module DA_table_3(table_in_3 , table_out_3);
input unsigned [15:0]table_in_3;
output [31:0]table_out_3;
wire  [31:0]LUT_3[65535:0]; 
wire [31:0]table_out_3; 
assign table_out_3 = LUT_3[table_in_3];
assign LUT_3[0] = 32'b00000000000000000000000000000000;
assign LUT_3[1] = 32'b00000000000000000110101011011101;
assign LUT_3[2] = 32'b00000000000000000010000111100100;
assign LUT_3[3] = 32'b00000000000000001000110011000001;
assign LUT_3[4] = 32'b11111111111111111101001101110110;
assign LUT_3[5] = 32'b00000000000000000011111001010011;
assign LUT_3[6] = 32'b11111111111111111111010101011010;
assign LUT_3[7] = 32'b00000000000000000110000000110111;
assign LUT_3[8] = 32'b00000000000000000101011001000110;
assign LUT_3[9] = 32'b00000000000000001100000100100011;
assign LUT_3[10] = 32'b00000000000000000111100000101010;
assign LUT_3[11] = 32'b00000000000000001110001100000111;
assign LUT_3[12] = 32'b00000000000000000010100110111100;
assign LUT_3[13] = 32'b00000000000000001001010010011001;
assign LUT_3[14] = 32'b00000000000000000100101110100000;
assign LUT_3[15] = 32'b00000000000000001011011001111101;
assign LUT_3[16] = 32'b00000000000000000011010011000011;
assign LUT_3[17] = 32'b00000000000000001001111110100000;
assign LUT_3[18] = 32'b00000000000000000101011010100111;
assign LUT_3[19] = 32'b00000000000000001100000110000100;
assign LUT_3[20] = 32'b00000000000000000000100000111001;
assign LUT_3[21] = 32'b00000000000000000111001100010110;
assign LUT_3[22] = 32'b00000000000000000010101000011101;
assign LUT_3[23] = 32'b00000000000000001001010011111010;
assign LUT_3[24] = 32'b00000000000000001000101100001001;
assign LUT_3[25] = 32'b00000000000000001111010111100110;
assign LUT_3[26] = 32'b00000000000000001010110011101101;
assign LUT_3[27] = 32'b00000000000000010001011111001010;
assign LUT_3[28] = 32'b00000000000000000101111001111111;
assign LUT_3[29] = 32'b00000000000000001100100101011100;
assign LUT_3[30] = 32'b00000000000000001000000001100011;
assign LUT_3[31] = 32'b00000000000000001110101101000000;
assign LUT_3[32] = 32'b00000000000000000001001110100000;
assign LUT_3[33] = 32'b00000000000000000111111001111101;
assign LUT_3[34] = 32'b00000000000000000011010110000100;
assign LUT_3[35] = 32'b00000000000000001010000001100001;
assign LUT_3[36] = 32'b11111111111111111110011100010110;
assign LUT_3[37] = 32'b00000000000000000101000111110011;
assign LUT_3[38] = 32'b00000000000000000000100011111010;
assign LUT_3[39] = 32'b00000000000000000111001111010111;
assign LUT_3[40] = 32'b00000000000000000110100111100110;
assign LUT_3[41] = 32'b00000000000000001101010011000011;
assign LUT_3[42] = 32'b00000000000000001000101111001010;
assign LUT_3[43] = 32'b00000000000000001111011010100111;
assign LUT_3[44] = 32'b00000000000000000011110101011100;
assign LUT_3[45] = 32'b00000000000000001010100000111001;
assign LUT_3[46] = 32'b00000000000000000101111101000000;
assign LUT_3[47] = 32'b00000000000000001100101000011101;
assign LUT_3[48] = 32'b00000000000000000100100001100011;
assign LUT_3[49] = 32'b00000000000000001011001101000000;
assign LUT_3[50] = 32'b00000000000000000110101001000111;
assign LUT_3[51] = 32'b00000000000000001101010100100100;
assign LUT_3[52] = 32'b00000000000000000001101111011001;
assign LUT_3[53] = 32'b00000000000000001000011010110110;
assign LUT_3[54] = 32'b00000000000000000011110110111101;
assign LUT_3[55] = 32'b00000000000000001010100010011010;
assign LUT_3[56] = 32'b00000000000000001001111010101001;
assign LUT_3[57] = 32'b00000000000000010000100110000110;
assign LUT_3[58] = 32'b00000000000000001100000010001101;
assign LUT_3[59] = 32'b00000000000000010010101101101010;
assign LUT_3[60] = 32'b00000000000000000111001000011111;
assign LUT_3[61] = 32'b00000000000000001101110011111100;
assign LUT_3[62] = 32'b00000000000000001001010000000011;
assign LUT_3[63] = 32'b00000000000000001111111011100000;
assign LUT_3[64] = 32'b11111111111111111111111000101011;
assign LUT_3[65] = 32'b00000000000000000110100100001000;
assign LUT_3[66] = 32'b00000000000000000010000000001111;
assign LUT_3[67] = 32'b00000000000000001000101011101100;
assign LUT_3[68] = 32'b11111111111111111101000110100001;
assign LUT_3[69] = 32'b00000000000000000011110001111110;
assign LUT_3[70] = 32'b11111111111111111111001110000101;
assign LUT_3[71] = 32'b00000000000000000101111001100010;
assign LUT_3[72] = 32'b00000000000000000101010001110001;
assign LUT_3[73] = 32'b00000000000000001011111101001110;
assign LUT_3[74] = 32'b00000000000000000111011001010101;
assign LUT_3[75] = 32'b00000000000000001110000100110010;
assign LUT_3[76] = 32'b00000000000000000010011111100111;
assign LUT_3[77] = 32'b00000000000000001001001011000100;
assign LUT_3[78] = 32'b00000000000000000100100111001011;
assign LUT_3[79] = 32'b00000000000000001011010010101000;
assign LUT_3[80] = 32'b00000000000000000011001011101110;
assign LUT_3[81] = 32'b00000000000000001001110111001011;
assign LUT_3[82] = 32'b00000000000000000101010011010010;
assign LUT_3[83] = 32'b00000000000000001011111110101111;
assign LUT_3[84] = 32'b00000000000000000000011001100100;
assign LUT_3[85] = 32'b00000000000000000111000101000001;
assign LUT_3[86] = 32'b00000000000000000010100001001000;
assign LUT_3[87] = 32'b00000000000000001001001100100101;
assign LUT_3[88] = 32'b00000000000000001000100100110100;
assign LUT_3[89] = 32'b00000000000000001111010000010001;
assign LUT_3[90] = 32'b00000000000000001010101100011000;
assign LUT_3[91] = 32'b00000000000000010001010111110101;
assign LUT_3[92] = 32'b00000000000000000101110010101010;
assign LUT_3[93] = 32'b00000000000000001100011110000111;
assign LUT_3[94] = 32'b00000000000000000111111010001110;
assign LUT_3[95] = 32'b00000000000000001110100101101011;
assign LUT_3[96] = 32'b00000000000000000001000111001011;
assign LUT_3[97] = 32'b00000000000000000111110010101000;
assign LUT_3[98] = 32'b00000000000000000011001110101111;
assign LUT_3[99] = 32'b00000000000000001001111010001100;
assign LUT_3[100] = 32'b11111111111111111110010101000001;
assign LUT_3[101] = 32'b00000000000000000101000000011110;
assign LUT_3[102] = 32'b00000000000000000000011100100101;
assign LUT_3[103] = 32'b00000000000000000111001000000010;
assign LUT_3[104] = 32'b00000000000000000110100000010001;
assign LUT_3[105] = 32'b00000000000000001101001011101110;
assign LUT_3[106] = 32'b00000000000000001000100111110101;
assign LUT_3[107] = 32'b00000000000000001111010011010010;
assign LUT_3[108] = 32'b00000000000000000011101110000111;
assign LUT_3[109] = 32'b00000000000000001010011001100100;
assign LUT_3[110] = 32'b00000000000000000101110101101011;
assign LUT_3[111] = 32'b00000000000000001100100001001000;
assign LUT_3[112] = 32'b00000000000000000100011010001110;
assign LUT_3[113] = 32'b00000000000000001011000101101011;
assign LUT_3[114] = 32'b00000000000000000110100001110010;
assign LUT_3[115] = 32'b00000000000000001101001101001111;
assign LUT_3[116] = 32'b00000000000000000001101000000100;
assign LUT_3[117] = 32'b00000000000000001000010011100001;
assign LUT_3[118] = 32'b00000000000000000011101111101000;
assign LUT_3[119] = 32'b00000000000000001010011011000101;
assign LUT_3[120] = 32'b00000000000000001001110011010100;
assign LUT_3[121] = 32'b00000000000000010000011110110001;
assign LUT_3[122] = 32'b00000000000000001011111010111000;
assign LUT_3[123] = 32'b00000000000000010010100110010101;
assign LUT_3[124] = 32'b00000000000000000111000001001010;
assign LUT_3[125] = 32'b00000000000000001101101100100111;
assign LUT_3[126] = 32'b00000000000000001001001000101110;
assign LUT_3[127] = 32'b00000000000000001111110100001011;
assign LUT_3[128] = 32'b00000000000000000010001010111110;
assign LUT_3[129] = 32'b00000000000000001000110110011011;
assign LUT_3[130] = 32'b00000000000000000100010010100010;
assign LUT_3[131] = 32'b00000000000000001010111101111111;
assign LUT_3[132] = 32'b11111111111111111111011000110100;
assign LUT_3[133] = 32'b00000000000000000110000100010001;
assign LUT_3[134] = 32'b00000000000000000001100000011000;
assign LUT_3[135] = 32'b00000000000000001000001011110101;
assign LUT_3[136] = 32'b00000000000000000111100100000100;
assign LUT_3[137] = 32'b00000000000000001110001111100001;
assign LUT_3[138] = 32'b00000000000000001001101011101000;
assign LUT_3[139] = 32'b00000000000000010000010111000101;
assign LUT_3[140] = 32'b00000000000000000100110001111010;
assign LUT_3[141] = 32'b00000000000000001011011101010111;
assign LUT_3[142] = 32'b00000000000000000110111001011110;
assign LUT_3[143] = 32'b00000000000000001101100100111011;
assign LUT_3[144] = 32'b00000000000000000101011110000001;
assign LUT_3[145] = 32'b00000000000000001100001001011110;
assign LUT_3[146] = 32'b00000000000000000111100101100101;
assign LUT_3[147] = 32'b00000000000000001110010001000010;
assign LUT_3[148] = 32'b00000000000000000010101011110111;
assign LUT_3[149] = 32'b00000000000000001001010111010100;
assign LUT_3[150] = 32'b00000000000000000100110011011011;
assign LUT_3[151] = 32'b00000000000000001011011110111000;
assign LUT_3[152] = 32'b00000000000000001010110111000111;
assign LUT_3[153] = 32'b00000000000000010001100010100100;
assign LUT_3[154] = 32'b00000000000000001100111110101011;
assign LUT_3[155] = 32'b00000000000000010011101010001000;
assign LUT_3[156] = 32'b00000000000000001000000100111101;
assign LUT_3[157] = 32'b00000000000000001110110000011010;
assign LUT_3[158] = 32'b00000000000000001010001100100001;
assign LUT_3[159] = 32'b00000000000000010000110111111110;
assign LUT_3[160] = 32'b00000000000000000011011001011110;
assign LUT_3[161] = 32'b00000000000000001010000100111011;
assign LUT_3[162] = 32'b00000000000000000101100001000010;
assign LUT_3[163] = 32'b00000000000000001100001100011111;
assign LUT_3[164] = 32'b00000000000000000000100111010100;
assign LUT_3[165] = 32'b00000000000000000111010010110001;
assign LUT_3[166] = 32'b00000000000000000010101110111000;
assign LUT_3[167] = 32'b00000000000000001001011010010101;
assign LUT_3[168] = 32'b00000000000000001000110010100100;
assign LUT_3[169] = 32'b00000000000000001111011110000001;
assign LUT_3[170] = 32'b00000000000000001010111010001000;
assign LUT_3[171] = 32'b00000000000000010001100101100101;
assign LUT_3[172] = 32'b00000000000000000110000000011010;
assign LUT_3[173] = 32'b00000000000000001100101011110111;
assign LUT_3[174] = 32'b00000000000000001000000111111110;
assign LUT_3[175] = 32'b00000000000000001110110011011011;
assign LUT_3[176] = 32'b00000000000000000110101100100001;
assign LUT_3[177] = 32'b00000000000000001101010111111110;
assign LUT_3[178] = 32'b00000000000000001000110100000101;
assign LUT_3[179] = 32'b00000000000000001111011111100010;
assign LUT_3[180] = 32'b00000000000000000011111010010111;
assign LUT_3[181] = 32'b00000000000000001010100101110100;
assign LUT_3[182] = 32'b00000000000000000110000001111011;
assign LUT_3[183] = 32'b00000000000000001100101101011000;
assign LUT_3[184] = 32'b00000000000000001100000101100111;
assign LUT_3[185] = 32'b00000000000000010010110001000100;
assign LUT_3[186] = 32'b00000000000000001110001101001011;
assign LUT_3[187] = 32'b00000000000000010100111000101000;
assign LUT_3[188] = 32'b00000000000000001001010011011101;
assign LUT_3[189] = 32'b00000000000000001111111110111010;
assign LUT_3[190] = 32'b00000000000000001011011011000001;
assign LUT_3[191] = 32'b00000000000000010010000110011110;
assign LUT_3[192] = 32'b00000000000000000010000011101001;
assign LUT_3[193] = 32'b00000000000000001000101111000110;
assign LUT_3[194] = 32'b00000000000000000100001011001101;
assign LUT_3[195] = 32'b00000000000000001010110110101010;
assign LUT_3[196] = 32'b11111111111111111111010001011111;
assign LUT_3[197] = 32'b00000000000000000101111100111100;
assign LUT_3[198] = 32'b00000000000000000001011001000011;
assign LUT_3[199] = 32'b00000000000000001000000100100000;
assign LUT_3[200] = 32'b00000000000000000111011100101111;
assign LUT_3[201] = 32'b00000000000000001110001000001100;
assign LUT_3[202] = 32'b00000000000000001001100100010011;
assign LUT_3[203] = 32'b00000000000000010000001111110000;
assign LUT_3[204] = 32'b00000000000000000100101010100101;
assign LUT_3[205] = 32'b00000000000000001011010110000010;
assign LUT_3[206] = 32'b00000000000000000110110010001001;
assign LUT_3[207] = 32'b00000000000000001101011101100110;
assign LUT_3[208] = 32'b00000000000000000101010110101100;
assign LUT_3[209] = 32'b00000000000000001100000010001001;
assign LUT_3[210] = 32'b00000000000000000111011110010000;
assign LUT_3[211] = 32'b00000000000000001110001001101101;
assign LUT_3[212] = 32'b00000000000000000010100100100010;
assign LUT_3[213] = 32'b00000000000000001001001111111111;
assign LUT_3[214] = 32'b00000000000000000100101100000110;
assign LUT_3[215] = 32'b00000000000000001011010111100011;
assign LUT_3[216] = 32'b00000000000000001010101111110010;
assign LUT_3[217] = 32'b00000000000000010001011011001111;
assign LUT_3[218] = 32'b00000000000000001100110111010110;
assign LUT_3[219] = 32'b00000000000000010011100010110011;
assign LUT_3[220] = 32'b00000000000000000111111101101000;
assign LUT_3[221] = 32'b00000000000000001110101001000101;
assign LUT_3[222] = 32'b00000000000000001010000101001100;
assign LUT_3[223] = 32'b00000000000000010000110000101001;
assign LUT_3[224] = 32'b00000000000000000011010010001001;
assign LUT_3[225] = 32'b00000000000000001001111101100110;
assign LUT_3[226] = 32'b00000000000000000101011001101101;
assign LUT_3[227] = 32'b00000000000000001100000101001010;
assign LUT_3[228] = 32'b00000000000000000000011111111111;
assign LUT_3[229] = 32'b00000000000000000111001011011100;
assign LUT_3[230] = 32'b00000000000000000010100111100011;
assign LUT_3[231] = 32'b00000000000000001001010011000000;
assign LUT_3[232] = 32'b00000000000000001000101011001111;
assign LUT_3[233] = 32'b00000000000000001111010110101100;
assign LUT_3[234] = 32'b00000000000000001010110010110011;
assign LUT_3[235] = 32'b00000000000000010001011110010000;
assign LUT_3[236] = 32'b00000000000000000101111001000101;
assign LUT_3[237] = 32'b00000000000000001100100100100010;
assign LUT_3[238] = 32'b00000000000000001000000000101001;
assign LUT_3[239] = 32'b00000000000000001110101100000110;
assign LUT_3[240] = 32'b00000000000000000110100101001100;
assign LUT_3[241] = 32'b00000000000000001101010000101001;
assign LUT_3[242] = 32'b00000000000000001000101100110000;
assign LUT_3[243] = 32'b00000000000000001111011000001101;
assign LUT_3[244] = 32'b00000000000000000011110011000010;
assign LUT_3[245] = 32'b00000000000000001010011110011111;
assign LUT_3[246] = 32'b00000000000000000101111010100110;
assign LUT_3[247] = 32'b00000000000000001100100110000011;
assign LUT_3[248] = 32'b00000000000000001011111110010010;
assign LUT_3[249] = 32'b00000000000000010010101001101111;
assign LUT_3[250] = 32'b00000000000000001110000101110110;
assign LUT_3[251] = 32'b00000000000000010100110001010011;
assign LUT_3[252] = 32'b00000000000000001001001100001000;
assign LUT_3[253] = 32'b00000000000000001111110111100101;
assign LUT_3[254] = 32'b00000000000000001011010011101100;
assign LUT_3[255] = 32'b00000000000000010001111111001001;
assign LUT_3[256] = 32'b11111111111111111100001111100001;
assign LUT_3[257] = 32'b00000000000000000010111010111110;
assign LUT_3[258] = 32'b11111111111111111110010111000101;
assign LUT_3[259] = 32'b00000000000000000101000010100010;
assign LUT_3[260] = 32'b11111111111111111001011101010111;
assign LUT_3[261] = 32'b00000000000000000000001000110100;
assign LUT_3[262] = 32'b11111111111111111011100100111011;
assign LUT_3[263] = 32'b00000000000000000010010000011000;
assign LUT_3[264] = 32'b00000000000000000001101000100111;
assign LUT_3[265] = 32'b00000000000000001000010100000100;
assign LUT_3[266] = 32'b00000000000000000011110000001011;
assign LUT_3[267] = 32'b00000000000000001010011011101000;
assign LUT_3[268] = 32'b11111111111111111110110110011101;
assign LUT_3[269] = 32'b00000000000000000101100001111010;
assign LUT_3[270] = 32'b00000000000000000000111110000001;
assign LUT_3[271] = 32'b00000000000000000111101001011110;
assign LUT_3[272] = 32'b11111111111111111111100010100100;
assign LUT_3[273] = 32'b00000000000000000110001110000001;
assign LUT_3[274] = 32'b00000000000000000001101010001000;
assign LUT_3[275] = 32'b00000000000000001000010101100101;
assign LUT_3[276] = 32'b11111111111111111100110000011010;
assign LUT_3[277] = 32'b00000000000000000011011011110111;
assign LUT_3[278] = 32'b11111111111111111110110111111110;
assign LUT_3[279] = 32'b00000000000000000101100011011011;
assign LUT_3[280] = 32'b00000000000000000100111011101010;
assign LUT_3[281] = 32'b00000000000000001011100111000111;
assign LUT_3[282] = 32'b00000000000000000111000011001110;
assign LUT_3[283] = 32'b00000000000000001101101110101011;
assign LUT_3[284] = 32'b00000000000000000010001001100000;
assign LUT_3[285] = 32'b00000000000000001000110100111101;
assign LUT_3[286] = 32'b00000000000000000100010001000100;
assign LUT_3[287] = 32'b00000000000000001010111100100001;
assign LUT_3[288] = 32'b11111111111111111101011110000001;
assign LUT_3[289] = 32'b00000000000000000100001001011110;
assign LUT_3[290] = 32'b11111111111111111111100101100101;
assign LUT_3[291] = 32'b00000000000000000110010001000010;
assign LUT_3[292] = 32'b11111111111111111010101011110111;
assign LUT_3[293] = 32'b00000000000000000001010111010100;
assign LUT_3[294] = 32'b11111111111111111100110011011011;
assign LUT_3[295] = 32'b00000000000000000011011110111000;
assign LUT_3[296] = 32'b00000000000000000010110111000111;
assign LUT_3[297] = 32'b00000000000000001001100010100100;
assign LUT_3[298] = 32'b00000000000000000100111110101011;
assign LUT_3[299] = 32'b00000000000000001011101010001000;
assign LUT_3[300] = 32'b00000000000000000000000100111101;
assign LUT_3[301] = 32'b00000000000000000110110000011010;
assign LUT_3[302] = 32'b00000000000000000010001100100001;
assign LUT_3[303] = 32'b00000000000000001000110111111110;
assign LUT_3[304] = 32'b00000000000000000000110001000100;
assign LUT_3[305] = 32'b00000000000000000111011100100001;
assign LUT_3[306] = 32'b00000000000000000010111000101000;
assign LUT_3[307] = 32'b00000000000000001001100100000101;
assign LUT_3[308] = 32'b11111111111111111101111110111010;
assign LUT_3[309] = 32'b00000000000000000100101010010111;
assign LUT_3[310] = 32'b00000000000000000000000110011110;
assign LUT_3[311] = 32'b00000000000000000110110001111011;
assign LUT_3[312] = 32'b00000000000000000110001010001010;
assign LUT_3[313] = 32'b00000000000000001100110101100111;
assign LUT_3[314] = 32'b00000000000000001000010001101110;
assign LUT_3[315] = 32'b00000000000000001110111101001011;
assign LUT_3[316] = 32'b00000000000000000011011000000000;
assign LUT_3[317] = 32'b00000000000000001010000011011101;
assign LUT_3[318] = 32'b00000000000000000101011111100100;
assign LUT_3[319] = 32'b00000000000000001100001011000001;
assign LUT_3[320] = 32'b11111111111111111100001000001100;
assign LUT_3[321] = 32'b00000000000000000010110011101001;
assign LUT_3[322] = 32'b11111111111111111110001111110000;
assign LUT_3[323] = 32'b00000000000000000100111011001101;
assign LUT_3[324] = 32'b11111111111111111001010110000010;
assign LUT_3[325] = 32'b00000000000000000000000001011111;
assign LUT_3[326] = 32'b11111111111111111011011101100110;
assign LUT_3[327] = 32'b00000000000000000010001001000011;
assign LUT_3[328] = 32'b00000000000000000001100001010010;
assign LUT_3[329] = 32'b00000000000000001000001100101111;
assign LUT_3[330] = 32'b00000000000000000011101000110110;
assign LUT_3[331] = 32'b00000000000000001010010100010011;
assign LUT_3[332] = 32'b11111111111111111110101111001000;
assign LUT_3[333] = 32'b00000000000000000101011010100101;
assign LUT_3[334] = 32'b00000000000000000000110110101100;
assign LUT_3[335] = 32'b00000000000000000111100010001001;
assign LUT_3[336] = 32'b11111111111111111111011011001111;
assign LUT_3[337] = 32'b00000000000000000110000110101100;
assign LUT_3[338] = 32'b00000000000000000001100010110011;
assign LUT_3[339] = 32'b00000000000000001000001110010000;
assign LUT_3[340] = 32'b11111111111111111100101001000101;
assign LUT_3[341] = 32'b00000000000000000011010100100010;
assign LUT_3[342] = 32'b11111111111111111110110000101001;
assign LUT_3[343] = 32'b00000000000000000101011100000110;
assign LUT_3[344] = 32'b00000000000000000100110100010101;
assign LUT_3[345] = 32'b00000000000000001011011111110010;
assign LUT_3[346] = 32'b00000000000000000110111011111001;
assign LUT_3[347] = 32'b00000000000000001101100111010110;
assign LUT_3[348] = 32'b00000000000000000010000010001011;
assign LUT_3[349] = 32'b00000000000000001000101101101000;
assign LUT_3[350] = 32'b00000000000000000100001001101111;
assign LUT_3[351] = 32'b00000000000000001010110101001100;
assign LUT_3[352] = 32'b11111111111111111101010110101100;
assign LUT_3[353] = 32'b00000000000000000100000010001001;
assign LUT_3[354] = 32'b11111111111111111111011110010000;
assign LUT_3[355] = 32'b00000000000000000110001001101101;
assign LUT_3[356] = 32'b11111111111111111010100100100010;
assign LUT_3[357] = 32'b00000000000000000001001111111111;
assign LUT_3[358] = 32'b11111111111111111100101100000110;
assign LUT_3[359] = 32'b00000000000000000011010111100011;
assign LUT_3[360] = 32'b00000000000000000010101111110010;
assign LUT_3[361] = 32'b00000000000000001001011011001111;
assign LUT_3[362] = 32'b00000000000000000100110111010110;
assign LUT_3[363] = 32'b00000000000000001011100010110011;
assign LUT_3[364] = 32'b11111111111111111111111101101000;
assign LUT_3[365] = 32'b00000000000000000110101001000101;
assign LUT_3[366] = 32'b00000000000000000010000101001100;
assign LUT_3[367] = 32'b00000000000000001000110000101001;
assign LUT_3[368] = 32'b00000000000000000000101001101111;
assign LUT_3[369] = 32'b00000000000000000111010101001100;
assign LUT_3[370] = 32'b00000000000000000010110001010011;
assign LUT_3[371] = 32'b00000000000000001001011100110000;
assign LUT_3[372] = 32'b11111111111111111101110111100101;
assign LUT_3[373] = 32'b00000000000000000100100011000010;
assign LUT_3[374] = 32'b11111111111111111111111111001001;
assign LUT_3[375] = 32'b00000000000000000110101010100110;
assign LUT_3[376] = 32'b00000000000000000110000010110101;
assign LUT_3[377] = 32'b00000000000000001100101110010010;
assign LUT_3[378] = 32'b00000000000000001000001010011001;
assign LUT_3[379] = 32'b00000000000000001110110101110110;
assign LUT_3[380] = 32'b00000000000000000011010000101011;
assign LUT_3[381] = 32'b00000000000000001001111100001000;
assign LUT_3[382] = 32'b00000000000000000101011000001111;
assign LUT_3[383] = 32'b00000000000000001100000011101100;
assign LUT_3[384] = 32'b11111111111111111110011010011111;
assign LUT_3[385] = 32'b00000000000000000101000101111100;
assign LUT_3[386] = 32'b00000000000000000000100010000011;
assign LUT_3[387] = 32'b00000000000000000111001101100000;
assign LUT_3[388] = 32'b11111111111111111011101000010101;
assign LUT_3[389] = 32'b00000000000000000010010011110010;
assign LUT_3[390] = 32'b11111111111111111101101111111001;
assign LUT_3[391] = 32'b00000000000000000100011011010110;
assign LUT_3[392] = 32'b00000000000000000011110011100101;
assign LUT_3[393] = 32'b00000000000000001010011111000010;
assign LUT_3[394] = 32'b00000000000000000101111011001001;
assign LUT_3[395] = 32'b00000000000000001100100110100110;
assign LUT_3[396] = 32'b00000000000000000001000001011011;
assign LUT_3[397] = 32'b00000000000000000111101100111000;
assign LUT_3[398] = 32'b00000000000000000011001000111111;
assign LUT_3[399] = 32'b00000000000000001001110100011100;
assign LUT_3[400] = 32'b00000000000000000001101101100010;
assign LUT_3[401] = 32'b00000000000000001000011000111111;
assign LUT_3[402] = 32'b00000000000000000011110101000110;
assign LUT_3[403] = 32'b00000000000000001010100000100011;
assign LUT_3[404] = 32'b11111111111111111110111011011000;
assign LUT_3[405] = 32'b00000000000000000101100110110101;
assign LUT_3[406] = 32'b00000000000000000001000010111100;
assign LUT_3[407] = 32'b00000000000000000111101110011001;
assign LUT_3[408] = 32'b00000000000000000111000110101000;
assign LUT_3[409] = 32'b00000000000000001101110010000101;
assign LUT_3[410] = 32'b00000000000000001001001110001100;
assign LUT_3[411] = 32'b00000000000000001111111001101001;
assign LUT_3[412] = 32'b00000000000000000100010100011110;
assign LUT_3[413] = 32'b00000000000000001010111111111011;
assign LUT_3[414] = 32'b00000000000000000110011100000010;
assign LUT_3[415] = 32'b00000000000000001101000111011111;
assign LUT_3[416] = 32'b11111111111111111111101000111111;
assign LUT_3[417] = 32'b00000000000000000110010100011100;
assign LUT_3[418] = 32'b00000000000000000001110000100011;
assign LUT_3[419] = 32'b00000000000000001000011100000000;
assign LUT_3[420] = 32'b11111111111111111100110110110101;
assign LUT_3[421] = 32'b00000000000000000011100010010010;
assign LUT_3[422] = 32'b11111111111111111110111110011001;
assign LUT_3[423] = 32'b00000000000000000101101001110110;
assign LUT_3[424] = 32'b00000000000000000101000010000101;
assign LUT_3[425] = 32'b00000000000000001011101101100010;
assign LUT_3[426] = 32'b00000000000000000111001001101001;
assign LUT_3[427] = 32'b00000000000000001101110101000110;
assign LUT_3[428] = 32'b00000000000000000010001111111011;
assign LUT_3[429] = 32'b00000000000000001000111011011000;
assign LUT_3[430] = 32'b00000000000000000100010111011111;
assign LUT_3[431] = 32'b00000000000000001011000010111100;
assign LUT_3[432] = 32'b00000000000000000010111100000010;
assign LUT_3[433] = 32'b00000000000000001001100111011111;
assign LUT_3[434] = 32'b00000000000000000101000011100110;
assign LUT_3[435] = 32'b00000000000000001011101111000011;
assign LUT_3[436] = 32'b00000000000000000000001001111000;
assign LUT_3[437] = 32'b00000000000000000110110101010101;
assign LUT_3[438] = 32'b00000000000000000010010001011100;
assign LUT_3[439] = 32'b00000000000000001000111100111001;
assign LUT_3[440] = 32'b00000000000000001000010101001000;
assign LUT_3[441] = 32'b00000000000000001111000000100101;
assign LUT_3[442] = 32'b00000000000000001010011100101100;
assign LUT_3[443] = 32'b00000000000000010001001000001001;
assign LUT_3[444] = 32'b00000000000000000101100010111110;
assign LUT_3[445] = 32'b00000000000000001100001110011011;
assign LUT_3[446] = 32'b00000000000000000111101010100010;
assign LUT_3[447] = 32'b00000000000000001110010101111111;
assign LUT_3[448] = 32'b11111111111111111110010011001010;
assign LUT_3[449] = 32'b00000000000000000100111110100111;
assign LUT_3[450] = 32'b00000000000000000000011010101110;
assign LUT_3[451] = 32'b00000000000000000111000110001011;
assign LUT_3[452] = 32'b11111111111111111011100001000000;
assign LUT_3[453] = 32'b00000000000000000010001100011101;
assign LUT_3[454] = 32'b11111111111111111101101000100100;
assign LUT_3[455] = 32'b00000000000000000100010100000001;
assign LUT_3[456] = 32'b00000000000000000011101100010000;
assign LUT_3[457] = 32'b00000000000000001010010111101101;
assign LUT_3[458] = 32'b00000000000000000101110011110100;
assign LUT_3[459] = 32'b00000000000000001100011111010001;
assign LUT_3[460] = 32'b00000000000000000000111010000110;
assign LUT_3[461] = 32'b00000000000000000111100101100011;
assign LUT_3[462] = 32'b00000000000000000011000001101010;
assign LUT_3[463] = 32'b00000000000000001001101101000111;
assign LUT_3[464] = 32'b00000000000000000001100110001101;
assign LUT_3[465] = 32'b00000000000000001000010001101010;
assign LUT_3[466] = 32'b00000000000000000011101101110001;
assign LUT_3[467] = 32'b00000000000000001010011001001110;
assign LUT_3[468] = 32'b11111111111111111110110100000011;
assign LUT_3[469] = 32'b00000000000000000101011111100000;
assign LUT_3[470] = 32'b00000000000000000000111011100111;
assign LUT_3[471] = 32'b00000000000000000111100111000100;
assign LUT_3[472] = 32'b00000000000000000110111111010011;
assign LUT_3[473] = 32'b00000000000000001101101010110000;
assign LUT_3[474] = 32'b00000000000000001001000110110111;
assign LUT_3[475] = 32'b00000000000000001111110010010100;
assign LUT_3[476] = 32'b00000000000000000100001101001001;
assign LUT_3[477] = 32'b00000000000000001010111000100110;
assign LUT_3[478] = 32'b00000000000000000110010100101101;
assign LUT_3[479] = 32'b00000000000000001101000000001010;
assign LUT_3[480] = 32'b11111111111111111111100001101010;
assign LUT_3[481] = 32'b00000000000000000110001101000111;
assign LUT_3[482] = 32'b00000000000000000001101001001110;
assign LUT_3[483] = 32'b00000000000000001000010100101011;
assign LUT_3[484] = 32'b11111111111111111100101111100000;
assign LUT_3[485] = 32'b00000000000000000011011010111101;
assign LUT_3[486] = 32'b11111111111111111110110111000100;
assign LUT_3[487] = 32'b00000000000000000101100010100001;
assign LUT_3[488] = 32'b00000000000000000100111010110000;
assign LUT_3[489] = 32'b00000000000000001011100110001101;
assign LUT_3[490] = 32'b00000000000000000111000010010100;
assign LUT_3[491] = 32'b00000000000000001101101101110001;
assign LUT_3[492] = 32'b00000000000000000010001000100110;
assign LUT_3[493] = 32'b00000000000000001000110100000011;
assign LUT_3[494] = 32'b00000000000000000100010000001010;
assign LUT_3[495] = 32'b00000000000000001010111011100111;
assign LUT_3[496] = 32'b00000000000000000010110100101101;
assign LUT_3[497] = 32'b00000000000000001001100000001010;
assign LUT_3[498] = 32'b00000000000000000100111100010001;
assign LUT_3[499] = 32'b00000000000000001011100111101110;
assign LUT_3[500] = 32'b00000000000000000000000010100011;
assign LUT_3[501] = 32'b00000000000000000110101110000000;
assign LUT_3[502] = 32'b00000000000000000010001010000111;
assign LUT_3[503] = 32'b00000000000000001000110101100100;
assign LUT_3[504] = 32'b00000000000000001000001101110011;
assign LUT_3[505] = 32'b00000000000000001110111001010000;
assign LUT_3[506] = 32'b00000000000000001010010101010111;
assign LUT_3[507] = 32'b00000000000000010001000000110100;
assign LUT_3[508] = 32'b00000000000000000101011011101001;
assign LUT_3[509] = 32'b00000000000000001100000111000110;
assign LUT_3[510] = 32'b00000000000000000111100011001101;
assign LUT_3[511] = 32'b00000000000000001110001110101010;
assign LUT_3[512] = 32'b00000000000000000011010101001100;
assign LUT_3[513] = 32'b00000000000000001010000000101001;
assign LUT_3[514] = 32'b00000000000000000101011100110000;
assign LUT_3[515] = 32'b00000000000000001100001000001101;
assign LUT_3[516] = 32'b00000000000000000000100011000010;
assign LUT_3[517] = 32'b00000000000000000111001110011111;
assign LUT_3[518] = 32'b00000000000000000010101010100110;
assign LUT_3[519] = 32'b00000000000000001001010110000011;
assign LUT_3[520] = 32'b00000000000000001000101110010010;
assign LUT_3[521] = 32'b00000000000000001111011001101111;
assign LUT_3[522] = 32'b00000000000000001010110101110110;
assign LUT_3[523] = 32'b00000000000000010001100001010011;
assign LUT_3[524] = 32'b00000000000000000101111100001000;
assign LUT_3[525] = 32'b00000000000000001100100111100101;
assign LUT_3[526] = 32'b00000000000000001000000011101100;
assign LUT_3[527] = 32'b00000000000000001110101111001001;
assign LUT_3[528] = 32'b00000000000000000110101000001111;
assign LUT_3[529] = 32'b00000000000000001101010011101100;
assign LUT_3[530] = 32'b00000000000000001000101111110011;
assign LUT_3[531] = 32'b00000000000000001111011011010000;
assign LUT_3[532] = 32'b00000000000000000011110110000101;
assign LUT_3[533] = 32'b00000000000000001010100001100010;
assign LUT_3[534] = 32'b00000000000000000101111101101001;
assign LUT_3[535] = 32'b00000000000000001100101001000110;
assign LUT_3[536] = 32'b00000000000000001100000001010101;
assign LUT_3[537] = 32'b00000000000000010010101100110010;
assign LUT_3[538] = 32'b00000000000000001110001000111001;
assign LUT_3[539] = 32'b00000000000000010100110100010110;
assign LUT_3[540] = 32'b00000000000000001001001111001011;
assign LUT_3[541] = 32'b00000000000000001111111010101000;
assign LUT_3[542] = 32'b00000000000000001011010110101111;
assign LUT_3[543] = 32'b00000000000000010010000010001100;
assign LUT_3[544] = 32'b00000000000000000100100011101100;
assign LUT_3[545] = 32'b00000000000000001011001111001001;
assign LUT_3[546] = 32'b00000000000000000110101011010000;
assign LUT_3[547] = 32'b00000000000000001101010110101101;
assign LUT_3[548] = 32'b00000000000000000001110001100010;
assign LUT_3[549] = 32'b00000000000000001000011100111111;
assign LUT_3[550] = 32'b00000000000000000011111001000110;
assign LUT_3[551] = 32'b00000000000000001010100100100011;
assign LUT_3[552] = 32'b00000000000000001001111100110010;
assign LUT_3[553] = 32'b00000000000000010000101000001111;
assign LUT_3[554] = 32'b00000000000000001100000100010110;
assign LUT_3[555] = 32'b00000000000000010010101111110011;
assign LUT_3[556] = 32'b00000000000000000111001010101000;
assign LUT_3[557] = 32'b00000000000000001101110110000101;
assign LUT_3[558] = 32'b00000000000000001001010010001100;
assign LUT_3[559] = 32'b00000000000000001111111101101001;
assign LUT_3[560] = 32'b00000000000000000111110110101111;
assign LUT_3[561] = 32'b00000000000000001110100010001100;
assign LUT_3[562] = 32'b00000000000000001001111110010011;
assign LUT_3[563] = 32'b00000000000000010000101001110000;
assign LUT_3[564] = 32'b00000000000000000101000100100101;
assign LUT_3[565] = 32'b00000000000000001011110000000010;
assign LUT_3[566] = 32'b00000000000000000111001100001001;
assign LUT_3[567] = 32'b00000000000000001101110111100110;
assign LUT_3[568] = 32'b00000000000000001101001111110101;
assign LUT_3[569] = 32'b00000000000000010011111011010010;
assign LUT_3[570] = 32'b00000000000000001111010111011001;
assign LUT_3[571] = 32'b00000000000000010110000010110110;
assign LUT_3[572] = 32'b00000000000000001010011101101011;
assign LUT_3[573] = 32'b00000000000000010001001001001000;
assign LUT_3[574] = 32'b00000000000000001100100101001111;
assign LUT_3[575] = 32'b00000000000000010011010000101100;
assign LUT_3[576] = 32'b00000000000000000011001101110111;
assign LUT_3[577] = 32'b00000000000000001001111001010100;
assign LUT_3[578] = 32'b00000000000000000101010101011011;
assign LUT_3[579] = 32'b00000000000000001100000000111000;
assign LUT_3[580] = 32'b00000000000000000000011011101101;
assign LUT_3[581] = 32'b00000000000000000111000111001010;
assign LUT_3[582] = 32'b00000000000000000010100011010001;
assign LUT_3[583] = 32'b00000000000000001001001110101110;
assign LUT_3[584] = 32'b00000000000000001000100110111101;
assign LUT_3[585] = 32'b00000000000000001111010010011010;
assign LUT_3[586] = 32'b00000000000000001010101110100001;
assign LUT_3[587] = 32'b00000000000000010001011001111110;
assign LUT_3[588] = 32'b00000000000000000101110100110011;
assign LUT_3[589] = 32'b00000000000000001100100000010000;
assign LUT_3[590] = 32'b00000000000000000111111100010111;
assign LUT_3[591] = 32'b00000000000000001110100111110100;
assign LUT_3[592] = 32'b00000000000000000110100000111010;
assign LUT_3[593] = 32'b00000000000000001101001100010111;
assign LUT_3[594] = 32'b00000000000000001000101000011110;
assign LUT_3[595] = 32'b00000000000000001111010011111011;
assign LUT_3[596] = 32'b00000000000000000011101110110000;
assign LUT_3[597] = 32'b00000000000000001010011010001101;
assign LUT_3[598] = 32'b00000000000000000101110110010100;
assign LUT_3[599] = 32'b00000000000000001100100001110001;
assign LUT_3[600] = 32'b00000000000000001011111010000000;
assign LUT_3[601] = 32'b00000000000000010010100101011101;
assign LUT_3[602] = 32'b00000000000000001110000001100100;
assign LUT_3[603] = 32'b00000000000000010100101101000001;
assign LUT_3[604] = 32'b00000000000000001001000111110110;
assign LUT_3[605] = 32'b00000000000000001111110011010011;
assign LUT_3[606] = 32'b00000000000000001011001111011010;
assign LUT_3[607] = 32'b00000000000000010001111010110111;
assign LUT_3[608] = 32'b00000000000000000100011100010111;
assign LUT_3[609] = 32'b00000000000000001011000111110100;
assign LUT_3[610] = 32'b00000000000000000110100011111011;
assign LUT_3[611] = 32'b00000000000000001101001111011000;
assign LUT_3[612] = 32'b00000000000000000001101010001101;
assign LUT_3[613] = 32'b00000000000000001000010101101010;
assign LUT_3[614] = 32'b00000000000000000011110001110001;
assign LUT_3[615] = 32'b00000000000000001010011101001110;
assign LUT_3[616] = 32'b00000000000000001001110101011101;
assign LUT_3[617] = 32'b00000000000000010000100000111010;
assign LUT_3[618] = 32'b00000000000000001011111101000001;
assign LUT_3[619] = 32'b00000000000000010010101000011110;
assign LUT_3[620] = 32'b00000000000000000111000011010011;
assign LUT_3[621] = 32'b00000000000000001101101110110000;
assign LUT_3[622] = 32'b00000000000000001001001010110111;
assign LUT_3[623] = 32'b00000000000000001111110110010100;
assign LUT_3[624] = 32'b00000000000000000111101111011010;
assign LUT_3[625] = 32'b00000000000000001110011010110111;
assign LUT_3[626] = 32'b00000000000000001001110110111110;
assign LUT_3[627] = 32'b00000000000000010000100010011011;
assign LUT_3[628] = 32'b00000000000000000100111101010000;
assign LUT_3[629] = 32'b00000000000000001011101000101101;
assign LUT_3[630] = 32'b00000000000000000111000100110100;
assign LUT_3[631] = 32'b00000000000000001101110000010001;
assign LUT_3[632] = 32'b00000000000000001101001000100000;
assign LUT_3[633] = 32'b00000000000000010011110011111101;
assign LUT_3[634] = 32'b00000000000000001111010000000100;
assign LUT_3[635] = 32'b00000000000000010101111011100001;
assign LUT_3[636] = 32'b00000000000000001010010110010110;
assign LUT_3[637] = 32'b00000000000000010001000001110011;
assign LUT_3[638] = 32'b00000000000000001100011101111010;
assign LUT_3[639] = 32'b00000000000000010011001001010111;
assign LUT_3[640] = 32'b00000000000000000101100000001010;
assign LUT_3[641] = 32'b00000000000000001100001011100111;
assign LUT_3[642] = 32'b00000000000000000111100111101110;
assign LUT_3[643] = 32'b00000000000000001110010011001011;
assign LUT_3[644] = 32'b00000000000000000010101110000000;
assign LUT_3[645] = 32'b00000000000000001001011001011101;
assign LUT_3[646] = 32'b00000000000000000100110101100100;
assign LUT_3[647] = 32'b00000000000000001011100001000001;
assign LUT_3[648] = 32'b00000000000000001010111001010000;
assign LUT_3[649] = 32'b00000000000000010001100100101101;
assign LUT_3[650] = 32'b00000000000000001101000000110100;
assign LUT_3[651] = 32'b00000000000000010011101100010001;
assign LUT_3[652] = 32'b00000000000000001000000111000110;
assign LUT_3[653] = 32'b00000000000000001110110010100011;
assign LUT_3[654] = 32'b00000000000000001010001110101010;
assign LUT_3[655] = 32'b00000000000000010000111010000111;
assign LUT_3[656] = 32'b00000000000000001000110011001101;
assign LUT_3[657] = 32'b00000000000000001111011110101010;
assign LUT_3[658] = 32'b00000000000000001010111010110001;
assign LUT_3[659] = 32'b00000000000000010001100110001110;
assign LUT_3[660] = 32'b00000000000000000110000001000011;
assign LUT_3[661] = 32'b00000000000000001100101100100000;
assign LUT_3[662] = 32'b00000000000000001000001000100111;
assign LUT_3[663] = 32'b00000000000000001110110100000100;
assign LUT_3[664] = 32'b00000000000000001110001100010011;
assign LUT_3[665] = 32'b00000000000000010100110111110000;
assign LUT_3[666] = 32'b00000000000000010000010011110111;
assign LUT_3[667] = 32'b00000000000000010110111111010100;
assign LUT_3[668] = 32'b00000000000000001011011010001001;
assign LUT_3[669] = 32'b00000000000000010010000101100110;
assign LUT_3[670] = 32'b00000000000000001101100001101101;
assign LUT_3[671] = 32'b00000000000000010100001101001010;
assign LUT_3[672] = 32'b00000000000000000110101110101010;
assign LUT_3[673] = 32'b00000000000000001101011010000111;
assign LUT_3[674] = 32'b00000000000000001000110110001110;
assign LUT_3[675] = 32'b00000000000000001111100001101011;
assign LUT_3[676] = 32'b00000000000000000011111100100000;
assign LUT_3[677] = 32'b00000000000000001010100111111101;
assign LUT_3[678] = 32'b00000000000000000110000100000100;
assign LUT_3[679] = 32'b00000000000000001100101111100001;
assign LUT_3[680] = 32'b00000000000000001100000111110000;
assign LUT_3[681] = 32'b00000000000000010010110011001101;
assign LUT_3[682] = 32'b00000000000000001110001111010100;
assign LUT_3[683] = 32'b00000000000000010100111010110001;
assign LUT_3[684] = 32'b00000000000000001001010101100110;
assign LUT_3[685] = 32'b00000000000000010000000001000011;
assign LUT_3[686] = 32'b00000000000000001011011101001010;
assign LUT_3[687] = 32'b00000000000000010010001000100111;
assign LUT_3[688] = 32'b00000000000000001010000001101101;
assign LUT_3[689] = 32'b00000000000000010000101101001010;
assign LUT_3[690] = 32'b00000000000000001100001001010001;
assign LUT_3[691] = 32'b00000000000000010010110100101110;
assign LUT_3[692] = 32'b00000000000000000111001111100011;
assign LUT_3[693] = 32'b00000000000000001101111011000000;
assign LUT_3[694] = 32'b00000000000000001001010111000111;
assign LUT_3[695] = 32'b00000000000000010000000010100100;
assign LUT_3[696] = 32'b00000000000000001111011010110011;
assign LUT_3[697] = 32'b00000000000000010110000110010000;
assign LUT_3[698] = 32'b00000000000000010001100010010111;
assign LUT_3[699] = 32'b00000000000000011000001101110100;
assign LUT_3[700] = 32'b00000000000000001100101000101001;
assign LUT_3[701] = 32'b00000000000000010011010100000110;
assign LUT_3[702] = 32'b00000000000000001110110000001101;
assign LUT_3[703] = 32'b00000000000000010101011011101010;
assign LUT_3[704] = 32'b00000000000000000101011000110101;
assign LUT_3[705] = 32'b00000000000000001100000100010010;
assign LUT_3[706] = 32'b00000000000000000111100000011001;
assign LUT_3[707] = 32'b00000000000000001110001011110110;
assign LUT_3[708] = 32'b00000000000000000010100110101011;
assign LUT_3[709] = 32'b00000000000000001001010010001000;
assign LUT_3[710] = 32'b00000000000000000100101110001111;
assign LUT_3[711] = 32'b00000000000000001011011001101100;
assign LUT_3[712] = 32'b00000000000000001010110001111011;
assign LUT_3[713] = 32'b00000000000000010001011101011000;
assign LUT_3[714] = 32'b00000000000000001100111001011111;
assign LUT_3[715] = 32'b00000000000000010011100100111100;
assign LUT_3[716] = 32'b00000000000000000111111111110001;
assign LUT_3[717] = 32'b00000000000000001110101011001110;
assign LUT_3[718] = 32'b00000000000000001010000111010101;
assign LUT_3[719] = 32'b00000000000000010000110010110010;
assign LUT_3[720] = 32'b00000000000000001000101011111000;
assign LUT_3[721] = 32'b00000000000000001111010111010101;
assign LUT_3[722] = 32'b00000000000000001010110011011100;
assign LUT_3[723] = 32'b00000000000000010001011110111001;
assign LUT_3[724] = 32'b00000000000000000101111001101110;
assign LUT_3[725] = 32'b00000000000000001100100101001011;
assign LUT_3[726] = 32'b00000000000000001000000001010010;
assign LUT_3[727] = 32'b00000000000000001110101100101111;
assign LUT_3[728] = 32'b00000000000000001110000100111110;
assign LUT_3[729] = 32'b00000000000000010100110000011011;
assign LUT_3[730] = 32'b00000000000000010000001100100010;
assign LUT_3[731] = 32'b00000000000000010110110111111111;
assign LUT_3[732] = 32'b00000000000000001011010010110100;
assign LUT_3[733] = 32'b00000000000000010001111110010001;
assign LUT_3[734] = 32'b00000000000000001101011010011000;
assign LUT_3[735] = 32'b00000000000000010100000101110101;
assign LUT_3[736] = 32'b00000000000000000110100111010101;
assign LUT_3[737] = 32'b00000000000000001101010010110010;
assign LUT_3[738] = 32'b00000000000000001000101110111001;
assign LUT_3[739] = 32'b00000000000000001111011010010110;
assign LUT_3[740] = 32'b00000000000000000011110101001011;
assign LUT_3[741] = 32'b00000000000000001010100000101000;
assign LUT_3[742] = 32'b00000000000000000101111100101111;
assign LUT_3[743] = 32'b00000000000000001100101000001100;
assign LUT_3[744] = 32'b00000000000000001100000000011011;
assign LUT_3[745] = 32'b00000000000000010010101011111000;
assign LUT_3[746] = 32'b00000000000000001110000111111111;
assign LUT_3[747] = 32'b00000000000000010100110011011100;
assign LUT_3[748] = 32'b00000000000000001001001110010001;
assign LUT_3[749] = 32'b00000000000000001111111001101110;
assign LUT_3[750] = 32'b00000000000000001011010101110101;
assign LUT_3[751] = 32'b00000000000000010010000001010010;
assign LUT_3[752] = 32'b00000000000000001001111010011000;
assign LUT_3[753] = 32'b00000000000000010000100101110101;
assign LUT_3[754] = 32'b00000000000000001100000001111100;
assign LUT_3[755] = 32'b00000000000000010010101101011001;
assign LUT_3[756] = 32'b00000000000000000111001000001110;
assign LUT_3[757] = 32'b00000000000000001101110011101011;
assign LUT_3[758] = 32'b00000000000000001001001111110010;
assign LUT_3[759] = 32'b00000000000000001111111011001111;
assign LUT_3[760] = 32'b00000000000000001111010011011110;
assign LUT_3[761] = 32'b00000000000000010101111110111011;
assign LUT_3[762] = 32'b00000000000000010001011011000010;
assign LUT_3[763] = 32'b00000000000000011000000110011111;
assign LUT_3[764] = 32'b00000000000000001100100001010100;
assign LUT_3[765] = 32'b00000000000000010011001100110001;
assign LUT_3[766] = 32'b00000000000000001110101000111000;
assign LUT_3[767] = 32'b00000000000000010101010100010101;
assign LUT_3[768] = 32'b11111111111111111111100100101101;
assign LUT_3[769] = 32'b00000000000000000110010000001010;
assign LUT_3[770] = 32'b00000000000000000001101100010001;
assign LUT_3[771] = 32'b00000000000000001000010111101110;
assign LUT_3[772] = 32'b11111111111111111100110010100011;
assign LUT_3[773] = 32'b00000000000000000011011110000000;
assign LUT_3[774] = 32'b11111111111111111110111010000111;
assign LUT_3[775] = 32'b00000000000000000101100101100100;
assign LUT_3[776] = 32'b00000000000000000100111101110011;
assign LUT_3[777] = 32'b00000000000000001011101001010000;
assign LUT_3[778] = 32'b00000000000000000111000101010111;
assign LUT_3[779] = 32'b00000000000000001101110000110100;
assign LUT_3[780] = 32'b00000000000000000010001011101001;
assign LUT_3[781] = 32'b00000000000000001000110111000110;
assign LUT_3[782] = 32'b00000000000000000100010011001101;
assign LUT_3[783] = 32'b00000000000000001010111110101010;
assign LUT_3[784] = 32'b00000000000000000010110111110000;
assign LUT_3[785] = 32'b00000000000000001001100011001101;
assign LUT_3[786] = 32'b00000000000000000100111111010100;
assign LUT_3[787] = 32'b00000000000000001011101010110001;
assign LUT_3[788] = 32'b00000000000000000000000101100110;
assign LUT_3[789] = 32'b00000000000000000110110001000011;
assign LUT_3[790] = 32'b00000000000000000010001101001010;
assign LUT_3[791] = 32'b00000000000000001000111000100111;
assign LUT_3[792] = 32'b00000000000000001000010000110110;
assign LUT_3[793] = 32'b00000000000000001110111100010011;
assign LUT_3[794] = 32'b00000000000000001010011000011010;
assign LUT_3[795] = 32'b00000000000000010001000011110111;
assign LUT_3[796] = 32'b00000000000000000101011110101100;
assign LUT_3[797] = 32'b00000000000000001100001010001001;
assign LUT_3[798] = 32'b00000000000000000111100110010000;
assign LUT_3[799] = 32'b00000000000000001110010001101101;
assign LUT_3[800] = 32'b00000000000000000000110011001101;
assign LUT_3[801] = 32'b00000000000000000111011110101010;
assign LUT_3[802] = 32'b00000000000000000010111010110001;
assign LUT_3[803] = 32'b00000000000000001001100110001110;
assign LUT_3[804] = 32'b11111111111111111110000001000011;
assign LUT_3[805] = 32'b00000000000000000100101100100000;
assign LUT_3[806] = 32'b00000000000000000000001000100111;
assign LUT_3[807] = 32'b00000000000000000110110100000100;
assign LUT_3[808] = 32'b00000000000000000110001100010011;
assign LUT_3[809] = 32'b00000000000000001100110111110000;
assign LUT_3[810] = 32'b00000000000000001000010011110111;
assign LUT_3[811] = 32'b00000000000000001110111111010100;
assign LUT_3[812] = 32'b00000000000000000011011010001001;
assign LUT_3[813] = 32'b00000000000000001010000101100110;
assign LUT_3[814] = 32'b00000000000000000101100001101101;
assign LUT_3[815] = 32'b00000000000000001100001101001010;
assign LUT_3[816] = 32'b00000000000000000100000110010000;
assign LUT_3[817] = 32'b00000000000000001010110001101101;
assign LUT_3[818] = 32'b00000000000000000110001101110100;
assign LUT_3[819] = 32'b00000000000000001100111001010001;
assign LUT_3[820] = 32'b00000000000000000001010100000110;
assign LUT_3[821] = 32'b00000000000000000111111111100011;
assign LUT_3[822] = 32'b00000000000000000011011011101010;
assign LUT_3[823] = 32'b00000000000000001010000111000111;
assign LUT_3[824] = 32'b00000000000000001001011111010110;
assign LUT_3[825] = 32'b00000000000000010000001010110011;
assign LUT_3[826] = 32'b00000000000000001011100110111010;
assign LUT_3[827] = 32'b00000000000000010010010010010111;
assign LUT_3[828] = 32'b00000000000000000110101101001100;
assign LUT_3[829] = 32'b00000000000000001101011000101001;
assign LUT_3[830] = 32'b00000000000000001000110100110000;
assign LUT_3[831] = 32'b00000000000000001111100000001101;
assign LUT_3[832] = 32'b11111111111111111111011101011000;
assign LUT_3[833] = 32'b00000000000000000110001000110101;
assign LUT_3[834] = 32'b00000000000000000001100100111100;
assign LUT_3[835] = 32'b00000000000000001000010000011001;
assign LUT_3[836] = 32'b11111111111111111100101011001110;
assign LUT_3[837] = 32'b00000000000000000011010110101011;
assign LUT_3[838] = 32'b11111111111111111110110010110010;
assign LUT_3[839] = 32'b00000000000000000101011110001111;
assign LUT_3[840] = 32'b00000000000000000100110110011110;
assign LUT_3[841] = 32'b00000000000000001011100001111011;
assign LUT_3[842] = 32'b00000000000000000110111110000010;
assign LUT_3[843] = 32'b00000000000000001101101001011111;
assign LUT_3[844] = 32'b00000000000000000010000100010100;
assign LUT_3[845] = 32'b00000000000000001000101111110001;
assign LUT_3[846] = 32'b00000000000000000100001011111000;
assign LUT_3[847] = 32'b00000000000000001010110111010101;
assign LUT_3[848] = 32'b00000000000000000010110000011011;
assign LUT_3[849] = 32'b00000000000000001001011011111000;
assign LUT_3[850] = 32'b00000000000000000100110111111111;
assign LUT_3[851] = 32'b00000000000000001011100011011100;
assign LUT_3[852] = 32'b11111111111111111111111110010001;
assign LUT_3[853] = 32'b00000000000000000110101001101110;
assign LUT_3[854] = 32'b00000000000000000010000101110101;
assign LUT_3[855] = 32'b00000000000000001000110001010010;
assign LUT_3[856] = 32'b00000000000000001000001001100001;
assign LUT_3[857] = 32'b00000000000000001110110100111110;
assign LUT_3[858] = 32'b00000000000000001010010001000101;
assign LUT_3[859] = 32'b00000000000000010000111100100010;
assign LUT_3[860] = 32'b00000000000000000101010111010111;
assign LUT_3[861] = 32'b00000000000000001100000010110100;
assign LUT_3[862] = 32'b00000000000000000111011110111011;
assign LUT_3[863] = 32'b00000000000000001110001010011000;
assign LUT_3[864] = 32'b00000000000000000000101011111000;
assign LUT_3[865] = 32'b00000000000000000111010111010101;
assign LUT_3[866] = 32'b00000000000000000010110011011100;
assign LUT_3[867] = 32'b00000000000000001001011110111001;
assign LUT_3[868] = 32'b11111111111111111101111001101110;
assign LUT_3[869] = 32'b00000000000000000100100101001011;
assign LUT_3[870] = 32'b00000000000000000000000001010010;
assign LUT_3[871] = 32'b00000000000000000110101100101111;
assign LUT_3[872] = 32'b00000000000000000110000100111110;
assign LUT_3[873] = 32'b00000000000000001100110000011011;
assign LUT_3[874] = 32'b00000000000000001000001100100010;
assign LUT_3[875] = 32'b00000000000000001110110111111111;
assign LUT_3[876] = 32'b00000000000000000011010010110100;
assign LUT_3[877] = 32'b00000000000000001001111110010001;
assign LUT_3[878] = 32'b00000000000000000101011010011000;
assign LUT_3[879] = 32'b00000000000000001100000101110101;
assign LUT_3[880] = 32'b00000000000000000011111110111011;
assign LUT_3[881] = 32'b00000000000000001010101010011000;
assign LUT_3[882] = 32'b00000000000000000110000110011111;
assign LUT_3[883] = 32'b00000000000000001100110001111100;
assign LUT_3[884] = 32'b00000000000000000001001100110001;
assign LUT_3[885] = 32'b00000000000000000111111000001110;
assign LUT_3[886] = 32'b00000000000000000011010100010101;
assign LUT_3[887] = 32'b00000000000000001001111111110010;
assign LUT_3[888] = 32'b00000000000000001001011000000001;
assign LUT_3[889] = 32'b00000000000000010000000011011110;
assign LUT_3[890] = 32'b00000000000000001011011111100101;
assign LUT_3[891] = 32'b00000000000000010010001011000010;
assign LUT_3[892] = 32'b00000000000000000110100101110111;
assign LUT_3[893] = 32'b00000000000000001101010001010100;
assign LUT_3[894] = 32'b00000000000000001000101101011011;
assign LUT_3[895] = 32'b00000000000000001111011000111000;
assign LUT_3[896] = 32'b00000000000000000001101111101011;
assign LUT_3[897] = 32'b00000000000000001000011011001000;
assign LUT_3[898] = 32'b00000000000000000011110111001111;
assign LUT_3[899] = 32'b00000000000000001010100010101100;
assign LUT_3[900] = 32'b11111111111111111110111101100001;
assign LUT_3[901] = 32'b00000000000000000101101000111110;
assign LUT_3[902] = 32'b00000000000000000001000101000101;
assign LUT_3[903] = 32'b00000000000000000111110000100010;
assign LUT_3[904] = 32'b00000000000000000111001000110001;
assign LUT_3[905] = 32'b00000000000000001101110100001110;
assign LUT_3[906] = 32'b00000000000000001001010000010101;
assign LUT_3[907] = 32'b00000000000000001111111011110010;
assign LUT_3[908] = 32'b00000000000000000100010110100111;
assign LUT_3[909] = 32'b00000000000000001011000010000100;
assign LUT_3[910] = 32'b00000000000000000110011110001011;
assign LUT_3[911] = 32'b00000000000000001101001001101000;
assign LUT_3[912] = 32'b00000000000000000101000010101110;
assign LUT_3[913] = 32'b00000000000000001011101110001011;
assign LUT_3[914] = 32'b00000000000000000111001010010010;
assign LUT_3[915] = 32'b00000000000000001101110101101111;
assign LUT_3[916] = 32'b00000000000000000010010000100100;
assign LUT_3[917] = 32'b00000000000000001000111100000001;
assign LUT_3[918] = 32'b00000000000000000100011000001000;
assign LUT_3[919] = 32'b00000000000000001011000011100101;
assign LUT_3[920] = 32'b00000000000000001010011011110100;
assign LUT_3[921] = 32'b00000000000000010001000111010001;
assign LUT_3[922] = 32'b00000000000000001100100011011000;
assign LUT_3[923] = 32'b00000000000000010011001110110101;
assign LUT_3[924] = 32'b00000000000000000111101001101010;
assign LUT_3[925] = 32'b00000000000000001110010101000111;
assign LUT_3[926] = 32'b00000000000000001001110001001110;
assign LUT_3[927] = 32'b00000000000000010000011100101011;
assign LUT_3[928] = 32'b00000000000000000010111110001011;
assign LUT_3[929] = 32'b00000000000000001001101001101000;
assign LUT_3[930] = 32'b00000000000000000101000101101111;
assign LUT_3[931] = 32'b00000000000000001011110001001100;
assign LUT_3[932] = 32'b00000000000000000000001100000001;
assign LUT_3[933] = 32'b00000000000000000110110111011110;
assign LUT_3[934] = 32'b00000000000000000010010011100101;
assign LUT_3[935] = 32'b00000000000000001000111111000010;
assign LUT_3[936] = 32'b00000000000000001000010111010001;
assign LUT_3[937] = 32'b00000000000000001111000010101110;
assign LUT_3[938] = 32'b00000000000000001010011110110101;
assign LUT_3[939] = 32'b00000000000000010001001010010010;
assign LUT_3[940] = 32'b00000000000000000101100101000111;
assign LUT_3[941] = 32'b00000000000000001100010000100100;
assign LUT_3[942] = 32'b00000000000000000111101100101011;
assign LUT_3[943] = 32'b00000000000000001110011000001000;
assign LUT_3[944] = 32'b00000000000000000110010001001110;
assign LUT_3[945] = 32'b00000000000000001100111100101011;
assign LUT_3[946] = 32'b00000000000000001000011000110010;
assign LUT_3[947] = 32'b00000000000000001111000100001111;
assign LUT_3[948] = 32'b00000000000000000011011111000100;
assign LUT_3[949] = 32'b00000000000000001010001010100001;
assign LUT_3[950] = 32'b00000000000000000101100110101000;
assign LUT_3[951] = 32'b00000000000000001100010010000101;
assign LUT_3[952] = 32'b00000000000000001011101010010100;
assign LUT_3[953] = 32'b00000000000000010010010101110001;
assign LUT_3[954] = 32'b00000000000000001101110001111000;
assign LUT_3[955] = 32'b00000000000000010100011101010101;
assign LUT_3[956] = 32'b00000000000000001000111000001010;
assign LUT_3[957] = 32'b00000000000000001111100011100111;
assign LUT_3[958] = 32'b00000000000000001010111111101110;
assign LUT_3[959] = 32'b00000000000000010001101011001011;
assign LUT_3[960] = 32'b00000000000000000001101000010110;
assign LUT_3[961] = 32'b00000000000000001000010011110011;
assign LUT_3[962] = 32'b00000000000000000011101111111010;
assign LUT_3[963] = 32'b00000000000000001010011011010111;
assign LUT_3[964] = 32'b11111111111111111110110110001100;
assign LUT_3[965] = 32'b00000000000000000101100001101001;
assign LUT_3[966] = 32'b00000000000000000000111101110000;
assign LUT_3[967] = 32'b00000000000000000111101001001101;
assign LUT_3[968] = 32'b00000000000000000111000001011100;
assign LUT_3[969] = 32'b00000000000000001101101100111001;
assign LUT_3[970] = 32'b00000000000000001001001001000000;
assign LUT_3[971] = 32'b00000000000000001111110100011101;
assign LUT_3[972] = 32'b00000000000000000100001111010010;
assign LUT_3[973] = 32'b00000000000000001010111010101111;
assign LUT_3[974] = 32'b00000000000000000110010110110110;
assign LUT_3[975] = 32'b00000000000000001101000010010011;
assign LUT_3[976] = 32'b00000000000000000100111011011001;
assign LUT_3[977] = 32'b00000000000000001011100110110110;
assign LUT_3[978] = 32'b00000000000000000111000010111101;
assign LUT_3[979] = 32'b00000000000000001101101110011010;
assign LUT_3[980] = 32'b00000000000000000010001001001111;
assign LUT_3[981] = 32'b00000000000000001000110100101100;
assign LUT_3[982] = 32'b00000000000000000100010000110011;
assign LUT_3[983] = 32'b00000000000000001010111100010000;
assign LUT_3[984] = 32'b00000000000000001010010100011111;
assign LUT_3[985] = 32'b00000000000000010000111111111100;
assign LUT_3[986] = 32'b00000000000000001100011100000011;
assign LUT_3[987] = 32'b00000000000000010011000111100000;
assign LUT_3[988] = 32'b00000000000000000111100010010101;
assign LUT_3[989] = 32'b00000000000000001110001101110010;
assign LUT_3[990] = 32'b00000000000000001001101001111001;
assign LUT_3[991] = 32'b00000000000000010000010101010110;
assign LUT_3[992] = 32'b00000000000000000010110110110110;
assign LUT_3[993] = 32'b00000000000000001001100010010011;
assign LUT_3[994] = 32'b00000000000000000100111110011010;
assign LUT_3[995] = 32'b00000000000000001011101001110111;
assign LUT_3[996] = 32'b00000000000000000000000100101100;
assign LUT_3[997] = 32'b00000000000000000110110000001001;
assign LUT_3[998] = 32'b00000000000000000010001100010000;
assign LUT_3[999] = 32'b00000000000000001000110111101101;
assign LUT_3[1000] = 32'b00000000000000001000001111111100;
assign LUT_3[1001] = 32'b00000000000000001110111011011001;
assign LUT_3[1002] = 32'b00000000000000001010010111100000;
assign LUT_3[1003] = 32'b00000000000000010001000010111101;
assign LUT_3[1004] = 32'b00000000000000000101011101110010;
assign LUT_3[1005] = 32'b00000000000000001100001001001111;
assign LUT_3[1006] = 32'b00000000000000000111100101010110;
assign LUT_3[1007] = 32'b00000000000000001110010000110011;
assign LUT_3[1008] = 32'b00000000000000000110001001111001;
assign LUT_3[1009] = 32'b00000000000000001100110101010110;
assign LUT_3[1010] = 32'b00000000000000001000010001011101;
assign LUT_3[1011] = 32'b00000000000000001110111100111010;
assign LUT_3[1012] = 32'b00000000000000000011010111101111;
assign LUT_3[1013] = 32'b00000000000000001010000011001100;
assign LUT_3[1014] = 32'b00000000000000000101011111010011;
assign LUT_3[1015] = 32'b00000000000000001100001010110000;
assign LUT_3[1016] = 32'b00000000000000001011100010111111;
assign LUT_3[1017] = 32'b00000000000000010010001110011100;
assign LUT_3[1018] = 32'b00000000000000001101101010100011;
assign LUT_3[1019] = 32'b00000000000000010100010110000000;
assign LUT_3[1020] = 32'b00000000000000001000110000110101;
assign LUT_3[1021] = 32'b00000000000000001111011100010010;
assign LUT_3[1022] = 32'b00000000000000001010111000011001;
assign LUT_3[1023] = 32'b00000000000000010001100011110110;
assign LUT_3[1024] = 32'b00000000000000000110100100111101;
assign LUT_3[1025] = 32'b00000000000000001101010000011010;
assign LUT_3[1026] = 32'b00000000000000001000101100100001;
assign LUT_3[1027] = 32'b00000000000000001111010111111110;
assign LUT_3[1028] = 32'b00000000000000000011110010110011;
assign LUT_3[1029] = 32'b00000000000000001010011110010000;
assign LUT_3[1030] = 32'b00000000000000000101111010010111;
assign LUT_3[1031] = 32'b00000000000000001100100101110100;
assign LUT_3[1032] = 32'b00000000000000001011111110000011;
assign LUT_3[1033] = 32'b00000000000000010010101001100000;
assign LUT_3[1034] = 32'b00000000000000001110000101100111;
assign LUT_3[1035] = 32'b00000000000000010100110001000100;
assign LUT_3[1036] = 32'b00000000000000001001001011111001;
assign LUT_3[1037] = 32'b00000000000000001111110111010110;
assign LUT_3[1038] = 32'b00000000000000001011010011011101;
assign LUT_3[1039] = 32'b00000000000000010001111110111010;
assign LUT_3[1040] = 32'b00000000000000001001111000000000;
assign LUT_3[1041] = 32'b00000000000000010000100011011101;
assign LUT_3[1042] = 32'b00000000000000001011111111100100;
assign LUT_3[1043] = 32'b00000000000000010010101011000001;
assign LUT_3[1044] = 32'b00000000000000000111000101110110;
assign LUT_3[1045] = 32'b00000000000000001101110001010011;
assign LUT_3[1046] = 32'b00000000000000001001001101011010;
assign LUT_3[1047] = 32'b00000000000000001111111000110111;
assign LUT_3[1048] = 32'b00000000000000001111010001000110;
assign LUT_3[1049] = 32'b00000000000000010101111100100011;
assign LUT_3[1050] = 32'b00000000000000010001011000101010;
assign LUT_3[1051] = 32'b00000000000000011000000100000111;
assign LUT_3[1052] = 32'b00000000000000001100011110111100;
assign LUT_3[1053] = 32'b00000000000000010011001010011001;
assign LUT_3[1054] = 32'b00000000000000001110100110100000;
assign LUT_3[1055] = 32'b00000000000000010101010001111101;
assign LUT_3[1056] = 32'b00000000000000000111110011011101;
assign LUT_3[1057] = 32'b00000000000000001110011110111010;
assign LUT_3[1058] = 32'b00000000000000001001111011000001;
assign LUT_3[1059] = 32'b00000000000000010000100110011110;
assign LUT_3[1060] = 32'b00000000000000000101000001010011;
assign LUT_3[1061] = 32'b00000000000000001011101100110000;
assign LUT_3[1062] = 32'b00000000000000000111001000110111;
assign LUT_3[1063] = 32'b00000000000000001101110100010100;
assign LUT_3[1064] = 32'b00000000000000001101001100100011;
assign LUT_3[1065] = 32'b00000000000000010011111000000000;
assign LUT_3[1066] = 32'b00000000000000001111010100000111;
assign LUT_3[1067] = 32'b00000000000000010101111111100100;
assign LUT_3[1068] = 32'b00000000000000001010011010011001;
assign LUT_3[1069] = 32'b00000000000000010001000101110110;
assign LUT_3[1070] = 32'b00000000000000001100100001111101;
assign LUT_3[1071] = 32'b00000000000000010011001101011010;
assign LUT_3[1072] = 32'b00000000000000001011000110100000;
assign LUT_3[1073] = 32'b00000000000000010001110001111101;
assign LUT_3[1074] = 32'b00000000000000001101001110000100;
assign LUT_3[1075] = 32'b00000000000000010011111001100001;
assign LUT_3[1076] = 32'b00000000000000001000010100010110;
assign LUT_3[1077] = 32'b00000000000000001110111111110011;
assign LUT_3[1078] = 32'b00000000000000001010011011111010;
assign LUT_3[1079] = 32'b00000000000000010001000111010111;
assign LUT_3[1080] = 32'b00000000000000010000011111100110;
assign LUT_3[1081] = 32'b00000000000000010111001011000011;
assign LUT_3[1082] = 32'b00000000000000010010100111001010;
assign LUT_3[1083] = 32'b00000000000000011001010010100111;
assign LUT_3[1084] = 32'b00000000000000001101101101011100;
assign LUT_3[1085] = 32'b00000000000000010100011000111001;
assign LUT_3[1086] = 32'b00000000000000001111110101000000;
assign LUT_3[1087] = 32'b00000000000000010110100000011101;
assign LUT_3[1088] = 32'b00000000000000000110011101101000;
assign LUT_3[1089] = 32'b00000000000000001101001001000101;
assign LUT_3[1090] = 32'b00000000000000001000100101001100;
assign LUT_3[1091] = 32'b00000000000000001111010000101001;
assign LUT_3[1092] = 32'b00000000000000000011101011011110;
assign LUT_3[1093] = 32'b00000000000000001010010110111011;
assign LUT_3[1094] = 32'b00000000000000000101110011000010;
assign LUT_3[1095] = 32'b00000000000000001100011110011111;
assign LUT_3[1096] = 32'b00000000000000001011110110101110;
assign LUT_3[1097] = 32'b00000000000000010010100010001011;
assign LUT_3[1098] = 32'b00000000000000001101111110010010;
assign LUT_3[1099] = 32'b00000000000000010100101001101111;
assign LUT_3[1100] = 32'b00000000000000001001000100100100;
assign LUT_3[1101] = 32'b00000000000000001111110000000001;
assign LUT_3[1102] = 32'b00000000000000001011001100001000;
assign LUT_3[1103] = 32'b00000000000000010001110111100101;
assign LUT_3[1104] = 32'b00000000000000001001110000101011;
assign LUT_3[1105] = 32'b00000000000000010000011100001000;
assign LUT_3[1106] = 32'b00000000000000001011111000001111;
assign LUT_3[1107] = 32'b00000000000000010010100011101100;
assign LUT_3[1108] = 32'b00000000000000000110111110100001;
assign LUT_3[1109] = 32'b00000000000000001101101001111110;
assign LUT_3[1110] = 32'b00000000000000001001000110000101;
assign LUT_3[1111] = 32'b00000000000000001111110001100010;
assign LUT_3[1112] = 32'b00000000000000001111001001110001;
assign LUT_3[1113] = 32'b00000000000000010101110101001110;
assign LUT_3[1114] = 32'b00000000000000010001010001010101;
assign LUT_3[1115] = 32'b00000000000000010111111100110010;
assign LUT_3[1116] = 32'b00000000000000001100010111100111;
assign LUT_3[1117] = 32'b00000000000000010011000011000100;
assign LUT_3[1118] = 32'b00000000000000001110011111001011;
assign LUT_3[1119] = 32'b00000000000000010101001010101000;
assign LUT_3[1120] = 32'b00000000000000000111101100001000;
assign LUT_3[1121] = 32'b00000000000000001110010111100101;
assign LUT_3[1122] = 32'b00000000000000001001110011101100;
assign LUT_3[1123] = 32'b00000000000000010000011111001001;
assign LUT_3[1124] = 32'b00000000000000000100111001111110;
assign LUT_3[1125] = 32'b00000000000000001011100101011011;
assign LUT_3[1126] = 32'b00000000000000000111000001100010;
assign LUT_3[1127] = 32'b00000000000000001101101100111111;
assign LUT_3[1128] = 32'b00000000000000001101000101001110;
assign LUT_3[1129] = 32'b00000000000000010011110000101011;
assign LUT_3[1130] = 32'b00000000000000001111001100110010;
assign LUT_3[1131] = 32'b00000000000000010101111000001111;
assign LUT_3[1132] = 32'b00000000000000001010010011000100;
assign LUT_3[1133] = 32'b00000000000000010000111110100001;
assign LUT_3[1134] = 32'b00000000000000001100011010101000;
assign LUT_3[1135] = 32'b00000000000000010011000110000101;
assign LUT_3[1136] = 32'b00000000000000001010111111001011;
assign LUT_3[1137] = 32'b00000000000000010001101010101000;
assign LUT_3[1138] = 32'b00000000000000001101000110101111;
assign LUT_3[1139] = 32'b00000000000000010011110010001100;
assign LUT_3[1140] = 32'b00000000000000001000001101000001;
assign LUT_3[1141] = 32'b00000000000000001110111000011110;
assign LUT_3[1142] = 32'b00000000000000001010010100100101;
assign LUT_3[1143] = 32'b00000000000000010001000000000010;
assign LUT_3[1144] = 32'b00000000000000010000011000010001;
assign LUT_3[1145] = 32'b00000000000000010111000011101110;
assign LUT_3[1146] = 32'b00000000000000010010011111110101;
assign LUT_3[1147] = 32'b00000000000000011001001011010010;
assign LUT_3[1148] = 32'b00000000000000001101100110000111;
assign LUT_3[1149] = 32'b00000000000000010100010001100100;
assign LUT_3[1150] = 32'b00000000000000001111101101101011;
assign LUT_3[1151] = 32'b00000000000000010110011001001000;
assign LUT_3[1152] = 32'b00000000000000001000101111111011;
assign LUT_3[1153] = 32'b00000000000000001111011011011000;
assign LUT_3[1154] = 32'b00000000000000001010110111011111;
assign LUT_3[1155] = 32'b00000000000000010001100010111100;
assign LUT_3[1156] = 32'b00000000000000000101111101110001;
assign LUT_3[1157] = 32'b00000000000000001100101001001110;
assign LUT_3[1158] = 32'b00000000000000001000000101010101;
assign LUT_3[1159] = 32'b00000000000000001110110000110010;
assign LUT_3[1160] = 32'b00000000000000001110001001000001;
assign LUT_3[1161] = 32'b00000000000000010100110100011110;
assign LUT_3[1162] = 32'b00000000000000010000010000100101;
assign LUT_3[1163] = 32'b00000000000000010110111100000010;
assign LUT_3[1164] = 32'b00000000000000001011010110110111;
assign LUT_3[1165] = 32'b00000000000000010010000010010100;
assign LUT_3[1166] = 32'b00000000000000001101011110011011;
assign LUT_3[1167] = 32'b00000000000000010100001001111000;
assign LUT_3[1168] = 32'b00000000000000001100000010111110;
assign LUT_3[1169] = 32'b00000000000000010010101110011011;
assign LUT_3[1170] = 32'b00000000000000001110001010100010;
assign LUT_3[1171] = 32'b00000000000000010100110101111111;
assign LUT_3[1172] = 32'b00000000000000001001010000110100;
assign LUT_3[1173] = 32'b00000000000000001111111100010001;
assign LUT_3[1174] = 32'b00000000000000001011011000011000;
assign LUT_3[1175] = 32'b00000000000000010010000011110101;
assign LUT_3[1176] = 32'b00000000000000010001011100000100;
assign LUT_3[1177] = 32'b00000000000000011000000111100001;
assign LUT_3[1178] = 32'b00000000000000010011100011101000;
assign LUT_3[1179] = 32'b00000000000000011010001111000101;
assign LUT_3[1180] = 32'b00000000000000001110101001111010;
assign LUT_3[1181] = 32'b00000000000000010101010101010111;
assign LUT_3[1182] = 32'b00000000000000010000110001011110;
assign LUT_3[1183] = 32'b00000000000000010111011100111011;
assign LUT_3[1184] = 32'b00000000000000001001111110011011;
assign LUT_3[1185] = 32'b00000000000000010000101001111000;
assign LUT_3[1186] = 32'b00000000000000001100000101111111;
assign LUT_3[1187] = 32'b00000000000000010010110001011100;
assign LUT_3[1188] = 32'b00000000000000000111001100010001;
assign LUT_3[1189] = 32'b00000000000000001101110111101110;
assign LUT_3[1190] = 32'b00000000000000001001010011110101;
assign LUT_3[1191] = 32'b00000000000000001111111111010010;
assign LUT_3[1192] = 32'b00000000000000001111010111100001;
assign LUT_3[1193] = 32'b00000000000000010110000010111110;
assign LUT_3[1194] = 32'b00000000000000010001011111000101;
assign LUT_3[1195] = 32'b00000000000000011000001010100010;
assign LUT_3[1196] = 32'b00000000000000001100100101010111;
assign LUT_3[1197] = 32'b00000000000000010011010000110100;
assign LUT_3[1198] = 32'b00000000000000001110101100111011;
assign LUT_3[1199] = 32'b00000000000000010101011000011000;
assign LUT_3[1200] = 32'b00000000000000001101010001011110;
assign LUT_3[1201] = 32'b00000000000000010011111100111011;
assign LUT_3[1202] = 32'b00000000000000001111011001000010;
assign LUT_3[1203] = 32'b00000000000000010110000100011111;
assign LUT_3[1204] = 32'b00000000000000001010011111010100;
assign LUT_3[1205] = 32'b00000000000000010001001010110001;
assign LUT_3[1206] = 32'b00000000000000001100100110111000;
assign LUT_3[1207] = 32'b00000000000000010011010010010101;
assign LUT_3[1208] = 32'b00000000000000010010101010100100;
assign LUT_3[1209] = 32'b00000000000000011001010110000001;
assign LUT_3[1210] = 32'b00000000000000010100110010001000;
assign LUT_3[1211] = 32'b00000000000000011011011101100101;
assign LUT_3[1212] = 32'b00000000000000001111111000011010;
assign LUT_3[1213] = 32'b00000000000000010110100011110111;
assign LUT_3[1214] = 32'b00000000000000010001111111111110;
assign LUT_3[1215] = 32'b00000000000000011000101011011011;
assign LUT_3[1216] = 32'b00000000000000001000101000100110;
assign LUT_3[1217] = 32'b00000000000000001111010100000011;
assign LUT_3[1218] = 32'b00000000000000001010110000001010;
assign LUT_3[1219] = 32'b00000000000000010001011011100111;
assign LUT_3[1220] = 32'b00000000000000000101110110011100;
assign LUT_3[1221] = 32'b00000000000000001100100001111001;
assign LUT_3[1222] = 32'b00000000000000000111111110000000;
assign LUT_3[1223] = 32'b00000000000000001110101001011101;
assign LUT_3[1224] = 32'b00000000000000001110000001101100;
assign LUT_3[1225] = 32'b00000000000000010100101101001001;
assign LUT_3[1226] = 32'b00000000000000010000001001010000;
assign LUT_3[1227] = 32'b00000000000000010110110100101101;
assign LUT_3[1228] = 32'b00000000000000001011001111100010;
assign LUT_3[1229] = 32'b00000000000000010001111010111111;
assign LUT_3[1230] = 32'b00000000000000001101010111000110;
assign LUT_3[1231] = 32'b00000000000000010100000010100011;
assign LUT_3[1232] = 32'b00000000000000001011111011101001;
assign LUT_3[1233] = 32'b00000000000000010010100111000110;
assign LUT_3[1234] = 32'b00000000000000001110000011001101;
assign LUT_3[1235] = 32'b00000000000000010100101110101010;
assign LUT_3[1236] = 32'b00000000000000001001001001011111;
assign LUT_3[1237] = 32'b00000000000000001111110100111100;
assign LUT_3[1238] = 32'b00000000000000001011010001000011;
assign LUT_3[1239] = 32'b00000000000000010001111100100000;
assign LUT_3[1240] = 32'b00000000000000010001010100101111;
assign LUT_3[1241] = 32'b00000000000000011000000000001100;
assign LUT_3[1242] = 32'b00000000000000010011011100010011;
assign LUT_3[1243] = 32'b00000000000000011010000111110000;
assign LUT_3[1244] = 32'b00000000000000001110100010100101;
assign LUT_3[1245] = 32'b00000000000000010101001110000010;
assign LUT_3[1246] = 32'b00000000000000010000101010001001;
assign LUT_3[1247] = 32'b00000000000000010111010101100110;
assign LUT_3[1248] = 32'b00000000000000001001110111000110;
assign LUT_3[1249] = 32'b00000000000000010000100010100011;
assign LUT_3[1250] = 32'b00000000000000001011111110101010;
assign LUT_3[1251] = 32'b00000000000000010010101010000111;
assign LUT_3[1252] = 32'b00000000000000000111000100111100;
assign LUT_3[1253] = 32'b00000000000000001101110000011001;
assign LUT_3[1254] = 32'b00000000000000001001001100100000;
assign LUT_3[1255] = 32'b00000000000000001111110111111101;
assign LUT_3[1256] = 32'b00000000000000001111010000001100;
assign LUT_3[1257] = 32'b00000000000000010101111011101001;
assign LUT_3[1258] = 32'b00000000000000010001010111110000;
assign LUT_3[1259] = 32'b00000000000000011000000011001101;
assign LUT_3[1260] = 32'b00000000000000001100011110000010;
assign LUT_3[1261] = 32'b00000000000000010011001001011111;
assign LUT_3[1262] = 32'b00000000000000001110100101100110;
assign LUT_3[1263] = 32'b00000000000000010101010001000011;
assign LUT_3[1264] = 32'b00000000000000001101001010001001;
assign LUT_3[1265] = 32'b00000000000000010011110101100110;
assign LUT_3[1266] = 32'b00000000000000001111010001101101;
assign LUT_3[1267] = 32'b00000000000000010101111101001010;
assign LUT_3[1268] = 32'b00000000000000001010010111111111;
assign LUT_3[1269] = 32'b00000000000000010001000011011100;
assign LUT_3[1270] = 32'b00000000000000001100011111100011;
assign LUT_3[1271] = 32'b00000000000000010011001011000000;
assign LUT_3[1272] = 32'b00000000000000010010100011001111;
assign LUT_3[1273] = 32'b00000000000000011001001110101100;
assign LUT_3[1274] = 32'b00000000000000010100101010110011;
assign LUT_3[1275] = 32'b00000000000000011011010110010000;
assign LUT_3[1276] = 32'b00000000000000001111110001000101;
assign LUT_3[1277] = 32'b00000000000000010110011100100010;
assign LUT_3[1278] = 32'b00000000000000010001111000101001;
assign LUT_3[1279] = 32'b00000000000000011000100100000110;
assign LUT_3[1280] = 32'b00000000000000000010110100011110;
assign LUT_3[1281] = 32'b00000000000000001001011111111011;
assign LUT_3[1282] = 32'b00000000000000000100111100000010;
assign LUT_3[1283] = 32'b00000000000000001011100111011111;
assign LUT_3[1284] = 32'b00000000000000000000000010010100;
assign LUT_3[1285] = 32'b00000000000000000110101101110001;
assign LUT_3[1286] = 32'b00000000000000000010001001111000;
assign LUT_3[1287] = 32'b00000000000000001000110101010101;
assign LUT_3[1288] = 32'b00000000000000001000001101100100;
assign LUT_3[1289] = 32'b00000000000000001110111001000001;
assign LUT_3[1290] = 32'b00000000000000001010010101001000;
assign LUT_3[1291] = 32'b00000000000000010001000000100101;
assign LUT_3[1292] = 32'b00000000000000000101011011011010;
assign LUT_3[1293] = 32'b00000000000000001100000110110111;
assign LUT_3[1294] = 32'b00000000000000000111100010111110;
assign LUT_3[1295] = 32'b00000000000000001110001110011011;
assign LUT_3[1296] = 32'b00000000000000000110000111100001;
assign LUT_3[1297] = 32'b00000000000000001100110010111110;
assign LUT_3[1298] = 32'b00000000000000001000001111000101;
assign LUT_3[1299] = 32'b00000000000000001110111010100010;
assign LUT_3[1300] = 32'b00000000000000000011010101010111;
assign LUT_3[1301] = 32'b00000000000000001010000000110100;
assign LUT_3[1302] = 32'b00000000000000000101011100111011;
assign LUT_3[1303] = 32'b00000000000000001100001000011000;
assign LUT_3[1304] = 32'b00000000000000001011100000100111;
assign LUT_3[1305] = 32'b00000000000000010010001100000100;
assign LUT_3[1306] = 32'b00000000000000001101101000001011;
assign LUT_3[1307] = 32'b00000000000000010100010011101000;
assign LUT_3[1308] = 32'b00000000000000001000101110011101;
assign LUT_3[1309] = 32'b00000000000000001111011001111010;
assign LUT_3[1310] = 32'b00000000000000001010110110000001;
assign LUT_3[1311] = 32'b00000000000000010001100001011110;
assign LUT_3[1312] = 32'b00000000000000000100000010111110;
assign LUT_3[1313] = 32'b00000000000000001010101110011011;
assign LUT_3[1314] = 32'b00000000000000000110001010100010;
assign LUT_3[1315] = 32'b00000000000000001100110101111111;
assign LUT_3[1316] = 32'b00000000000000000001010000110100;
assign LUT_3[1317] = 32'b00000000000000000111111100010001;
assign LUT_3[1318] = 32'b00000000000000000011011000011000;
assign LUT_3[1319] = 32'b00000000000000001010000011110101;
assign LUT_3[1320] = 32'b00000000000000001001011100000100;
assign LUT_3[1321] = 32'b00000000000000010000000111100001;
assign LUT_3[1322] = 32'b00000000000000001011100011101000;
assign LUT_3[1323] = 32'b00000000000000010010001111000101;
assign LUT_3[1324] = 32'b00000000000000000110101001111010;
assign LUT_3[1325] = 32'b00000000000000001101010101010111;
assign LUT_3[1326] = 32'b00000000000000001000110001011110;
assign LUT_3[1327] = 32'b00000000000000001111011100111011;
assign LUT_3[1328] = 32'b00000000000000000111010110000001;
assign LUT_3[1329] = 32'b00000000000000001110000001011110;
assign LUT_3[1330] = 32'b00000000000000001001011101100101;
assign LUT_3[1331] = 32'b00000000000000010000001001000010;
assign LUT_3[1332] = 32'b00000000000000000100100011110111;
assign LUT_3[1333] = 32'b00000000000000001011001111010100;
assign LUT_3[1334] = 32'b00000000000000000110101011011011;
assign LUT_3[1335] = 32'b00000000000000001101010110111000;
assign LUT_3[1336] = 32'b00000000000000001100101111000111;
assign LUT_3[1337] = 32'b00000000000000010011011010100100;
assign LUT_3[1338] = 32'b00000000000000001110110110101011;
assign LUT_3[1339] = 32'b00000000000000010101100010001000;
assign LUT_3[1340] = 32'b00000000000000001001111100111101;
assign LUT_3[1341] = 32'b00000000000000010000101000011010;
assign LUT_3[1342] = 32'b00000000000000001100000100100001;
assign LUT_3[1343] = 32'b00000000000000010010101111111110;
assign LUT_3[1344] = 32'b00000000000000000010101101001001;
assign LUT_3[1345] = 32'b00000000000000001001011000100110;
assign LUT_3[1346] = 32'b00000000000000000100110100101101;
assign LUT_3[1347] = 32'b00000000000000001011100000001010;
assign LUT_3[1348] = 32'b11111111111111111111111010111111;
assign LUT_3[1349] = 32'b00000000000000000110100110011100;
assign LUT_3[1350] = 32'b00000000000000000010000010100011;
assign LUT_3[1351] = 32'b00000000000000001000101110000000;
assign LUT_3[1352] = 32'b00000000000000001000000110001111;
assign LUT_3[1353] = 32'b00000000000000001110110001101100;
assign LUT_3[1354] = 32'b00000000000000001010001101110011;
assign LUT_3[1355] = 32'b00000000000000010000111001010000;
assign LUT_3[1356] = 32'b00000000000000000101010100000101;
assign LUT_3[1357] = 32'b00000000000000001011111111100010;
assign LUT_3[1358] = 32'b00000000000000000111011011101001;
assign LUT_3[1359] = 32'b00000000000000001110000111000110;
assign LUT_3[1360] = 32'b00000000000000000110000000001100;
assign LUT_3[1361] = 32'b00000000000000001100101011101001;
assign LUT_3[1362] = 32'b00000000000000001000000111110000;
assign LUT_3[1363] = 32'b00000000000000001110110011001101;
assign LUT_3[1364] = 32'b00000000000000000011001110000010;
assign LUT_3[1365] = 32'b00000000000000001001111001011111;
assign LUT_3[1366] = 32'b00000000000000000101010101100110;
assign LUT_3[1367] = 32'b00000000000000001100000001000011;
assign LUT_3[1368] = 32'b00000000000000001011011001010010;
assign LUT_3[1369] = 32'b00000000000000010010000100101111;
assign LUT_3[1370] = 32'b00000000000000001101100000110110;
assign LUT_3[1371] = 32'b00000000000000010100001100010011;
assign LUT_3[1372] = 32'b00000000000000001000100111001000;
assign LUT_3[1373] = 32'b00000000000000001111010010100101;
assign LUT_3[1374] = 32'b00000000000000001010101110101100;
assign LUT_3[1375] = 32'b00000000000000010001011010001001;
assign LUT_3[1376] = 32'b00000000000000000011111011101001;
assign LUT_3[1377] = 32'b00000000000000001010100111000110;
assign LUT_3[1378] = 32'b00000000000000000110000011001101;
assign LUT_3[1379] = 32'b00000000000000001100101110101010;
assign LUT_3[1380] = 32'b00000000000000000001001001011111;
assign LUT_3[1381] = 32'b00000000000000000111110100111100;
assign LUT_3[1382] = 32'b00000000000000000011010001000011;
assign LUT_3[1383] = 32'b00000000000000001001111100100000;
assign LUT_3[1384] = 32'b00000000000000001001010100101111;
assign LUT_3[1385] = 32'b00000000000000010000000000001100;
assign LUT_3[1386] = 32'b00000000000000001011011100010011;
assign LUT_3[1387] = 32'b00000000000000010010000111110000;
assign LUT_3[1388] = 32'b00000000000000000110100010100101;
assign LUT_3[1389] = 32'b00000000000000001101001110000010;
assign LUT_3[1390] = 32'b00000000000000001000101010001001;
assign LUT_3[1391] = 32'b00000000000000001111010101100110;
assign LUT_3[1392] = 32'b00000000000000000111001110101100;
assign LUT_3[1393] = 32'b00000000000000001101111010001001;
assign LUT_3[1394] = 32'b00000000000000001001010110010000;
assign LUT_3[1395] = 32'b00000000000000010000000001101101;
assign LUT_3[1396] = 32'b00000000000000000100011100100010;
assign LUT_3[1397] = 32'b00000000000000001011000111111111;
assign LUT_3[1398] = 32'b00000000000000000110100100000110;
assign LUT_3[1399] = 32'b00000000000000001101001111100011;
assign LUT_3[1400] = 32'b00000000000000001100100111110010;
assign LUT_3[1401] = 32'b00000000000000010011010011001111;
assign LUT_3[1402] = 32'b00000000000000001110101111010110;
assign LUT_3[1403] = 32'b00000000000000010101011010110011;
assign LUT_3[1404] = 32'b00000000000000001001110101101000;
assign LUT_3[1405] = 32'b00000000000000010000100001000101;
assign LUT_3[1406] = 32'b00000000000000001011111101001100;
assign LUT_3[1407] = 32'b00000000000000010010101000101001;
assign LUT_3[1408] = 32'b00000000000000000100111111011100;
assign LUT_3[1409] = 32'b00000000000000001011101010111001;
assign LUT_3[1410] = 32'b00000000000000000111000111000000;
assign LUT_3[1411] = 32'b00000000000000001101110010011101;
assign LUT_3[1412] = 32'b00000000000000000010001101010010;
assign LUT_3[1413] = 32'b00000000000000001000111000101111;
assign LUT_3[1414] = 32'b00000000000000000100010100110110;
assign LUT_3[1415] = 32'b00000000000000001011000000010011;
assign LUT_3[1416] = 32'b00000000000000001010011000100010;
assign LUT_3[1417] = 32'b00000000000000010001000011111111;
assign LUT_3[1418] = 32'b00000000000000001100100000000110;
assign LUT_3[1419] = 32'b00000000000000010011001011100011;
assign LUT_3[1420] = 32'b00000000000000000111100110011000;
assign LUT_3[1421] = 32'b00000000000000001110010001110101;
assign LUT_3[1422] = 32'b00000000000000001001101101111100;
assign LUT_3[1423] = 32'b00000000000000010000011001011001;
assign LUT_3[1424] = 32'b00000000000000001000010010011111;
assign LUT_3[1425] = 32'b00000000000000001110111101111100;
assign LUT_3[1426] = 32'b00000000000000001010011010000011;
assign LUT_3[1427] = 32'b00000000000000010001000101100000;
assign LUT_3[1428] = 32'b00000000000000000101100000010101;
assign LUT_3[1429] = 32'b00000000000000001100001011110010;
assign LUT_3[1430] = 32'b00000000000000000111100111111001;
assign LUT_3[1431] = 32'b00000000000000001110010011010110;
assign LUT_3[1432] = 32'b00000000000000001101101011100101;
assign LUT_3[1433] = 32'b00000000000000010100010111000010;
assign LUT_3[1434] = 32'b00000000000000001111110011001001;
assign LUT_3[1435] = 32'b00000000000000010110011110100110;
assign LUT_3[1436] = 32'b00000000000000001010111001011011;
assign LUT_3[1437] = 32'b00000000000000010001100100111000;
assign LUT_3[1438] = 32'b00000000000000001101000000111111;
assign LUT_3[1439] = 32'b00000000000000010011101100011100;
assign LUT_3[1440] = 32'b00000000000000000110001101111100;
assign LUT_3[1441] = 32'b00000000000000001100111001011001;
assign LUT_3[1442] = 32'b00000000000000001000010101100000;
assign LUT_3[1443] = 32'b00000000000000001111000000111101;
assign LUT_3[1444] = 32'b00000000000000000011011011110010;
assign LUT_3[1445] = 32'b00000000000000001010000111001111;
assign LUT_3[1446] = 32'b00000000000000000101100011010110;
assign LUT_3[1447] = 32'b00000000000000001100001110110011;
assign LUT_3[1448] = 32'b00000000000000001011100111000010;
assign LUT_3[1449] = 32'b00000000000000010010010010011111;
assign LUT_3[1450] = 32'b00000000000000001101101110100110;
assign LUT_3[1451] = 32'b00000000000000010100011010000011;
assign LUT_3[1452] = 32'b00000000000000001000110100111000;
assign LUT_3[1453] = 32'b00000000000000001111100000010101;
assign LUT_3[1454] = 32'b00000000000000001010111100011100;
assign LUT_3[1455] = 32'b00000000000000010001100111111001;
assign LUT_3[1456] = 32'b00000000000000001001100000111111;
assign LUT_3[1457] = 32'b00000000000000010000001100011100;
assign LUT_3[1458] = 32'b00000000000000001011101000100011;
assign LUT_3[1459] = 32'b00000000000000010010010100000000;
assign LUT_3[1460] = 32'b00000000000000000110101110110101;
assign LUT_3[1461] = 32'b00000000000000001101011010010010;
assign LUT_3[1462] = 32'b00000000000000001000110110011001;
assign LUT_3[1463] = 32'b00000000000000001111100001110110;
assign LUT_3[1464] = 32'b00000000000000001110111010000101;
assign LUT_3[1465] = 32'b00000000000000010101100101100010;
assign LUT_3[1466] = 32'b00000000000000010001000001101001;
assign LUT_3[1467] = 32'b00000000000000010111101101000110;
assign LUT_3[1468] = 32'b00000000000000001100000111111011;
assign LUT_3[1469] = 32'b00000000000000010010110011011000;
assign LUT_3[1470] = 32'b00000000000000001110001111011111;
assign LUT_3[1471] = 32'b00000000000000010100111010111100;
assign LUT_3[1472] = 32'b00000000000000000100111000000111;
assign LUT_3[1473] = 32'b00000000000000001011100011100100;
assign LUT_3[1474] = 32'b00000000000000000110111111101011;
assign LUT_3[1475] = 32'b00000000000000001101101011001000;
assign LUT_3[1476] = 32'b00000000000000000010000101111101;
assign LUT_3[1477] = 32'b00000000000000001000110001011010;
assign LUT_3[1478] = 32'b00000000000000000100001101100001;
assign LUT_3[1479] = 32'b00000000000000001010111000111110;
assign LUT_3[1480] = 32'b00000000000000001010010001001101;
assign LUT_3[1481] = 32'b00000000000000010000111100101010;
assign LUT_3[1482] = 32'b00000000000000001100011000110001;
assign LUT_3[1483] = 32'b00000000000000010011000100001110;
assign LUT_3[1484] = 32'b00000000000000000111011111000011;
assign LUT_3[1485] = 32'b00000000000000001110001010100000;
assign LUT_3[1486] = 32'b00000000000000001001100110100111;
assign LUT_3[1487] = 32'b00000000000000010000010010000100;
assign LUT_3[1488] = 32'b00000000000000001000001011001010;
assign LUT_3[1489] = 32'b00000000000000001110110110100111;
assign LUT_3[1490] = 32'b00000000000000001010010010101110;
assign LUT_3[1491] = 32'b00000000000000010000111110001011;
assign LUT_3[1492] = 32'b00000000000000000101011001000000;
assign LUT_3[1493] = 32'b00000000000000001100000100011101;
assign LUT_3[1494] = 32'b00000000000000000111100000100100;
assign LUT_3[1495] = 32'b00000000000000001110001100000001;
assign LUT_3[1496] = 32'b00000000000000001101100100010000;
assign LUT_3[1497] = 32'b00000000000000010100001111101101;
assign LUT_3[1498] = 32'b00000000000000001111101011110100;
assign LUT_3[1499] = 32'b00000000000000010110010111010001;
assign LUT_3[1500] = 32'b00000000000000001010110010000110;
assign LUT_3[1501] = 32'b00000000000000010001011101100011;
assign LUT_3[1502] = 32'b00000000000000001100111001101010;
assign LUT_3[1503] = 32'b00000000000000010011100101000111;
assign LUT_3[1504] = 32'b00000000000000000110000110100111;
assign LUT_3[1505] = 32'b00000000000000001100110010000100;
assign LUT_3[1506] = 32'b00000000000000001000001110001011;
assign LUT_3[1507] = 32'b00000000000000001110111001101000;
assign LUT_3[1508] = 32'b00000000000000000011010100011101;
assign LUT_3[1509] = 32'b00000000000000001001111111111010;
assign LUT_3[1510] = 32'b00000000000000000101011100000001;
assign LUT_3[1511] = 32'b00000000000000001100000111011110;
assign LUT_3[1512] = 32'b00000000000000001011011111101101;
assign LUT_3[1513] = 32'b00000000000000010010001011001010;
assign LUT_3[1514] = 32'b00000000000000001101100111010001;
assign LUT_3[1515] = 32'b00000000000000010100010010101110;
assign LUT_3[1516] = 32'b00000000000000001000101101100011;
assign LUT_3[1517] = 32'b00000000000000001111011001000000;
assign LUT_3[1518] = 32'b00000000000000001010110101000111;
assign LUT_3[1519] = 32'b00000000000000010001100000100100;
assign LUT_3[1520] = 32'b00000000000000001001011001101010;
assign LUT_3[1521] = 32'b00000000000000010000000101000111;
assign LUT_3[1522] = 32'b00000000000000001011100001001110;
assign LUT_3[1523] = 32'b00000000000000010010001100101011;
assign LUT_3[1524] = 32'b00000000000000000110100111100000;
assign LUT_3[1525] = 32'b00000000000000001101010010111101;
assign LUT_3[1526] = 32'b00000000000000001000101111000100;
assign LUT_3[1527] = 32'b00000000000000001111011010100001;
assign LUT_3[1528] = 32'b00000000000000001110110010110000;
assign LUT_3[1529] = 32'b00000000000000010101011110001101;
assign LUT_3[1530] = 32'b00000000000000010000111010010100;
assign LUT_3[1531] = 32'b00000000000000010111100101110001;
assign LUT_3[1532] = 32'b00000000000000001100000000100110;
assign LUT_3[1533] = 32'b00000000000000010010101100000011;
assign LUT_3[1534] = 32'b00000000000000001110001000001010;
assign LUT_3[1535] = 32'b00000000000000010100110011100111;
assign LUT_3[1536] = 32'b00000000000000001001111010001001;
assign LUT_3[1537] = 32'b00000000000000010000100101100110;
assign LUT_3[1538] = 32'b00000000000000001100000001101101;
assign LUT_3[1539] = 32'b00000000000000010010101101001010;
assign LUT_3[1540] = 32'b00000000000000000111000111111111;
assign LUT_3[1541] = 32'b00000000000000001101110011011100;
assign LUT_3[1542] = 32'b00000000000000001001001111100011;
assign LUT_3[1543] = 32'b00000000000000001111111011000000;
assign LUT_3[1544] = 32'b00000000000000001111010011001111;
assign LUT_3[1545] = 32'b00000000000000010101111110101100;
assign LUT_3[1546] = 32'b00000000000000010001011010110011;
assign LUT_3[1547] = 32'b00000000000000011000000110010000;
assign LUT_3[1548] = 32'b00000000000000001100100001000101;
assign LUT_3[1549] = 32'b00000000000000010011001100100010;
assign LUT_3[1550] = 32'b00000000000000001110101000101001;
assign LUT_3[1551] = 32'b00000000000000010101010100000110;
assign LUT_3[1552] = 32'b00000000000000001101001101001100;
assign LUT_3[1553] = 32'b00000000000000010011111000101001;
assign LUT_3[1554] = 32'b00000000000000001111010100110000;
assign LUT_3[1555] = 32'b00000000000000010110000000001101;
assign LUT_3[1556] = 32'b00000000000000001010011011000010;
assign LUT_3[1557] = 32'b00000000000000010001000110011111;
assign LUT_3[1558] = 32'b00000000000000001100100010100110;
assign LUT_3[1559] = 32'b00000000000000010011001110000011;
assign LUT_3[1560] = 32'b00000000000000010010100110010010;
assign LUT_3[1561] = 32'b00000000000000011001010001101111;
assign LUT_3[1562] = 32'b00000000000000010100101101110110;
assign LUT_3[1563] = 32'b00000000000000011011011001010011;
assign LUT_3[1564] = 32'b00000000000000001111110100001000;
assign LUT_3[1565] = 32'b00000000000000010110011111100101;
assign LUT_3[1566] = 32'b00000000000000010001111011101100;
assign LUT_3[1567] = 32'b00000000000000011000100111001001;
assign LUT_3[1568] = 32'b00000000000000001011001000101001;
assign LUT_3[1569] = 32'b00000000000000010001110100000110;
assign LUT_3[1570] = 32'b00000000000000001101010000001101;
assign LUT_3[1571] = 32'b00000000000000010011111011101010;
assign LUT_3[1572] = 32'b00000000000000001000010110011111;
assign LUT_3[1573] = 32'b00000000000000001111000001111100;
assign LUT_3[1574] = 32'b00000000000000001010011110000011;
assign LUT_3[1575] = 32'b00000000000000010001001001100000;
assign LUT_3[1576] = 32'b00000000000000010000100001101111;
assign LUT_3[1577] = 32'b00000000000000010111001101001100;
assign LUT_3[1578] = 32'b00000000000000010010101001010011;
assign LUT_3[1579] = 32'b00000000000000011001010100110000;
assign LUT_3[1580] = 32'b00000000000000001101101111100101;
assign LUT_3[1581] = 32'b00000000000000010100011011000010;
assign LUT_3[1582] = 32'b00000000000000001111110111001001;
assign LUT_3[1583] = 32'b00000000000000010110100010100110;
assign LUT_3[1584] = 32'b00000000000000001110011011101100;
assign LUT_3[1585] = 32'b00000000000000010101000111001001;
assign LUT_3[1586] = 32'b00000000000000010000100011010000;
assign LUT_3[1587] = 32'b00000000000000010111001110101101;
assign LUT_3[1588] = 32'b00000000000000001011101001100010;
assign LUT_3[1589] = 32'b00000000000000010010010100111111;
assign LUT_3[1590] = 32'b00000000000000001101110001000110;
assign LUT_3[1591] = 32'b00000000000000010100011100100011;
assign LUT_3[1592] = 32'b00000000000000010011110100110010;
assign LUT_3[1593] = 32'b00000000000000011010100000001111;
assign LUT_3[1594] = 32'b00000000000000010101111100010110;
assign LUT_3[1595] = 32'b00000000000000011100100111110011;
assign LUT_3[1596] = 32'b00000000000000010001000010101000;
assign LUT_3[1597] = 32'b00000000000000010111101110000101;
assign LUT_3[1598] = 32'b00000000000000010011001010001100;
assign LUT_3[1599] = 32'b00000000000000011001110101101001;
assign LUT_3[1600] = 32'b00000000000000001001110010110100;
assign LUT_3[1601] = 32'b00000000000000010000011110010001;
assign LUT_3[1602] = 32'b00000000000000001011111010011000;
assign LUT_3[1603] = 32'b00000000000000010010100101110101;
assign LUT_3[1604] = 32'b00000000000000000111000000101010;
assign LUT_3[1605] = 32'b00000000000000001101101100000111;
assign LUT_3[1606] = 32'b00000000000000001001001000001110;
assign LUT_3[1607] = 32'b00000000000000001111110011101011;
assign LUT_3[1608] = 32'b00000000000000001111001011111010;
assign LUT_3[1609] = 32'b00000000000000010101110111010111;
assign LUT_3[1610] = 32'b00000000000000010001010011011110;
assign LUT_3[1611] = 32'b00000000000000010111111110111011;
assign LUT_3[1612] = 32'b00000000000000001100011001110000;
assign LUT_3[1613] = 32'b00000000000000010011000101001101;
assign LUT_3[1614] = 32'b00000000000000001110100001010100;
assign LUT_3[1615] = 32'b00000000000000010101001100110001;
assign LUT_3[1616] = 32'b00000000000000001101000101110111;
assign LUT_3[1617] = 32'b00000000000000010011110001010100;
assign LUT_3[1618] = 32'b00000000000000001111001101011011;
assign LUT_3[1619] = 32'b00000000000000010101111000111000;
assign LUT_3[1620] = 32'b00000000000000001010010011101101;
assign LUT_3[1621] = 32'b00000000000000010000111111001010;
assign LUT_3[1622] = 32'b00000000000000001100011011010001;
assign LUT_3[1623] = 32'b00000000000000010011000110101110;
assign LUT_3[1624] = 32'b00000000000000010010011110111101;
assign LUT_3[1625] = 32'b00000000000000011001001010011010;
assign LUT_3[1626] = 32'b00000000000000010100100110100001;
assign LUT_3[1627] = 32'b00000000000000011011010001111110;
assign LUT_3[1628] = 32'b00000000000000001111101100110011;
assign LUT_3[1629] = 32'b00000000000000010110011000010000;
assign LUT_3[1630] = 32'b00000000000000010001110100010111;
assign LUT_3[1631] = 32'b00000000000000011000011111110100;
assign LUT_3[1632] = 32'b00000000000000001011000001010100;
assign LUT_3[1633] = 32'b00000000000000010001101100110001;
assign LUT_3[1634] = 32'b00000000000000001101001000111000;
assign LUT_3[1635] = 32'b00000000000000010011110100010101;
assign LUT_3[1636] = 32'b00000000000000001000001111001010;
assign LUT_3[1637] = 32'b00000000000000001110111010100111;
assign LUT_3[1638] = 32'b00000000000000001010010110101110;
assign LUT_3[1639] = 32'b00000000000000010001000010001011;
assign LUT_3[1640] = 32'b00000000000000010000011010011010;
assign LUT_3[1641] = 32'b00000000000000010111000101110111;
assign LUT_3[1642] = 32'b00000000000000010010100001111110;
assign LUT_3[1643] = 32'b00000000000000011001001101011011;
assign LUT_3[1644] = 32'b00000000000000001101101000010000;
assign LUT_3[1645] = 32'b00000000000000010100010011101101;
assign LUT_3[1646] = 32'b00000000000000001111101111110100;
assign LUT_3[1647] = 32'b00000000000000010110011011010001;
assign LUT_3[1648] = 32'b00000000000000001110010100010111;
assign LUT_3[1649] = 32'b00000000000000010100111111110100;
assign LUT_3[1650] = 32'b00000000000000010000011011111011;
assign LUT_3[1651] = 32'b00000000000000010111000111011000;
assign LUT_3[1652] = 32'b00000000000000001011100010001101;
assign LUT_3[1653] = 32'b00000000000000010010001101101010;
assign LUT_3[1654] = 32'b00000000000000001101101001110001;
assign LUT_3[1655] = 32'b00000000000000010100010101001110;
assign LUT_3[1656] = 32'b00000000000000010011101101011101;
assign LUT_3[1657] = 32'b00000000000000011010011000111010;
assign LUT_3[1658] = 32'b00000000000000010101110101000001;
assign LUT_3[1659] = 32'b00000000000000011100100000011110;
assign LUT_3[1660] = 32'b00000000000000010000111011010011;
assign LUT_3[1661] = 32'b00000000000000010111100110110000;
assign LUT_3[1662] = 32'b00000000000000010011000010110111;
assign LUT_3[1663] = 32'b00000000000000011001101110010100;
assign LUT_3[1664] = 32'b00000000000000001100000101000111;
assign LUT_3[1665] = 32'b00000000000000010010110000100100;
assign LUT_3[1666] = 32'b00000000000000001110001100101011;
assign LUT_3[1667] = 32'b00000000000000010100111000001000;
assign LUT_3[1668] = 32'b00000000000000001001010010111101;
assign LUT_3[1669] = 32'b00000000000000001111111110011010;
assign LUT_3[1670] = 32'b00000000000000001011011010100001;
assign LUT_3[1671] = 32'b00000000000000010010000101111110;
assign LUT_3[1672] = 32'b00000000000000010001011110001101;
assign LUT_3[1673] = 32'b00000000000000011000001001101010;
assign LUT_3[1674] = 32'b00000000000000010011100101110001;
assign LUT_3[1675] = 32'b00000000000000011010010001001110;
assign LUT_3[1676] = 32'b00000000000000001110101100000011;
assign LUT_3[1677] = 32'b00000000000000010101010111100000;
assign LUT_3[1678] = 32'b00000000000000010000110011100111;
assign LUT_3[1679] = 32'b00000000000000010111011111000100;
assign LUT_3[1680] = 32'b00000000000000001111011000001010;
assign LUT_3[1681] = 32'b00000000000000010110000011100111;
assign LUT_3[1682] = 32'b00000000000000010001011111101110;
assign LUT_3[1683] = 32'b00000000000000011000001011001011;
assign LUT_3[1684] = 32'b00000000000000001100100110000000;
assign LUT_3[1685] = 32'b00000000000000010011010001011101;
assign LUT_3[1686] = 32'b00000000000000001110101101100100;
assign LUT_3[1687] = 32'b00000000000000010101011001000001;
assign LUT_3[1688] = 32'b00000000000000010100110001010000;
assign LUT_3[1689] = 32'b00000000000000011011011100101101;
assign LUT_3[1690] = 32'b00000000000000010110111000110100;
assign LUT_3[1691] = 32'b00000000000000011101100100010001;
assign LUT_3[1692] = 32'b00000000000000010001111111000110;
assign LUT_3[1693] = 32'b00000000000000011000101010100011;
assign LUT_3[1694] = 32'b00000000000000010100000110101010;
assign LUT_3[1695] = 32'b00000000000000011010110010000111;
assign LUT_3[1696] = 32'b00000000000000001101010011100111;
assign LUT_3[1697] = 32'b00000000000000010011111111000100;
assign LUT_3[1698] = 32'b00000000000000001111011011001011;
assign LUT_3[1699] = 32'b00000000000000010110000110101000;
assign LUT_3[1700] = 32'b00000000000000001010100001011101;
assign LUT_3[1701] = 32'b00000000000000010001001100111010;
assign LUT_3[1702] = 32'b00000000000000001100101001000001;
assign LUT_3[1703] = 32'b00000000000000010011010100011110;
assign LUT_3[1704] = 32'b00000000000000010010101100101101;
assign LUT_3[1705] = 32'b00000000000000011001011000001010;
assign LUT_3[1706] = 32'b00000000000000010100110100010001;
assign LUT_3[1707] = 32'b00000000000000011011011111101110;
assign LUT_3[1708] = 32'b00000000000000001111111010100011;
assign LUT_3[1709] = 32'b00000000000000010110100110000000;
assign LUT_3[1710] = 32'b00000000000000010010000010000111;
assign LUT_3[1711] = 32'b00000000000000011000101101100100;
assign LUT_3[1712] = 32'b00000000000000010000100110101010;
assign LUT_3[1713] = 32'b00000000000000010111010010000111;
assign LUT_3[1714] = 32'b00000000000000010010101110001110;
assign LUT_3[1715] = 32'b00000000000000011001011001101011;
assign LUT_3[1716] = 32'b00000000000000001101110100100000;
assign LUT_3[1717] = 32'b00000000000000010100011111111101;
assign LUT_3[1718] = 32'b00000000000000001111111100000100;
assign LUT_3[1719] = 32'b00000000000000010110100111100001;
assign LUT_3[1720] = 32'b00000000000000010101111111110000;
assign LUT_3[1721] = 32'b00000000000000011100101011001101;
assign LUT_3[1722] = 32'b00000000000000011000000111010100;
assign LUT_3[1723] = 32'b00000000000000011110110010110001;
assign LUT_3[1724] = 32'b00000000000000010011001101100110;
assign LUT_3[1725] = 32'b00000000000000011001111001000011;
assign LUT_3[1726] = 32'b00000000000000010101010101001010;
assign LUT_3[1727] = 32'b00000000000000011100000000100111;
assign LUT_3[1728] = 32'b00000000000000001011111101110010;
assign LUT_3[1729] = 32'b00000000000000010010101001001111;
assign LUT_3[1730] = 32'b00000000000000001110000101010110;
assign LUT_3[1731] = 32'b00000000000000010100110000110011;
assign LUT_3[1732] = 32'b00000000000000001001001011101000;
assign LUT_3[1733] = 32'b00000000000000001111110111000101;
assign LUT_3[1734] = 32'b00000000000000001011010011001100;
assign LUT_3[1735] = 32'b00000000000000010001111110101001;
assign LUT_3[1736] = 32'b00000000000000010001010110111000;
assign LUT_3[1737] = 32'b00000000000000011000000010010101;
assign LUT_3[1738] = 32'b00000000000000010011011110011100;
assign LUT_3[1739] = 32'b00000000000000011010001001111001;
assign LUT_3[1740] = 32'b00000000000000001110100100101110;
assign LUT_3[1741] = 32'b00000000000000010101010000001011;
assign LUT_3[1742] = 32'b00000000000000010000101100010010;
assign LUT_3[1743] = 32'b00000000000000010111010111101111;
assign LUT_3[1744] = 32'b00000000000000001111010000110101;
assign LUT_3[1745] = 32'b00000000000000010101111100010010;
assign LUT_3[1746] = 32'b00000000000000010001011000011001;
assign LUT_3[1747] = 32'b00000000000000011000000011110110;
assign LUT_3[1748] = 32'b00000000000000001100011110101011;
assign LUT_3[1749] = 32'b00000000000000010011001010001000;
assign LUT_3[1750] = 32'b00000000000000001110100110001111;
assign LUT_3[1751] = 32'b00000000000000010101010001101100;
assign LUT_3[1752] = 32'b00000000000000010100101001111011;
assign LUT_3[1753] = 32'b00000000000000011011010101011000;
assign LUT_3[1754] = 32'b00000000000000010110110001011111;
assign LUT_3[1755] = 32'b00000000000000011101011100111100;
assign LUT_3[1756] = 32'b00000000000000010001110111110001;
assign LUT_3[1757] = 32'b00000000000000011000100011001110;
assign LUT_3[1758] = 32'b00000000000000010011111111010101;
assign LUT_3[1759] = 32'b00000000000000011010101010110010;
assign LUT_3[1760] = 32'b00000000000000001101001100010010;
assign LUT_3[1761] = 32'b00000000000000010011110111101111;
assign LUT_3[1762] = 32'b00000000000000001111010011110110;
assign LUT_3[1763] = 32'b00000000000000010101111111010011;
assign LUT_3[1764] = 32'b00000000000000001010011010001000;
assign LUT_3[1765] = 32'b00000000000000010001000101100101;
assign LUT_3[1766] = 32'b00000000000000001100100001101100;
assign LUT_3[1767] = 32'b00000000000000010011001101001001;
assign LUT_3[1768] = 32'b00000000000000010010100101011000;
assign LUT_3[1769] = 32'b00000000000000011001010000110101;
assign LUT_3[1770] = 32'b00000000000000010100101100111100;
assign LUT_3[1771] = 32'b00000000000000011011011000011001;
assign LUT_3[1772] = 32'b00000000000000001111110011001110;
assign LUT_3[1773] = 32'b00000000000000010110011110101011;
assign LUT_3[1774] = 32'b00000000000000010001111010110010;
assign LUT_3[1775] = 32'b00000000000000011000100110001111;
assign LUT_3[1776] = 32'b00000000000000010000011111010101;
assign LUT_3[1777] = 32'b00000000000000010111001010110010;
assign LUT_3[1778] = 32'b00000000000000010010100110111001;
assign LUT_3[1779] = 32'b00000000000000011001010010010110;
assign LUT_3[1780] = 32'b00000000000000001101101101001011;
assign LUT_3[1781] = 32'b00000000000000010100011000101000;
assign LUT_3[1782] = 32'b00000000000000001111110100101111;
assign LUT_3[1783] = 32'b00000000000000010110100000001100;
assign LUT_3[1784] = 32'b00000000000000010101111000011011;
assign LUT_3[1785] = 32'b00000000000000011100100011111000;
assign LUT_3[1786] = 32'b00000000000000010111111111111111;
assign LUT_3[1787] = 32'b00000000000000011110101011011100;
assign LUT_3[1788] = 32'b00000000000000010011000110010001;
assign LUT_3[1789] = 32'b00000000000000011001110001101110;
assign LUT_3[1790] = 32'b00000000000000010101001101110101;
assign LUT_3[1791] = 32'b00000000000000011011111001010010;
assign LUT_3[1792] = 32'b00000000000000000110001001101010;
assign LUT_3[1793] = 32'b00000000000000001100110101000111;
assign LUT_3[1794] = 32'b00000000000000001000010001001110;
assign LUT_3[1795] = 32'b00000000000000001110111100101011;
assign LUT_3[1796] = 32'b00000000000000000011010111100000;
assign LUT_3[1797] = 32'b00000000000000001010000010111101;
assign LUT_3[1798] = 32'b00000000000000000101011111000100;
assign LUT_3[1799] = 32'b00000000000000001100001010100001;
assign LUT_3[1800] = 32'b00000000000000001011100010110000;
assign LUT_3[1801] = 32'b00000000000000010010001110001101;
assign LUT_3[1802] = 32'b00000000000000001101101010010100;
assign LUT_3[1803] = 32'b00000000000000010100010101110001;
assign LUT_3[1804] = 32'b00000000000000001000110000100110;
assign LUT_3[1805] = 32'b00000000000000001111011100000011;
assign LUT_3[1806] = 32'b00000000000000001010111000001010;
assign LUT_3[1807] = 32'b00000000000000010001100011100111;
assign LUT_3[1808] = 32'b00000000000000001001011100101101;
assign LUT_3[1809] = 32'b00000000000000010000001000001010;
assign LUT_3[1810] = 32'b00000000000000001011100100010001;
assign LUT_3[1811] = 32'b00000000000000010010001111101110;
assign LUT_3[1812] = 32'b00000000000000000110101010100011;
assign LUT_3[1813] = 32'b00000000000000001101010110000000;
assign LUT_3[1814] = 32'b00000000000000001000110010000111;
assign LUT_3[1815] = 32'b00000000000000001111011101100100;
assign LUT_3[1816] = 32'b00000000000000001110110101110011;
assign LUT_3[1817] = 32'b00000000000000010101100001010000;
assign LUT_3[1818] = 32'b00000000000000010000111101010111;
assign LUT_3[1819] = 32'b00000000000000010111101000110100;
assign LUT_3[1820] = 32'b00000000000000001100000011101001;
assign LUT_3[1821] = 32'b00000000000000010010101111000110;
assign LUT_3[1822] = 32'b00000000000000001110001011001101;
assign LUT_3[1823] = 32'b00000000000000010100110110101010;
assign LUT_3[1824] = 32'b00000000000000000111011000001010;
assign LUT_3[1825] = 32'b00000000000000001110000011100111;
assign LUT_3[1826] = 32'b00000000000000001001011111101110;
assign LUT_3[1827] = 32'b00000000000000010000001011001011;
assign LUT_3[1828] = 32'b00000000000000000100100110000000;
assign LUT_3[1829] = 32'b00000000000000001011010001011101;
assign LUT_3[1830] = 32'b00000000000000000110101101100100;
assign LUT_3[1831] = 32'b00000000000000001101011001000001;
assign LUT_3[1832] = 32'b00000000000000001100110001010000;
assign LUT_3[1833] = 32'b00000000000000010011011100101101;
assign LUT_3[1834] = 32'b00000000000000001110111000110100;
assign LUT_3[1835] = 32'b00000000000000010101100100010001;
assign LUT_3[1836] = 32'b00000000000000001001111111000110;
assign LUT_3[1837] = 32'b00000000000000010000101010100011;
assign LUT_3[1838] = 32'b00000000000000001100000110101010;
assign LUT_3[1839] = 32'b00000000000000010010110010000111;
assign LUT_3[1840] = 32'b00000000000000001010101011001101;
assign LUT_3[1841] = 32'b00000000000000010001010110101010;
assign LUT_3[1842] = 32'b00000000000000001100110010110001;
assign LUT_3[1843] = 32'b00000000000000010011011110001110;
assign LUT_3[1844] = 32'b00000000000000000111111001000011;
assign LUT_3[1845] = 32'b00000000000000001110100100100000;
assign LUT_3[1846] = 32'b00000000000000001010000000100111;
assign LUT_3[1847] = 32'b00000000000000010000101100000100;
assign LUT_3[1848] = 32'b00000000000000010000000100010011;
assign LUT_3[1849] = 32'b00000000000000010110101111110000;
assign LUT_3[1850] = 32'b00000000000000010010001011110111;
assign LUT_3[1851] = 32'b00000000000000011000110111010100;
assign LUT_3[1852] = 32'b00000000000000001101010010001001;
assign LUT_3[1853] = 32'b00000000000000010011111101100110;
assign LUT_3[1854] = 32'b00000000000000001111011001101101;
assign LUT_3[1855] = 32'b00000000000000010110000101001010;
assign LUT_3[1856] = 32'b00000000000000000110000010010101;
assign LUT_3[1857] = 32'b00000000000000001100101101110010;
assign LUT_3[1858] = 32'b00000000000000001000001001111001;
assign LUT_3[1859] = 32'b00000000000000001110110101010110;
assign LUT_3[1860] = 32'b00000000000000000011010000001011;
assign LUT_3[1861] = 32'b00000000000000001001111011101000;
assign LUT_3[1862] = 32'b00000000000000000101010111101111;
assign LUT_3[1863] = 32'b00000000000000001100000011001100;
assign LUT_3[1864] = 32'b00000000000000001011011011011011;
assign LUT_3[1865] = 32'b00000000000000010010000110111000;
assign LUT_3[1866] = 32'b00000000000000001101100010111111;
assign LUT_3[1867] = 32'b00000000000000010100001110011100;
assign LUT_3[1868] = 32'b00000000000000001000101001010001;
assign LUT_3[1869] = 32'b00000000000000001111010100101110;
assign LUT_3[1870] = 32'b00000000000000001010110000110101;
assign LUT_3[1871] = 32'b00000000000000010001011100010010;
assign LUT_3[1872] = 32'b00000000000000001001010101011000;
assign LUT_3[1873] = 32'b00000000000000010000000000110101;
assign LUT_3[1874] = 32'b00000000000000001011011100111100;
assign LUT_3[1875] = 32'b00000000000000010010001000011001;
assign LUT_3[1876] = 32'b00000000000000000110100011001110;
assign LUT_3[1877] = 32'b00000000000000001101001110101011;
assign LUT_3[1878] = 32'b00000000000000001000101010110010;
assign LUT_3[1879] = 32'b00000000000000001111010110001111;
assign LUT_3[1880] = 32'b00000000000000001110101110011110;
assign LUT_3[1881] = 32'b00000000000000010101011001111011;
assign LUT_3[1882] = 32'b00000000000000010000110110000010;
assign LUT_3[1883] = 32'b00000000000000010111100001011111;
assign LUT_3[1884] = 32'b00000000000000001011111100010100;
assign LUT_3[1885] = 32'b00000000000000010010100111110001;
assign LUT_3[1886] = 32'b00000000000000001110000011111000;
assign LUT_3[1887] = 32'b00000000000000010100101111010101;
assign LUT_3[1888] = 32'b00000000000000000111010000110101;
assign LUT_3[1889] = 32'b00000000000000001101111100010010;
assign LUT_3[1890] = 32'b00000000000000001001011000011001;
assign LUT_3[1891] = 32'b00000000000000010000000011110110;
assign LUT_3[1892] = 32'b00000000000000000100011110101011;
assign LUT_3[1893] = 32'b00000000000000001011001010001000;
assign LUT_3[1894] = 32'b00000000000000000110100110001111;
assign LUT_3[1895] = 32'b00000000000000001101010001101100;
assign LUT_3[1896] = 32'b00000000000000001100101001111011;
assign LUT_3[1897] = 32'b00000000000000010011010101011000;
assign LUT_3[1898] = 32'b00000000000000001110110001011111;
assign LUT_3[1899] = 32'b00000000000000010101011100111100;
assign LUT_3[1900] = 32'b00000000000000001001110111110001;
assign LUT_3[1901] = 32'b00000000000000010000100011001110;
assign LUT_3[1902] = 32'b00000000000000001011111111010101;
assign LUT_3[1903] = 32'b00000000000000010010101010110010;
assign LUT_3[1904] = 32'b00000000000000001010100011111000;
assign LUT_3[1905] = 32'b00000000000000010001001111010101;
assign LUT_3[1906] = 32'b00000000000000001100101011011100;
assign LUT_3[1907] = 32'b00000000000000010011010110111001;
assign LUT_3[1908] = 32'b00000000000000000111110001101110;
assign LUT_3[1909] = 32'b00000000000000001110011101001011;
assign LUT_3[1910] = 32'b00000000000000001001111001010010;
assign LUT_3[1911] = 32'b00000000000000010000100100101111;
assign LUT_3[1912] = 32'b00000000000000001111111100111110;
assign LUT_3[1913] = 32'b00000000000000010110101000011011;
assign LUT_3[1914] = 32'b00000000000000010010000100100010;
assign LUT_3[1915] = 32'b00000000000000011000101111111111;
assign LUT_3[1916] = 32'b00000000000000001101001010110100;
assign LUT_3[1917] = 32'b00000000000000010011110110010001;
assign LUT_3[1918] = 32'b00000000000000001111010010011000;
assign LUT_3[1919] = 32'b00000000000000010101111101110101;
assign LUT_3[1920] = 32'b00000000000000001000010100101000;
assign LUT_3[1921] = 32'b00000000000000001111000000000101;
assign LUT_3[1922] = 32'b00000000000000001010011100001100;
assign LUT_3[1923] = 32'b00000000000000010001000111101001;
assign LUT_3[1924] = 32'b00000000000000000101100010011110;
assign LUT_3[1925] = 32'b00000000000000001100001101111011;
assign LUT_3[1926] = 32'b00000000000000000111101010000010;
assign LUT_3[1927] = 32'b00000000000000001110010101011111;
assign LUT_3[1928] = 32'b00000000000000001101101101101110;
assign LUT_3[1929] = 32'b00000000000000010100011001001011;
assign LUT_3[1930] = 32'b00000000000000001111110101010010;
assign LUT_3[1931] = 32'b00000000000000010110100000101111;
assign LUT_3[1932] = 32'b00000000000000001010111011100100;
assign LUT_3[1933] = 32'b00000000000000010001100111000001;
assign LUT_3[1934] = 32'b00000000000000001101000011001000;
assign LUT_3[1935] = 32'b00000000000000010011101110100101;
assign LUT_3[1936] = 32'b00000000000000001011100111101011;
assign LUT_3[1937] = 32'b00000000000000010010010011001000;
assign LUT_3[1938] = 32'b00000000000000001101101111001111;
assign LUT_3[1939] = 32'b00000000000000010100011010101100;
assign LUT_3[1940] = 32'b00000000000000001000110101100001;
assign LUT_3[1941] = 32'b00000000000000001111100000111110;
assign LUT_3[1942] = 32'b00000000000000001010111101000101;
assign LUT_3[1943] = 32'b00000000000000010001101000100010;
assign LUT_3[1944] = 32'b00000000000000010001000000110001;
assign LUT_3[1945] = 32'b00000000000000010111101100001110;
assign LUT_3[1946] = 32'b00000000000000010011001000010101;
assign LUT_3[1947] = 32'b00000000000000011001110011110010;
assign LUT_3[1948] = 32'b00000000000000001110001110100111;
assign LUT_3[1949] = 32'b00000000000000010100111010000100;
assign LUT_3[1950] = 32'b00000000000000010000010110001011;
assign LUT_3[1951] = 32'b00000000000000010111000001101000;
assign LUT_3[1952] = 32'b00000000000000001001100011001000;
assign LUT_3[1953] = 32'b00000000000000010000001110100101;
assign LUT_3[1954] = 32'b00000000000000001011101010101100;
assign LUT_3[1955] = 32'b00000000000000010010010110001001;
assign LUT_3[1956] = 32'b00000000000000000110110000111110;
assign LUT_3[1957] = 32'b00000000000000001101011100011011;
assign LUT_3[1958] = 32'b00000000000000001000111000100010;
assign LUT_3[1959] = 32'b00000000000000001111100011111111;
assign LUT_3[1960] = 32'b00000000000000001110111100001110;
assign LUT_3[1961] = 32'b00000000000000010101100111101011;
assign LUT_3[1962] = 32'b00000000000000010001000011110010;
assign LUT_3[1963] = 32'b00000000000000010111101111001111;
assign LUT_3[1964] = 32'b00000000000000001100001010000100;
assign LUT_3[1965] = 32'b00000000000000010010110101100001;
assign LUT_3[1966] = 32'b00000000000000001110010001101000;
assign LUT_3[1967] = 32'b00000000000000010100111101000101;
assign LUT_3[1968] = 32'b00000000000000001100110110001011;
assign LUT_3[1969] = 32'b00000000000000010011100001101000;
assign LUT_3[1970] = 32'b00000000000000001110111101101111;
assign LUT_3[1971] = 32'b00000000000000010101101001001100;
assign LUT_3[1972] = 32'b00000000000000001010000100000001;
assign LUT_3[1973] = 32'b00000000000000010000101111011110;
assign LUT_3[1974] = 32'b00000000000000001100001011100101;
assign LUT_3[1975] = 32'b00000000000000010010110111000010;
assign LUT_3[1976] = 32'b00000000000000010010001111010001;
assign LUT_3[1977] = 32'b00000000000000011000111010101110;
assign LUT_3[1978] = 32'b00000000000000010100010110110101;
assign LUT_3[1979] = 32'b00000000000000011011000010010010;
assign LUT_3[1980] = 32'b00000000000000001111011101000111;
assign LUT_3[1981] = 32'b00000000000000010110001000100100;
assign LUT_3[1982] = 32'b00000000000000010001100100101011;
assign LUT_3[1983] = 32'b00000000000000011000010000001000;
assign LUT_3[1984] = 32'b00000000000000001000001101010011;
assign LUT_3[1985] = 32'b00000000000000001110111000110000;
assign LUT_3[1986] = 32'b00000000000000001010010100110111;
assign LUT_3[1987] = 32'b00000000000000010001000000010100;
assign LUT_3[1988] = 32'b00000000000000000101011011001001;
assign LUT_3[1989] = 32'b00000000000000001100000110100110;
assign LUT_3[1990] = 32'b00000000000000000111100010101101;
assign LUT_3[1991] = 32'b00000000000000001110001110001010;
assign LUT_3[1992] = 32'b00000000000000001101100110011001;
assign LUT_3[1993] = 32'b00000000000000010100010001110110;
assign LUT_3[1994] = 32'b00000000000000001111101101111101;
assign LUT_3[1995] = 32'b00000000000000010110011001011010;
assign LUT_3[1996] = 32'b00000000000000001010110100001111;
assign LUT_3[1997] = 32'b00000000000000010001011111101100;
assign LUT_3[1998] = 32'b00000000000000001100111011110011;
assign LUT_3[1999] = 32'b00000000000000010011100111010000;
assign LUT_3[2000] = 32'b00000000000000001011100000010110;
assign LUT_3[2001] = 32'b00000000000000010010001011110011;
assign LUT_3[2002] = 32'b00000000000000001101100111111010;
assign LUT_3[2003] = 32'b00000000000000010100010011010111;
assign LUT_3[2004] = 32'b00000000000000001000101110001100;
assign LUT_3[2005] = 32'b00000000000000001111011001101001;
assign LUT_3[2006] = 32'b00000000000000001010110101110000;
assign LUT_3[2007] = 32'b00000000000000010001100001001101;
assign LUT_3[2008] = 32'b00000000000000010000111001011100;
assign LUT_3[2009] = 32'b00000000000000010111100100111001;
assign LUT_3[2010] = 32'b00000000000000010011000001000000;
assign LUT_3[2011] = 32'b00000000000000011001101100011101;
assign LUT_3[2012] = 32'b00000000000000001110000111010010;
assign LUT_3[2013] = 32'b00000000000000010100110010101111;
assign LUT_3[2014] = 32'b00000000000000010000001110110110;
assign LUT_3[2015] = 32'b00000000000000010110111010010011;
assign LUT_3[2016] = 32'b00000000000000001001011011110011;
assign LUT_3[2017] = 32'b00000000000000010000000111010000;
assign LUT_3[2018] = 32'b00000000000000001011100011010111;
assign LUT_3[2019] = 32'b00000000000000010010001110110100;
assign LUT_3[2020] = 32'b00000000000000000110101001101001;
assign LUT_3[2021] = 32'b00000000000000001101010101000110;
assign LUT_3[2022] = 32'b00000000000000001000110001001101;
assign LUT_3[2023] = 32'b00000000000000001111011100101010;
assign LUT_3[2024] = 32'b00000000000000001110110100111001;
assign LUT_3[2025] = 32'b00000000000000010101100000010110;
assign LUT_3[2026] = 32'b00000000000000010000111100011101;
assign LUT_3[2027] = 32'b00000000000000010111100111111010;
assign LUT_3[2028] = 32'b00000000000000001100000010101111;
assign LUT_3[2029] = 32'b00000000000000010010101110001100;
assign LUT_3[2030] = 32'b00000000000000001110001010010011;
assign LUT_3[2031] = 32'b00000000000000010100110101110000;
assign LUT_3[2032] = 32'b00000000000000001100101110110110;
assign LUT_3[2033] = 32'b00000000000000010011011010010011;
assign LUT_3[2034] = 32'b00000000000000001110110110011010;
assign LUT_3[2035] = 32'b00000000000000010101100001110111;
assign LUT_3[2036] = 32'b00000000000000001001111100101100;
assign LUT_3[2037] = 32'b00000000000000010000101000001001;
assign LUT_3[2038] = 32'b00000000000000001100000100010000;
assign LUT_3[2039] = 32'b00000000000000010010101111101101;
assign LUT_3[2040] = 32'b00000000000000010010000111111100;
assign LUT_3[2041] = 32'b00000000000000011000110011011001;
assign LUT_3[2042] = 32'b00000000000000010100001111100000;
assign LUT_3[2043] = 32'b00000000000000011010111010111101;
assign LUT_3[2044] = 32'b00000000000000001111010101110010;
assign LUT_3[2045] = 32'b00000000000000010110000001001111;
assign LUT_3[2046] = 32'b00000000000000010001011101010110;
assign LUT_3[2047] = 32'b00000000000000011000001000110011;
assign LUT_3[2048] = 32'b00000000000000000001110110001110;
assign LUT_3[2049] = 32'b00000000000000001000100001101011;
assign LUT_3[2050] = 32'b00000000000000000011111101110010;
assign LUT_3[2051] = 32'b00000000000000001010101001001111;
assign LUT_3[2052] = 32'b11111111111111111111000100000100;
assign LUT_3[2053] = 32'b00000000000000000101101111100001;
assign LUT_3[2054] = 32'b00000000000000000001001011101000;
assign LUT_3[2055] = 32'b00000000000000000111110111000101;
assign LUT_3[2056] = 32'b00000000000000000111001111010100;
assign LUT_3[2057] = 32'b00000000000000001101111010110001;
assign LUT_3[2058] = 32'b00000000000000001001010110111000;
assign LUT_3[2059] = 32'b00000000000000010000000010010101;
assign LUT_3[2060] = 32'b00000000000000000100011101001010;
assign LUT_3[2061] = 32'b00000000000000001011001000100111;
assign LUT_3[2062] = 32'b00000000000000000110100100101110;
assign LUT_3[2063] = 32'b00000000000000001101010000001011;
assign LUT_3[2064] = 32'b00000000000000000101001001010001;
assign LUT_3[2065] = 32'b00000000000000001011110100101110;
assign LUT_3[2066] = 32'b00000000000000000111010000110101;
assign LUT_3[2067] = 32'b00000000000000001101111100010010;
assign LUT_3[2068] = 32'b00000000000000000010010111000111;
assign LUT_3[2069] = 32'b00000000000000001001000010100100;
assign LUT_3[2070] = 32'b00000000000000000100011110101011;
assign LUT_3[2071] = 32'b00000000000000001011001010001000;
assign LUT_3[2072] = 32'b00000000000000001010100010010111;
assign LUT_3[2073] = 32'b00000000000000010001001101110100;
assign LUT_3[2074] = 32'b00000000000000001100101001111011;
assign LUT_3[2075] = 32'b00000000000000010011010101011000;
assign LUT_3[2076] = 32'b00000000000000000111110000001101;
assign LUT_3[2077] = 32'b00000000000000001110011011101010;
assign LUT_3[2078] = 32'b00000000000000001001110111110001;
assign LUT_3[2079] = 32'b00000000000000010000100011001110;
assign LUT_3[2080] = 32'b00000000000000000011000100101110;
assign LUT_3[2081] = 32'b00000000000000001001110000001011;
assign LUT_3[2082] = 32'b00000000000000000101001100010010;
assign LUT_3[2083] = 32'b00000000000000001011110111101111;
assign LUT_3[2084] = 32'b00000000000000000000010010100100;
assign LUT_3[2085] = 32'b00000000000000000110111110000001;
assign LUT_3[2086] = 32'b00000000000000000010011010001000;
assign LUT_3[2087] = 32'b00000000000000001001000101100101;
assign LUT_3[2088] = 32'b00000000000000001000011101110100;
assign LUT_3[2089] = 32'b00000000000000001111001001010001;
assign LUT_3[2090] = 32'b00000000000000001010100101011000;
assign LUT_3[2091] = 32'b00000000000000010001010000110101;
assign LUT_3[2092] = 32'b00000000000000000101101011101010;
assign LUT_3[2093] = 32'b00000000000000001100010111000111;
assign LUT_3[2094] = 32'b00000000000000000111110011001110;
assign LUT_3[2095] = 32'b00000000000000001110011110101011;
assign LUT_3[2096] = 32'b00000000000000000110010111110001;
assign LUT_3[2097] = 32'b00000000000000001101000011001110;
assign LUT_3[2098] = 32'b00000000000000001000011111010101;
assign LUT_3[2099] = 32'b00000000000000001111001010110010;
assign LUT_3[2100] = 32'b00000000000000000011100101100111;
assign LUT_3[2101] = 32'b00000000000000001010010001000100;
assign LUT_3[2102] = 32'b00000000000000000101101101001011;
assign LUT_3[2103] = 32'b00000000000000001100011000101000;
assign LUT_3[2104] = 32'b00000000000000001011110000110111;
assign LUT_3[2105] = 32'b00000000000000010010011100010100;
assign LUT_3[2106] = 32'b00000000000000001101111000011011;
assign LUT_3[2107] = 32'b00000000000000010100100011111000;
assign LUT_3[2108] = 32'b00000000000000001000111110101101;
assign LUT_3[2109] = 32'b00000000000000001111101010001010;
assign LUT_3[2110] = 32'b00000000000000001011000110010001;
assign LUT_3[2111] = 32'b00000000000000010001110001101110;
assign LUT_3[2112] = 32'b00000000000000000001101110111001;
assign LUT_3[2113] = 32'b00000000000000001000011010010110;
assign LUT_3[2114] = 32'b00000000000000000011110110011101;
assign LUT_3[2115] = 32'b00000000000000001010100001111010;
assign LUT_3[2116] = 32'b11111111111111111110111100101111;
assign LUT_3[2117] = 32'b00000000000000000101101000001100;
assign LUT_3[2118] = 32'b00000000000000000001000100010011;
assign LUT_3[2119] = 32'b00000000000000000111101111110000;
assign LUT_3[2120] = 32'b00000000000000000111000111111111;
assign LUT_3[2121] = 32'b00000000000000001101110011011100;
assign LUT_3[2122] = 32'b00000000000000001001001111100011;
assign LUT_3[2123] = 32'b00000000000000001111111011000000;
assign LUT_3[2124] = 32'b00000000000000000100010101110101;
assign LUT_3[2125] = 32'b00000000000000001011000001010010;
assign LUT_3[2126] = 32'b00000000000000000110011101011001;
assign LUT_3[2127] = 32'b00000000000000001101001000110110;
assign LUT_3[2128] = 32'b00000000000000000101000001111100;
assign LUT_3[2129] = 32'b00000000000000001011101101011001;
assign LUT_3[2130] = 32'b00000000000000000111001001100000;
assign LUT_3[2131] = 32'b00000000000000001101110100111101;
assign LUT_3[2132] = 32'b00000000000000000010001111110010;
assign LUT_3[2133] = 32'b00000000000000001000111011001111;
assign LUT_3[2134] = 32'b00000000000000000100010111010110;
assign LUT_3[2135] = 32'b00000000000000001011000010110011;
assign LUT_3[2136] = 32'b00000000000000001010011011000010;
assign LUT_3[2137] = 32'b00000000000000010001000110011111;
assign LUT_3[2138] = 32'b00000000000000001100100010100110;
assign LUT_3[2139] = 32'b00000000000000010011001110000011;
assign LUT_3[2140] = 32'b00000000000000000111101000111000;
assign LUT_3[2141] = 32'b00000000000000001110010100010101;
assign LUT_3[2142] = 32'b00000000000000001001110000011100;
assign LUT_3[2143] = 32'b00000000000000010000011011111001;
assign LUT_3[2144] = 32'b00000000000000000010111101011001;
assign LUT_3[2145] = 32'b00000000000000001001101000110110;
assign LUT_3[2146] = 32'b00000000000000000101000100111101;
assign LUT_3[2147] = 32'b00000000000000001011110000011010;
assign LUT_3[2148] = 32'b00000000000000000000001011001111;
assign LUT_3[2149] = 32'b00000000000000000110110110101100;
assign LUT_3[2150] = 32'b00000000000000000010010010110011;
assign LUT_3[2151] = 32'b00000000000000001000111110010000;
assign LUT_3[2152] = 32'b00000000000000001000010110011111;
assign LUT_3[2153] = 32'b00000000000000001111000001111100;
assign LUT_3[2154] = 32'b00000000000000001010011110000011;
assign LUT_3[2155] = 32'b00000000000000010001001001100000;
assign LUT_3[2156] = 32'b00000000000000000101100100010101;
assign LUT_3[2157] = 32'b00000000000000001100001111110010;
assign LUT_3[2158] = 32'b00000000000000000111101011111001;
assign LUT_3[2159] = 32'b00000000000000001110010111010110;
assign LUT_3[2160] = 32'b00000000000000000110010000011100;
assign LUT_3[2161] = 32'b00000000000000001100111011111001;
assign LUT_3[2162] = 32'b00000000000000001000011000000000;
assign LUT_3[2163] = 32'b00000000000000001111000011011101;
assign LUT_3[2164] = 32'b00000000000000000011011110010010;
assign LUT_3[2165] = 32'b00000000000000001010001001101111;
assign LUT_3[2166] = 32'b00000000000000000101100101110110;
assign LUT_3[2167] = 32'b00000000000000001100010001010011;
assign LUT_3[2168] = 32'b00000000000000001011101001100010;
assign LUT_3[2169] = 32'b00000000000000010010010100111111;
assign LUT_3[2170] = 32'b00000000000000001101110001000110;
assign LUT_3[2171] = 32'b00000000000000010100011100100011;
assign LUT_3[2172] = 32'b00000000000000001000110111011000;
assign LUT_3[2173] = 32'b00000000000000001111100010110101;
assign LUT_3[2174] = 32'b00000000000000001010111110111100;
assign LUT_3[2175] = 32'b00000000000000010001101010011001;
assign LUT_3[2176] = 32'b00000000000000000100000001001100;
assign LUT_3[2177] = 32'b00000000000000001010101100101001;
assign LUT_3[2178] = 32'b00000000000000000110001000110000;
assign LUT_3[2179] = 32'b00000000000000001100110100001101;
assign LUT_3[2180] = 32'b00000000000000000001001111000010;
assign LUT_3[2181] = 32'b00000000000000000111111010011111;
assign LUT_3[2182] = 32'b00000000000000000011010110100110;
assign LUT_3[2183] = 32'b00000000000000001010000010000011;
assign LUT_3[2184] = 32'b00000000000000001001011010010010;
assign LUT_3[2185] = 32'b00000000000000010000000101101111;
assign LUT_3[2186] = 32'b00000000000000001011100001110110;
assign LUT_3[2187] = 32'b00000000000000010010001101010011;
assign LUT_3[2188] = 32'b00000000000000000110101000001000;
assign LUT_3[2189] = 32'b00000000000000001101010011100101;
assign LUT_3[2190] = 32'b00000000000000001000101111101100;
assign LUT_3[2191] = 32'b00000000000000001111011011001001;
assign LUT_3[2192] = 32'b00000000000000000111010100001111;
assign LUT_3[2193] = 32'b00000000000000001101111111101100;
assign LUT_3[2194] = 32'b00000000000000001001011011110011;
assign LUT_3[2195] = 32'b00000000000000010000000111010000;
assign LUT_3[2196] = 32'b00000000000000000100100010000101;
assign LUT_3[2197] = 32'b00000000000000001011001101100010;
assign LUT_3[2198] = 32'b00000000000000000110101001101001;
assign LUT_3[2199] = 32'b00000000000000001101010101000110;
assign LUT_3[2200] = 32'b00000000000000001100101101010101;
assign LUT_3[2201] = 32'b00000000000000010011011000110010;
assign LUT_3[2202] = 32'b00000000000000001110110100111001;
assign LUT_3[2203] = 32'b00000000000000010101100000010110;
assign LUT_3[2204] = 32'b00000000000000001001111011001011;
assign LUT_3[2205] = 32'b00000000000000010000100110101000;
assign LUT_3[2206] = 32'b00000000000000001100000010101111;
assign LUT_3[2207] = 32'b00000000000000010010101110001100;
assign LUT_3[2208] = 32'b00000000000000000101001111101100;
assign LUT_3[2209] = 32'b00000000000000001011111011001001;
assign LUT_3[2210] = 32'b00000000000000000111010111010000;
assign LUT_3[2211] = 32'b00000000000000001110000010101101;
assign LUT_3[2212] = 32'b00000000000000000010011101100010;
assign LUT_3[2213] = 32'b00000000000000001001001000111111;
assign LUT_3[2214] = 32'b00000000000000000100100101000110;
assign LUT_3[2215] = 32'b00000000000000001011010000100011;
assign LUT_3[2216] = 32'b00000000000000001010101000110010;
assign LUT_3[2217] = 32'b00000000000000010001010100001111;
assign LUT_3[2218] = 32'b00000000000000001100110000010110;
assign LUT_3[2219] = 32'b00000000000000010011011011110011;
assign LUT_3[2220] = 32'b00000000000000000111110110101000;
assign LUT_3[2221] = 32'b00000000000000001110100010000101;
assign LUT_3[2222] = 32'b00000000000000001001111110001100;
assign LUT_3[2223] = 32'b00000000000000010000101001101001;
assign LUT_3[2224] = 32'b00000000000000001000100010101111;
assign LUT_3[2225] = 32'b00000000000000001111001110001100;
assign LUT_3[2226] = 32'b00000000000000001010101010010011;
assign LUT_3[2227] = 32'b00000000000000010001010101110000;
assign LUT_3[2228] = 32'b00000000000000000101110000100101;
assign LUT_3[2229] = 32'b00000000000000001100011100000010;
assign LUT_3[2230] = 32'b00000000000000000111111000001001;
assign LUT_3[2231] = 32'b00000000000000001110100011100110;
assign LUT_3[2232] = 32'b00000000000000001101111011110101;
assign LUT_3[2233] = 32'b00000000000000010100100111010010;
assign LUT_3[2234] = 32'b00000000000000010000000011011001;
assign LUT_3[2235] = 32'b00000000000000010110101110110110;
assign LUT_3[2236] = 32'b00000000000000001011001001101011;
assign LUT_3[2237] = 32'b00000000000000010001110101001000;
assign LUT_3[2238] = 32'b00000000000000001101010001001111;
assign LUT_3[2239] = 32'b00000000000000010011111100101100;
assign LUT_3[2240] = 32'b00000000000000000011111001110111;
assign LUT_3[2241] = 32'b00000000000000001010100101010100;
assign LUT_3[2242] = 32'b00000000000000000110000001011011;
assign LUT_3[2243] = 32'b00000000000000001100101100111000;
assign LUT_3[2244] = 32'b00000000000000000001000111101101;
assign LUT_3[2245] = 32'b00000000000000000111110011001010;
assign LUT_3[2246] = 32'b00000000000000000011001111010001;
assign LUT_3[2247] = 32'b00000000000000001001111010101110;
assign LUT_3[2248] = 32'b00000000000000001001010010111101;
assign LUT_3[2249] = 32'b00000000000000001111111110011010;
assign LUT_3[2250] = 32'b00000000000000001011011010100001;
assign LUT_3[2251] = 32'b00000000000000010010000101111110;
assign LUT_3[2252] = 32'b00000000000000000110100000110011;
assign LUT_3[2253] = 32'b00000000000000001101001100010000;
assign LUT_3[2254] = 32'b00000000000000001000101000010111;
assign LUT_3[2255] = 32'b00000000000000001111010011110100;
assign LUT_3[2256] = 32'b00000000000000000111001100111010;
assign LUT_3[2257] = 32'b00000000000000001101111000010111;
assign LUT_3[2258] = 32'b00000000000000001001010100011110;
assign LUT_3[2259] = 32'b00000000000000001111111111111011;
assign LUT_3[2260] = 32'b00000000000000000100011010110000;
assign LUT_3[2261] = 32'b00000000000000001011000110001101;
assign LUT_3[2262] = 32'b00000000000000000110100010010100;
assign LUT_3[2263] = 32'b00000000000000001101001101110001;
assign LUT_3[2264] = 32'b00000000000000001100100110000000;
assign LUT_3[2265] = 32'b00000000000000010011010001011101;
assign LUT_3[2266] = 32'b00000000000000001110101101100100;
assign LUT_3[2267] = 32'b00000000000000010101011001000001;
assign LUT_3[2268] = 32'b00000000000000001001110011110110;
assign LUT_3[2269] = 32'b00000000000000010000011111010011;
assign LUT_3[2270] = 32'b00000000000000001011111011011010;
assign LUT_3[2271] = 32'b00000000000000010010100110110111;
assign LUT_3[2272] = 32'b00000000000000000101001000010111;
assign LUT_3[2273] = 32'b00000000000000001011110011110100;
assign LUT_3[2274] = 32'b00000000000000000111001111111011;
assign LUT_3[2275] = 32'b00000000000000001101111011011000;
assign LUT_3[2276] = 32'b00000000000000000010010110001101;
assign LUT_3[2277] = 32'b00000000000000001001000001101010;
assign LUT_3[2278] = 32'b00000000000000000100011101110001;
assign LUT_3[2279] = 32'b00000000000000001011001001001110;
assign LUT_3[2280] = 32'b00000000000000001010100001011101;
assign LUT_3[2281] = 32'b00000000000000010001001100111010;
assign LUT_3[2282] = 32'b00000000000000001100101001000001;
assign LUT_3[2283] = 32'b00000000000000010011010100011110;
assign LUT_3[2284] = 32'b00000000000000000111101111010011;
assign LUT_3[2285] = 32'b00000000000000001110011010110000;
assign LUT_3[2286] = 32'b00000000000000001001110110110111;
assign LUT_3[2287] = 32'b00000000000000010000100010010100;
assign LUT_3[2288] = 32'b00000000000000001000011011011010;
assign LUT_3[2289] = 32'b00000000000000001111000110110111;
assign LUT_3[2290] = 32'b00000000000000001010100010111110;
assign LUT_3[2291] = 32'b00000000000000010001001110011011;
assign LUT_3[2292] = 32'b00000000000000000101101001010000;
assign LUT_3[2293] = 32'b00000000000000001100010100101101;
assign LUT_3[2294] = 32'b00000000000000000111110000110100;
assign LUT_3[2295] = 32'b00000000000000001110011100010001;
assign LUT_3[2296] = 32'b00000000000000001101110100100000;
assign LUT_3[2297] = 32'b00000000000000010100011111111101;
assign LUT_3[2298] = 32'b00000000000000001111111100000100;
assign LUT_3[2299] = 32'b00000000000000010110100111100001;
assign LUT_3[2300] = 32'b00000000000000001011000010010110;
assign LUT_3[2301] = 32'b00000000000000010001101101110011;
assign LUT_3[2302] = 32'b00000000000000001101001001111010;
assign LUT_3[2303] = 32'b00000000000000010011110101010111;
assign LUT_3[2304] = 32'b11111111111111111110000101101111;
assign LUT_3[2305] = 32'b00000000000000000100110001001100;
assign LUT_3[2306] = 32'b00000000000000000000001101010011;
assign LUT_3[2307] = 32'b00000000000000000110111000110000;
assign LUT_3[2308] = 32'b11111111111111111011010011100101;
assign LUT_3[2309] = 32'b00000000000000000001111111000010;
assign LUT_3[2310] = 32'b11111111111111111101011011001001;
assign LUT_3[2311] = 32'b00000000000000000100000110100110;
assign LUT_3[2312] = 32'b00000000000000000011011110110101;
assign LUT_3[2313] = 32'b00000000000000001010001010010010;
assign LUT_3[2314] = 32'b00000000000000000101100110011001;
assign LUT_3[2315] = 32'b00000000000000001100010001110110;
assign LUT_3[2316] = 32'b00000000000000000000101100101011;
assign LUT_3[2317] = 32'b00000000000000000111011000001000;
assign LUT_3[2318] = 32'b00000000000000000010110100001111;
assign LUT_3[2319] = 32'b00000000000000001001011111101100;
assign LUT_3[2320] = 32'b00000000000000000001011000110010;
assign LUT_3[2321] = 32'b00000000000000001000000100001111;
assign LUT_3[2322] = 32'b00000000000000000011100000010110;
assign LUT_3[2323] = 32'b00000000000000001010001011110011;
assign LUT_3[2324] = 32'b11111111111111111110100110101000;
assign LUT_3[2325] = 32'b00000000000000000101010010000101;
assign LUT_3[2326] = 32'b00000000000000000000101110001100;
assign LUT_3[2327] = 32'b00000000000000000111011001101001;
assign LUT_3[2328] = 32'b00000000000000000110110001111000;
assign LUT_3[2329] = 32'b00000000000000001101011101010101;
assign LUT_3[2330] = 32'b00000000000000001000111001011100;
assign LUT_3[2331] = 32'b00000000000000001111100100111001;
assign LUT_3[2332] = 32'b00000000000000000011111111101110;
assign LUT_3[2333] = 32'b00000000000000001010101011001011;
assign LUT_3[2334] = 32'b00000000000000000110000111010010;
assign LUT_3[2335] = 32'b00000000000000001100110010101111;
assign LUT_3[2336] = 32'b11111111111111111111010100001111;
assign LUT_3[2337] = 32'b00000000000000000101111111101100;
assign LUT_3[2338] = 32'b00000000000000000001011011110011;
assign LUT_3[2339] = 32'b00000000000000001000000111010000;
assign LUT_3[2340] = 32'b11111111111111111100100010000101;
assign LUT_3[2341] = 32'b00000000000000000011001101100010;
assign LUT_3[2342] = 32'b11111111111111111110101001101001;
assign LUT_3[2343] = 32'b00000000000000000101010101000110;
assign LUT_3[2344] = 32'b00000000000000000100101101010101;
assign LUT_3[2345] = 32'b00000000000000001011011000110010;
assign LUT_3[2346] = 32'b00000000000000000110110100111001;
assign LUT_3[2347] = 32'b00000000000000001101100000010110;
assign LUT_3[2348] = 32'b00000000000000000001111011001011;
assign LUT_3[2349] = 32'b00000000000000001000100110101000;
assign LUT_3[2350] = 32'b00000000000000000100000010101111;
assign LUT_3[2351] = 32'b00000000000000001010101110001100;
assign LUT_3[2352] = 32'b00000000000000000010100111010010;
assign LUT_3[2353] = 32'b00000000000000001001010010101111;
assign LUT_3[2354] = 32'b00000000000000000100101110110110;
assign LUT_3[2355] = 32'b00000000000000001011011010010011;
assign LUT_3[2356] = 32'b11111111111111111111110101001000;
assign LUT_3[2357] = 32'b00000000000000000110100000100101;
assign LUT_3[2358] = 32'b00000000000000000001111100101100;
assign LUT_3[2359] = 32'b00000000000000001000101000001001;
assign LUT_3[2360] = 32'b00000000000000001000000000011000;
assign LUT_3[2361] = 32'b00000000000000001110101011110101;
assign LUT_3[2362] = 32'b00000000000000001010000111111100;
assign LUT_3[2363] = 32'b00000000000000010000110011011001;
assign LUT_3[2364] = 32'b00000000000000000101001110001110;
assign LUT_3[2365] = 32'b00000000000000001011111001101011;
assign LUT_3[2366] = 32'b00000000000000000111010101110010;
assign LUT_3[2367] = 32'b00000000000000001110000001001111;
assign LUT_3[2368] = 32'b11111111111111111101111110011010;
assign LUT_3[2369] = 32'b00000000000000000100101001110111;
assign LUT_3[2370] = 32'b00000000000000000000000101111110;
assign LUT_3[2371] = 32'b00000000000000000110110001011011;
assign LUT_3[2372] = 32'b11111111111111111011001100010000;
assign LUT_3[2373] = 32'b00000000000000000001110111101101;
assign LUT_3[2374] = 32'b11111111111111111101010011110100;
assign LUT_3[2375] = 32'b00000000000000000011111111010001;
assign LUT_3[2376] = 32'b00000000000000000011010111100000;
assign LUT_3[2377] = 32'b00000000000000001010000010111101;
assign LUT_3[2378] = 32'b00000000000000000101011111000100;
assign LUT_3[2379] = 32'b00000000000000001100001010100001;
assign LUT_3[2380] = 32'b00000000000000000000100101010110;
assign LUT_3[2381] = 32'b00000000000000000111010000110011;
assign LUT_3[2382] = 32'b00000000000000000010101100111010;
assign LUT_3[2383] = 32'b00000000000000001001011000010111;
assign LUT_3[2384] = 32'b00000000000000000001010001011101;
assign LUT_3[2385] = 32'b00000000000000000111111100111010;
assign LUT_3[2386] = 32'b00000000000000000011011001000001;
assign LUT_3[2387] = 32'b00000000000000001010000100011110;
assign LUT_3[2388] = 32'b11111111111111111110011111010011;
assign LUT_3[2389] = 32'b00000000000000000101001010110000;
assign LUT_3[2390] = 32'b00000000000000000000100110110111;
assign LUT_3[2391] = 32'b00000000000000000111010010010100;
assign LUT_3[2392] = 32'b00000000000000000110101010100011;
assign LUT_3[2393] = 32'b00000000000000001101010110000000;
assign LUT_3[2394] = 32'b00000000000000001000110010000111;
assign LUT_3[2395] = 32'b00000000000000001111011101100100;
assign LUT_3[2396] = 32'b00000000000000000011111000011001;
assign LUT_3[2397] = 32'b00000000000000001010100011110110;
assign LUT_3[2398] = 32'b00000000000000000101111111111101;
assign LUT_3[2399] = 32'b00000000000000001100101011011010;
assign LUT_3[2400] = 32'b11111111111111111111001100111010;
assign LUT_3[2401] = 32'b00000000000000000101111000010111;
assign LUT_3[2402] = 32'b00000000000000000001010100011110;
assign LUT_3[2403] = 32'b00000000000000000111111111111011;
assign LUT_3[2404] = 32'b11111111111111111100011010110000;
assign LUT_3[2405] = 32'b00000000000000000011000110001101;
assign LUT_3[2406] = 32'b11111111111111111110100010010100;
assign LUT_3[2407] = 32'b00000000000000000101001101110001;
assign LUT_3[2408] = 32'b00000000000000000100100110000000;
assign LUT_3[2409] = 32'b00000000000000001011010001011101;
assign LUT_3[2410] = 32'b00000000000000000110101101100100;
assign LUT_3[2411] = 32'b00000000000000001101011001000001;
assign LUT_3[2412] = 32'b00000000000000000001110011110110;
assign LUT_3[2413] = 32'b00000000000000001000011111010011;
assign LUT_3[2414] = 32'b00000000000000000011111011011010;
assign LUT_3[2415] = 32'b00000000000000001010100110110111;
assign LUT_3[2416] = 32'b00000000000000000010011111111101;
assign LUT_3[2417] = 32'b00000000000000001001001011011010;
assign LUT_3[2418] = 32'b00000000000000000100100111100001;
assign LUT_3[2419] = 32'b00000000000000001011010010111110;
assign LUT_3[2420] = 32'b11111111111111111111101101110011;
assign LUT_3[2421] = 32'b00000000000000000110011001010000;
assign LUT_3[2422] = 32'b00000000000000000001110101010111;
assign LUT_3[2423] = 32'b00000000000000001000100000110100;
assign LUT_3[2424] = 32'b00000000000000000111111001000011;
assign LUT_3[2425] = 32'b00000000000000001110100100100000;
assign LUT_3[2426] = 32'b00000000000000001010000000100111;
assign LUT_3[2427] = 32'b00000000000000010000101100000100;
assign LUT_3[2428] = 32'b00000000000000000101000110111001;
assign LUT_3[2429] = 32'b00000000000000001011110010010110;
assign LUT_3[2430] = 32'b00000000000000000111001110011101;
assign LUT_3[2431] = 32'b00000000000000001101111001111010;
assign LUT_3[2432] = 32'b00000000000000000000010000101101;
assign LUT_3[2433] = 32'b00000000000000000110111100001010;
assign LUT_3[2434] = 32'b00000000000000000010011000010001;
assign LUT_3[2435] = 32'b00000000000000001001000011101110;
assign LUT_3[2436] = 32'b11111111111111111101011110100011;
assign LUT_3[2437] = 32'b00000000000000000100001010000000;
assign LUT_3[2438] = 32'b11111111111111111111100110000111;
assign LUT_3[2439] = 32'b00000000000000000110010001100100;
assign LUT_3[2440] = 32'b00000000000000000101101001110011;
assign LUT_3[2441] = 32'b00000000000000001100010101010000;
assign LUT_3[2442] = 32'b00000000000000000111110001010111;
assign LUT_3[2443] = 32'b00000000000000001110011100110100;
assign LUT_3[2444] = 32'b00000000000000000010110111101001;
assign LUT_3[2445] = 32'b00000000000000001001100011000110;
assign LUT_3[2446] = 32'b00000000000000000100111111001101;
assign LUT_3[2447] = 32'b00000000000000001011101010101010;
assign LUT_3[2448] = 32'b00000000000000000011100011110000;
assign LUT_3[2449] = 32'b00000000000000001010001111001101;
assign LUT_3[2450] = 32'b00000000000000000101101011010100;
assign LUT_3[2451] = 32'b00000000000000001100010110110001;
assign LUT_3[2452] = 32'b00000000000000000000110001100110;
assign LUT_3[2453] = 32'b00000000000000000111011101000011;
assign LUT_3[2454] = 32'b00000000000000000010111001001010;
assign LUT_3[2455] = 32'b00000000000000001001100100100111;
assign LUT_3[2456] = 32'b00000000000000001000111100110110;
assign LUT_3[2457] = 32'b00000000000000001111101000010011;
assign LUT_3[2458] = 32'b00000000000000001011000100011010;
assign LUT_3[2459] = 32'b00000000000000010001101111110111;
assign LUT_3[2460] = 32'b00000000000000000110001010101100;
assign LUT_3[2461] = 32'b00000000000000001100110110001001;
assign LUT_3[2462] = 32'b00000000000000001000010010010000;
assign LUT_3[2463] = 32'b00000000000000001110111101101101;
assign LUT_3[2464] = 32'b00000000000000000001011111001101;
assign LUT_3[2465] = 32'b00000000000000001000001010101010;
assign LUT_3[2466] = 32'b00000000000000000011100110110001;
assign LUT_3[2467] = 32'b00000000000000001010010010001110;
assign LUT_3[2468] = 32'b11111111111111111110101101000011;
assign LUT_3[2469] = 32'b00000000000000000101011000100000;
assign LUT_3[2470] = 32'b00000000000000000000110100100111;
assign LUT_3[2471] = 32'b00000000000000000111100000000100;
assign LUT_3[2472] = 32'b00000000000000000110111000010011;
assign LUT_3[2473] = 32'b00000000000000001101100011110000;
assign LUT_3[2474] = 32'b00000000000000001000111111110111;
assign LUT_3[2475] = 32'b00000000000000001111101011010100;
assign LUT_3[2476] = 32'b00000000000000000100000110001001;
assign LUT_3[2477] = 32'b00000000000000001010110001100110;
assign LUT_3[2478] = 32'b00000000000000000110001101101101;
assign LUT_3[2479] = 32'b00000000000000001100111001001010;
assign LUT_3[2480] = 32'b00000000000000000100110010010000;
assign LUT_3[2481] = 32'b00000000000000001011011101101101;
assign LUT_3[2482] = 32'b00000000000000000110111001110100;
assign LUT_3[2483] = 32'b00000000000000001101100101010001;
assign LUT_3[2484] = 32'b00000000000000000010000000000110;
assign LUT_3[2485] = 32'b00000000000000001000101011100011;
assign LUT_3[2486] = 32'b00000000000000000100000111101010;
assign LUT_3[2487] = 32'b00000000000000001010110011000111;
assign LUT_3[2488] = 32'b00000000000000001010001011010110;
assign LUT_3[2489] = 32'b00000000000000010000110110110011;
assign LUT_3[2490] = 32'b00000000000000001100010010111010;
assign LUT_3[2491] = 32'b00000000000000010010111110010111;
assign LUT_3[2492] = 32'b00000000000000000111011001001100;
assign LUT_3[2493] = 32'b00000000000000001110000100101001;
assign LUT_3[2494] = 32'b00000000000000001001100000110000;
assign LUT_3[2495] = 32'b00000000000000010000001100001101;
assign LUT_3[2496] = 32'b00000000000000000000001001011000;
assign LUT_3[2497] = 32'b00000000000000000110110100110101;
assign LUT_3[2498] = 32'b00000000000000000010010000111100;
assign LUT_3[2499] = 32'b00000000000000001000111100011001;
assign LUT_3[2500] = 32'b11111111111111111101010111001110;
assign LUT_3[2501] = 32'b00000000000000000100000010101011;
assign LUT_3[2502] = 32'b11111111111111111111011110110010;
assign LUT_3[2503] = 32'b00000000000000000110001010001111;
assign LUT_3[2504] = 32'b00000000000000000101100010011110;
assign LUT_3[2505] = 32'b00000000000000001100001101111011;
assign LUT_3[2506] = 32'b00000000000000000111101010000010;
assign LUT_3[2507] = 32'b00000000000000001110010101011111;
assign LUT_3[2508] = 32'b00000000000000000010110000010100;
assign LUT_3[2509] = 32'b00000000000000001001011011110001;
assign LUT_3[2510] = 32'b00000000000000000100110111111000;
assign LUT_3[2511] = 32'b00000000000000001011100011010101;
assign LUT_3[2512] = 32'b00000000000000000011011100011011;
assign LUT_3[2513] = 32'b00000000000000001010000111111000;
assign LUT_3[2514] = 32'b00000000000000000101100011111111;
assign LUT_3[2515] = 32'b00000000000000001100001111011100;
assign LUT_3[2516] = 32'b00000000000000000000101010010001;
assign LUT_3[2517] = 32'b00000000000000000111010101101110;
assign LUT_3[2518] = 32'b00000000000000000010110001110101;
assign LUT_3[2519] = 32'b00000000000000001001011101010010;
assign LUT_3[2520] = 32'b00000000000000001000110101100001;
assign LUT_3[2521] = 32'b00000000000000001111100000111110;
assign LUT_3[2522] = 32'b00000000000000001010111101000101;
assign LUT_3[2523] = 32'b00000000000000010001101000100010;
assign LUT_3[2524] = 32'b00000000000000000110000011010111;
assign LUT_3[2525] = 32'b00000000000000001100101110110100;
assign LUT_3[2526] = 32'b00000000000000001000001010111011;
assign LUT_3[2527] = 32'b00000000000000001110110110011000;
assign LUT_3[2528] = 32'b00000000000000000001010111111000;
assign LUT_3[2529] = 32'b00000000000000001000000011010101;
assign LUT_3[2530] = 32'b00000000000000000011011111011100;
assign LUT_3[2531] = 32'b00000000000000001010001010111001;
assign LUT_3[2532] = 32'b11111111111111111110100101101110;
assign LUT_3[2533] = 32'b00000000000000000101010001001011;
assign LUT_3[2534] = 32'b00000000000000000000101101010010;
assign LUT_3[2535] = 32'b00000000000000000111011000101111;
assign LUT_3[2536] = 32'b00000000000000000110110000111110;
assign LUT_3[2537] = 32'b00000000000000001101011100011011;
assign LUT_3[2538] = 32'b00000000000000001000111000100010;
assign LUT_3[2539] = 32'b00000000000000001111100011111111;
assign LUT_3[2540] = 32'b00000000000000000011111110110100;
assign LUT_3[2541] = 32'b00000000000000001010101010010001;
assign LUT_3[2542] = 32'b00000000000000000110000110011000;
assign LUT_3[2543] = 32'b00000000000000001100110001110101;
assign LUT_3[2544] = 32'b00000000000000000100101010111011;
assign LUT_3[2545] = 32'b00000000000000001011010110011000;
assign LUT_3[2546] = 32'b00000000000000000110110010011111;
assign LUT_3[2547] = 32'b00000000000000001101011101111100;
assign LUT_3[2548] = 32'b00000000000000000001111000110001;
assign LUT_3[2549] = 32'b00000000000000001000100100001110;
assign LUT_3[2550] = 32'b00000000000000000100000000010101;
assign LUT_3[2551] = 32'b00000000000000001010101011110010;
assign LUT_3[2552] = 32'b00000000000000001010000100000001;
assign LUT_3[2553] = 32'b00000000000000010000101111011110;
assign LUT_3[2554] = 32'b00000000000000001100001011100101;
assign LUT_3[2555] = 32'b00000000000000010010110111000010;
assign LUT_3[2556] = 32'b00000000000000000111010001110111;
assign LUT_3[2557] = 32'b00000000000000001101111101010100;
assign LUT_3[2558] = 32'b00000000000000001001011001011011;
assign LUT_3[2559] = 32'b00000000000000010000000100111000;
assign LUT_3[2560] = 32'b00000000000000000101001011011010;
assign LUT_3[2561] = 32'b00000000000000001011110110110111;
assign LUT_3[2562] = 32'b00000000000000000111010010111110;
assign LUT_3[2563] = 32'b00000000000000001101111110011011;
assign LUT_3[2564] = 32'b00000000000000000010011001010000;
assign LUT_3[2565] = 32'b00000000000000001001000100101101;
assign LUT_3[2566] = 32'b00000000000000000100100000110100;
assign LUT_3[2567] = 32'b00000000000000001011001100010001;
assign LUT_3[2568] = 32'b00000000000000001010100100100000;
assign LUT_3[2569] = 32'b00000000000000010001001111111101;
assign LUT_3[2570] = 32'b00000000000000001100101100000100;
assign LUT_3[2571] = 32'b00000000000000010011010111100001;
assign LUT_3[2572] = 32'b00000000000000000111110010010110;
assign LUT_3[2573] = 32'b00000000000000001110011101110011;
assign LUT_3[2574] = 32'b00000000000000001001111001111010;
assign LUT_3[2575] = 32'b00000000000000010000100101010111;
assign LUT_3[2576] = 32'b00000000000000001000011110011101;
assign LUT_3[2577] = 32'b00000000000000001111001001111010;
assign LUT_3[2578] = 32'b00000000000000001010100110000001;
assign LUT_3[2579] = 32'b00000000000000010001010001011110;
assign LUT_3[2580] = 32'b00000000000000000101101100010011;
assign LUT_3[2581] = 32'b00000000000000001100010111110000;
assign LUT_3[2582] = 32'b00000000000000000111110011110111;
assign LUT_3[2583] = 32'b00000000000000001110011111010100;
assign LUT_3[2584] = 32'b00000000000000001101110111100011;
assign LUT_3[2585] = 32'b00000000000000010100100011000000;
assign LUT_3[2586] = 32'b00000000000000001111111111000111;
assign LUT_3[2587] = 32'b00000000000000010110101010100100;
assign LUT_3[2588] = 32'b00000000000000001011000101011001;
assign LUT_3[2589] = 32'b00000000000000010001110000110110;
assign LUT_3[2590] = 32'b00000000000000001101001100111101;
assign LUT_3[2591] = 32'b00000000000000010011111000011010;
assign LUT_3[2592] = 32'b00000000000000000110011001111010;
assign LUT_3[2593] = 32'b00000000000000001101000101010111;
assign LUT_3[2594] = 32'b00000000000000001000100001011110;
assign LUT_3[2595] = 32'b00000000000000001111001100111011;
assign LUT_3[2596] = 32'b00000000000000000011100111110000;
assign LUT_3[2597] = 32'b00000000000000001010010011001101;
assign LUT_3[2598] = 32'b00000000000000000101101111010100;
assign LUT_3[2599] = 32'b00000000000000001100011010110001;
assign LUT_3[2600] = 32'b00000000000000001011110011000000;
assign LUT_3[2601] = 32'b00000000000000010010011110011101;
assign LUT_3[2602] = 32'b00000000000000001101111010100100;
assign LUT_3[2603] = 32'b00000000000000010100100110000001;
assign LUT_3[2604] = 32'b00000000000000001001000000110110;
assign LUT_3[2605] = 32'b00000000000000001111101100010011;
assign LUT_3[2606] = 32'b00000000000000001011001000011010;
assign LUT_3[2607] = 32'b00000000000000010001110011110111;
assign LUT_3[2608] = 32'b00000000000000001001101100111101;
assign LUT_3[2609] = 32'b00000000000000010000011000011010;
assign LUT_3[2610] = 32'b00000000000000001011110100100001;
assign LUT_3[2611] = 32'b00000000000000010010011111111110;
assign LUT_3[2612] = 32'b00000000000000000110111010110011;
assign LUT_3[2613] = 32'b00000000000000001101100110010000;
assign LUT_3[2614] = 32'b00000000000000001001000010010111;
assign LUT_3[2615] = 32'b00000000000000001111101101110100;
assign LUT_3[2616] = 32'b00000000000000001111000110000011;
assign LUT_3[2617] = 32'b00000000000000010101110001100000;
assign LUT_3[2618] = 32'b00000000000000010001001101100111;
assign LUT_3[2619] = 32'b00000000000000010111111001000100;
assign LUT_3[2620] = 32'b00000000000000001100010011111001;
assign LUT_3[2621] = 32'b00000000000000010010111111010110;
assign LUT_3[2622] = 32'b00000000000000001110011011011101;
assign LUT_3[2623] = 32'b00000000000000010101000110111010;
assign LUT_3[2624] = 32'b00000000000000000101000100000101;
assign LUT_3[2625] = 32'b00000000000000001011101111100010;
assign LUT_3[2626] = 32'b00000000000000000111001011101001;
assign LUT_3[2627] = 32'b00000000000000001101110111000110;
assign LUT_3[2628] = 32'b00000000000000000010010001111011;
assign LUT_3[2629] = 32'b00000000000000001000111101011000;
assign LUT_3[2630] = 32'b00000000000000000100011001011111;
assign LUT_3[2631] = 32'b00000000000000001011000100111100;
assign LUT_3[2632] = 32'b00000000000000001010011101001011;
assign LUT_3[2633] = 32'b00000000000000010001001000101000;
assign LUT_3[2634] = 32'b00000000000000001100100100101111;
assign LUT_3[2635] = 32'b00000000000000010011010000001100;
assign LUT_3[2636] = 32'b00000000000000000111101011000001;
assign LUT_3[2637] = 32'b00000000000000001110010110011110;
assign LUT_3[2638] = 32'b00000000000000001001110010100101;
assign LUT_3[2639] = 32'b00000000000000010000011110000010;
assign LUT_3[2640] = 32'b00000000000000001000010111001000;
assign LUT_3[2641] = 32'b00000000000000001111000010100101;
assign LUT_3[2642] = 32'b00000000000000001010011110101100;
assign LUT_3[2643] = 32'b00000000000000010001001010001001;
assign LUT_3[2644] = 32'b00000000000000000101100100111110;
assign LUT_3[2645] = 32'b00000000000000001100010000011011;
assign LUT_3[2646] = 32'b00000000000000000111101100100010;
assign LUT_3[2647] = 32'b00000000000000001110010111111111;
assign LUT_3[2648] = 32'b00000000000000001101110000001110;
assign LUT_3[2649] = 32'b00000000000000010100011011101011;
assign LUT_3[2650] = 32'b00000000000000001111110111110010;
assign LUT_3[2651] = 32'b00000000000000010110100011001111;
assign LUT_3[2652] = 32'b00000000000000001010111110000100;
assign LUT_3[2653] = 32'b00000000000000010001101001100001;
assign LUT_3[2654] = 32'b00000000000000001101000101101000;
assign LUT_3[2655] = 32'b00000000000000010011110001000101;
assign LUT_3[2656] = 32'b00000000000000000110010010100101;
assign LUT_3[2657] = 32'b00000000000000001100111110000010;
assign LUT_3[2658] = 32'b00000000000000001000011010001001;
assign LUT_3[2659] = 32'b00000000000000001111000101100110;
assign LUT_3[2660] = 32'b00000000000000000011100000011011;
assign LUT_3[2661] = 32'b00000000000000001010001011111000;
assign LUT_3[2662] = 32'b00000000000000000101100111111111;
assign LUT_3[2663] = 32'b00000000000000001100010011011100;
assign LUT_3[2664] = 32'b00000000000000001011101011101011;
assign LUT_3[2665] = 32'b00000000000000010010010111001000;
assign LUT_3[2666] = 32'b00000000000000001101110011001111;
assign LUT_3[2667] = 32'b00000000000000010100011110101100;
assign LUT_3[2668] = 32'b00000000000000001000111001100001;
assign LUT_3[2669] = 32'b00000000000000001111100100111110;
assign LUT_3[2670] = 32'b00000000000000001011000001000101;
assign LUT_3[2671] = 32'b00000000000000010001101100100010;
assign LUT_3[2672] = 32'b00000000000000001001100101101000;
assign LUT_3[2673] = 32'b00000000000000010000010001000101;
assign LUT_3[2674] = 32'b00000000000000001011101101001100;
assign LUT_3[2675] = 32'b00000000000000010010011000101001;
assign LUT_3[2676] = 32'b00000000000000000110110011011110;
assign LUT_3[2677] = 32'b00000000000000001101011110111011;
assign LUT_3[2678] = 32'b00000000000000001000111011000010;
assign LUT_3[2679] = 32'b00000000000000001111100110011111;
assign LUT_3[2680] = 32'b00000000000000001110111110101110;
assign LUT_3[2681] = 32'b00000000000000010101101010001011;
assign LUT_3[2682] = 32'b00000000000000010001000110010010;
assign LUT_3[2683] = 32'b00000000000000010111110001101111;
assign LUT_3[2684] = 32'b00000000000000001100001100100100;
assign LUT_3[2685] = 32'b00000000000000010010111000000001;
assign LUT_3[2686] = 32'b00000000000000001110010100001000;
assign LUT_3[2687] = 32'b00000000000000010100111111100101;
assign LUT_3[2688] = 32'b00000000000000000111010110011000;
assign LUT_3[2689] = 32'b00000000000000001110000001110101;
assign LUT_3[2690] = 32'b00000000000000001001011101111100;
assign LUT_3[2691] = 32'b00000000000000010000001001011001;
assign LUT_3[2692] = 32'b00000000000000000100100100001110;
assign LUT_3[2693] = 32'b00000000000000001011001111101011;
assign LUT_3[2694] = 32'b00000000000000000110101011110010;
assign LUT_3[2695] = 32'b00000000000000001101010111001111;
assign LUT_3[2696] = 32'b00000000000000001100101111011110;
assign LUT_3[2697] = 32'b00000000000000010011011010111011;
assign LUT_3[2698] = 32'b00000000000000001110110111000010;
assign LUT_3[2699] = 32'b00000000000000010101100010011111;
assign LUT_3[2700] = 32'b00000000000000001001111101010100;
assign LUT_3[2701] = 32'b00000000000000010000101000110001;
assign LUT_3[2702] = 32'b00000000000000001100000100111000;
assign LUT_3[2703] = 32'b00000000000000010010110000010101;
assign LUT_3[2704] = 32'b00000000000000001010101001011011;
assign LUT_3[2705] = 32'b00000000000000010001010100111000;
assign LUT_3[2706] = 32'b00000000000000001100110000111111;
assign LUT_3[2707] = 32'b00000000000000010011011100011100;
assign LUT_3[2708] = 32'b00000000000000000111110111010001;
assign LUT_3[2709] = 32'b00000000000000001110100010101110;
assign LUT_3[2710] = 32'b00000000000000001001111110110101;
assign LUT_3[2711] = 32'b00000000000000010000101010010010;
assign LUT_3[2712] = 32'b00000000000000010000000010100001;
assign LUT_3[2713] = 32'b00000000000000010110101101111110;
assign LUT_3[2714] = 32'b00000000000000010010001010000101;
assign LUT_3[2715] = 32'b00000000000000011000110101100010;
assign LUT_3[2716] = 32'b00000000000000001101010000010111;
assign LUT_3[2717] = 32'b00000000000000010011111011110100;
assign LUT_3[2718] = 32'b00000000000000001111010111111011;
assign LUT_3[2719] = 32'b00000000000000010110000011011000;
assign LUT_3[2720] = 32'b00000000000000001000100100111000;
assign LUT_3[2721] = 32'b00000000000000001111010000010101;
assign LUT_3[2722] = 32'b00000000000000001010101100011100;
assign LUT_3[2723] = 32'b00000000000000010001010111111001;
assign LUT_3[2724] = 32'b00000000000000000101110010101110;
assign LUT_3[2725] = 32'b00000000000000001100011110001011;
assign LUT_3[2726] = 32'b00000000000000000111111010010010;
assign LUT_3[2727] = 32'b00000000000000001110100101101111;
assign LUT_3[2728] = 32'b00000000000000001101111101111110;
assign LUT_3[2729] = 32'b00000000000000010100101001011011;
assign LUT_3[2730] = 32'b00000000000000010000000101100010;
assign LUT_3[2731] = 32'b00000000000000010110110000111111;
assign LUT_3[2732] = 32'b00000000000000001011001011110100;
assign LUT_3[2733] = 32'b00000000000000010001110111010001;
assign LUT_3[2734] = 32'b00000000000000001101010011011000;
assign LUT_3[2735] = 32'b00000000000000010011111110110101;
assign LUT_3[2736] = 32'b00000000000000001011110111111011;
assign LUT_3[2737] = 32'b00000000000000010010100011011000;
assign LUT_3[2738] = 32'b00000000000000001101111111011111;
assign LUT_3[2739] = 32'b00000000000000010100101010111100;
assign LUT_3[2740] = 32'b00000000000000001001000101110001;
assign LUT_3[2741] = 32'b00000000000000001111110001001110;
assign LUT_3[2742] = 32'b00000000000000001011001101010101;
assign LUT_3[2743] = 32'b00000000000000010001111000110010;
assign LUT_3[2744] = 32'b00000000000000010001010001000001;
assign LUT_3[2745] = 32'b00000000000000010111111100011110;
assign LUT_3[2746] = 32'b00000000000000010011011000100101;
assign LUT_3[2747] = 32'b00000000000000011010000100000010;
assign LUT_3[2748] = 32'b00000000000000001110011110110111;
assign LUT_3[2749] = 32'b00000000000000010101001010010100;
assign LUT_3[2750] = 32'b00000000000000010000100110011011;
assign LUT_3[2751] = 32'b00000000000000010111010001111000;
assign LUT_3[2752] = 32'b00000000000000000111001111000011;
assign LUT_3[2753] = 32'b00000000000000001101111010100000;
assign LUT_3[2754] = 32'b00000000000000001001010110100111;
assign LUT_3[2755] = 32'b00000000000000010000000010000100;
assign LUT_3[2756] = 32'b00000000000000000100011100111001;
assign LUT_3[2757] = 32'b00000000000000001011001000010110;
assign LUT_3[2758] = 32'b00000000000000000110100100011101;
assign LUT_3[2759] = 32'b00000000000000001101001111111010;
assign LUT_3[2760] = 32'b00000000000000001100101000001001;
assign LUT_3[2761] = 32'b00000000000000010011010011100110;
assign LUT_3[2762] = 32'b00000000000000001110101111101101;
assign LUT_3[2763] = 32'b00000000000000010101011011001010;
assign LUT_3[2764] = 32'b00000000000000001001110101111111;
assign LUT_3[2765] = 32'b00000000000000010000100001011100;
assign LUT_3[2766] = 32'b00000000000000001011111101100011;
assign LUT_3[2767] = 32'b00000000000000010010101001000000;
assign LUT_3[2768] = 32'b00000000000000001010100010000110;
assign LUT_3[2769] = 32'b00000000000000010001001101100011;
assign LUT_3[2770] = 32'b00000000000000001100101001101010;
assign LUT_3[2771] = 32'b00000000000000010011010101000111;
assign LUT_3[2772] = 32'b00000000000000000111101111111100;
assign LUT_3[2773] = 32'b00000000000000001110011011011001;
assign LUT_3[2774] = 32'b00000000000000001001110111100000;
assign LUT_3[2775] = 32'b00000000000000010000100010111101;
assign LUT_3[2776] = 32'b00000000000000001111111011001100;
assign LUT_3[2777] = 32'b00000000000000010110100110101001;
assign LUT_3[2778] = 32'b00000000000000010010000010110000;
assign LUT_3[2779] = 32'b00000000000000011000101110001101;
assign LUT_3[2780] = 32'b00000000000000001101001001000010;
assign LUT_3[2781] = 32'b00000000000000010011110100011111;
assign LUT_3[2782] = 32'b00000000000000001111010000100110;
assign LUT_3[2783] = 32'b00000000000000010101111100000011;
assign LUT_3[2784] = 32'b00000000000000001000011101100011;
assign LUT_3[2785] = 32'b00000000000000001111001001000000;
assign LUT_3[2786] = 32'b00000000000000001010100101000111;
assign LUT_3[2787] = 32'b00000000000000010001010000100100;
assign LUT_3[2788] = 32'b00000000000000000101101011011001;
assign LUT_3[2789] = 32'b00000000000000001100010110110110;
assign LUT_3[2790] = 32'b00000000000000000111110010111101;
assign LUT_3[2791] = 32'b00000000000000001110011110011010;
assign LUT_3[2792] = 32'b00000000000000001101110110101001;
assign LUT_3[2793] = 32'b00000000000000010100100010000110;
assign LUT_3[2794] = 32'b00000000000000001111111110001101;
assign LUT_3[2795] = 32'b00000000000000010110101001101010;
assign LUT_3[2796] = 32'b00000000000000001011000100011111;
assign LUT_3[2797] = 32'b00000000000000010001101111111100;
assign LUT_3[2798] = 32'b00000000000000001101001100000011;
assign LUT_3[2799] = 32'b00000000000000010011110111100000;
assign LUT_3[2800] = 32'b00000000000000001011110000100110;
assign LUT_3[2801] = 32'b00000000000000010010011100000011;
assign LUT_3[2802] = 32'b00000000000000001101111000001010;
assign LUT_3[2803] = 32'b00000000000000010100100011100111;
assign LUT_3[2804] = 32'b00000000000000001000111110011100;
assign LUT_3[2805] = 32'b00000000000000001111101001111001;
assign LUT_3[2806] = 32'b00000000000000001011000110000000;
assign LUT_3[2807] = 32'b00000000000000010001110001011101;
assign LUT_3[2808] = 32'b00000000000000010001001001101100;
assign LUT_3[2809] = 32'b00000000000000010111110101001001;
assign LUT_3[2810] = 32'b00000000000000010011010001010000;
assign LUT_3[2811] = 32'b00000000000000011001111100101101;
assign LUT_3[2812] = 32'b00000000000000001110010111100010;
assign LUT_3[2813] = 32'b00000000000000010101000010111111;
assign LUT_3[2814] = 32'b00000000000000010000011111000110;
assign LUT_3[2815] = 32'b00000000000000010111001010100011;
assign LUT_3[2816] = 32'b00000000000000000001011010111011;
assign LUT_3[2817] = 32'b00000000000000001000000110011000;
assign LUT_3[2818] = 32'b00000000000000000011100010011111;
assign LUT_3[2819] = 32'b00000000000000001010001101111100;
assign LUT_3[2820] = 32'b11111111111111111110101000110001;
assign LUT_3[2821] = 32'b00000000000000000101010100001110;
assign LUT_3[2822] = 32'b00000000000000000000110000010101;
assign LUT_3[2823] = 32'b00000000000000000111011011110010;
assign LUT_3[2824] = 32'b00000000000000000110110100000001;
assign LUT_3[2825] = 32'b00000000000000001101011111011110;
assign LUT_3[2826] = 32'b00000000000000001000111011100101;
assign LUT_3[2827] = 32'b00000000000000001111100111000010;
assign LUT_3[2828] = 32'b00000000000000000100000001110111;
assign LUT_3[2829] = 32'b00000000000000001010101101010100;
assign LUT_3[2830] = 32'b00000000000000000110001001011011;
assign LUT_3[2831] = 32'b00000000000000001100110100111000;
assign LUT_3[2832] = 32'b00000000000000000100101101111110;
assign LUT_3[2833] = 32'b00000000000000001011011001011011;
assign LUT_3[2834] = 32'b00000000000000000110110101100010;
assign LUT_3[2835] = 32'b00000000000000001101100000111111;
assign LUT_3[2836] = 32'b00000000000000000001111011110100;
assign LUT_3[2837] = 32'b00000000000000001000100111010001;
assign LUT_3[2838] = 32'b00000000000000000100000011011000;
assign LUT_3[2839] = 32'b00000000000000001010101110110101;
assign LUT_3[2840] = 32'b00000000000000001010000111000100;
assign LUT_3[2841] = 32'b00000000000000010000110010100001;
assign LUT_3[2842] = 32'b00000000000000001100001110101000;
assign LUT_3[2843] = 32'b00000000000000010010111010000101;
assign LUT_3[2844] = 32'b00000000000000000111010100111010;
assign LUT_3[2845] = 32'b00000000000000001110000000010111;
assign LUT_3[2846] = 32'b00000000000000001001011100011110;
assign LUT_3[2847] = 32'b00000000000000010000000111111011;
assign LUT_3[2848] = 32'b00000000000000000010101001011011;
assign LUT_3[2849] = 32'b00000000000000001001010100111000;
assign LUT_3[2850] = 32'b00000000000000000100110000111111;
assign LUT_3[2851] = 32'b00000000000000001011011100011100;
assign LUT_3[2852] = 32'b11111111111111111111110111010001;
assign LUT_3[2853] = 32'b00000000000000000110100010101110;
assign LUT_3[2854] = 32'b00000000000000000001111110110101;
assign LUT_3[2855] = 32'b00000000000000001000101010010010;
assign LUT_3[2856] = 32'b00000000000000001000000010100001;
assign LUT_3[2857] = 32'b00000000000000001110101101111110;
assign LUT_3[2858] = 32'b00000000000000001010001010000101;
assign LUT_3[2859] = 32'b00000000000000010000110101100010;
assign LUT_3[2860] = 32'b00000000000000000101010000010111;
assign LUT_3[2861] = 32'b00000000000000001011111011110100;
assign LUT_3[2862] = 32'b00000000000000000111010111111011;
assign LUT_3[2863] = 32'b00000000000000001110000011011000;
assign LUT_3[2864] = 32'b00000000000000000101111100011110;
assign LUT_3[2865] = 32'b00000000000000001100100111111011;
assign LUT_3[2866] = 32'b00000000000000001000000100000010;
assign LUT_3[2867] = 32'b00000000000000001110101111011111;
assign LUT_3[2868] = 32'b00000000000000000011001010010100;
assign LUT_3[2869] = 32'b00000000000000001001110101110001;
assign LUT_3[2870] = 32'b00000000000000000101010001111000;
assign LUT_3[2871] = 32'b00000000000000001011111101010101;
assign LUT_3[2872] = 32'b00000000000000001011010101100100;
assign LUT_3[2873] = 32'b00000000000000010010000001000001;
assign LUT_3[2874] = 32'b00000000000000001101011101001000;
assign LUT_3[2875] = 32'b00000000000000010100001000100101;
assign LUT_3[2876] = 32'b00000000000000001000100011011010;
assign LUT_3[2877] = 32'b00000000000000001111001110110111;
assign LUT_3[2878] = 32'b00000000000000001010101010111110;
assign LUT_3[2879] = 32'b00000000000000010001010110011011;
assign LUT_3[2880] = 32'b00000000000000000001010011100110;
assign LUT_3[2881] = 32'b00000000000000000111111111000011;
assign LUT_3[2882] = 32'b00000000000000000011011011001010;
assign LUT_3[2883] = 32'b00000000000000001010000110100111;
assign LUT_3[2884] = 32'b11111111111111111110100001011100;
assign LUT_3[2885] = 32'b00000000000000000101001100111001;
assign LUT_3[2886] = 32'b00000000000000000000101001000000;
assign LUT_3[2887] = 32'b00000000000000000111010100011101;
assign LUT_3[2888] = 32'b00000000000000000110101100101100;
assign LUT_3[2889] = 32'b00000000000000001101011000001001;
assign LUT_3[2890] = 32'b00000000000000001000110100010000;
assign LUT_3[2891] = 32'b00000000000000001111011111101101;
assign LUT_3[2892] = 32'b00000000000000000011111010100010;
assign LUT_3[2893] = 32'b00000000000000001010100101111111;
assign LUT_3[2894] = 32'b00000000000000000110000010000110;
assign LUT_3[2895] = 32'b00000000000000001100101101100011;
assign LUT_3[2896] = 32'b00000000000000000100100110101001;
assign LUT_3[2897] = 32'b00000000000000001011010010000110;
assign LUT_3[2898] = 32'b00000000000000000110101110001101;
assign LUT_3[2899] = 32'b00000000000000001101011001101010;
assign LUT_3[2900] = 32'b00000000000000000001110100011111;
assign LUT_3[2901] = 32'b00000000000000001000011111111100;
assign LUT_3[2902] = 32'b00000000000000000011111100000011;
assign LUT_3[2903] = 32'b00000000000000001010100111100000;
assign LUT_3[2904] = 32'b00000000000000001001111111101111;
assign LUT_3[2905] = 32'b00000000000000010000101011001100;
assign LUT_3[2906] = 32'b00000000000000001100000111010011;
assign LUT_3[2907] = 32'b00000000000000010010110010110000;
assign LUT_3[2908] = 32'b00000000000000000111001101100101;
assign LUT_3[2909] = 32'b00000000000000001101111001000010;
assign LUT_3[2910] = 32'b00000000000000001001010101001001;
assign LUT_3[2911] = 32'b00000000000000010000000000100110;
assign LUT_3[2912] = 32'b00000000000000000010100010000110;
assign LUT_3[2913] = 32'b00000000000000001001001101100011;
assign LUT_3[2914] = 32'b00000000000000000100101001101010;
assign LUT_3[2915] = 32'b00000000000000001011010101000111;
assign LUT_3[2916] = 32'b11111111111111111111101111111100;
assign LUT_3[2917] = 32'b00000000000000000110011011011001;
assign LUT_3[2918] = 32'b00000000000000000001110111100000;
assign LUT_3[2919] = 32'b00000000000000001000100010111101;
assign LUT_3[2920] = 32'b00000000000000000111111011001100;
assign LUT_3[2921] = 32'b00000000000000001110100110101001;
assign LUT_3[2922] = 32'b00000000000000001010000010110000;
assign LUT_3[2923] = 32'b00000000000000010000101110001101;
assign LUT_3[2924] = 32'b00000000000000000101001001000010;
assign LUT_3[2925] = 32'b00000000000000001011110100011111;
assign LUT_3[2926] = 32'b00000000000000000111010000100110;
assign LUT_3[2927] = 32'b00000000000000001101111100000011;
assign LUT_3[2928] = 32'b00000000000000000101110101001001;
assign LUT_3[2929] = 32'b00000000000000001100100000100110;
assign LUT_3[2930] = 32'b00000000000000000111111100101101;
assign LUT_3[2931] = 32'b00000000000000001110101000001010;
assign LUT_3[2932] = 32'b00000000000000000011000010111111;
assign LUT_3[2933] = 32'b00000000000000001001101110011100;
assign LUT_3[2934] = 32'b00000000000000000101001010100011;
assign LUT_3[2935] = 32'b00000000000000001011110110000000;
assign LUT_3[2936] = 32'b00000000000000001011001110001111;
assign LUT_3[2937] = 32'b00000000000000010001111001101100;
assign LUT_3[2938] = 32'b00000000000000001101010101110011;
assign LUT_3[2939] = 32'b00000000000000010100000001010000;
assign LUT_3[2940] = 32'b00000000000000001000011100000101;
assign LUT_3[2941] = 32'b00000000000000001111000111100010;
assign LUT_3[2942] = 32'b00000000000000001010100011101001;
assign LUT_3[2943] = 32'b00000000000000010001001111000110;
assign LUT_3[2944] = 32'b00000000000000000011100101111001;
assign LUT_3[2945] = 32'b00000000000000001010010001010110;
assign LUT_3[2946] = 32'b00000000000000000101101101011101;
assign LUT_3[2947] = 32'b00000000000000001100011000111010;
assign LUT_3[2948] = 32'b00000000000000000000110011101111;
assign LUT_3[2949] = 32'b00000000000000000111011111001100;
assign LUT_3[2950] = 32'b00000000000000000010111011010011;
assign LUT_3[2951] = 32'b00000000000000001001100110110000;
assign LUT_3[2952] = 32'b00000000000000001000111110111111;
assign LUT_3[2953] = 32'b00000000000000001111101010011100;
assign LUT_3[2954] = 32'b00000000000000001011000110100011;
assign LUT_3[2955] = 32'b00000000000000010001110010000000;
assign LUT_3[2956] = 32'b00000000000000000110001100110101;
assign LUT_3[2957] = 32'b00000000000000001100111000010010;
assign LUT_3[2958] = 32'b00000000000000001000010100011001;
assign LUT_3[2959] = 32'b00000000000000001110111111110110;
assign LUT_3[2960] = 32'b00000000000000000110111000111100;
assign LUT_3[2961] = 32'b00000000000000001101100100011001;
assign LUT_3[2962] = 32'b00000000000000001001000000100000;
assign LUT_3[2963] = 32'b00000000000000001111101011111101;
assign LUT_3[2964] = 32'b00000000000000000100000110110010;
assign LUT_3[2965] = 32'b00000000000000001010110010001111;
assign LUT_3[2966] = 32'b00000000000000000110001110010110;
assign LUT_3[2967] = 32'b00000000000000001100111001110011;
assign LUT_3[2968] = 32'b00000000000000001100010010000010;
assign LUT_3[2969] = 32'b00000000000000010010111101011111;
assign LUT_3[2970] = 32'b00000000000000001110011001100110;
assign LUT_3[2971] = 32'b00000000000000010101000101000011;
assign LUT_3[2972] = 32'b00000000000000001001011111111000;
assign LUT_3[2973] = 32'b00000000000000010000001011010101;
assign LUT_3[2974] = 32'b00000000000000001011100111011100;
assign LUT_3[2975] = 32'b00000000000000010010010010111001;
assign LUT_3[2976] = 32'b00000000000000000100110100011001;
assign LUT_3[2977] = 32'b00000000000000001011011111110110;
assign LUT_3[2978] = 32'b00000000000000000110111011111101;
assign LUT_3[2979] = 32'b00000000000000001101100111011010;
assign LUT_3[2980] = 32'b00000000000000000010000010001111;
assign LUT_3[2981] = 32'b00000000000000001000101101101100;
assign LUT_3[2982] = 32'b00000000000000000100001001110011;
assign LUT_3[2983] = 32'b00000000000000001010110101010000;
assign LUT_3[2984] = 32'b00000000000000001010001101011111;
assign LUT_3[2985] = 32'b00000000000000010000111000111100;
assign LUT_3[2986] = 32'b00000000000000001100010101000011;
assign LUT_3[2987] = 32'b00000000000000010011000000100000;
assign LUT_3[2988] = 32'b00000000000000000111011011010101;
assign LUT_3[2989] = 32'b00000000000000001110000110110010;
assign LUT_3[2990] = 32'b00000000000000001001100010111001;
assign LUT_3[2991] = 32'b00000000000000010000001110010110;
assign LUT_3[2992] = 32'b00000000000000001000000111011100;
assign LUT_3[2993] = 32'b00000000000000001110110010111001;
assign LUT_3[2994] = 32'b00000000000000001010001111000000;
assign LUT_3[2995] = 32'b00000000000000010000111010011101;
assign LUT_3[2996] = 32'b00000000000000000101010101010010;
assign LUT_3[2997] = 32'b00000000000000001100000000101111;
assign LUT_3[2998] = 32'b00000000000000000111011100110110;
assign LUT_3[2999] = 32'b00000000000000001110001000010011;
assign LUT_3[3000] = 32'b00000000000000001101100000100010;
assign LUT_3[3001] = 32'b00000000000000010100001011111111;
assign LUT_3[3002] = 32'b00000000000000001111101000000110;
assign LUT_3[3003] = 32'b00000000000000010110010011100011;
assign LUT_3[3004] = 32'b00000000000000001010101110011000;
assign LUT_3[3005] = 32'b00000000000000010001011001110101;
assign LUT_3[3006] = 32'b00000000000000001100110101111100;
assign LUT_3[3007] = 32'b00000000000000010011100001011001;
assign LUT_3[3008] = 32'b00000000000000000011011110100100;
assign LUT_3[3009] = 32'b00000000000000001010001010000001;
assign LUT_3[3010] = 32'b00000000000000000101100110001000;
assign LUT_3[3011] = 32'b00000000000000001100010001100101;
assign LUT_3[3012] = 32'b00000000000000000000101100011010;
assign LUT_3[3013] = 32'b00000000000000000111010111110111;
assign LUT_3[3014] = 32'b00000000000000000010110011111110;
assign LUT_3[3015] = 32'b00000000000000001001011111011011;
assign LUT_3[3016] = 32'b00000000000000001000110111101010;
assign LUT_3[3017] = 32'b00000000000000001111100011000111;
assign LUT_3[3018] = 32'b00000000000000001010111111001110;
assign LUT_3[3019] = 32'b00000000000000010001101010101011;
assign LUT_3[3020] = 32'b00000000000000000110000101100000;
assign LUT_3[3021] = 32'b00000000000000001100110000111101;
assign LUT_3[3022] = 32'b00000000000000001000001101000100;
assign LUT_3[3023] = 32'b00000000000000001110111000100001;
assign LUT_3[3024] = 32'b00000000000000000110110001100111;
assign LUT_3[3025] = 32'b00000000000000001101011101000100;
assign LUT_3[3026] = 32'b00000000000000001000111001001011;
assign LUT_3[3027] = 32'b00000000000000001111100100101000;
assign LUT_3[3028] = 32'b00000000000000000011111111011101;
assign LUT_3[3029] = 32'b00000000000000001010101010111010;
assign LUT_3[3030] = 32'b00000000000000000110000111000001;
assign LUT_3[3031] = 32'b00000000000000001100110010011110;
assign LUT_3[3032] = 32'b00000000000000001100001010101101;
assign LUT_3[3033] = 32'b00000000000000010010110110001010;
assign LUT_3[3034] = 32'b00000000000000001110010010010001;
assign LUT_3[3035] = 32'b00000000000000010100111101101110;
assign LUT_3[3036] = 32'b00000000000000001001011000100011;
assign LUT_3[3037] = 32'b00000000000000010000000100000000;
assign LUT_3[3038] = 32'b00000000000000001011100000000111;
assign LUT_3[3039] = 32'b00000000000000010010001011100100;
assign LUT_3[3040] = 32'b00000000000000000100101101000100;
assign LUT_3[3041] = 32'b00000000000000001011011000100001;
assign LUT_3[3042] = 32'b00000000000000000110110100101000;
assign LUT_3[3043] = 32'b00000000000000001101100000000101;
assign LUT_3[3044] = 32'b00000000000000000001111010111010;
assign LUT_3[3045] = 32'b00000000000000001000100110010111;
assign LUT_3[3046] = 32'b00000000000000000100000010011110;
assign LUT_3[3047] = 32'b00000000000000001010101101111011;
assign LUT_3[3048] = 32'b00000000000000001010000110001010;
assign LUT_3[3049] = 32'b00000000000000010000110001100111;
assign LUT_3[3050] = 32'b00000000000000001100001101101110;
assign LUT_3[3051] = 32'b00000000000000010010111001001011;
assign LUT_3[3052] = 32'b00000000000000000111010100000000;
assign LUT_3[3053] = 32'b00000000000000001101111111011101;
assign LUT_3[3054] = 32'b00000000000000001001011011100100;
assign LUT_3[3055] = 32'b00000000000000010000000111000001;
assign LUT_3[3056] = 32'b00000000000000001000000000000111;
assign LUT_3[3057] = 32'b00000000000000001110101011100100;
assign LUT_3[3058] = 32'b00000000000000001010000111101011;
assign LUT_3[3059] = 32'b00000000000000010000110011001000;
assign LUT_3[3060] = 32'b00000000000000000101001101111101;
assign LUT_3[3061] = 32'b00000000000000001011111001011010;
assign LUT_3[3062] = 32'b00000000000000000111010101100001;
assign LUT_3[3063] = 32'b00000000000000001110000000111110;
assign LUT_3[3064] = 32'b00000000000000001101011001001101;
assign LUT_3[3065] = 32'b00000000000000010100000100101010;
assign LUT_3[3066] = 32'b00000000000000001111100000110001;
assign LUT_3[3067] = 32'b00000000000000010110001100001110;
assign LUT_3[3068] = 32'b00000000000000001010100111000011;
assign LUT_3[3069] = 32'b00000000000000010001010010100000;
assign LUT_3[3070] = 32'b00000000000000001100101110100111;
assign LUT_3[3071] = 32'b00000000000000010011011010000100;
assign LUT_3[3072] = 32'b00000000000000001000011011001011;
assign LUT_3[3073] = 32'b00000000000000001111000110101000;
assign LUT_3[3074] = 32'b00000000000000001010100010101111;
assign LUT_3[3075] = 32'b00000000000000010001001110001100;
assign LUT_3[3076] = 32'b00000000000000000101101001000001;
assign LUT_3[3077] = 32'b00000000000000001100010100011110;
assign LUT_3[3078] = 32'b00000000000000000111110000100101;
assign LUT_3[3079] = 32'b00000000000000001110011100000010;
assign LUT_3[3080] = 32'b00000000000000001101110100010001;
assign LUT_3[3081] = 32'b00000000000000010100011111101110;
assign LUT_3[3082] = 32'b00000000000000001111111011110101;
assign LUT_3[3083] = 32'b00000000000000010110100111010010;
assign LUT_3[3084] = 32'b00000000000000001011000010000111;
assign LUT_3[3085] = 32'b00000000000000010001101101100100;
assign LUT_3[3086] = 32'b00000000000000001101001001101011;
assign LUT_3[3087] = 32'b00000000000000010011110101001000;
assign LUT_3[3088] = 32'b00000000000000001011101110001110;
assign LUT_3[3089] = 32'b00000000000000010010011001101011;
assign LUT_3[3090] = 32'b00000000000000001101110101110010;
assign LUT_3[3091] = 32'b00000000000000010100100001001111;
assign LUT_3[3092] = 32'b00000000000000001000111100000100;
assign LUT_3[3093] = 32'b00000000000000001111100111100001;
assign LUT_3[3094] = 32'b00000000000000001011000011101000;
assign LUT_3[3095] = 32'b00000000000000010001101111000101;
assign LUT_3[3096] = 32'b00000000000000010001000111010100;
assign LUT_3[3097] = 32'b00000000000000010111110010110001;
assign LUT_3[3098] = 32'b00000000000000010011001110111000;
assign LUT_3[3099] = 32'b00000000000000011001111010010101;
assign LUT_3[3100] = 32'b00000000000000001110010101001010;
assign LUT_3[3101] = 32'b00000000000000010101000000100111;
assign LUT_3[3102] = 32'b00000000000000010000011100101110;
assign LUT_3[3103] = 32'b00000000000000010111001000001011;
assign LUT_3[3104] = 32'b00000000000000001001101001101011;
assign LUT_3[3105] = 32'b00000000000000010000010101001000;
assign LUT_3[3106] = 32'b00000000000000001011110001001111;
assign LUT_3[3107] = 32'b00000000000000010010011100101100;
assign LUT_3[3108] = 32'b00000000000000000110110111100001;
assign LUT_3[3109] = 32'b00000000000000001101100010111110;
assign LUT_3[3110] = 32'b00000000000000001000111111000101;
assign LUT_3[3111] = 32'b00000000000000001111101010100010;
assign LUT_3[3112] = 32'b00000000000000001111000010110001;
assign LUT_3[3113] = 32'b00000000000000010101101110001110;
assign LUT_3[3114] = 32'b00000000000000010001001010010101;
assign LUT_3[3115] = 32'b00000000000000010111110101110010;
assign LUT_3[3116] = 32'b00000000000000001100010000100111;
assign LUT_3[3117] = 32'b00000000000000010010111100000100;
assign LUT_3[3118] = 32'b00000000000000001110011000001011;
assign LUT_3[3119] = 32'b00000000000000010101000011101000;
assign LUT_3[3120] = 32'b00000000000000001100111100101110;
assign LUT_3[3121] = 32'b00000000000000010011101000001011;
assign LUT_3[3122] = 32'b00000000000000001111000100010010;
assign LUT_3[3123] = 32'b00000000000000010101101111101111;
assign LUT_3[3124] = 32'b00000000000000001010001010100100;
assign LUT_3[3125] = 32'b00000000000000010000110110000001;
assign LUT_3[3126] = 32'b00000000000000001100010010001000;
assign LUT_3[3127] = 32'b00000000000000010010111101100101;
assign LUT_3[3128] = 32'b00000000000000010010010101110100;
assign LUT_3[3129] = 32'b00000000000000011001000001010001;
assign LUT_3[3130] = 32'b00000000000000010100011101011000;
assign LUT_3[3131] = 32'b00000000000000011011001000110101;
assign LUT_3[3132] = 32'b00000000000000001111100011101010;
assign LUT_3[3133] = 32'b00000000000000010110001111000111;
assign LUT_3[3134] = 32'b00000000000000010001101011001110;
assign LUT_3[3135] = 32'b00000000000000011000010110101011;
assign LUT_3[3136] = 32'b00000000000000001000010011110110;
assign LUT_3[3137] = 32'b00000000000000001110111111010011;
assign LUT_3[3138] = 32'b00000000000000001010011011011010;
assign LUT_3[3139] = 32'b00000000000000010001000110110111;
assign LUT_3[3140] = 32'b00000000000000000101100001101100;
assign LUT_3[3141] = 32'b00000000000000001100001101001001;
assign LUT_3[3142] = 32'b00000000000000000111101001010000;
assign LUT_3[3143] = 32'b00000000000000001110010100101101;
assign LUT_3[3144] = 32'b00000000000000001101101100111100;
assign LUT_3[3145] = 32'b00000000000000010100011000011001;
assign LUT_3[3146] = 32'b00000000000000001111110100100000;
assign LUT_3[3147] = 32'b00000000000000010110011111111101;
assign LUT_3[3148] = 32'b00000000000000001010111010110010;
assign LUT_3[3149] = 32'b00000000000000010001100110001111;
assign LUT_3[3150] = 32'b00000000000000001101000010010110;
assign LUT_3[3151] = 32'b00000000000000010011101101110011;
assign LUT_3[3152] = 32'b00000000000000001011100110111001;
assign LUT_3[3153] = 32'b00000000000000010010010010010110;
assign LUT_3[3154] = 32'b00000000000000001101101110011101;
assign LUT_3[3155] = 32'b00000000000000010100011001111010;
assign LUT_3[3156] = 32'b00000000000000001000110100101111;
assign LUT_3[3157] = 32'b00000000000000001111100000001100;
assign LUT_3[3158] = 32'b00000000000000001010111100010011;
assign LUT_3[3159] = 32'b00000000000000010001100111110000;
assign LUT_3[3160] = 32'b00000000000000010000111111111111;
assign LUT_3[3161] = 32'b00000000000000010111101011011100;
assign LUT_3[3162] = 32'b00000000000000010011000111100011;
assign LUT_3[3163] = 32'b00000000000000011001110011000000;
assign LUT_3[3164] = 32'b00000000000000001110001101110101;
assign LUT_3[3165] = 32'b00000000000000010100111001010010;
assign LUT_3[3166] = 32'b00000000000000010000010101011001;
assign LUT_3[3167] = 32'b00000000000000010111000000110110;
assign LUT_3[3168] = 32'b00000000000000001001100010010110;
assign LUT_3[3169] = 32'b00000000000000010000001101110011;
assign LUT_3[3170] = 32'b00000000000000001011101001111010;
assign LUT_3[3171] = 32'b00000000000000010010010101010111;
assign LUT_3[3172] = 32'b00000000000000000110110000001100;
assign LUT_3[3173] = 32'b00000000000000001101011011101001;
assign LUT_3[3174] = 32'b00000000000000001000110111110000;
assign LUT_3[3175] = 32'b00000000000000001111100011001101;
assign LUT_3[3176] = 32'b00000000000000001110111011011100;
assign LUT_3[3177] = 32'b00000000000000010101100110111001;
assign LUT_3[3178] = 32'b00000000000000010001000011000000;
assign LUT_3[3179] = 32'b00000000000000010111101110011101;
assign LUT_3[3180] = 32'b00000000000000001100001001010010;
assign LUT_3[3181] = 32'b00000000000000010010110100101111;
assign LUT_3[3182] = 32'b00000000000000001110010000110110;
assign LUT_3[3183] = 32'b00000000000000010100111100010011;
assign LUT_3[3184] = 32'b00000000000000001100110101011001;
assign LUT_3[3185] = 32'b00000000000000010011100000110110;
assign LUT_3[3186] = 32'b00000000000000001110111100111101;
assign LUT_3[3187] = 32'b00000000000000010101101000011010;
assign LUT_3[3188] = 32'b00000000000000001010000011001111;
assign LUT_3[3189] = 32'b00000000000000010000101110101100;
assign LUT_3[3190] = 32'b00000000000000001100001010110011;
assign LUT_3[3191] = 32'b00000000000000010010110110010000;
assign LUT_3[3192] = 32'b00000000000000010010001110011111;
assign LUT_3[3193] = 32'b00000000000000011000111001111100;
assign LUT_3[3194] = 32'b00000000000000010100010110000011;
assign LUT_3[3195] = 32'b00000000000000011011000001100000;
assign LUT_3[3196] = 32'b00000000000000001111011100010101;
assign LUT_3[3197] = 32'b00000000000000010110000111110010;
assign LUT_3[3198] = 32'b00000000000000010001100011111001;
assign LUT_3[3199] = 32'b00000000000000011000001111010110;
assign LUT_3[3200] = 32'b00000000000000001010100110001001;
assign LUT_3[3201] = 32'b00000000000000010001010001100110;
assign LUT_3[3202] = 32'b00000000000000001100101101101101;
assign LUT_3[3203] = 32'b00000000000000010011011001001010;
assign LUT_3[3204] = 32'b00000000000000000111110011111111;
assign LUT_3[3205] = 32'b00000000000000001110011111011100;
assign LUT_3[3206] = 32'b00000000000000001001111011100011;
assign LUT_3[3207] = 32'b00000000000000010000100111000000;
assign LUT_3[3208] = 32'b00000000000000001111111111001111;
assign LUT_3[3209] = 32'b00000000000000010110101010101100;
assign LUT_3[3210] = 32'b00000000000000010010000110110011;
assign LUT_3[3211] = 32'b00000000000000011000110010010000;
assign LUT_3[3212] = 32'b00000000000000001101001101000101;
assign LUT_3[3213] = 32'b00000000000000010011111000100010;
assign LUT_3[3214] = 32'b00000000000000001111010100101001;
assign LUT_3[3215] = 32'b00000000000000010110000000000110;
assign LUT_3[3216] = 32'b00000000000000001101111001001100;
assign LUT_3[3217] = 32'b00000000000000010100100100101001;
assign LUT_3[3218] = 32'b00000000000000010000000000110000;
assign LUT_3[3219] = 32'b00000000000000010110101100001101;
assign LUT_3[3220] = 32'b00000000000000001011000111000010;
assign LUT_3[3221] = 32'b00000000000000010001110010011111;
assign LUT_3[3222] = 32'b00000000000000001101001110100110;
assign LUT_3[3223] = 32'b00000000000000010011111010000011;
assign LUT_3[3224] = 32'b00000000000000010011010010010010;
assign LUT_3[3225] = 32'b00000000000000011001111101101111;
assign LUT_3[3226] = 32'b00000000000000010101011001110110;
assign LUT_3[3227] = 32'b00000000000000011100000101010011;
assign LUT_3[3228] = 32'b00000000000000010000100000001000;
assign LUT_3[3229] = 32'b00000000000000010111001011100101;
assign LUT_3[3230] = 32'b00000000000000010010100111101100;
assign LUT_3[3231] = 32'b00000000000000011001010011001001;
assign LUT_3[3232] = 32'b00000000000000001011110100101001;
assign LUT_3[3233] = 32'b00000000000000010010100000000110;
assign LUT_3[3234] = 32'b00000000000000001101111100001101;
assign LUT_3[3235] = 32'b00000000000000010100100111101010;
assign LUT_3[3236] = 32'b00000000000000001001000010011111;
assign LUT_3[3237] = 32'b00000000000000001111101101111100;
assign LUT_3[3238] = 32'b00000000000000001011001010000011;
assign LUT_3[3239] = 32'b00000000000000010001110101100000;
assign LUT_3[3240] = 32'b00000000000000010001001101101111;
assign LUT_3[3241] = 32'b00000000000000010111111001001100;
assign LUT_3[3242] = 32'b00000000000000010011010101010011;
assign LUT_3[3243] = 32'b00000000000000011010000000110000;
assign LUT_3[3244] = 32'b00000000000000001110011011100101;
assign LUT_3[3245] = 32'b00000000000000010101000111000010;
assign LUT_3[3246] = 32'b00000000000000010000100011001001;
assign LUT_3[3247] = 32'b00000000000000010111001110100110;
assign LUT_3[3248] = 32'b00000000000000001111000111101100;
assign LUT_3[3249] = 32'b00000000000000010101110011001001;
assign LUT_3[3250] = 32'b00000000000000010001001111010000;
assign LUT_3[3251] = 32'b00000000000000010111111010101101;
assign LUT_3[3252] = 32'b00000000000000001100010101100010;
assign LUT_3[3253] = 32'b00000000000000010011000000111111;
assign LUT_3[3254] = 32'b00000000000000001110011101000110;
assign LUT_3[3255] = 32'b00000000000000010101001000100011;
assign LUT_3[3256] = 32'b00000000000000010100100000110010;
assign LUT_3[3257] = 32'b00000000000000011011001100001111;
assign LUT_3[3258] = 32'b00000000000000010110101000010110;
assign LUT_3[3259] = 32'b00000000000000011101010011110011;
assign LUT_3[3260] = 32'b00000000000000010001101110101000;
assign LUT_3[3261] = 32'b00000000000000011000011010000101;
assign LUT_3[3262] = 32'b00000000000000010011110110001100;
assign LUT_3[3263] = 32'b00000000000000011010100001101001;
assign LUT_3[3264] = 32'b00000000000000001010011110110100;
assign LUT_3[3265] = 32'b00000000000000010001001010010001;
assign LUT_3[3266] = 32'b00000000000000001100100110011000;
assign LUT_3[3267] = 32'b00000000000000010011010001110101;
assign LUT_3[3268] = 32'b00000000000000000111101100101010;
assign LUT_3[3269] = 32'b00000000000000001110011000000111;
assign LUT_3[3270] = 32'b00000000000000001001110100001110;
assign LUT_3[3271] = 32'b00000000000000010000011111101011;
assign LUT_3[3272] = 32'b00000000000000001111110111111010;
assign LUT_3[3273] = 32'b00000000000000010110100011010111;
assign LUT_3[3274] = 32'b00000000000000010001111111011110;
assign LUT_3[3275] = 32'b00000000000000011000101010111011;
assign LUT_3[3276] = 32'b00000000000000001101000101110000;
assign LUT_3[3277] = 32'b00000000000000010011110001001101;
assign LUT_3[3278] = 32'b00000000000000001111001101010100;
assign LUT_3[3279] = 32'b00000000000000010101111000110001;
assign LUT_3[3280] = 32'b00000000000000001101110001110111;
assign LUT_3[3281] = 32'b00000000000000010100011101010100;
assign LUT_3[3282] = 32'b00000000000000001111111001011011;
assign LUT_3[3283] = 32'b00000000000000010110100100111000;
assign LUT_3[3284] = 32'b00000000000000001010111111101101;
assign LUT_3[3285] = 32'b00000000000000010001101011001010;
assign LUT_3[3286] = 32'b00000000000000001101000111010001;
assign LUT_3[3287] = 32'b00000000000000010011110010101110;
assign LUT_3[3288] = 32'b00000000000000010011001010111101;
assign LUT_3[3289] = 32'b00000000000000011001110110011010;
assign LUT_3[3290] = 32'b00000000000000010101010010100001;
assign LUT_3[3291] = 32'b00000000000000011011111101111110;
assign LUT_3[3292] = 32'b00000000000000010000011000110011;
assign LUT_3[3293] = 32'b00000000000000010111000100010000;
assign LUT_3[3294] = 32'b00000000000000010010100000010111;
assign LUT_3[3295] = 32'b00000000000000011001001011110100;
assign LUT_3[3296] = 32'b00000000000000001011101101010100;
assign LUT_3[3297] = 32'b00000000000000010010011000110001;
assign LUT_3[3298] = 32'b00000000000000001101110100111000;
assign LUT_3[3299] = 32'b00000000000000010100100000010101;
assign LUT_3[3300] = 32'b00000000000000001000111011001010;
assign LUT_3[3301] = 32'b00000000000000001111100110100111;
assign LUT_3[3302] = 32'b00000000000000001011000010101110;
assign LUT_3[3303] = 32'b00000000000000010001101110001011;
assign LUT_3[3304] = 32'b00000000000000010001000110011010;
assign LUT_3[3305] = 32'b00000000000000010111110001110111;
assign LUT_3[3306] = 32'b00000000000000010011001101111110;
assign LUT_3[3307] = 32'b00000000000000011001111001011011;
assign LUT_3[3308] = 32'b00000000000000001110010100010000;
assign LUT_3[3309] = 32'b00000000000000010100111111101101;
assign LUT_3[3310] = 32'b00000000000000010000011011110100;
assign LUT_3[3311] = 32'b00000000000000010111000111010001;
assign LUT_3[3312] = 32'b00000000000000001111000000010111;
assign LUT_3[3313] = 32'b00000000000000010101101011110100;
assign LUT_3[3314] = 32'b00000000000000010001000111111011;
assign LUT_3[3315] = 32'b00000000000000010111110011011000;
assign LUT_3[3316] = 32'b00000000000000001100001110001101;
assign LUT_3[3317] = 32'b00000000000000010010111001101010;
assign LUT_3[3318] = 32'b00000000000000001110010101110001;
assign LUT_3[3319] = 32'b00000000000000010101000001001110;
assign LUT_3[3320] = 32'b00000000000000010100011001011101;
assign LUT_3[3321] = 32'b00000000000000011011000100111010;
assign LUT_3[3322] = 32'b00000000000000010110100001000001;
assign LUT_3[3323] = 32'b00000000000000011101001100011110;
assign LUT_3[3324] = 32'b00000000000000010001100111010011;
assign LUT_3[3325] = 32'b00000000000000011000010010110000;
assign LUT_3[3326] = 32'b00000000000000010011101110110111;
assign LUT_3[3327] = 32'b00000000000000011010011010010100;
assign LUT_3[3328] = 32'b00000000000000000100101010101100;
assign LUT_3[3329] = 32'b00000000000000001011010110001001;
assign LUT_3[3330] = 32'b00000000000000000110110010010000;
assign LUT_3[3331] = 32'b00000000000000001101011101101101;
assign LUT_3[3332] = 32'b00000000000000000001111000100010;
assign LUT_3[3333] = 32'b00000000000000001000100011111111;
assign LUT_3[3334] = 32'b00000000000000000100000000000110;
assign LUT_3[3335] = 32'b00000000000000001010101011100011;
assign LUT_3[3336] = 32'b00000000000000001010000011110010;
assign LUT_3[3337] = 32'b00000000000000010000101111001111;
assign LUT_3[3338] = 32'b00000000000000001100001011010110;
assign LUT_3[3339] = 32'b00000000000000010010110110110011;
assign LUT_3[3340] = 32'b00000000000000000111010001101000;
assign LUT_3[3341] = 32'b00000000000000001101111101000101;
assign LUT_3[3342] = 32'b00000000000000001001011001001100;
assign LUT_3[3343] = 32'b00000000000000010000000100101001;
assign LUT_3[3344] = 32'b00000000000000000111111101101111;
assign LUT_3[3345] = 32'b00000000000000001110101001001100;
assign LUT_3[3346] = 32'b00000000000000001010000101010011;
assign LUT_3[3347] = 32'b00000000000000010000110000110000;
assign LUT_3[3348] = 32'b00000000000000000101001011100101;
assign LUT_3[3349] = 32'b00000000000000001011110111000010;
assign LUT_3[3350] = 32'b00000000000000000111010011001001;
assign LUT_3[3351] = 32'b00000000000000001101111110100110;
assign LUT_3[3352] = 32'b00000000000000001101010110110101;
assign LUT_3[3353] = 32'b00000000000000010100000010010010;
assign LUT_3[3354] = 32'b00000000000000001111011110011001;
assign LUT_3[3355] = 32'b00000000000000010110001001110110;
assign LUT_3[3356] = 32'b00000000000000001010100100101011;
assign LUT_3[3357] = 32'b00000000000000010001010000001000;
assign LUT_3[3358] = 32'b00000000000000001100101100001111;
assign LUT_3[3359] = 32'b00000000000000010011010111101100;
assign LUT_3[3360] = 32'b00000000000000000101111001001100;
assign LUT_3[3361] = 32'b00000000000000001100100100101001;
assign LUT_3[3362] = 32'b00000000000000001000000000110000;
assign LUT_3[3363] = 32'b00000000000000001110101100001101;
assign LUT_3[3364] = 32'b00000000000000000011000111000010;
assign LUT_3[3365] = 32'b00000000000000001001110010011111;
assign LUT_3[3366] = 32'b00000000000000000101001110100110;
assign LUT_3[3367] = 32'b00000000000000001011111010000011;
assign LUT_3[3368] = 32'b00000000000000001011010010010010;
assign LUT_3[3369] = 32'b00000000000000010001111101101111;
assign LUT_3[3370] = 32'b00000000000000001101011001110110;
assign LUT_3[3371] = 32'b00000000000000010100000101010011;
assign LUT_3[3372] = 32'b00000000000000001000100000001000;
assign LUT_3[3373] = 32'b00000000000000001111001011100101;
assign LUT_3[3374] = 32'b00000000000000001010100111101100;
assign LUT_3[3375] = 32'b00000000000000010001010011001001;
assign LUT_3[3376] = 32'b00000000000000001001001100001111;
assign LUT_3[3377] = 32'b00000000000000001111110111101100;
assign LUT_3[3378] = 32'b00000000000000001011010011110011;
assign LUT_3[3379] = 32'b00000000000000010001111111010000;
assign LUT_3[3380] = 32'b00000000000000000110011010000101;
assign LUT_3[3381] = 32'b00000000000000001101000101100010;
assign LUT_3[3382] = 32'b00000000000000001000100001101001;
assign LUT_3[3383] = 32'b00000000000000001111001101000110;
assign LUT_3[3384] = 32'b00000000000000001110100101010101;
assign LUT_3[3385] = 32'b00000000000000010101010000110010;
assign LUT_3[3386] = 32'b00000000000000010000101100111001;
assign LUT_3[3387] = 32'b00000000000000010111011000010110;
assign LUT_3[3388] = 32'b00000000000000001011110011001011;
assign LUT_3[3389] = 32'b00000000000000010010011110101000;
assign LUT_3[3390] = 32'b00000000000000001101111010101111;
assign LUT_3[3391] = 32'b00000000000000010100100110001100;
assign LUT_3[3392] = 32'b00000000000000000100100011010111;
assign LUT_3[3393] = 32'b00000000000000001011001110110100;
assign LUT_3[3394] = 32'b00000000000000000110101010111011;
assign LUT_3[3395] = 32'b00000000000000001101010110011000;
assign LUT_3[3396] = 32'b00000000000000000001110001001101;
assign LUT_3[3397] = 32'b00000000000000001000011100101010;
assign LUT_3[3398] = 32'b00000000000000000011111000110001;
assign LUT_3[3399] = 32'b00000000000000001010100100001110;
assign LUT_3[3400] = 32'b00000000000000001001111100011101;
assign LUT_3[3401] = 32'b00000000000000010000100111111010;
assign LUT_3[3402] = 32'b00000000000000001100000100000001;
assign LUT_3[3403] = 32'b00000000000000010010101111011110;
assign LUT_3[3404] = 32'b00000000000000000111001010010011;
assign LUT_3[3405] = 32'b00000000000000001101110101110000;
assign LUT_3[3406] = 32'b00000000000000001001010001110111;
assign LUT_3[3407] = 32'b00000000000000001111111101010100;
assign LUT_3[3408] = 32'b00000000000000000111110110011010;
assign LUT_3[3409] = 32'b00000000000000001110100001110111;
assign LUT_3[3410] = 32'b00000000000000001001111101111110;
assign LUT_3[3411] = 32'b00000000000000010000101001011011;
assign LUT_3[3412] = 32'b00000000000000000101000100010000;
assign LUT_3[3413] = 32'b00000000000000001011101111101101;
assign LUT_3[3414] = 32'b00000000000000000111001011110100;
assign LUT_3[3415] = 32'b00000000000000001101110111010001;
assign LUT_3[3416] = 32'b00000000000000001101001111100000;
assign LUT_3[3417] = 32'b00000000000000010011111010111101;
assign LUT_3[3418] = 32'b00000000000000001111010111000100;
assign LUT_3[3419] = 32'b00000000000000010110000010100001;
assign LUT_3[3420] = 32'b00000000000000001010011101010110;
assign LUT_3[3421] = 32'b00000000000000010001001000110011;
assign LUT_3[3422] = 32'b00000000000000001100100100111010;
assign LUT_3[3423] = 32'b00000000000000010011010000010111;
assign LUT_3[3424] = 32'b00000000000000000101110001110111;
assign LUT_3[3425] = 32'b00000000000000001100011101010100;
assign LUT_3[3426] = 32'b00000000000000000111111001011011;
assign LUT_3[3427] = 32'b00000000000000001110100100111000;
assign LUT_3[3428] = 32'b00000000000000000010111111101101;
assign LUT_3[3429] = 32'b00000000000000001001101011001010;
assign LUT_3[3430] = 32'b00000000000000000101000111010001;
assign LUT_3[3431] = 32'b00000000000000001011110010101110;
assign LUT_3[3432] = 32'b00000000000000001011001010111101;
assign LUT_3[3433] = 32'b00000000000000010001110110011010;
assign LUT_3[3434] = 32'b00000000000000001101010010100001;
assign LUT_3[3435] = 32'b00000000000000010011111101111110;
assign LUT_3[3436] = 32'b00000000000000001000011000110011;
assign LUT_3[3437] = 32'b00000000000000001111000100010000;
assign LUT_3[3438] = 32'b00000000000000001010100000010111;
assign LUT_3[3439] = 32'b00000000000000010001001011110100;
assign LUT_3[3440] = 32'b00000000000000001001000100111010;
assign LUT_3[3441] = 32'b00000000000000001111110000010111;
assign LUT_3[3442] = 32'b00000000000000001011001100011110;
assign LUT_3[3443] = 32'b00000000000000010001110111111011;
assign LUT_3[3444] = 32'b00000000000000000110010010110000;
assign LUT_3[3445] = 32'b00000000000000001100111110001101;
assign LUT_3[3446] = 32'b00000000000000001000011010010100;
assign LUT_3[3447] = 32'b00000000000000001111000101110001;
assign LUT_3[3448] = 32'b00000000000000001110011110000000;
assign LUT_3[3449] = 32'b00000000000000010101001001011101;
assign LUT_3[3450] = 32'b00000000000000010000100101100100;
assign LUT_3[3451] = 32'b00000000000000010111010001000001;
assign LUT_3[3452] = 32'b00000000000000001011101011110110;
assign LUT_3[3453] = 32'b00000000000000010010010111010011;
assign LUT_3[3454] = 32'b00000000000000001101110011011010;
assign LUT_3[3455] = 32'b00000000000000010100011110110111;
assign LUT_3[3456] = 32'b00000000000000000110110101101010;
assign LUT_3[3457] = 32'b00000000000000001101100001000111;
assign LUT_3[3458] = 32'b00000000000000001000111101001110;
assign LUT_3[3459] = 32'b00000000000000001111101000101011;
assign LUT_3[3460] = 32'b00000000000000000100000011100000;
assign LUT_3[3461] = 32'b00000000000000001010101110111101;
assign LUT_3[3462] = 32'b00000000000000000110001011000100;
assign LUT_3[3463] = 32'b00000000000000001100110110100001;
assign LUT_3[3464] = 32'b00000000000000001100001110110000;
assign LUT_3[3465] = 32'b00000000000000010010111010001101;
assign LUT_3[3466] = 32'b00000000000000001110010110010100;
assign LUT_3[3467] = 32'b00000000000000010101000001110001;
assign LUT_3[3468] = 32'b00000000000000001001011100100110;
assign LUT_3[3469] = 32'b00000000000000010000001000000011;
assign LUT_3[3470] = 32'b00000000000000001011100100001010;
assign LUT_3[3471] = 32'b00000000000000010010001111100111;
assign LUT_3[3472] = 32'b00000000000000001010001000101101;
assign LUT_3[3473] = 32'b00000000000000010000110100001010;
assign LUT_3[3474] = 32'b00000000000000001100010000010001;
assign LUT_3[3475] = 32'b00000000000000010010111011101110;
assign LUT_3[3476] = 32'b00000000000000000111010110100011;
assign LUT_3[3477] = 32'b00000000000000001110000010000000;
assign LUT_3[3478] = 32'b00000000000000001001011110000111;
assign LUT_3[3479] = 32'b00000000000000010000001001100100;
assign LUT_3[3480] = 32'b00000000000000001111100001110011;
assign LUT_3[3481] = 32'b00000000000000010110001101010000;
assign LUT_3[3482] = 32'b00000000000000010001101001010111;
assign LUT_3[3483] = 32'b00000000000000011000010100110100;
assign LUT_3[3484] = 32'b00000000000000001100101111101001;
assign LUT_3[3485] = 32'b00000000000000010011011011000110;
assign LUT_3[3486] = 32'b00000000000000001110110111001101;
assign LUT_3[3487] = 32'b00000000000000010101100010101010;
assign LUT_3[3488] = 32'b00000000000000001000000100001010;
assign LUT_3[3489] = 32'b00000000000000001110101111100111;
assign LUT_3[3490] = 32'b00000000000000001010001011101110;
assign LUT_3[3491] = 32'b00000000000000010000110111001011;
assign LUT_3[3492] = 32'b00000000000000000101010010000000;
assign LUT_3[3493] = 32'b00000000000000001011111101011101;
assign LUT_3[3494] = 32'b00000000000000000111011001100100;
assign LUT_3[3495] = 32'b00000000000000001110000101000001;
assign LUT_3[3496] = 32'b00000000000000001101011101010000;
assign LUT_3[3497] = 32'b00000000000000010100001000101101;
assign LUT_3[3498] = 32'b00000000000000001111100100110100;
assign LUT_3[3499] = 32'b00000000000000010110010000010001;
assign LUT_3[3500] = 32'b00000000000000001010101011000110;
assign LUT_3[3501] = 32'b00000000000000010001010110100011;
assign LUT_3[3502] = 32'b00000000000000001100110010101010;
assign LUT_3[3503] = 32'b00000000000000010011011110000111;
assign LUT_3[3504] = 32'b00000000000000001011010111001101;
assign LUT_3[3505] = 32'b00000000000000010010000010101010;
assign LUT_3[3506] = 32'b00000000000000001101011110110001;
assign LUT_3[3507] = 32'b00000000000000010100001010001110;
assign LUT_3[3508] = 32'b00000000000000001000100101000011;
assign LUT_3[3509] = 32'b00000000000000001111010000100000;
assign LUT_3[3510] = 32'b00000000000000001010101100100111;
assign LUT_3[3511] = 32'b00000000000000010001011000000100;
assign LUT_3[3512] = 32'b00000000000000010000110000010011;
assign LUT_3[3513] = 32'b00000000000000010111011011110000;
assign LUT_3[3514] = 32'b00000000000000010010110111110111;
assign LUT_3[3515] = 32'b00000000000000011001100011010100;
assign LUT_3[3516] = 32'b00000000000000001101111110001001;
assign LUT_3[3517] = 32'b00000000000000010100101001100110;
assign LUT_3[3518] = 32'b00000000000000010000000101101101;
assign LUT_3[3519] = 32'b00000000000000010110110001001010;
assign LUT_3[3520] = 32'b00000000000000000110101110010101;
assign LUT_3[3521] = 32'b00000000000000001101011001110010;
assign LUT_3[3522] = 32'b00000000000000001000110101111001;
assign LUT_3[3523] = 32'b00000000000000001111100001010110;
assign LUT_3[3524] = 32'b00000000000000000011111100001011;
assign LUT_3[3525] = 32'b00000000000000001010100111101000;
assign LUT_3[3526] = 32'b00000000000000000110000011101111;
assign LUT_3[3527] = 32'b00000000000000001100101111001100;
assign LUT_3[3528] = 32'b00000000000000001100000111011011;
assign LUT_3[3529] = 32'b00000000000000010010110010111000;
assign LUT_3[3530] = 32'b00000000000000001110001110111111;
assign LUT_3[3531] = 32'b00000000000000010100111010011100;
assign LUT_3[3532] = 32'b00000000000000001001010101010001;
assign LUT_3[3533] = 32'b00000000000000010000000000101110;
assign LUT_3[3534] = 32'b00000000000000001011011100110101;
assign LUT_3[3535] = 32'b00000000000000010010001000010010;
assign LUT_3[3536] = 32'b00000000000000001010000001011000;
assign LUT_3[3537] = 32'b00000000000000010000101100110101;
assign LUT_3[3538] = 32'b00000000000000001100001000111100;
assign LUT_3[3539] = 32'b00000000000000010010110100011001;
assign LUT_3[3540] = 32'b00000000000000000111001111001110;
assign LUT_3[3541] = 32'b00000000000000001101111010101011;
assign LUT_3[3542] = 32'b00000000000000001001010110110010;
assign LUT_3[3543] = 32'b00000000000000010000000010001111;
assign LUT_3[3544] = 32'b00000000000000001111011010011110;
assign LUT_3[3545] = 32'b00000000000000010110000101111011;
assign LUT_3[3546] = 32'b00000000000000010001100010000010;
assign LUT_3[3547] = 32'b00000000000000011000001101011111;
assign LUT_3[3548] = 32'b00000000000000001100101000010100;
assign LUT_3[3549] = 32'b00000000000000010011010011110001;
assign LUT_3[3550] = 32'b00000000000000001110101111111000;
assign LUT_3[3551] = 32'b00000000000000010101011011010101;
assign LUT_3[3552] = 32'b00000000000000000111111100110101;
assign LUT_3[3553] = 32'b00000000000000001110101000010010;
assign LUT_3[3554] = 32'b00000000000000001010000100011001;
assign LUT_3[3555] = 32'b00000000000000010000101111110110;
assign LUT_3[3556] = 32'b00000000000000000101001010101011;
assign LUT_3[3557] = 32'b00000000000000001011110110001000;
assign LUT_3[3558] = 32'b00000000000000000111010010001111;
assign LUT_3[3559] = 32'b00000000000000001101111101101100;
assign LUT_3[3560] = 32'b00000000000000001101010101111011;
assign LUT_3[3561] = 32'b00000000000000010100000001011000;
assign LUT_3[3562] = 32'b00000000000000001111011101011111;
assign LUT_3[3563] = 32'b00000000000000010110001000111100;
assign LUT_3[3564] = 32'b00000000000000001010100011110001;
assign LUT_3[3565] = 32'b00000000000000010001001111001110;
assign LUT_3[3566] = 32'b00000000000000001100101011010101;
assign LUT_3[3567] = 32'b00000000000000010011010110110010;
assign LUT_3[3568] = 32'b00000000000000001011001111111000;
assign LUT_3[3569] = 32'b00000000000000010001111011010101;
assign LUT_3[3570] = 32'b00000000000000001101010111011100;
assign LUT_3[3571] = 32'b00000000000000010100000010111001;
assign LUT_3[3572] = 32'b00000000000000001000011101101110;
assign LUT_3[3573] = 32'b00000000000000001111001001001011;
assign LUT_3[3574] = 32'b00000000000000001010100101010010;
assign LUT_3[3575] = 32'b00000000000000010001010000101111;
assign LUT_3[3576] = 32'b00000000000000010000101000111110;
assign LUT_3[3577] = 32'b00000000000000010111010100011011;
assign LUT_3[3578] = 32'b00000000000000010010110000100010;
assign LUT_3[3579] = 32'b00000000000000011001011011111111;
assign LUT_3[3580] = 32'b00000000000000001101110110110100;
assign LUT_3[3581] = 32'b00000000000000010100100010010001;
assign LUT_3[3582] = 32'b00000000000000001111111110011000;
assign LUT_3[3583] = 32'b00000000000000010110101001110101;
assign LUT_3[3584] = 32'b00000000000000001011110000010111;
assign LUT_3[3585] = 32'b00000000000000010010011011110100;
assign LUT_3[3586] = 32'b00000000000000001101110111111011;
assign LUT_3[3587] = 32'b00000000000000010100100011011000;
assign LUT_3[3588] = 32'b00000000000000001000111110001101;
assign LUT_3[3589] = 32'b00000000000000001111101001101010;
assign LUT_3[3590] = 32'b00000000000000001011000101110001;
assign LUT_3[3591] = 32'b00000000000000010001110001001110;
assign LUT_3[3592] = 32'b00000000000000010001001001011101;
assign LUT_3[3593] = 32'b00000000000000010111110100111010;
assign LUT_3[3594] = 32'b00000000000000010011010001000001;
assign LUT_3[3595] = 32'b00000000000000011001111100011110;
assign LUT_3[3596] = 32'b00000000000000001110010111010011;
assign LUT_3[3597] = 32'b00000000000000010101000010110000;
assign LUT_3[3598] = 32'b00000000000000010000011110110111;
assign LUT_3[3599] = 32'b00000000000000010111001010010100;
assign LUT_3[3600] = 32'b00000000000000001111000011011010;
assign LUT_3[3601] = 32'b00000000000000010101101110110111;
assign LUT_3[3602] = 32'b00000000000000010001001010111110;
assign LUT_3[3603] = 32'b00000000000000010111110110011011;
assign LUT_3[3604] = 32'b00000000000000001100010001010000;
assign LUT_3[3605] = 32'b00000000000000010010111100101101;
assign LUT_3[3606] = 32'b00000000000000001110011000110100;
assign LUT_3[3607] = 32'b00000000000000010101000100010001;
assign LUT_3[3608] = 32'b00000000000000010100011100100000;
assign LUT_3[3609] = 32'b00000000000000011011000111111101;
assign LUT_3[3610] = 32'b00000000000000010110100100000100;
assign LUT_3[3611] = 32'b00000000000000011101001111100001;
assign LUT_3[3612] = 32'b00000000000000010001101010010110;
assign LUT_3[3613] = 32'b00000000000000011000010101110011;
assign LUT_3[3614] = 32'b00000000000000010011110001111010;
assign LUT_3[3615] = 32'b00000000000000011010011101010111;
assign LUT_3[3616] = 32'b00000000000000001100111110110111;
assign LUT_3[3617] = 32'b00000000000000010011101010010100;
assign LUT_3[3618] = 32'b00000000000000001111000110011011;
assign LUT_3[3619] = 32'b00000000000000010101110001111000;
assign LUT_3[3620] = 32'b00000000000000001010001100101101;
assign LUT_3[3621] = 32'b00000000000000010000111000001010;
assign LUT_3[3622] = 32'b00000000000000001100010100010001;
assign LUT_3[3623] = 32'b00000000000000010010111111101110;
assign LUT_3[3624] = 32'b00000000000000010010010111111101;
assign LUT_3[3625] = 32'b00000000000000011001000011011010;
assign LUT_3[3626] = 32'b00000000000000010100011111100001;
assign LUT_3[3627] = 32'b00000000000000011011001010111110;
assign LUT_3[3628] = 32'b00000000000000001111100101110011;
assign LUT_3[3629] = 32'b00000000000000010110010001010000;
assign LUT_3[3630] = 32'b00000000000000010001101101010111;
assign LUT_3[3631] = 32'b00000000000000011000011000110100;
assign LUT_3[3632] = 32'b00000000000000010000010001111010;
assign LUT_3[3633] = 32'b00000000000000010110111101010111;
assign LUT_3[3634] = 32'b00000000000000010010011001011110;
assign LUT_3[3635] = 32'b00000000000000011001000100111011;
assign LUT_3[3636] = 32'b00000000000000001101011111110000;
assign LUT_3[3637] = 32'b00000000000000010100001011001101;
assign LUT_3[3638] = 32'b00000000000000001111100111010100;
assign LUT_3[3639] = 32'b00000000000000010110010010110001;
assign LUT_3[3640] = 32'b00000000000000010101101011000000;
assign LUT_3[3641] = 32'b00000000000000011100010110011101;
assign LUT_3[3642] = 32'b00000000000000010111110010100100;
assign LUT_3[3643] = 32'b00000000000000011110011110000001;
assign LUT_3[3644] = 32'b00000000000000010010111000110110;
assign LUT_3[3645] = 32'b00000000000000011001100100010011;
assign LUT_3[3646] = 32'b00000000000000010101000000011010;
assign LUT_3[3647] = 32'b00000000000000011011101011110111;
assign LUT_3[3648] = 32'b00000000000000001011101001000010;
assign LUT_3[3649] = 32'b00000000000000010010010100011111;
assign LUT_3[3650] = 32'b00000000000000001101110000100110;
assign LUT_3[3651] = 32'b00000000000000010100011100000011;
assign LUT_3[3652] = 32'b00000000000000001000110110111000;
assign LUT_3[3653] = 32'b00000000000000001111100010010101;
assign LUT_3[3654] = 32'b00000000000000001010111110011100;
assign LUT_3[3655] = 32'b00000000000000010001101001111001;
assign LUT_3[3656] = 32'b00000000000000010001000010001000;
assign LUT_3[3657] = 32'b00000000000000010111101101100101;
assign LUT_3[3658] = 32'b00000000000000010011001001101100;
assign LUT_3[3659] = 32'b00000000000000011001110101001001;
assign LUT_3[3660] = 32'b00000000000000001110001111111110;
assign LUT_3[3661] = 32'b00000000000000010100111011011011;
assign LUT_3[3662] = 32'b00000000000000010000010111100010;
assign LUT_3[3663] = 32'b00000000000000010111000010111111;
assign LUT_3[3664] = 32'b00000000000000001110111100000101;
assign LUT_3[3665] = 32'b00000000000000010101100111100010;
assign LUT_3[3666] = 32'b00000000000000010001000011101001;
assign LUT_3[3667] = 32'b00000000000000010111101111000110;
assign LUT_3[3668] = 32'b00000000000000001100001001111011;
assign LUT_3[3669] = 32'b00000000000000010010110101011000;
assign LUT_3[3670] = 32'b00000000000000001110010001011111;
assign LUT_3[3671] = 32'b00000000000000010100111100111100;
assign LUT_3[3672] = 32'b00000000000000010100010101001011;
assign LUT_3[3673] = 32'b00000000000000011011000000101000;
assign LUT_3[3674] = 32'b00000000000000010110011100101111;
assign LUT_3[3675] = 32'b00000000000000011101001000001100;
assign LUT_3[3676] = 32'b00000000000000010001100011000001;
assign LUT_3[3677] = 32'b00000000000000011000001110011110;
assign LUT_3[3678] = 32'b00000000000000010011101010100101;
assign LUT_3[3679] = 32'b00000000000000011010010110000010;
assign LUT_3[3680] = 32'b00000000000000001100110111100010;
assign LUT_3[3681] = 32'b00000000000000010011100010111111;
assign LUT_3[3682] = 32'b00000000000000001110111111000110;
assign LUT_3[3683] = 32'b00000000000000010101101010100011;
assign LUT_3[3684] = 32'b00000000000000001010000101011000;
assign LUT_3[3685] = 32'b00000000000000010000110000110101;
assign LUT_3[3686] = 32'b00000000000000001100001100111100;
assign LUT_3[3687] = 32'b00000000000000010010111000011001;
assign LUT_3[3688] = 32'b00000000000000010010010000101000;
assign LUT_3[3689] = 32'b00000000000000011000111100000101;
assign LUT_3[3690] = 32'b00000000000000010100011000001100;
assign LUT_3[3691] = 32'b00000000000000011011000011101001;
assign LUT_3[3692] = 32'b00000000000000001111011110011110;
assign LUT_3[3693] = 32'b00000000000000010110001001111011;
assign LUT_3[3694] = 32'b00000000000000010001100110000010;
assign LUT_3[3695] = 32'b00000000000000011000010001011111;
assign LUT_3[3696] = 32'b00000000000000010000001010100101;
assign LUT_3[3697] = 32'b00000000000000010110110110000010;
assign LUT_3[3698] = 32'b00000000000000010010010010001001;
assign LUT_3[3699] = 32'b00000000000000011000111101100110;
assign LUT_3[3700] = 32'b00000000000000001101011000011011;
assign LUT_3[3701] = 32'b00000000000000010100000011111000;
assign LUT_3[3702] = 32'b00000000000000001111011111111111;
assign LUT_3[3703] = 32'b00000000000000010110001011011100;
assign LUT_3[3704] = 32'b00000000000000010101100011101011;
assign LUT_3[3705] = 32'b00000000000000011100001111001000;
assign LUT_3[3706] = 32'b00000000000000010111101011001111;
assign LUT_3[3707] = 32'b00000000000000011110010110101100;
assign LUT_3[3708] = 32'b00000000000000010010110001100001;
assign LUT_3[3709] = 32'b00000000000000011001011100111110;
assign LUT_3[3710] = 32'b00000000000000010100111001000101;
assign LUT_3[3711] = 32'b00000000000000011011100100100010;
assign LUT_3[3712] = 32'b00000000000000001101111011010101;
assign LUT_3[3713] = 32'b00000000000000010100100110110010;
assign LUT_3[3714] = 32'b00000000000000010000000010111001;
assign LUT_3[3715] = 32'b00000000000000010110101110010110;
assign LUT_3[3716] = 32'b00000000000000001011001001001011;
assign LUT_3[3717] = 32'b00000000000000010001110100101000;
assign LUT_3[3718] = 32'b00000000000000001101010000101111;
assign LUT_3[3719] = 32'b00000000000000010011111100001100;
assign LUT_3[3720] = 32'b00000000000000010011010100011011;
assign LUT_3[3721] = 32'b00000000000000011001111111111000;
assign LUT_3[3722] = 32'b00000000000000010101011011111111;
assign LUT_3[3723] = 32'b00000000000000011100000111011100;
assign LUT_3[3724] = 32'b00000000000000010000100010010001;
assign LUT_3[3725] = 32'b00000000000000010111001101101110;
assign LUT_3[3726] = 32'b00000000000000010010101001110101;
assign LUT_3[3727] = 32'b00000000000000011001010101010010;
assign LUT_3[3728] = 32'b00000000000000010001001110011000;
assign LUT_3[3729] = 32'b00000000000000010111111001110101;
assign LUT_3[3730] = 32'b00000000000000010011010101111100;
assign LUT_3[3731] = 32'b00000000000000011010000001011001;
assign LUT_3[3732] = 32'b00000000000000001110011100001110;
assign LUT_3[3733] = 32'b00000000000000010101000111101011;
assign LUT_3[3734] = 32'b00000000000000010000100011110010;
assign LUT_3[3735] = 32'b00000000000000010111001111001111;
assign LUT_3[3736] = 32'b00000000000000010110100111011110;
assign LUT_3[3737] = 32'b00000000000000011101010010111011;
assign LUT_3[3738] = 32'b00000000000000011000101111000010;
assign LUT_3[3739] = 32'b00000000000000011111011010011111;
assign LUT_3[3740] = 32'b00000000000000010011110101010100;
assign LUT_3[3741] = 32'b00000000000000011010100000110001;
assign LUT_3[3742] = 32'b00000000000000010101111100111000;
assign LUT_3[3743] = 32'b00000000000000011100101000010101;
assign LUT_3[3744] = 32'b00000000000000001111001001110101;
assign LUT_3[3745] = 32'b00000000000000010101110101010010;
assign LUT_3[3746] = 32'b00000000000000010001010001011001;
assign LUT_3[3747] = 32'b00000000000000010111111100110110;
assign LUT_3[3748] = 32'b00000000000000001100010111101011;
assign LUT_3[3749] = 32'b00000000000000010011000011001000;
assign LUT_3[3750] = 32'b00000000000000001110011111001111;
assign LUT_3[3751] = 32'b00000000000000010101001010101100;
assign LUT_3[3752] = 32'b00000000000000010100100010111011;
assign LUT_3[3753] = 32'b00000000000000011011001110011000;
assign LUT_3[3754] = 32'b00000000000000010110101010011111;
assign LUT_3[3755] = 32'b00000000000000011101010101111100;
assign LUT_3[3756] = 32'b00000000000000010001110000110001;
assign LUT_3[3757] = 32'b00000000000000011000011100001110;
assign LUT_3[3758] = 32'b00000000000000010011111000010101;
assign LUT_3[3759] = 32'b00000000000000011010100011110010;
assign LUT_3[3760] = 32'b00000000000000010010011100111000;
assign LUT_3[3761] = 32'b00000000000000011001001000010101;
assign LUT_3[3762] = 32'b00000000000000010100100100011100;
assign LUT_3[3763] = 32'b00000000000000011011001111111001;
assign LUT_3[3764] = 32'b00000000000000001111101010101110;
assign LUT_3[3765] = 32'b00000000000000010110010110001011;
assign LUT_3[3766] = 32'b00000000000000010001110010010010;
assign LUT_3[3767] = 32'b00000000000000011000011101101111;
assign LUT_3[3768] = 32'b00000000000000010111110101111110;
assign LUT_3[3769] = 32'b00000000000000011110100001011011;
assign LUT_3[3770] = 32'b00000000000000011001111101100010;
assign LUT_3[3771] = 32'b00000000000000100000101000111111;
assign LUT_3[3772] = 32'b00000000000000010101000011110100;
assign LUT_3[3773] = 32'b00000000000000011011101111010001;
assign LUT_3[3774] = 32'b00000000000000010111001011011000;
assign LUT_3[3775] = 32'b00000000000000011101110110110101;
assign LUT_3[3776] = 32'b00000000000000001101110100000000;
assign LUT_3[3777] = 32'b00000000000000010100011111011101;
assign LUT_3[3778] = 32'b00000000000000001111111011100100;
assign LUT_3[3779] = 32'b00000000000000010110100111000001;
assign LUT_3[3780] = 32'b00000000000000001011000001110110;
assign LUT_3[3781] = 32'b00000000000000010001101101010011;
assign LUT_3[3782] = 32'b00000000000000001101001001011010;
assign LUT_3[3783] = 32'b00000000000000010011110100110111;
assign LUT_3[3784] = 32'b00000000000000010011001101000110;
assign LUT_3[3785] = 32'b00000000000000011001111000100011;
assign LUT_3[3786] = 32'b00000000000000010101010100101010;
assign LUT_3[3787] = 32'b00000000000000011100000000000111;
assign LUT_3[3788] = 32'b00000000000000010000011010111100;
assign LUT_3[3789] = 32'b00000000000000010111000110011001;
assign LUT_3[3790] = 32'b00000000000000010010100010100000;
assign LUT_3[3791] = 32'b00000000000000011001001101111101;
assign LUT_3[3792] = 32'b00000000000000010001000111000011;
assign LUT_3[3793] = 32'b00000000000000010111110010100000;
assign LUT_3[3794] = 32'b00000000000000010011001110100111;
assign LUT_3[3795] = 32'b00000000000000011001111010000100;
assign LUT_3[3796] = 32'b00000000000000001110010100111001;
assign LUT_3[3797] = 32'b00000000000000010101000000010110;
assign LUT_3[3798] = 32'b00000000000000010000011100011101;
assign LUT_3[3799] = 32'b00000000000000010111000111111010;
assign LUT_3[3800] = 32'b00000000000000010110100000001001;
assign LUT_3[3801] = 32'b00000000000000011101001011100110;
assign LUT_3[3802] = 32'b00000000000000011000100111101101;
assign LUT_3[3803] = 32'b00000000000000011111010011001010;
assign LUT_3[3804] = 32'b00000000000000010011101101111111;
assign LUT_3[3805] = 32'b00000000000000011010011001011100;
assign LUT_3[3806] = 32'b00000000000000010101110101100011;
assign LUT_3[3807] = 32'b00000000000000011100100001000000;
assign LUT_3[3808] = 32'b00000000000000001111000010100000;
assign LUT_3[3809] = 32'b00000000000000010101101101111101;
assign LUT_3[3810] = 32'b00000000000000010001001010000100;
assign LUT_3[3811] = 32'b00000000000000010111110101100001;
assign LUT_3[3812] = 32'b00000000000000001100010000010110;
assign LUT_3[3813] = 32'b00000000000000010010111011110011;
assign LUT_3[3814] = 32'b00000000000000001110010111111010;
assign LUT_3[3815] = 32'b00000000000000010101000011010111;
assign LUT_3[3816] = 32'b00000000000000010100011011100110;
assign LUT_3[3817] = 32'b00000000000000011011000111000011;
assign LUT_3[3818] = 32'b00000000000000010110100011001010;
assign LUT_3[3819] = 32'b00000000000000011101001110100111;
assign LUT_3[3820] = 32'b00000000000000010001101001011100;
assign LUT_3[3821] = 32'b00000000000000011000010100111001;
assign LUT_3[3822] = 32'b00000000000000010011110001000000;
assign LUT_3[3823] = 32'b00000000000000011010011100011101;
assign LUT_3[3824] = 32'b00000000000000010010010101100011;
assign LUT_3[3825] = 32'b00000000000000011001000001000000;
assign LUT_3[3826] = 32'b00000000000000010100011101000111;
assign LUT_3[3827] = 32'b00000000000000011011001000100100;
assign LUT_3[3828] = 32'b00000000000000001111100011011001;
assign LUT_3[3829] = 32'b00000000000000010110001110110110;
assign LUT_3[3830] = 32'b00000000000000010001101010111101;
assign LUT_3[3831] = 32'b00000000000000011000010110011010;
assign LUT_3[3832] = 32'b00000000000000010111101110101001;
assign LUT_3[3833] = 32'b00000000000000011110011010000110;
assign LUT_3[3834] = 32'b00000000000000011001110110001101;
assign LUT_3[3835] = 32'b00000000000000100000100001101010;
assign LUT_3[3836] = 32'b00000000000000010100111100011111;
assign LUT_3[3837] = 32'b00000000000000011011100111111100;
assign LUT_3[3838] = 32'b00000000000000010111000100000011;
assign LUT_3[3839] = 32'b00000000000000011101101111100000;
assign LUT_3[3840] = 32'b00000000000000000111111111111000;
assign LUT_3[3841] = 32'b00000000000000001110101011010101;
assign LUT_3[3842] = 32'b00000000000000001010000111011100;
assign LUT_3[3843] = 32'b00000000000000010000110010111001;
assign LUT_3[3844] = 32'b00000000000000000101001101101110;
assign LUT_3[3845] = 32'b00000000000000001011111001001011;
assign LUT_3[3846] = 32'b00000000000000000111010101010010;
assign LUT_3[3847] = 32'b00000000000000001110000000101111;
assign LUT_3[3848] = 32'b00000000000000001101011000111110;
assign LUT_3[3849] = 32'b00000000000000010100000100011011;
assign LUT_3[3850] = 32'b00000000000000001111100000100010;
assign LUT_3[3851] = 32'b00000000000000010110001011111111;
assign LUT_3[3852] = 32'b00000000000000001010100110110100;
assign LUT_3[3853] = 32'b00000000000000010001010010010001;
assign LUT_3[3854] = 32'b00000000000000001100101110011000;
assign LUT_3[3855] = 32'b00000000000000010011011001110101;
assign LUT_3[3856] = 32'b00000000000000001011010010111011;
assign LUT_3[3857] = 32'b00000000000000010001111110011000;
assign LUT_3[3858] = 32'b00000000000000001101011010011111;
assign LUT_3[3859] = 32'b00000000000000010100000101111100;
assign LUT_3[3860] = 32'b00000000000000001000100000110001;
assign LUT_3[3861] = 32'b00000000000000001111001100001110;
assign LUT_3[3862] = 32'b00000000000000001010101000010101;
assign LUT_3[3863] = 32'b00000000000000010001010011110010;
assign LUT_3[3864] = 32'b00000000000000010000101100000001;
assign LUT_3[3865] = 32'b00000000000000010111010111011110;
assign LUT_3[3866] = 32'b00000000000000010010110011100101;
assign LUT_3[3867] = 32'b00000000000000011001011111000010;
assign LUT_3[3868] = 32'b00000000000000001101111001110111;
assign LUT_3[3869] = 32'b00000000000000010100100101010100;
assign LUT_3[3870] = 32'b00000000000000010000000001011011;
assign LUT_3[3871] = 32'b00000000000000010110101100111000;
assign LUT_3[3872] = 32'b00000000000000001001001110011000;
assign LUT_3[3873] = 32'b00000000000000001111111001110101;
assign LUT_3[3874] = 32'b00000000000000001011010101111100;
assign LUT_3[3875] = 32'b00000000000000010010000001011001;
assign LUT_3[3876] = 32'b00000000000000000110011100001110;
assign LUT_3[3877] = 32'b00000000000000001101000111101011;
assign LUT_3[3878] = 32'b00000000000000001000100011110010;
assign LUT_3[3879] = 32'b00000000000000001111001111001111;
assign LUT_3[3880] = 32'b00000000000000001110100111011110;
assign LUT_3[3881] = 32'b00000000000000010101010010111011;
assign LUT_3[3882] = 32'b00000000000000010000101111000010;
assign LUT_3[3883] = 32'b00000000000000010111011010011111;
assign LUT_3[3884] = 32'b00000000000000001011110101010100;
assign LUT_3[3885] = 32'b00000000000000010010100000110001;
assign LUT_3[3886] = 32'b00000000000000001101111100111000;
assign LUT_3[3887] = 32'b00000000000000010100101000010101;
assign LUT_3[3888] = 32'b00000000000000001100100001011011;
assign LUT_3[3889] = 32'b00000000000000010011001100111000;
assign LUT_3[3890] = 32'b00000000000000001110101000111111;
assign LUT_3[3891] = 32'b00000000000000010101010100011100;
assign LUT_3[3892] = 32'b00000000000000001001101111010001;
assign LUT_3[3893] = 32'b00000000000000010000011010101110;
assign LUT_3[3894] = 32'b00000000000000001011110110110101;
assign LUT_3[3895] = 32'b00000000000000010010100010010010;
assign LUT_3[3896] = 32'b00000000000000010001111010100001;
assign LUT_3[3897] = 32'b00000000000000011000100101111110;
assign LUT_3[3898] = 32'b00000000000000010100000010000101;
assign LUT_3[3899] = 32'b00000000000000011010101101100010;
assign LUT_3[3900] = 32'b00000000000000001111001000010111;
assign LUT_3[3901] = 32'b00000000000000010101110011110100;
assign LUT_3[3902] = 32'b00000000000000010001001111111011;
assign LUT_3[3903] = 32'b00000000000000010111111011011000;
assign LUT_3[3904] = 32'b00000000000000000111111000100011;
assign LUT_3[3905] = 32'b00000000000000001110100100000000;
assign LUT_3[3906] = 32'b00000000000000001010000000000111;
assign LUT_3[3907] = 32'b00000000000000010000101011100100;
assign LUT_3[3908] = 32'b00000000000000000101000110011001;
assign LUT_3[3909] = 32'b00000000000000001011110001110110;
assign LUT_3[3910] = 32'b00000000000000000111001101111101;
assign LUT_3[3911] = 32'b00000000000000001101111001011010;
assign LUT_3[3912] = 32'b00000000000000001101010001101001;
assign LUT_3[3913] = 32'b00000000000000010011111101000110;
assign LUT_3[3914] = 32'b00000000000000001111011001001101;
assign LUT_3[3915] = 32'b00000000000000010110000100101010;
assign LUT_3[3916] = 32'b00000000000000001010011111011111;
assign LUT_3[3917] = 32'b00000000000000010001001010111100;
assign LUT_3[3918] = 32'b00000000000000001100100111000011;
assign LUT_3[3919] = 32'b00000000000000010011010010100000;
assign LUT_3[3920] = 32'b00000000000000001011001011100110;
assign LUT_3[3921] = 32'b00000000000000010001110111000011;
assign LUT_3[3922] = 32'b00000000000000001101010011001010;
assign LUT_3[3923] = 32'b00000000000000010011111110100111;
assign LUT_3[3924] = 32'b00000000000000001000011001011100;
assign LUT_3[3925] = 32'b00000000000000001111000100111001;
assign LUT_3[3926] = 32'b00000000000000001010100001000000;
assign LUT_3[3927] = 32'b00000000000000010001001100011101;
assign LUT_3[3928] = 32'b00000000000000010000100100101100;
assign LUT_3[3929] = 32'b00000000000000010111010000001001;
assign LUT_3[3930] = 32'b00000000000000010010101100010000;
assign LUT_3[3931] = 32'b00000000000000011001010111101101;
assign LUT_3[3932] = 32'b00000000000000001101110010100010;
assign LUT_3[3933] = 32'b00000000000000010100011101111111;
assign LUT_3[3934] = 32'b00000000000000001111111010000110;
assign LUT_3[3935] = 32'b00000000000000010110100101100011;
assign LUT_3[3936] = 32'b00000000000000001001000111000011;
assign LUT_3[3937] = 32'b00000000000000001111110010100000;
assign LUT_3[3938] = 32'b00000000000000001011001110100111;
assign LUT_3[3939] = 32'b00000000000000010001111010000100;
assign LUT_3[3940] = 32'b00000000000000000110010100111001;
assign LUT_3[3941] = 32'b00000000000000001101000000010110;
assign LUT_3[3942] = 32'b00000000000000001000011100011101;
assign LUT_3[3943] = 32'b00000000000000001111000111111010;
assign LUT_3[3944] = 32'b00000000000000001110100000001001;
assign LUT_3[3945] = 32'b00000000000000010101001011100110;
assign LUT_3[3946] = 32'b00000000000000010000100111101101;
assign LUT_3[3947] = 32'b00000000000000010111010011001010;
assign LUT_3[3948] = 32'b00000000000000001011101101111111;
assign LUT_3[3949] = 32'b00000000000000010010011001011100;
assign LUT_3[3950] = 32'b00000000000000001101110101100011;
assign LUT_3[3951] = 32'b00000000000000010100100001000000;
assign LUT_3[3952] = 32'b00000000000000001100011010000110;
assign LUT_3[3953] = 32'b00000000000000010011000101100011;
assign LUT_3[3954] = 32'b00000000000000001110100001101010;
assign LUT_3[3955] = 32'b00000000000000010101001101000111;
assign LUT_3[3956] = 32'b00000000000000001001100111111100;
assign LUT_3[3957] = 32'b00000000000000010000010011011001;
assign LUT_3[3958] = 32'b00000000000000001011101111100000;
assign LUT_3[3959] = 32'b00000000000000010010011010111101;
assign LUT_3[3960] = 32'b00000000000000010001110011001100;
assign LUT_3[3961] = 32'b00000000000000011000011110101001;
assign LUT_3[3962] = 32'b00000000000000010011111010110000;
assign LUT_3[3963] = 32'b00000000000000011010100110001101;
assign LUT_3[3964] = 32'b00000000000000001111000001000010;
assign LUT_3[3965] = 32'b00000000000000010101101100011111;
assign LUT_3[3966] = 32'b00000000000000010001001000100110;
assign LUT_3[3967] = 32'b00000000000000010111110100000011;
assign LUT_3[3968] = 32'b00000000000000001010001010110110;
assign LUT_3[3969] = 32'b00000000000000010000110110010011;
assign LUT_3[3970] = 32'b00000000000000001100010010011010;
assign LUT_3[3971] = 32'b00000000000000010010111101110111;
assign LUT_3[3972] = 32'b00000000000000000111011000101100;
assign LUT_3[3973] = 32'b00000000000000001110000100001001;
assign LUT_3[3974] = 32'b00000000000000001001100000010000;
assign LUT_3[3975] = 32'b00000000000000010000001011101101;
assign LUT_3[3976] = 32'b00000000000000001111100011111100;
assign LUT_3[3977] = 32'b00000000000000010110001111011001;
assign LUT_3[3978] = 32'b00000000000000010001101011100000;
assign LUT_3[3979] = 32'b00000000000000011000010110111101;
assign LUT_3[3980] = 32'b00000000000000001100110001110010;
assign LUT_3[3981] = 32'b00000000000000010011011101001111;
assign LUT_3[3982] = 32'b00000000000000001110111001010110;
assign LUT_3[3983] = 32'b00000000000000010101100100110011;
assign LUT_3[3984] = 32'b00000000000000001101011101111001;
assign LUT_3[3985] = 32'b00000000000000010100001001010110;
assign LUT_3[3986] = 32'b00000000000000001111100101011101;
assign LUT_3[3987] = 32'b00000000000000010110010000111010;
assign LUT_3[3988] = 32'b00000000000000001010101011101111;
assign LUT_3[3989] = 32'b00000000000000010001010111001100;
assign LUT_3[3990] = 32'b00000000000000001100110011010011;
assign LUT_3[3991] = 32'b00000000000000010011011110110000;
assign LUT_3[3992] = 32'b00000000000000010010110110111111;
assign LUT_3[3993] = 32'b00000000000000011001100010011100;
assign LUT_3[3994] = 32'b00000000000000010100111110100011;
assign LUT_3[3995] = 32'b00000000000000011011101010000000;
assign LUT_3[3996] = 32'b00000000000000010000000100110101;
assign LUT_3[3997] = 32'b00000000000000010110110000010010;
assign LUT_3[3998] = 32'b00000000000000010010001100011001;
assign LUT_3[3999] = 32'b00000000000000011000110111110110;
assign LUT_3[4000] = 32'b00000000000000001011011001010110;
assign LUT_3[4001] = 32'b00000000000000010010000100110011;
assign LUT_3[4002] = 32'b00000000000000001101100000111010;
assign LUT_3[4003] = 32'b00000000000000010100001100010111;
assign LUT_3[4004] = 32'b00000000000000001000100111001100;
assign LUT_3[4005] = 32'b00000000000000001111010010101001;
assign LUT_3[4006] = 32'b00000000000000001010101110110000;
assign LUT_3[4007] = 32'b00000000000000010001011010001101;
assign LUT_3[4008] = 32'b00000000000000010000110010011100;
assign LUT_3[4009] = 32'b00000000000000010111011101111001;
assign LUT_3[4010] = 32'b00000000000000010010111010000000;
assign LUT_3[4011] = 32'b00000000000000011001100101011101;
assign LUT_3[4012] = 32'b00000000000000001110000000010010;
assign LUT_3[4013] = 32'b00000000000000010100101011101111;
assign LUT_3[4014] = 32'b00000000000000010000000111110110;
assign LUT_3[4015] = 32'b00000000000000010110110011010011;
assign LUT_3[4016] = 32'b00000000000000001110101100011001;
assign LUT_3[4017] = 32'b00000000000000010101010111110110;
assign LUT_3[4018] = 32'b00000000000000010000110011111101;
assign LUT_3[4019] = 32'b00000000000000010111011111011010;
assign LUT_3[4020] = 32'b00000000000000001011111010001111;
assign LUT_3[4021] = 32'b00000000000000010010100101101100;
assign LUT_3[4022] = 32'b00000000000000001110000001110011;
assign LUT_3[4023] = 32'b00000000000000010100101101010000;
assign LUT_3[4024] = 32'b00000000000000010100000101011111;
assign LUT_3[4025] = 32'b00000000000000011010110000111100;
assign LUT_3[4026] = 32'b00000000000000010110001101000011;
assign LUT_3[4027] = 32'b00000000000000011100111000100000;
assign LUT_3[4028] = 32'b00000000000000010001010011010101;
assign LUT_3[4029] = 32'b00000000000000010111111110110010;
assign LUT_3[4030] = 32'b00000000000000010011011010111001;
assign LUT_3[4031] = 32'b00000000000000011010000110010110;
assign LUT_3[4032] = 32'b00000000000000001010000011100001;
assign LUT_3[4033] = 32'b00000000000000010000101110111110;
assign LUT_3[4034] = 32'b00000000000000001100001011000101;
assign LUT_3[4035] = 32'b00000000000000010010110110100010;
assign LUT_3[4036] = 32'b00000000000000000111010001010111;
assign LUT_3[4037] = 32'b00000000000000001101111100110100;
assign LUT_3[4038] = 32'b00000000000000001001011000111011;
assign LUT_3[4039] = 32'b00000000000000010000000100011000;
assign LUT_3[4040] = 32'b00000000000000001111011100100111;
assign LUT_3[4041] = 32'b00000000000000010110001000000100;
assign LUT_3[4042] = 32'b00000000000000010001100100001011;
assign LUT_3[4043] = 32'b00000000000000011000001111101000;
assign LUT_3[4044] = 32'b00000000000000001100101010011101;
assign LUT_3[4045] = 32'b00000000000000010011010101111010;
assign LUT_3[4046] = 32'b00000000000000001110110010000001;
assign LUT_3[4047] = 32'b00000000000000010101011101011110;
assign LUT_3[4048] = 32'b00000000000000001101010110100100;
assign LUT_3[4049] = 32'b00000000000000010100000010000001;
assign LUT_3[4050] = 32'b00000000000000001111011110001000;
assign LUT_3[4051] = 32'b00000000000000010110001001100101;
assign LUT_3[4052] = 32'b00000000000000001010100100011010;
assign LUT_3[4053] = 32'b00000000000000010001001111110111;
assign LUT_3[4054] = 32'b00000000000000001100101011111110;
assign LUT_3[4055] = 32'b00000000000000010011010111011011;
assign LUT_3[4056] = 32'b00000000000000010010101111101010;
assign LUT_3[4057] = 32'b00000000000000011001011011000111;
assign LUT_3[4058] = 32'b00000000000000010100110111001110;
assign LUT_3[4059] = 32'b00000000000000011011100010101011;
assign LUT_3[4060] = 32'b00000000000000001111111101100000;
assign LUT_3[4061] = 32'b00000000000000010110101000111101;
assign LUT_3[4062] = 32'b00000000000000010010000101000100;
assign LUT_3[4063] = 32'b00000000000000011000110000100001;
assign LUT_3[4064] = 32'b00000000000000001011010010000001;
assign LUT_3[4065] = 32'b00000000000000010001111101011110;
assign LUT_3[4066] = 32'b00000000000000001101011001100101;
assign LUT_3[4067] = 32'b00000000000000010100000101000010;
assign LUT_3[4068] = 32'b00000000000000001000011111110111;
assign LUT_3[4069] = 32'b00000000000000001111001011010100;
assign LUT_3[4070] = 32'b00000000000000001010100111011011;
assign LUT_3[4071] = 32'b00000000000000010001010010111000;
assign LUT_3[4072] = 32'b00000000000000010000101011000111;
assign LUT_3[4073] = 32'b00000000000000010111010110100100;
assign LUT_3[4074] = 32'b00000000000000010010110010101011;
assign LUT_3[4075] = 32'b00000000000000011001011110001000;
assign LUT_3[4076] = 32'b00000000000000001101111000111101;
assign LUT_3[4077] = 32'b00000000000000010100100100011010;
assign LUT_3[4078] = 32'b00000000000000010000000000100001;
assign LUT_3[4079] = 32'b00000000000000010110101011111110;
assign LUT_3[4080] = 32'b00000000000000001110100101000100;
assign LUT_3[4081] = 32'b00000000000000010101010000100001;
assign LUT_3[4082] = 32'b00000000000000010000101100101000;
assign LUT_3[4083] = 32'b00000000000000010111011000000101;
assign LUT_3[4084] = 32'b00000000000000001011110010111010;
assign LUT_3[4085] = 32'b00000000000000010010011110010111;
assign LUT_3[4086] = 32'b00000000000000001101111010011110;
assign LUT_3[4087] = 32'b00000000000000010100100101111011;
assign LUT_3[4088] = 32'b00000000000000010011111110001010;
assign LUT_3[4089] = 32'b00000000000000011010101001100111;
assign LUT_3[4090] = 32'b00000000000000010110000101101110;
assign LUT_3[4091] = 32'b00000000000000011100110001001011;
assign LUT_3[4092] = 32'b00000000000000010001001100000000;
assign LUT_3[4093] = 32'b00000000000000010111110111011101;
assign LUT_3[4094] = 32'b00000000000000010011010011100100;
assign LUT_3[4095] = 32'b00000000000000011001111111000001;
assign LUT_3[4096] = 32'b00000000000000000100010001011011;
assign LUT_3[4097] = 32'b00000000000000001010111100111000;
assign LUT_3[4098] = 32'b00000000000000000110011000111111;
assign LUT_3[4099] = 32'b00000000000000001101000100011100;
assign LUT_3[4100] = 32'b00000000000000000001011111010001;
assign LUT_3[4101] = 32'b00000000000000001000001010101110;
assign LUT_3[4102] = 32'b00000000000000000011100110110101;
assign LUT_3[4103] = 32'b00000000000000001010010010010010;
assign LUT_3[4104] = 32'b00000000000000001001101010100001;
assign LUT_3[4105] = 32'b00000000000000010000010101111110;
assign LUT_3[4106] = 32'b00000000000000001011110010000101;
assign LUT_3[4107] = 32'b00000000000000010010011101100010;
assign LUT_3[4108] = 32'b00000000000000000110111000010111;
assign LUT_3[4109] = 32'b00000000000000001101100011110100;
assign LUT_3[4110] = 32'b00000000000000001000111111111011;
assign LUT_3[4111] = 32'b00000000000000001111101011011000;
assign LUT_3[4112] = 32'b00000000000000000111100100011110;
assign LUT_3[4113] = 32'b00000000000000001110001111111011;
assign LUT_3[4114] = 32'b00000000000000001001101100000010;
assign LUT_3[4115] = 32'b00000000000000010000010111011111;
assign LUT_3[4116] = 32'b00000000000000000100110010010100;
assign LUT_3[4117] = 32'b00000000000000001011011101110001;
assign LUT_3[4118] = 32'b00000000000000000110111001111000;
assign LUT_3[4119] = 32'b00000000000000001101100101010101;
assign LUT_3[4120] = 32'b00000000000000001100111101100100;
assign LUT_3[4121] = 32'b00000000000000010011101001000001;
assign LUT_3[4122] = 32'b00000000000000001111000101001000;
assign LUT_3[4123] = 32'b00000000000000010101110000100101;
assign LUT_3[4124] = 32'b00000000000000001010001011011010;
assign LUT_3[4125] = 32'b00000000000000010000110110110111;
assign LUT_3[4126] = 32'b00000000000000001100010010111110;
assign LUT_3[4127] = 32'b00000000000000010010111110011011;
assign LUT_3[4128] = 32'b00000000000000000101011111111011;
assign LUT_3[4129] = 32'b00000000000000001100001011011000;
assign LUT_3[4130] = 32'b00000000000000000111100111011111;
assign LUT_3[4131] = 32'b00000000000000001110010010111100;
assign LUT_3[4132] = 32'b00000000000000000010101101110001;
assign LUT_3[4133] = 32'b00000000000000001001011001001110;
assign LUT_3[4134] = 32'b00000000000000000100110101010101;
assign LUT_3[4135] = 32'b00000000000000001011100000110010;
assign LUT_3[4136] = 32'b00000000000000001010111001000001;
assign LUT_3[4137] = 32'b00000000000000010001100100011110;
assign LUT_3[4138] = 32'b00000000000000001101000000100101;
assign LUT_3[4139] = 32'b00000000000000010011101100000010;
assign LUT_3[4140] = 32'b00000000000000001000000110110111;
assign LUT_3[4141] = 32'b00000000000000001110110010010100;
assign LUT_3[4142] = 32'b00000000000000001010001110011011;
assign LUT_3[4143] = 32'b00000000000000010000111001111000;
assign LUT_3[4144] = 32'b00000000000000001000110010111110;
assign LUT_3[4145] = 32'b00000000000000001111011110011011;
assign LUT_3[4146] = 32'b00000000000000001010111010100010;
assign LUT_3[4147] = 32'b00000000000000010001100101111111;
assign LUT_3[4148] = 32'b00000000000000000110000000110100;
assign LUT_3[4149] = 32'b00000000000000001100101100010001;
assign LUT_3[4150] = 32'b00000000000000001000001000011000;
assign LUT_3[4151] = 32'b00000000000000001110110011110101;
assign LUT_3[4152] = 32'b00000000000000001110001100000100;
assign LUT_3[4153] = 32'b00000000000000010100110111100001;
assign LUT_3[4154] = 32'b00000000000000010000010011101000;
assign LUT_3[4155] = 32'b00000000000000010110111111000101;
assign LUT_3[4156] = 32'b00000000000000001011011001111010;
assign LUT_3[4157] = 32'b00000000000000010010000101010111;
assign LUT_3[4158] = 32'b00000000000000001101100001011110;
assign LUT_3[4159] = 32'b00000000000000010100001100111011;
assign LUT_3[4160] = 32'b00000000000000000100001010000110;
assign LUT_3[4161] = 32'b00000000000000001010110101100011;
assign LUT_3[4162] = 32'b00000000000000000110010001101010;
assign LUT_3[4163] = 32'b00000000000000001100111101000111;
assign LUT_3[4164] = 32'b00000000000000000001010111111100;
assign LUT_3[4165] = 32'b00000000000000001000000011011001;
assign LUT_3[4166] = 32'b00000000000000000011011111100000;
assign LUT_3[4167] = 32'b00000000000000001010001010111101;
assign LUT_3[4168] = 32'b00000000000000001001100011001100;
assign LUT_3[4169] = 32'b00000000000000010000001110101001;
assign LUT_3[4170] = 32'b00000000000000001011101010110000;
assign LUT_3[4171] = 32'b00000000000000010010010110001101;
assign LUT_3[4172] = 32'b00000000000000000110110001000010;
assign LUT_3[4173] = 32'b00000000000000001101011100011111;
assign LUT_3[4174] = 32'b00000000000000001000111000100110;
assign LUT_3[4175] = 32'b00000000000000001111100100000011;
assign LUT_3[4176] = 32'b00000000000000000111011101001001;
assign LUT_3[4177] = 32'b00000000000000001110001000100110;
assign LUT_3[4178] = 32'b00000000000000001001100100101101;
assign LUT_3[4179] = 32'b00000000000000010000010000001010;
assign LUT_3[4180] = 32'b00000000000000000100101010111111;
assign LUT_3[4181] = 32'b00000000000000001011010110011100;
assign LUT_3[4182] = 32'b00000000000000000110110010100011;
assign LUT_3[4183] = 32'b00000000000000001101011110000000;
assign LUT_3[4184] = 32'b00000000000000001100110110001111;
assign LUT_3[4185] = 32'b00000000000000010011100001101100;
assign LUT_3[4186] = 32'b00000000000000001110111101110011;
assign LUT_3[4187] = 32'b00000000000000010101101001010000;
assign LUT_3[4188] = 32'b00000000000000001010000100000101;
assign LUT_3[4189] = 32'b00000000000000010000101111100010;
assign LUT_3[4190] = 32'b00000000000000001100001011101001;
assign LUT_3[4191] = 32'b00000000000000010010110111000110;
assign LUT_3[4192] = 32'b00000000000000000101011000100110;
assign LUT_3[4193] = 32'b00000000000000001100000100000011;
assign LUT_3[4194] = 32'b00000000000000000111100000001010;
assign LUT_3[4195] = 32'b00000000000000001110001011100111;
assign LUT_3[4196] = 32'b00000000000000000010100110011100;
assign LUT_3[4197] = 32'b00000000000000001001010001111001;
assign LUT_3[4198] = 32'b00000000000000000100101110000000;
assign LUT_3[4199] = 32'b00000000000000001011011001011101;
assign LUT_3[4200] = 32'b00000000000000001010110001101100;
assign LUT_3[4201] = 32'b00000000000000010001011101001001;
assign LUT_3[4202] = 32'b00000000000000001100111001010000;
assign LUT_3[4203] = 32'b00000000000000010011100100101101;
assign LUT_3[4204] = 32'b00000000000000000111111111100010;
assign LUT_3[4205] = 32'b00000000000000001110101010111111;
assign LUT_3[4206] = 32'b00000000000000001010000111000110;
assign LUT_3[4207] = 32'b00000000000000010000110010100011;
assign LUT_3[4208] = 32'b00000000000000001000101011101001;
assign LUT_3[4209] = 32'b00000000000000001111010111000110;
assign LUT_3[4210] = 32'b00000000000000001010110011001101;
assign LUT_3[4211] = 32'b00000000000000010001011110101010;
assign LUT_3[4212] = 32'b00000000000000000101111001011111;
assign LUT_3[4213] = 32'b00000000000000001100100100111100;
assign LUT_3[4214] = 32'b00000000000000001000000001000011;
assign LUT_3[4215] = 32'b00000000000000001110101100100000;
assign LUT_3[4216] = 32'b00000000000000001110000100101111;
assign LUT_3[4217] = 32'b00000000000000010100110000001100;
assign LUT_3[4218] = 32'b00000000000000010000001100010011;
assign LUT_3[4219] = 32'b00000000000000010110110111110000;
assign LUT_3[4220] = 32'b00000000000000001011010010100101;
assign LUT_3[4221] = 32'b00000000000000010001111110000010;
assign LUT_3[4222] = 32'b00000000000000001101011010001001;
assign LUT_3[4223] = 32'b00000000000000010100000101100110;
assign LUT_3[4224] = 32'b00000000000000000110011100011001;
assign LUT_3[4225] = 32'b00000000000000001101000111110110;
assign LUT_3[4226] = 32'b00000000000000001000100011111101;
assign LUT_3[4227] = 32'b00000000000000001111001111011010;
assign LUT_3[4228] = 32'b00000000000000000011101010001111;
assign LUT_3[4229] = 32'b00000000000000001010010101101100;
assign LUT_3[4230] = 32'b00000000000000000101110001110011;
assign LUT_3[4231] = 32'b00000000000000001100011101010000;
assign LUT_3[4232] = 32'b00000000000000001011110101011111;
assign LUT_3[4233] = 32'b00000000000000010010100000111100;
assign LUT_3[4234] = 32'b00000000000000001101111101000011;
assign LUT_3[4235] = 32'b00000000000000010100101000100000;
assign LUT_3[4236] = 32'b00000000000000001001000011010101;
assign LUT_3[4237] = 32'b00000000000000001111101110110010;
assign LUT_3[4238] = 32'b00000000000000001011001010111001;
assign LUT_3[4239] = 32'b00000000000000010001110110010110;
assign LUT_3[4240] = 32'b00000000000000001001101111011100;
assign LUT_3[4241] = 32'b00000000000000010000011010111001;
assign LUT_3[4242] = 32'b00000000000000001011110111000000;
assign LUT_3[4243] = 32'b00000000000000010010100010011101;
assign LUT_3[4244] = 32'b00000000000000000110111101010010;
assign LUT_3[4245] = 32'b00000000000000001101101000101111;
assign LUT_3[4246] = 32'b00000000000000001001000100110110;
assign LUT_3[4247] = 32'b00000000000000001111110000010011;
assign LUT_3[4248] = 32'b00000000000000001111001000100010;
assign LUT_3[4249] = 32'b00000000000000010101110011111111;
assign LUT_3[4250] = 32'b00000000000000010001010000000110;
assign LUT_3[4251] = 32'b00000000000000010111111011100011;
assign LUT_3[4252] = 32'b00000000000000001100010110011000;
assign LUT_3[4253] = 32'b00000000000000010011000001110101;
assign LUT_3[4254] = 32'b00000000000000001110011101111100;
assign LUT_3[4255] = 32'b00000000000000010101001001011001;
assign LUT_3[4256] = 32'b00000000000000000111101010111001;
assign LUT_3[4257] = 32'b00000000000000001110010110010110;
assign LUT_3[4258] = 32'b00000000000000001001110010011101;
assign LUT_3[4259] = 32'b00000000000000010000011101111010;
assign LUT_3[4260] = 32'b00000000000000000100111000101111;
assign LUT_3[4261] = 32'b00000000000000001011100100001100;
assign LUT_3[4262] = 32'b00000000000000000111000000010011;
assign LUT_3[4263] = 32'b00000000000000001101101011110000;
assign LUT_3[4264] = 32'b00000000000000001101000011111111;
assign LUT_3[4265] = 32'b00000000000000010011101111011100;
assign LUT_3[4266] = 32'b00000000000000001111001011100011;
assign LUT_3[4267] = 32'b00000000000000010101110111000000;
assign LUT_3[4268] = 32'b00000000000000001010010001110101;
assign LUT_3[4269] = 32'b00000000000000010000111101010010;
assign LUT_3[4270] = 32'b00000000000000001100011001011001;
assign LUT_3[4271] = 32'b00000000000000010011000100110110;
assign LUT_3[4272] = 32'b00000000000000001010111101111100;
assign LUT_3[4273] = 32'b00000000000000010001101001011001;
assign LUT_3[4274] = 32'b00000000000000001101000101100000;
assign LUT_3[4275] = 32'b00000000000000010011110000111101;
assign LUT_3[4276] = 32'b00000000000000001000001011110010;
assign LUT_3[4277] = 32'b00000000000000001110110111001111;
assign LUT_3[4278] = 32'b00000000000000001010010011010110;
assign LUT_3[4279] = 32'b00000000000000010000111110110011;
assign LUT_3[4280] = 32'b00000000000000010000010111000010;
assign LUT_3[4281] = 32'b00000000000000010111000010011111;
assign LUT_3[4282] = 32'b00000000000000010010011110100110;
assign LUT_3[4283] = 32'b00000000000000011001001010000011;
assign LUT_3[4284] = 32'b00000000000000001101100100111000;
assign LUT_3[4285] = 32'b00000000000000010100010000010101;
assign LUT_3[4286] = 32'b00000000000000001111101100011100;
assign LUT_3[4287] = 32'b00000000000000010110010111111001;
assign LUT_3[4288] = 32'b00000000000000000110010101000100;
assign LUT_3[4289] = 32'b00000000000000001101000000100001;
assign LUT_3[4290] = 32'b00000000000000001000011100101000;
assign LUT_3[4291] = 32'b00000000000000001111001000000101;
assign LUT_3[4292] = 32'b00000000000000000011100010111010;
assign LUT_3[4293] = 32'b00000000000000001010001110010111;
assign LUT_3[4294] = 32'b00000000000000000101101010011110;
assign LUT_3[4295] = 32'b00000000000000001100010101111011;
assign LUT_3[4296] = 32'b00000000000000001011101110001010;
assign LUT_3[4297] = 32'b00000000000000010010011001100111;
assign LUT_3[4298] = 32'b00000000000000001101110101101110;
assign LUT_3[4299] = 32'b00000000000000010100100001001011;
assign LUT_3[4300] = 32'b00000000000000001000111100000000;
assign LUT_3[4301] = 32'b00000000000000001111100111011101;
assign LUT_3[4302] = 32'b00000000000000001011000011100100;
assign LUT_3[4303] = 32'b00000000000000010001101111000001;
assign LUT_3[4304] = 32'b00000000000000001001101000000111;
assign LUT_3[4305] = 32'b00000000000000010000010011100100;
assign LUT_3[4306] = 32'b00000000000000001011101111101011;
assign LUT_3[4307] = 32'b00000000000000010010011011001000;
assign LUT_3[4308] = 32'b00000000000000000110110101111101;
assign LUT_3[4309] = 32'b00000000000000001101100001011010;
assign LUT_3[4310] = 32'b00000000000000001000111101100001;
assign LUT_3[4311] = 32'b00000000000000001111101000111110;
assign LUT_3[4312] = 32'b00000000000000001111000001001101;
assign LUT_3[4313] = 32'b00000000000000010101101100101010;
assign LUT_3[4314] = 32'b00000000000000010001001000110001;
assign LUT_3[4315] = 32'b00000000000000010111110100001110;
assign LUT_3[4316] = 32'b00000000000000001100001111000011;
assign LUT_3[4317] = 32'b00000000000000010010111010100000;
assign LUT_3[4318] = 32'b00000000000000001110010110100111;
assign LUT_3[4319] = 32'b00000000000000010101000010000100;
assign LUT_3[4320] = 32'b00000000000000000111100011100100;
assign LUT_3[4321] = 32'b00000000000000001110001111000001;
assign LUT_3[4322] = 32'b00000000000000001001101011001000;
assign LUT_3[4323] = 32'b00000000000000010000010110100101;
assign LUT_3[4324] = 32'b00000000000000000100110001011010;
assign LUT_3[4325] = 32'b00000000000000001011011100110111;
assign LUT_3[4326] = 32'b00000000000000000110111000111110;
assign LUT_3[4327] = 32'b00000000000000001101100100011011;
assign LUT_3[4328] = 32'b00000000000000001100111100101010;
assign LUT_3[4329] = 32'b00000000000000010011101000000111;
assign LUT_3[4330] = 32'b00000000000000001111000100001110;
assign LUT_3[4331] = 32'b00000000000000010101101111101011;
assign LUT_3[4332] = 32'b00000000000000001010001010100000;
assign LUT_3[4333] = 32'b00000000000000010000110101111101;
assign LUT_3[4334] = 32'b00000000000000001100010010000100;
assign LUT_3[4335] = 32'b00000000000000010010111101100001;
assign LUT_3[4336] = 32'b00000000000000001010110110100111;
assign LUT_3[4337] = 32'b00000000000000010001100010000100;
assign LUT_3[4338] = 32'b00000000000000001100111110001011;
assign LUT_3[4339] = 32'b00000000000000010011101001101000;
assign LUT_3[4340] = 32'b00000000000000001000000100011101;
assign LUT_3[4341] = 32'b00000000000000001110101111111010;
assign LUT_3[4342] = 32'b00000000000000001010001100000001;
assign LUT_3[4343] = 32'b00000000000000010000110111011110;
assign LUT_3[4344] = 32'b00000000000000010000001111101101;
assign LUT_3[4345] = 32'b00000000000000010110111011001010;
assign LUT_3[4346] = 32'b00000000000000010010010111010001;
assign LUT_3[4347] = 32'b00000000000000011001000010101110;
assign LUT_3[4348] = 32'b00000000000000001101011101100011;
assign LUT_3[4349] = 32'b00000000000000010100001001000000;
assign LUT_3[4350] = 32'b00000000000000001111100101000111;
assign LUT_3[4351] = 32'b00000000000000010110010000100100;
assign LUT_3[4352] = 32'b00000000000000000000100000111100;
assign LUT_3[4353] = 32'b00000000000000000111001100011001;
assign LUT_3[4354] = 32'b00000000000000000010101000100000;
assign LUT_3[4355] = 32'b00000000000000001001010011111101;
assign LUT_3[4356] = 32'b11111111111111111101101110110010;
assign LUT_3[4357] = 32'b00000000000000000100011010001111;
assign LUT_3[4358] = 32'b11111111111111111111110110010110;
assign LUT_3[4359] = 32'b00000000000000000110100001110011;
assign LUT_3[4360] = 32'b00000000000000000101111010000010;
assign LUT_3[4361] = 32'b00000000000000001100100101011111;
assign LUT_3[4362] = 32'b00000000000000001000000001100110;
assign LUT_3[4363] = 32'b00000000000000001110101101000011;
assign LUT_3[4364] = 32'b00000000000000000011000111111000;
assign LUT_3[4365] = 32'b00000000000000001001110011010101;
assign LUT_3[4366] = 32'b00000000000000000101001111011100;
assign LUT_3[4367] = 32'b00000000000000001011111010111001;
assign LUT_3[4368] = 32'b00000000000000000011110011111111;
assign LUT_3[4369] = 32'b00000000000000001010011111011100;
assign LUT_3[4370] = 32'b00000000000000000101111011100011;
assign LUT_3[4371] = 32'b00000000000000001100100111000000;
assign LUT_3[4372] = 32'b00000000000000000001000001110101;
assign LUT_3[4373] = 32'b00000000000000000111101101010010;
assign LUT_3[4374] = 32'b00000000000000000011001001011001;
assign LUT_3[4375] = 32'b00000000000000001001110100110110;
assign LUT_3[4376] = 32'b00000000000000001001001101000101;
assign LUT_3[4377] = 32'b00000000000000001111111000100010;
assign LUT_3[4378] = 32'b00000000000000001011010100101001;
assign LUT_3[4379] = 32'b00000000000000010010000000000110;
assign LUT_3[4380] = 32'b00000000000000000110011010111011;
assign LUT_3[4381] = 32'b00000000000000001101000110011000;
assign LUT_3[4382] = 32'b00000000000000001000100010011111;
assign LUT_3[4383] = 32'b00000000000000001111001101111100;
assign LUT_3[4384] = 32'b00000000000000000001101111011100;
assign LUT_3[4385] = 32'b00000000000000001000011010111001;
assign LUT_3[4386] = 32'b00000000000000000011110111000000;
assign LUT_3[4387] = 32'b00000000000000001010100010011101;
assign LUT_3[4388] = 32'b11111111111111111110111101010010;
assign LUT_3[4389] = 32'b00000000000000000101101000101111;
assign LUT_3[4390] = 32'b00000000000000000001000100110110;
assign LUT_3[4391] = 32'b00000000000000000111110000010011;
assign LUT_3[4392] = 32'b00000000000000000111001000100010;
assign LUT_3[4393] = 32'b00000000000000001101110011111111;
assign LUT_3[4394] = 32'b00000000000000001001010000000110;
assign LUT_3[4395] = 32'b00000000000000001111111011100011;
assign LUT_3[4396] = 32'b00000000000000000100010110011000;
assign LUT_3[4397] = 32'b00000000000000001011000001110101;
assign LUT_3[4398] = 32'b00000000000000000110011101111100;
assign LUT_3[4399] = 32'b00000000000000001101001001011001;
assign LUT_3[4400] = 32'b00000000000000000101000010011111;
assign LUT_3[4401] = 32'b00000000000000001011101101111100;
assign LUT_3[4402] = 32'b00000000000000000111001010000011;
assign LUT_3[4403] = 32'b00000000000000001101110101100000;
assign LUT_3[4404] = 32'b00000000000000000010010000010101;
assign LUT_3[4405] = 32'b00000000000000001000111011110010;
assign LUT_3[4406] = 32'b00000000000000000100010111111001;
assign LUT_3[4407] = 32'b00000000000000001011000011010110;
assign LUT_3[4408] = 32'b00000000000000001010011011100101;
assign LUT_3[4409] = 32'b00000000000000010001000111000010;
assign LUT_3[4410] = 32'b00000000000000001100100011001001;
assign LUT_3[4411] = 32'b00000000000000010011001110100110;
assign LUT_3[4412] = 32'b00000000000000000111101001011011;
assign LUT_3[4413] = 32'b00000000000000001110010100111000;
assign LUT_3[4414] = 32'b00000000000000001001110000111111;
assign LUT_3[4415] = 32'b00000000000000010000011100011100;
assign LUT_3[4416] = 32'b00000000000000000000011001100111;
assign LUT_3[4417] = 32'b00000000000000000111000101000100;
assign LUT_3[4418] = 32'b00000000000000000010100001001011;
assign LUT_3[4419] = 32'b00000000000000001001001100101000;
assign LUT_3[4420] = 32'b11111111111111111101100111011101;
assign LUT_3[4421] = 32'b00000000000000000100010010111010;
assign LUT_3[4422] = 32'b11111111111111111111101111000001;
assign LUT_3[4423] = 32'b00000000000000000110011010011110;
assign LUT_3[4424] = 32'b00000000000000000101110010101101;
assign LUT_3[4425] = 32'b00000000000000001100011110001010;
assign LUT_3[4426] = 32'b00000000000000000111111010010001;
assign LUT_3[4427] = 32'b00000000000000001110100101101110;
assign LUT_3[4428] = 32'b00000000000000000011000000100011;
assign LUT_3[4429] = 32'b00000000000000001001101100000000;
assign LUT_3[4430] = 32'b00000000000000000101001000000111;
assign LUT_3[4431] = 32'b00000000000000001011110011100100;
assign LUT_3[4432] = 32'b00000000000000000011101100101010;
assign LUT_3[4433] = 32'b00000000000000001010011000000111;
assign LUT_3[4434] = 32'b00000000000000000101110100001110;
assign LUT_3[4435] = 32'b00000000000000001100011111101011;
assign LUT_3[4436] = 32'b00000000000000000000111010100000;
assign LUT_3[4437] = 32'b00000000000000000111100101111101;
assign LUT_3[4438] = 32'b00000000000000000011000010000100;
assign LUT_3[4439] = 32'b00000000000000001001101101100001;
assign LUT_3[4440] = 32'b00000000000000001001000101110000;
assign LUT_3[4441] = 32'b00000000000000001111110001001101;
assign LUT_3[4442] = 32'b00000000000000001011001101010100;
assign LUT_3[4443] = 32'b00000000000000010001111000110001;
assign LUT_3[4444] = 32'b00000000000000000110010011100110;
assign LUT_3[4445] = 32'b00000000000000001100111111000011;
assign LUT_3[4446] = 32'b00000000000000001000011011001010;
assign LUT_3[4447] = 32'b00000000000000001111000110100111;
assign LUT_3[4448] = 32'b00000000000000000001101000000111;
assign LUT_3[4449] = 32'b00000000000000001000010011100100;
assign LUT_3[4450] = 32'b00000000000000000011101111101011;
assign LUT_3[4451] = 32'b00000000000000001010011011001000;
assign LUT_3[4452] = 32'b11111111111111111110110101111101;
assign LUT_3[4453] = 32'b00000000000000000101100001011010;
assign LUT_3[4454] = 32'b00000000000000000000111101100001;
assign LUT_3[4455] = 32'b00000000000000000111101000111110;
assign LUT_3[4456] = 32'b00000000000000000111000001001101;
assign LUT_3[4457] = 32'b00000000000000001101101100101010;
assign LUT_3[4458] = 32'b00000000000000001001001000110001;
assign LUT_3[4459] = 32'b00000000000000001111110100001110;
assign LUT_3[4460] = 32'b00000000000000000100001111000011;
assign LUT_3[4461] = 32'b00000000000000001010111010100000;
assign LUT_3[4462] = 32'b00000000000000000110010110100111;
assign LUT_3[4463] = 32'b00000000000000001101000010000100;
assign LUT_3[4464] = 32'b00000000000000000100111011001010;
assign LUT_3[4465] = 32'b00000000000000001011100110100111;
assign LUT_3[4466] = 32'b00000000000000000111000010101110;
assign LUT_3[4467] = 32'b00000000000000001101101110001011;
assign LUT_3[4468] = 32'b00000000000000000010001001000000;
assign LUT_3[4469] = 32'b00000000000000001000110100011101;
assign LUT_3[4470] = 32'b00000000000000000100010000100100;
assign LUT_3[4471] = 32'b00000000000000001010111100000001;
assign LUT_3[4472] = 32'b00000000000000001010010100010000;
assign LUT_3[4473] = 32'b00000000000000010000111111101101;
assign LUT_3[4474] = 32'b00000000000000001100011011110100;
assign LUT_3[4475] = 32'b00000000000000010011000111010001;
assign LUT_3[4476] = 32'b00000000000000000111100010000110;
assign LUT_3[4477] = 32'b00000000000000001110001101100011;
assign LUT_3[4478] = 32'b00000000000000001001101001101010;
assign LUT_3[4479] = 32'b00000000000000010000010101000111;
assign LUT_3[4480] = 32'b00000000000000000010101011111010;
assign LUT_3[4481] = 32'b00000000000000001001010111010111;
assign LUT_3[4482] = 32'b00000000000000000100110011011110;
assign LUT_3[4483] = 32'b00000000000000001011011110111011;
assign LUT_3[4484] = 32'b11111111111111111111111001110000;
assign LUT_3[4485] = 32'b00000000000000000110100101001101;
assign LUT_3[4486] = 32'b00000000000000000010000001010100;
assign LUT_3[4487] = 32'b00000000000000001000101100110001;
assign LUT_3[4488] = 32'b00000000000000001000000101000000;
assign LUT_3[4489] = 32'b00000000000000001110110000011101;
assign LUT_3[4490] = 32'b00000000000000001010001100100100;
assign LUT_3[4491] = 32'b00000000000000010000111000000001;
assign LUT_3[4492] = 32'b00000000000000000101010010110110;
assign LUT_3[4493] = 32'b00000000000000001011111110010011;
assign LUT_3[4494] = 32'b00000000000000000111011010011010;
assign LUT_3[4495] = 32'b00000000000000001110000101110111;
assign LUT_3[4496] = 32'b00000000000000000101111110111101;
assign LUT_3[4497] = 32'b00000000000000001100101010011010;
assign LUT_3[4498] = 32'b00000000000000001000000110100001;
assign LUT_3[4499] = 32'b00000000000000001110110001111110;
assign LUT_3[4500] = 32'b00000000000000000011001100110011;
assign LUT_3[4501] = 32'b00000000000000001001111000010000;
assign LUT_3[4502] = 32'b00000000000000000101010100010111;
assign LUT_3[4503] = 32'b00000000000000001011111111110100;
assign LUT_3[4504] = 32'b00000000000000001011011000000011;
assign LUT_3[4505] = 32'b00000000000000010010000011100000;
assign LUT_3[4506] = 32'b00000000000000001101011111100111;
assign LUT_3[4507] = 32'b00000000000000010100001011000100;
assign LUT_3[4508] = 32'b00000000000000001000100101111001;
assign LUT_3[4509] = 32'b00000000000000001111010001010110;
assign LUT_3[4510] = 32'b00000000000000001010101101011101;
assign LUT_3[4511] = 32'b00000000000000010001011000111010;
assign LUT_3[4512] = 32'b00000000000000000011111010011010;
assign LUT_3[4513] = 32'b00000000000000001010100101110111;
assign LUT_3[4514] = 32'b00000000000000000110000001111110;
assign LUT_3[4515] = 32'b00000000000000001100101101011011;
assign LUT_3[4516] = 32'b00000000000000000001001000010000;
assign LUT_3[4517] = 32'b00000000000000000111110011101101;
assign LUT_3[4518] = 32'b00000000000000000011001111110100;
assign LUT_3[4519] = 32'b00000000000000001001111011010001;
assign LUT_3[4520] = 32'b00000000000000001001010011100000;
assign LUT_3[4521] = 32'b00000000000000001111111110111101;
assign LUT_3[4522] = 32'b00000000000000001011011011000100;
assign LUT_3[4523] = 32'b00000000000000010010000110100001;
assign LUT_3[4524] = 32'b00000000000000000110100001010110;
assign LUT_3[4525] = 32'b00000000000000001101001100110011;
assign LUT_3[4526] = 32'b00000000000000001000101000111010;
assign LUT_3[4527] = 32'b00000000000000001111010100010111;
assign LUT_3[4528] = 32'b00000000000000000111001101011101;
assign LUT_3[4529] = 32'b00000000000000001101111000111010;
assign LUT_3[4530] = 32'b00000000000000001001010101000001;
assign LUT_3[4531] = 32'b00000000000000010000000000011110;
assign LUT_3[4532] = 32'b00000000000000000100011011010011;
assign LUT_3[4533] = 32'b00000000000000001011000110110000;
assign LUT_3[4534] = 32'b00000000000000000110100010110111;
assign LUT_3[4535] = 32'b00000000000000001101001110010100;
assign LUT_3[4536] = 32'b00000000000000001100100110100011;
assign LUT_3[4537] = 32'b00000000000000010011010010000000;
assign LUT_3[4538] = 32'b00000000000000001110101110000111;
assign LUT_3[4539] = 32'b00000000000000010101011001100100;
assign LUT_3[4540] = 32'b00000000000000001001110100011001;
assign LUT_3[4541] = 32'b00000000000000010000011111110110;
assign LUT_3[4542] = 32'b00000000000000001011111011111101;
assign LUT_3[4543] = 32'b00000000000000010010100111011010;
assign LUT_3[4544] = 32'b00000000000000000010100100100101;
assign LUT_3[4545] = 32'b00000000000000001001010000000010;
assign LUT_3[4546] = 32'b00000000000000000100101100001001;
assign LUT_3[4547] = 32'b00000000000000001011010111100110;
assign LUT_3[4548] = 32'b11111111111111111111110010011011;
assign LUT_3[4549] = 32'b00000000000000000110011101111000;
assign LUT_3[4550] = 32'b00000000000000000001111001111111;
assign LUT_3[4551] = 32'b00000000000000001000100101011100;
assign LUT_3[4552] = 32'b00000000000000000111111101101011;
assign LUT_3[4553] = 32'b00000000000000001110101001001000;
assign LUT_3[4554] = 32'b00000000000000001010000101001111;
assign LUT_3[4555] = 32'b00000000000000010000110000101100;
assign LUT_3[4556] = 32'b00000000000000000101001011100001;
assign LUT_3[4557] = 32'b00000000000000001011110110111110;
assign LUT_3[4558] = 32'b00000000000000000111010011000101;
assign LUT_3[4559] = 32'b00000000000000001101111110100010;
assign LUT_3[4560] = 32'b00000000000000000101110111101000;
assign LUT_3[4561] = 32'b00000000000000001100100011000101;
assign LUT_3[4562] = 32'b00000000000000000111111111001100;
assign LUT_3[4563] = 32'b00000000000000001110101010101001;
assign LUT_3[4564] = 32'b00000000000000000011000101011110;
assign LUT_3[4565] = 32'b00000000000000001001110000111011;
assign LUT_3[4566] = 32'b00000000000000000101001101000010;
assign LUT_3[4567] = 32'b00000000000000001011111000011111;
assign LUT_3[4568] = 32'b00000000000000001011010000101110;
assign LUT_3[4569] = 32'b00000000000000010001111100001011;
assign LUT_3[4570] = 32'b00000000000000001101011000010010;
assign LUT_3[4571] = 32'b00000000000000010100000011101111;
assign LUT_3[4572] = 32'b00000000000000001000011110100100;
assign LUT_3[4573] = 32'b00000000000000001111001010000001;
assign LUT_3[4574] = 32'b00000000000000001010100110001000;
assign LUT_3[4575] = 32'b00000000000000010001010001100101;
assign LUT_3[4576] = 32'b00000000000000000011110011000101;
assign LUT_3[4577] = 32'b00000000000000001010011110100010;
assign LUT_3[4578] = 32'b00000000000000000101111010101001;
assign LUT_3[4579] = 32'b00000000000000001100100110000110;
assign LUT_3[4580] = 32'b00000000000000000001000000111011;
assign LUT_3[4581] = 32'b00000000000000000111101100011000;
assign LUT_3[4582] = 32'b00000000000000000011001000011111;
assign LUT_3[4583] = 32'b00000000000000001001110011111100;
assign LUT_3[4584] = 32'b00000000000000001001001100001011;
assign LUT_3[4585] = 32'b00000000000000001111110111101000;
assign LUT_3[4586] = 32'b00000000000000001011010011101111;
assign LUT_3[4587] = 32'b00000000000000010001111111001100;
assign LUT_3[4588] = 32'b00000000000000000110011010000001;
assign LUT_3[4589] = 32'b00000000000000001101000101011110;
assign LUT_3[4590] = 32'b00000000000000001000100001100101;
assign LUT_3[4591] = 32'b00000000000000001111001101000010;
assign LUT_3[4592] = 32'b00000000000000000111000110001000;
assign LUT_3[4593] = 32'b00000000000000001101110001100101;
assign LUT_3[4594] = 32'b00000000000000001001001101101100;
assign LUT_3[4595] = 32'b00000000000000001111111001001001;
assign LUT_3[4596] = 32'b00000000000000000100010011111110;
assign LUT_3[4597] = 32'b00000000000000001010111111011011;
assign LUT_3[4598] = 32'b00000000000000000110011011100010;
assign LUT_3[4599] = 32'b00000000000000001101000110111111;
assign LUT_3[4600] = 32'b00000000000000001100011111001110;
assign LUT_3[4601] = 32'b00000000000000010011001010101011;
assign LUT_3[4602] = 32'b00000000000000001110100110110010;
assign LUT_3[4603] = 32'b00000000000000010101010010001111;
assign LUT_3[4604] = 32'b00000000000000001001101101000100;
assign LUT_3[4605] = 32'b00000000000000010000011000100001;
assign LUT_3[4606] = 32'b00000000000000001011110100101000;
assign LUT_3[4607] = 32'b00000000000000010010100000000101;
assign LUT_3[4608] = 32'b00000000000000000111100110100111;
assign LUT_3[4609] = 32'b00000000000000001110010010000100;
assign LUT_3[4610] = 32'b00000000000000001001101110001011;
assign LUT_3[4611] = 32'b00000000000000010000011001101000;
assign LUT_3[4612] = 32'b00000000000000000100110100011101;
assign LUT_3[4613] = 32'b00000000000000001011011111111010;
assign LUT_3[4614] = 32'b00000000000000000110111100000001;
assign LUT_3[4615] = 32'b00000000000000001101100111011110;
assign LUT_3[4616] = 32'b00000000000000001100111111101101;
assign LUT_3[4617] = 32'b00000000000000010011101011001010;
assign LUT_3[4618] = 32'b00000000000000001111000111010001;
assign LUT_3[4619] = 32'b00000000000000010101110010101110;
assign LUT_3[4620] = 32'b00000000000000001010001101100011;
assign LUT_3[4621] = 32'b00000000000000010000111001000000;
assign LUT_3[4622] = 32'b00000000000000001100010101000111;
assign LUT_3[4623] = 32'b00000000000000010011000000100100;
assign LUT_3[4624] = 32'b00000000000000001010111001101010;
assign LUT_3[4625] = 32'b00000000000000010001100101000111;
assign LUT_3[4626] = 32'b00000000000000001101000001001110;
assign LUT_3[4627] = 32'b00000000000000010011101100101011;
assign LUT_3[4628] = 32'b00000000000000001000000111100000;
assign LUT_3[4629] = 32'b00000000000000001110110010111101;
assign LUT_3[4630] = 32'b00000000000000001010001111000100;
assign LUT_3[4631] = 32'b00000000000000010000111010100001;
assign LUT_3[4632] = 32'b00000000000000010000010010110000;
assign LUT_3[4633] = 32'b00000000000000010110111110001101;
assign LUT_3[4634] = 32'b00000000000000010010011010010100;
assign LUT_3[4635] = 32'b00000000000000011001000101110001;
assign LUT_3[4636] = 32'b00000000000000001101100000100110;
assign LUT_3[4637] = 32'b00000000000000010100001100000011;
assign LUT_3[4638] = 32'b00000000000000001111101000001010;
assign LUT_3[4639] = 32'b00000000000000010110010011100111;
assign LUT_3[4640] = 32'b00000000000000001000110101000111;
assign LUT_3[4641] = 32'b00000000000000001111100000100100;
assign LUT_3[4642] = 32'b00000000000000001010111100101011;
assign LUT_3[4643] = 32'b00000000000000010001101000001000;
assign LUT_3[4644] = 32'b00000000000000000110000010111101;
assign LUT_3[4645] = 32'b00000000000000001100101110011010;
assign LUT_3[4646] = 32'b00000000000000001000001010100001;
assign LUT_3[4647] = 32'b00000000000000001110110101111110;
assign LUT_3[4648] = 32'b00000000000000001110001110001101;
assign LUT_3[4649] = 32'b00000000000000010100111001101010;
assign LUT_3[4650] = 32'b00000000000000010000010101110001;
assign LUT_3[4651] = 32'b00000000000000010111000001001110;
assign LUT_3[4652] = 32'b00000000000000001011011100000011;
assign LUT_3[4653] = 32'b00000000000000010010000111100000;
assign LUT_3[4654] = 32'b00000000000000001101100011100111;
assign LUT_3[4655] = 32'b00000000000000010100001111000100;
assign LUT_3[4656] = 32'b00000000000000001100001000001010;
assign LUT_3[4657] = 32'b00000000000000010010110011100111;
assign LUT_3[4658] = 32'b00000000000000001110001111101110;
assign LUT_3[4659] = 32'b00000000000000010100111011001011;
assign LUT_3[4660] = 32'b00000000000000001001010110000000;
assign LUT_3[4661] = 32'b00000000000000010000000001011101;
assign LUT_3[4662] = 32'b00000000000000001011011101100100;
assign LUT_3[4663] = 32'b00000000000000010010001001000001;
assign LUT_3[4664] = 32'b00000000000000010001100001010000;
assign LUT_3[4665] = 32'b00000000000000011000001100101101;
assign LUT_3[4666] = 32'b00000000000000010011101000110100;
assign LUT_3[4667] = 32'b00000000000000011010010100010001;
assign LUT_3[4668] = 32'b00000000000000001110101111000110;
assign LUT_3[4669] = 32'b00000000000000010101011010100011;
assign LUT_3[4670] = 32'b00000000000000010000110110101010;
assign LUT_3[4671] = 32'b00000000000000010111100010000111;
assign LUT_3[4672] = 32'b00000000000000000111011111010010;
assign LUT_3[4673] = 32'b00000000000000001110001010101111;
assign LUT_3[4674] = 32'b00000000000000001001100110110110;
assign LUT_3[4675] = 32'b00000000000000010000010010010011;
assign LUT_3[4676] = 32'b00000000000000000100101101001000;
assign LUT_3[4677] = 32'b00000000000000001011011000100101;
assign LUT_3[4678] = 32'b00000000000000000110110100101100;
assign LUT_3[4679] = 32'b00000000000000001101100000001001;
assign LUT_3[4680] = 32'b00000000000000001100111000011000;
assign LUT_3[4681] = 32'b00000000000000010011100011110101;
assign LUT_3[4682] = 32'b00000000000000001110111111111100;
assign LUT_3[4683] = 32'b00000000000000010101101011011001;
assign LUT_3[4684] = 32'b00000000000000001010000110001110;
assign LUT_3[4685] = 32'b00000000000000010000110001101011;
assign LUT_3[4686] = 32'b00000000000000001100001101110010;
assign LUT_3[4687] = 32'b00000000000000010010111001001111;
assign LUT_3[4688] = 32'b00000000000000001010110010010101;
assign LUT_3[4689] = 32'b00000000000000010001011101110010;
assign LUT_3[4690] = 32'b00000000000000001100111001111001;
assign LUT_3[4691] = 32'b00000000000000010011100101010110;
assign LUT_3[4692] = 32'b00000000000000001000000000001011;
assign LUT_3[4693] = 32'b00000000000000001110101011101000;
assign LUT_3[4694] = 32'b00000000000000001010000111101111;
assign LUT_3[4695] = 32'b00000000000000010000110011001100;
assign LUT_3[4696] = 32'b00000000000000010000001011011011;
assign LUT_3[4697] = 32'b00000000000000010110110110111000;
assign LUT_3[4698] = 32'b00000000000000010010010010111111;
assign LUT_3[4699] = 32'b00000000000000011000111110011100;
assign LUT_3[4700] = 32'b00000000000000001101011001010001;
assign LUT_3[4701] = 32'b00000000000000010100000100101110;
assign LUT_3[4702] = 32'b00000000000000001111100000110101;
assign LUT_3[4703] = 32'b00000000000000010110001100010010;
assign LUT_3[4704] = 32'b00000000000000001000101101110010;
assign LUT_3[4705] = 32'b00000000000000001111011001001111;
assign LUT_3[4706] = 32'b00000000000000001010110101010110;
assign LUT_3[4707] = 32'b00000000000000010001100000110011;
assign LUT_3[4708] = 32'b00000000000000000101111011101000;
assign LUT_3[4709] = 32'b00000000000000001100100111000101;
assign LUT_3[4710] = 32'b00000000000000001000000011001100;
assign LUT_3[4711] = 32'b00000000000000001110101110101001;
assign LUT_3[4712] = 32'b00000000000000001110000110111000;
assign LUT_3[4713] = 32'b00000000000000010100110010010101;
assign LUT_3[4714] = 32'b00000000000000010000001110011100;
assign LUT_3[4715] = 32'b00000000000000010110111001111001;
assign LUT_3[4716] = 32'b00000000000000001011010100101110;
assign LUT_3[4717] = 32'b00000000000000010010000000001011;
assign LUT_3[4718] = 32'b00000000000000001101011100010010;
assign LUT_3[4719] = 32'b00000000000000010100000111101111;
assign LUT_3[4720] = 32'b00000000000000001100000000110101;
assign LUT_3[4721] = 32'b00000000000000010010101100010010;
assign LUT_3[4722] = 32'b00000000000000001110001000011001;
assign LUT_3[4723] = 32'b00000000000000010100110011110110;
assign LUT_3[4724] = 32'b00000000000000001001001110101011;
assign LUT_3[4725] = 32'b00000000000000001111111010001000;
assign LUT_3[4726] = 32'b00000000000000001011010110001111;
assign LUT_3[4727] = 32'b00000000000000010010000001101100;
assign LUT_3[4728] = 32'b00000000000000010001011001111011;
assign LUT_3[4729] = 32'b00000000000000011000000101011000;
assign LUT_3[4730] = 32'b00000000000000010011100001011111;
assign LUT_3[4731] = 32'b00000000000000011010001100111100;
assign LUT_3[4732] = 32'b00000000000000001110100111110001;
assign LUT_3[4733] = 32'b00000000000000010101010011001110;
assign LUT_3[4734] = 32'b00000000000000010000101111010101;
assign LUT_3[4735] = 32'b00000000000000010111011010110010;
assign LUT_3[4736] = 32'b00000000000000001001110001100101;
assign LUT_3[4737] = 32'b00000000000000010000011101000010;
assign LUT_3[4738] = 32'b00000000000000001011111001001001;
assign LUT_3[4739] = 32'b00000000000000010010100100100110;
assign LUT_3[4740] = 32'b00000000000000000110111111011011;
assign LUT_3[4741] = 32'b00000000000000001101101010111000;
assign LUT_3[4742] = 32'b00000000000000001001000110111111;
assign LUT_3[4743] = 32'b00000000000000001111110010011100;
assign LUT_3[4744] = 32'b00000000000000001111001010101011;
assign LUT_3[4745] = 32'b00000000000000010101110110001000;
assign LUT_3[4746] = 32'b00000000000000010001010010001111;
assign LUT_3[4747] = 32'b00000000000000010111111101101100;
assign LUT_3[4748] = 32'b00000000000000001100011000100001;
assign LUT_3[4749] = 32'b00000000000000010011000011111110;
assign LUT_3[4750] = 32'b00000000000000001110100000000101;
assign LUT_3[4751] = 32'b00000000000000010101001011100010;
assign LUT_3[4752] = 32'b00000000000000001101000100101000;
assign LUT_3[4753] = 32'b00000000000000010011110000000101;
assign LUT_3[4754] = 32'b00000000000000001111001100001100;
assign LUT_3[4755] = 32'b00000000000000010101110111101001;
assign LUT_3[4756] = 32'b00000000000000001010010010011110;
assign LUT_3[4757] = 32'b00000000000000010000111101111011;
assign LUT_3[4758] = 32'b00000000000000001100011010000010;
assign LUT_3[4759] = 32'b00000000000000010011000101011111;
assign LUT_3[4760] = 32'b00000000000000010010011101101110;
assign LUT_3[4761] = 32'b00000000000000011001001001001011;
assign LUT_3[4762] = 32'b00000000000000010100100101010010;
assign LUT_3[4763] = 32'b00000000000000011011010000101111;
assign LUT_3[4764] = 32'b00000000000000001111101011100100;
assign LUT_3[4765] = 32'b00000000000000010110010111000001;
assign LUT_3[4766] = 32'b00000000000000010001110011001000;
assign LUT_3[4767] = 32'b00000000000000011000011110100101;
assign LUT_3[4768] = 32'b00000000000000001011000000000101;
assign LUT_3[4769] = 32'b00000000000000010001101011100010;
assign LUT_3[4770] = 32'b00000000000000001101000111101001;
assign LUT_3[4771] = 32'b00000000000000010011110011000110;
assign LUT_3[4772] = 32'b00000000000000001000001101111011;
assign LUT_3[4773] = 32'b00000000000000001110111001011000;
assign LUT_3[4774] = 32'b00000000000000001010010101011111;
assign LUT_3[4775] = 32'b00000000000000010001000000111100;
assign LUT_3[4776] = 32'b00000000000000010000011001001011;
assign LUT_3[4777] = 32'b00000000000000010111000100101000;
assign LUT_3[4778] = 32'b00000000000000010010100000101111;
assign LUT_3[4779] = 32'b00000000000000011001001100001100;
assign LUT_3[4780] = 32'b00000000000000001101100111000001;
assign LUT_3[4781] = 32'b00000000000000010100010010011110;
assign LUT_3[4782] = 32'b00000000000000001111101110100101;
assign LUT_3[4783] = 32'b00000000000000010110011010000010;
assign LUT_3[4784] = 32'b00000000000000001110010011001000;
assign LUT_3[4785] = 32'b00000000000000010100111110100101;
assign LUT_3[4786] = 32'b00000000000000010000011010101100;
assign LUT_3[4787] = 32'b00000000000000010111000110001001;
assign LUT_3[4788] = 32'b00000000000000001011100000111110;
assign LUT_3[4789] = 32'b00000000000000010010001100011011;
assign LUT_3[4790] = 32'b00000000000000001101101000100010;
assign LUT_3[4791] = 32'b00000000000000010100010011111111;
assign LUT_3[4792] = 32'b00000000000000010011101100001110;
assign LUT_3[4793] = 32'b00000000000000011010010111101011;
assign LUT_3[4794] = 32'b00000000000000010101110011110010;
assign LUT_3[4795] = 32'b00000000000000011100011111001111;
assign LUT_3[4796] = 32'b00000000000000010000111010000100;
assign LUT_3[4797] = 32'b00000000000000010111100101100001;
assign LUT_3[4798] = 32'b00000000000000010011000001101000;
assign LUT_3[4799] = 32'b00000000000000011001101101000101;
assign LUT_3[4800] = 32'b00000000000000001001101010010000;
assign LUT_3[4801] = 32'b00000000000000010000010101101101;
assign LUT_3[4802] = 32'b00000000000000001011110001110100;
assign LUT_3[4803] = 32'b00000000000000010010011101010001;
assign LUT_3[4804] = 32'b00000000000000000110111000000110;
assign LUT_3[4805] = 32'b00000000000000001101100011100011;
assign LUT_3[4806] = 32'b00000000000000001000111111101010;
assign LUT_3[4807] = 32'b00000000000000001111101011000111;
assign LUT_3[4808] = 32'b00000000000000001111000011010110;
assign LUT_3[4809] = 32'b00000000000000010101101110110011;
assign LUT_3[4810] = 32'b00000000000000010001001010111010;
assign LUT_3[4811] = 32'b00000000000000010111110110010111;
assign LUT_3[4812] = 32'b00000000000000001100010001001100;
assign LUT_3[4813] = 32'b00000000000000010010111100101001;
assign LUT_3[4814] = 32'b00000000000000001110011000110000;
assign LUT_3[4815] = 32'b00000000000000010101000100001101;
assign LUT_3[4816] = 32'b00000000000000001100111101010011;
assign LUT_3[4817] = 32'b00000000000000010011101000110000;
assign LUT_3[4818] = 32'b00000000000000001111000100110111;
assign LUT_3[4819] = 32'b00000000000000010101110000010100;
assign LUT_3[4820] = 32'b00000000000000001010001011001001;
assign LUT_3[4821] = 32'b00000000000000010000110110100110;
assign LUT_3[4822] = 32'b00000000000000001100010010101101;
assign LUT_3[4823] = 32'b00000000000000010010111110001010;
assign LUT_3[4824] = 32'b00000000000000010010010110011001;
assign LUT_3[4825] = 32'b00000000000000011001000001110110;
assign LUT_3[4826] = 32'b00000000000000010100011101111101;
assign LUT_3[4827] = 32'b00000000000000011011001001011010;
assign LUT_3[4828] = 32'b00000000000000001111100100001111;
assign LUT_3[4829] = 32'b00000000000000010110001111101100;
assign LUT_3[4830] = 32'b00000000000000010001101011110011;
assign LUT_3[4831] = 32'b00000000000000011000010111010000;
assign LUT_3[4832] = 32'b00000000000000001010111000110000;
assign LUT_3[4833] = 32'b00000000000000010001100100001101;
assign LUT_3[4834] = 32'b00000000000000001101000000010100;
assign LUT_3[4835] = 32'b00000000000000010011101011110001;
assign LUT_3[4836] = 32'b00000000000000001000000110100110;
assign LUT_3[4837] = 32'b00000000000000001110110010000011;
assign LUT_3[4838] = 32'b00000000000000001010001110001010;
assign LUT_3[4839] = 32'b00000000000000010000111001100111;
assign LUT_3[4840] = 32'b00000000000000010000010001110110;
assign LUT_3[4841] = 32'b00000000000000010110111101010011;
assign LUT_3[4842] = 32'b00000000000000010010011001011010;
assign LUT_3[4843] = 32'b00000000000000011001000100110111;
assign LUT_3[4844] = 32'b00000000000000001101011111101100;
assign LUT_3[4845] = 32'b00000000000000010100001011001001;
assign LUT_3[4846] = 32'b00000000000000001111100111010000;
assign LUT_3[4847] = 32'b00000000000000010110010010101101;
assign LUT_3[4848] = 32'b00000000000000001110001011110011;
assign LUT_3[4849] = 32'b00000000000000010100110111010000;
assign LUT_3[4850] = 32'b00000000000000010000010011010111;
assign LUT_3[4851] = 32'b00000000000000010110111110110100;
assign LUT_3[4852] = 32'b00000000000000001011011001101001;
assign LUT_3[4853] = 32'b00000000000000010010000101000110;
assign LUT_3[4854] = 32'b00000000000000001101100001001101;
assign LUT_3[4855] = 32'b00000000000000010100001100101010;
assign LUT_3[4856] = 32'b00000000000000010011100100111001;
assign LUT_3[4857] = 32'b00000000000000011010010000010110;
assign LUT_3[4858] = 32'b00000000000000010101101100011101;
assign LUT_3[4859] = 32'b00000000000000011100010111111010;
assign LUT_3[4860] = 32'b00000000000000010000110010101111;
assign LUT_3[4861] = 32'b00000000000000010111011110001100;
assign LUT_3[4862] = 32'b00000000000000010010111010010011;
assign LUT_3[4863] = 32'b00000000000000011001100101110000;
assign LUT_3[4864] = 32'b00000000000000000011110110001000;
assign LUT_3[4865] = 32'b00000000000000001010100001100101;
assign LUT_3[4866] = 32'b00000000000000000101111101101100;
assign LUT_3[4867] = 32'b00000000000000001100101001001001;
assign LUT_3[4868] = 32'b00000000000000000001000011111110;
assign LUT_3[4869] = 32'b00000000000000000111101111011011;
assign LUT_3[4870] = 32'b00000000000000000011001011100010;
assign LUT_3[4871] = 32'b00000000000000001001110110111111;
assign LUT_3[4872] = 32'b00000000000000001001001111001110;
assign LUT_3[4873] = 32'b00000000000000001111111010101011;
assign LUT_3[4874] = 32'b00000000000000001011010110110010;
assign LUT_3[4875] = 32'b00000000000000010010000010001111;
assign LUT_3[4876] = 32'b00000000000000000110011101000100;
assign LUT_3[4877] = 32'b00000000000000001101001000100001;
assign LUT_3[4878] = 32'b00000000000000001000100100101000;
assign LUT_3[4879] = 32'b00000000000000001111010000000101;
assign LUT_3[4880] = 32'b00000000000000000111001001001011;
assign LUT_3[4881] = 32'b00000000000000001101110100101000;
assign LUT_3[4882] = 32'b00000000000000001001010000101111;
assign LUT_3[4883] = 32'b00000000000000001111111100001100;
assign LUT_3[4884] = 32'b00000000000000000100010111000001;
assign LUT_3[4885] = 32'b00000000000000001011000010011110;
assign LUT_3[4886] = 32'b00000000000000000110011110100101;
assign LUT_3[4887] = 32'b00000000000000001101001010000010;
assign LUT_3[4888] = 32'b00000000000000001100100010010001;
assign LUT_3[4889] = 32'b00000000000000010011001101101110;
assign LUT_3[4890] = 32'b00000000000000001110101001110101;
assign LUT_3[4891] = 32'b00000000000000010101010101010010;
assign LUT_3[4892] = 32'b00000000000000001001110000000111;
assign LUT_3[4893] = 32'b00000000000000010000011011100100;
assign LUT_3[4894] = 32'b00000000000000001011110111101011;
assign LUT_3[4895] = 32'b00000000000000010010100011001000;
assign LUT_3[4896] = 32'b00000000000000000101000100101000;
assign LUT_3[4897] = 32'b00000000000000001011110000000101;
assign LUT_3[4898] = 32'b00000000000000000111001100001100;
assign LUT_3[4899] = 32'b00000000000000001101110111101001;
assign LUT_3[4900] = 32'b00000000000000000010010010011110;
assign LUT_3[4901] = 32'b00000000000000001000111101111011;
assign LUT_3[4902] = 32'b00000000000000000100011010000010;
assign LUT_3[4903] = 32'b00000000000000001011000101011111;
assign LUT_3[4904] = 32'b00000000000000001010011101101110;
assign LUT_3[4905] = 32'b00000000000000010001001001001011;
assign LUT_3[4906] = 32'b00000000000000001100100101010010;
assign LUT_3[4907] = 32'b00000000000000010011010000101111;
assign LUT_3[4908] = 32'b00000000000000000111101011100100;
assign LUT_3[4909] = 32'b00000000000000001110010111000001;
assign LUT_3[4910] = 32'b00000000000000001001110011001000;
assign LUT_3[4911] = 32'b00000000000000010000011110100101;
assign LUT_3[4912] = 32'b00000000000000001000010111101011;
assign LUT_3[4913] = 32'b00000000000000001111000011001000;
assign LUT_3[4914] = 32'b00000000000000001010011111001111;
assign LUT_3[4915] = 32'b00000000000000010001001010101100;
assign LUT_3[4916] = 32'b00000000000000000101100101100001;
assign LUT_3[4917] = 32'b00000000000000001100010000111110;
assign LUT_3[4918] = 32'b00000000000000000111101101000101;
assign LUT_3[4919] = 32'b00000000000000001110011000100010;
assign LUT_3[4920] = 32'b00000000000000001101110000110001;
assign LUT_3[4921] = 32'b00000000000000010100011100001110;
assign LUT_3[4922] = 32'b00000000000000001111111000010101;
assign LUT_3[4923] = 32'b00000000000000010110100011110010;
assign LUT_3[4924] = 32'b00000000000000001010111110100111;
assign LUT_3[4925] = 32'b00000000000000010001101010000100;
assign LUT_3[4926] = 32'b00000000000000001101000110001011;
assign LUT_3[4927] = 32'b00000000000000010011110001101000;
assign LUT_3[4928] = 32'b00000000000000000011101110110011;
assign LUT_3[4929] = 32'b00000000000000001010011010010000;
assign LUT_3[4930] = 32'b00000000000000000101110110010111;
assign LUT_3[4931] = 32'b00000000000000001100100001110100;
assign LUT_3[4932] = 32'b00000000000000000000111100101001;
assign LUT_3[4933] = 32'b00000000000000000111101000000110;
assign LUT_3[4934] = 32'b00000000000000000011000100001101;
assign LUT_3[4935] = 32'b00000000000000001001101111101010;
assign LUT_3[4936] = 32'b00000000000000001001000111111001;
assign LUT_3[4937] = 32'b00000000000000001111110011010110;
assign LUT_3[4938] = 32'b00000000000000001011001111011101;
assign LUT_3[4939] = 32'b00000000000000010001111010111010;
assign LUT_3[4940] = 32'b00000000000000000110010101101111;
assign LUT_3[4941] = 32'b00000000000000001101000001001100;
assign LUT_3[4942] = 32'b00000000000000001000011101010011;
assign LUT_3[4943] = 32'b00000000000000001111001000110000;
assign LUT_3[4944] = 32'b00000000000000000111000001110110;
assign LUT_3[4945] = 32'b00000000000000001101101101010011;
assign LUT_3[4946] = 32'b00000000000000001001001001011010;
assign LUT_3[4947] = 32'b00000000000000001111110100110111;
assign LUT_3[4948] = 32'b00000000000000000100001111101100;
assign LUT_3[4949] = 32'b00000000000000001010111011001001;
assign LUT_3[4950] = 32'b00000000000000000110010111010000;
assign LUT_3[4951] = 32'b00000000000000001101000010101101;
assign LUT_3[4952] = 32'b00000000000000001100011010111100;
assign LUT_3[4953] = 32'b00000000000000010011000110011001;
assign LUT_3[4954] = 32'b00000000000000001110100010100000;
assign LUT_3[4955] = 32'b00000000000000010101001101111101;
assign LUT_3[4956] = 32'b00000000000000001001101000110010;
assign LUT_3[4957] = 32'b00000000000000010000010100001111;
assign LUT_3[4958] = 32'b00000000000000001011110000010110;
assign LUT_3[4959] = 32'b00000000000000010010011011110011;
assign LUT_3[4960] = 32'b00000000000000000100111101010011;
assign LUT_3[4961] = 32'b00000000000000001011101000110000;
assign LUT_3[4962] = 32'b00000000000000000111000100110111;
assign LUT_3[4963] = 32'b00000000000000001101110000010100;
assign LUT_3[4964] = 32'b00000000000000000010001011001001;
assign LUT_3[4965] = 32'b00000000000000001000110110100110;
assign LUT_3[4966] = 32'b00000000000000000100010010101101;
assign LUT_3[4967] = 32'b00000000000000001010111110001010;
assign LUT_3[4968] = 32'b00000000000000001010010110011001;
assign LUT_3[4969] = 32'b00000000000000010001000001110110;
assign LUT_3[4970] = 32'b00000000000000001100011101111101;
assign LUT_3[4971] = 32'b00000000000000010011001001011010;
assign LUT_3[4972] = 32'b00000000000000000111100100001111;
assign LUT_3[4973] = 32'b00000000000000001110001111101100;
assign LUT_3[4974] = 32'b00000000000000001001101011110011;
assign LUT_3[4975] = 32'b00000000000000010000010111010000;
assign LUT_3[4976] = 32'b00000000000000001000010000010110;
assign LUT_3[4977] = 32'b00000000000000001110111011110011;
assign LUT_3[4978] = 32'b00000000000000001010010111111010;
assign LUT_3[4979] = 32'b00000000000000010001000011010111;
assign LUT_3[4980] = 32'b00000000000000000101011110001100;
assign LUT_3[4981] = 32'b00000000000000001100001001101001;
assign LUT_3[4982] = 32'b00000000000000000111100101110000;
assign LUT_3[4983] = 32'b00000000000000001110010001001101;
assign LUT_3[4984] = 32'b00000000000000001101101001011100;
assign LUT_3[4985] = 32'b00000000000000010100010100111001;
assign LUT_3[4986] = 32'b00000000000000001111110001000000;
assign LUT_3[4987] = 32'b00000000000000010110011100011101;
assign LUT_3[4988] = 32'b00000000000000001010110111010010;
assign LUT_3[4989] = 32'b00000000000000010001100010101111;
assign LUT_3[4990] = 32'b00000000000000001100111110110110;
assign LUT_3[4991] = 32'b00000000000000010011101010010011;
assign LUT_3[4992] = 32'b00000000000000000110000001000110;
assign LUT_3[4993] = 32'b00000000000000001100101100100011;
assign LUT_3[4994] = 32'b00000000000000001000001000101010;
assign LUT_3[4995] = 32'b00000000000000001110110100000111;
assign LUT_3[4996] = 32'b00000000000000000011001110111100;
assign LUT_3[4997] = 32'b00000000000000001001111010011001;
assign LUT_3[4998] = 32'b00000000000000000101010110100000;
assign LUT_3[4999] = 32'b00000000000000001100000001111101;
assign LUT_3[5000] = 32'b00000000000000001011011010001100;
assign LUT_3[5001] = 32'b00000000000000010010000101101001;
assign LUT_3[5002] = 32'b00000000000000001101100001110000;
assign LUT_3[5003] = 32'b00000000000000010100001101001101;
assign LUT_3[5004] = 32'b00000000000000001000101000000010;
assign LUT_3[5005] = 32'b00000000000000001111010011011111;
assign LUT_3[5006] = 32'b00000000000000001010101111100110;
assign LUT_3[5007] = 32'b00000000000000010001011011000011;
assign LUT_3[5008] = 32'b00000000000000001001010100001001;
assign LUT_3[5009] = 32'b00000000000000001111111111100110;
assign LUT_3[5010] = 32'b00000000000000001011011011101101;
assign LUT_3[5011] = 32'b00000000000000010010000111001010;
assign LUT_3[5012] = 32'b00000000000000000110100001111111;
assign LUT_3[5013] = 32'b00000000000000001101001101011100;
assign LUT_3[5014] = 32'b00000000000000001000101001100011;
assign LUT_3[5015] = 32'b00000000000000001111010101000000;
assign LUT_3[5016] = 32'b00000000000000001110101101001111;
assign LUT_3[5017] = 32'b00000000000000010101011000101100;
assign LUT_3[5018] = 32'b00000000000000010000110100110011;
assign LUT_3[5019] = 32'b00000000000000010111100000010000;
assign LUT_3[5020] = 32'b00000000000000001011111011000101;
assign LUT_3[5021] = 32'b00000000000000010010100110100010;
assign LUT_3[5022] = 32'b00000000000000001110000010101001;
assign LUT_3[5023] = 32'b00000000000000010100101110000110;
assign LUT_3[5024] = 32'b00000000000000000111001111100110;
assign LUT_3[5025] = 32'b00000000000000001101111011000011;
assign LUT_3[5026] = 32'b00000000000000001001010111001010;
assign LUT_3[5027] = 32'b00000000000000010000000010100111;
assign LUT_3[5028] = 32'b00000000000000000100011101011100;
assign LUT_3[5029] = 32'b00000000000000001011001000111001;
assign LUT_3[5030] = 32'b00000000000000000110100101000000;
assign LUT_3[5031] = 32'b00000000000000001101010000011101;
assign LUT_3[5032] = 32'b00000000000000001100101000101100;
assign LUT_3[5033] = 32'b00000000000000010011010100001001;
assign LUT_3[5034] = 32'b00000000000000001110110000010000;
assign LUT_3[5035] = 32'b00000000000000010101011011101101;
assign LUT_3[5036] = 32'b00000000000000001001110110100010;
assign LUT_3[5037] = 32'b00000000000000010000100001111111;
assign LUT_3[5038] = 32'b00000000000000001011111110000110;
assign LUT_3[5039] = 32'b00000000000000010010101001100011;
assign LUT_3[5040] = 32'b00000000000000001010100010101001;
assign LUT_3[5041] = 32'b00000000000000010001001110000110;
assign LUT_3[5042] = 32'b00000000000000001100101010001101;
assign LUT_3[5043] = 32'b00000000000000010011010101101010;
assign LUT_3[5044] = 32'b00000000000000000111110000011111;
assign LUT_3[5045] = 32'b00000000000000001110011011111100;
assign LUT_3[5046] = 32'b00000000000000001001111000000011;
assign LUT_3[5047] = 32'b00000000000000010000100011100000;
assign LUT_3[5048] = 32'b00000000000000001111111011101111;
assign LUT_3[5049] = 32'b00000000000000010110100111001100;
assign LUT_3[5050] = 32'b00000000000000010010000011010011;
assign LUT_3[5051] = 32'b00000000000000011000101110110000;
assign LUT_3[5052] = 32'b00000000000000001101001001100101;
assign LUT_3[5053] = 32'b00000000000000010011110101000010;
assign LUT_3[5054] = 32'b00000000000000001111010001001001;
assign LUT_3[5055] = 32'b00000000000000010101111100100110;
assign LUT_3[5056] = 32'b00000000000000000101111001110001;
assign LUT_3[5057] = 32'b00000000000000001100100101001110;
assign LUT_3[5058] = 32'b00000000000000001000000001010101;
assign LUT_3[5059] = 32'b00000000000000001110101100110010;
assign LUT_3[5060] = 32'b00000000000000000011000111100111;
assign LUT_3[5061] = 32'b00000000000000001001110011000100;
assign LUT_3[5062] = 32'b00000000000000000101001111001011;
assign LUT_3[5063] = 32'b00000000000000001011111010101000;
assign LUT_3[5064] = 32'b00000000000000001011010010110111;
assign LUT_3[5065] = 32'b00000000000000010001111110010100;
assign LUT_3[5066] = 32'b00000000000000001101011010011011;
assign LUT_3[5067] = 32'b00000000000000010100000101111000;
assign LUT_3[5068] = 32'b00000000000000001000100000101101;
assign LUT_3[5069] = 32'b00000000000000001111001100001010;
assign LUT_3[5070] = 32'b00000000000000001010101000010001;
assign LUT_3[5071] = 32'b00000000000000010001010011101110;
assign LUT_3[5072] = 32'b00000000000000001001001100110100;
assign LUT_3[5073] = 32'b00000000000000001111111000010001;
assign LUT_3[5074] = 32'b00000000000000001011010100011000;
assign LUT_3[5075] = 32'b00000000000000010001111111110101;
assign LUT_3[5076] = 32'b00000000000000000110011010101010;
assign LUT_3[5077] = 32'b00000000000000001101000110000111;
assign LUT_3[5078] = 32'b00000000000000001000100010001110;
assign LUT_3[5079] = 32'b00000000000000001111001101101011;
assign LUT_3[5080] = 32'b00000000000000001110100101111010;
assign LUT_3[5081] = 32'b00000000000000010101010001010111;
assign LUT_3[5082] = 32'b00000000000000010000101101011110;
assign LUT_3[5083] = 32'b00000000000000010111011000111011;
assign LUT_3[5084] = 32'b00000000000000001011110011110000;
assign LUT_3[5085] = 32'b00000000000000010010011111001101;
assign LUT_3[5086] = 32'b00000000000000001101111011010100;
assign LUT_3[5087] = 32'b00000000000000010100100110110001;
assign LUT_3[5088] = 32'b00000000000000000111001000010001;
assign LUT_3[5089] = 32'b00000000000000001101110011101110;
assign LUT_3[5090] = 32'b00000000000000001001001111110101;
assign LUT_3[5091] = 32'b00000000000000001111111011010010;
assign LUT_3[5092] = 32'b00000000000000000100010110000111;
assign LUT_3[5093] = 32'b00000000000000001011000001100100;
assign LUT_3[5094] = 32'b00000000000000000110011101101011;
assign LUT_3[5095] = 32'b00000000000000001101001001001000;
assign LUT_3[5096] = 32'b00000000000000001100100001010111;
assign LUT_3[5097] = 32'b00000000000000010011001100110100;
assign LUT_3[5098] = 32'b00000000000000001110101000111011;
assign LUT_3[5099] = 32'b00000000000000010101010100011000;
assign LUT_3[5100] = 32'b00000000000000001001101111001101;
assign LUT_3[5101] = 32'b00000000000000010000011010101010;
assign LUT_3[5102] = 32'b00000000000000001011110110110001;
assign LUT_3[5103] = 32'b00000000000000010010100010001110;
assign LUT_3[5104] = 32'b00000000000000001010011011010100;
assign LUT_3[5105] = 32'b00000000000000010001000110110001;
assign LUT_3[5106] = 32'b00000000000000001100100010111000;
assign LUT_3[5107] = 32'b00000000000000010011001110010101;
assign LUT_3[5108] = 32'b00000000000000000111101001001010;
assign LUT_3[5109] = 32'b00000000000000001110010100100111;
assign LUT_3[5110] = 32'b00000000000000001001110000101110;
assign LUT_3[5111] = 32'b00000000000000010000011100001011;
assign LUT_3[5112] = 32'b00000000000000001111110100011010;
assign LUT_3[5113] = 32'b00000000000000010110011111110111;
assign LUT_3[5114] = 32'b00000000000000010001111011111110;
assign LUT_3[5115] = 32'b00000000000000011000100111011011;
assign LUT_3[5116] = 32'b00000000000000001101000010010000;
assign LUT_3[5117] = 32'b00000000000000010011101101101101;
assign LUT_3[5118] = 32'b00000000000000001111001001110100;
assign LUT_3[5119] = 32'b00000000000000010101110101010001;
assign LUT_3[5120] = 32'b00000000000000001010110110011000;
assign LUT_3[5121] = 32'b00000000000000010001100001110101;
assign LUT_3[5122] = 32'b00000000000000001100111101111100;
assign LUT_3[5123] = 32'b00000000000000010011101001011001;
assign LUT_3[5124] = 32'b00000000000000001000000100001110;
assign LUT_3[5125] = 32'b00000000000000001110101111101011;
assign LUT_3[5126] = 32'b00000000000000001010001011110010;
assign LUT_3[5127] = 32'b00000000000000010000110111001111;
assign LUT_3[5128] = 32'b00000000000000010000001111011110;
assign LUT_3[5129] = 32'b00000000000000010110111010111011;
assign LUT_3[5130] = 32'b00000000000000010010010111000010;
assign LUT_3[5131] = 32'b00000000000000011001000010011111;
assign LUT_3[5132] = 32'b00000000000000001101011101010100;
assign LUT_3[5133] = 32'b00000000000000010100001000110001;
assign LUT_3[5134] = 32'b00000000000000001111100100111000;
assign LUT_3[5135] = 32'b00000000000000010110010000010101;
assign LUT_3[5136] = 32'b00000000000000001110001001011011;
assign LUT_3[5137] = 32'b00000000000000010100110100111000;
assign LUT_3[5138] = 32'b00000000000000010000010000111111;
assign LUT_3[5139] = 32'b00000000000000010110111100011100;
assign LUT_3[5140] = 32'b00000000000000001011010111010001;
assign LUT_3[5141] = 32'b00000000000000010010000010101110;
assign LUT_3[5142] = 32'b00000000000000001101011110110101;
assign LUT_3[5143] = 32'b00000000000000010100001010010010;
assign LUT_3[5144] = 32'b00000000000000010011100010100001;
assign LUT_3[5145] = 32'b00000000000000011010001101111110;
assign LUT_3[5146] = 32'b00000000000000010101101010000101;
assign LUT_3[5147] = 32'b00000000000000011100010101100010;
assign LUT_3[5148] = 32'b00000000000000010000110000010111;
assign LUT_3[5149] = 32'b00000000000000010111011011110100;
assign LUT_3[5150] = 32'b00000000000000010010110111111011;
assign LUT_3[5151] = 32'b00000000000000011001100011011000;
assign LUT_3[5152] = 32'b00000000000000001100000100111000;
assign LUT_3[5153] = 32'b00000000000000010010110000010101;
assign LUT_3[5154] = 32'b00000000000000001110001100011100;
assign LUT_3[5155] = 32'b00000000000000010100110111111001;
assign LUT_3[5156] = 32'b00000000000000001001010010101110;
assign LUT_3[5157] = 32'b00000000000000001111111110001011;
assign LUT_3[5158] = 32'b00000000000000001011011010010010;
assign LUT_3[5159] = 32'b00000000000000010010000101101111;
assign LUT_3[5160] = 32'b00000000000000010001011101111110;
assign LUT_3[5161] = 32'b00000000000000011000001001011011;
assign LUT_3[5162] = 32'b00000000000000010011100101100010;
assign LUT_3[5163] = 32'b00000000000000011010010000111111;
assign LUT_3[5164] = 32'b00000000000000001110101011110100;
assign LUT_3[5165] = 32'b00000000000000010101010111010001;
assign LUT_3[5166] = 32'b00000000000000010000110011011000;
assign LUT_3[5167] = 32'b00000000000000010111011110110101;
assign LUT_3[5168] = 32'b00000000000000001111010111111011;
assign LUT_3[5169] = 32'b00000000000000010110000011011000;
assign LUT_3[5170] = 32'b00000000000000010001011111011111;
assign LUT_3[5171] = 32'b00000000000000011000001010111100;
assign LUT_3[5172] = 32'b00000000000000001100100101110001;
assign LUT_3[5173] = 32'b00000000000000010011010001001110;
assign LUT_3[5174] = 32'b00000000000000001110101101010101;
assign LUT_3[5175] = 32'b00000000000000010101011000110010;
assign LUT_3[5176] = 32'b00000000000000010100110001000001;
assign LUT_3[5177] = 32'b00000000000000011011011100011110;
assign LUT_3[5178] = 32'b00000000000000010110111000100101;
assign LUT_3[5179] = 32'b00000000000000011101100100000010;
assign LUT_3[5180] = 32'b00000000000000010001111110110111;
assign LUT_3[5181] = 32'b00000000000000011000101010010100;
assign LUT_3[5182] = 32'b00000000000000010100000110011011;
assign LUT_3[5183] = 32'b00000000000000011010110001111000;
assign LUT_3[5184] = 32'b00000000000000001010101111000011;
assign LUT_3[5185] = 32'b00000000000000010001011010100000;
assign LUT_3[5186] = 32'b00000000000000001100110110100111;
assign LUT_3[5187] = 32'b00000000000000010011100010000100;
assign LUT_3[5188] = 32'b00000000000000000111111100111001;
assign LUT_3[5189] = 32'b00000000000000001110101000010110;
assign LUT_3[5190] = 32'b00000000000000001010000100011101;
assign LUT_3[5191] = 32'b00000000000000010000101111111010;
assign LUT_3[5192] = 32'b00000000000000010000001000001001;
assign LUT_3[5193] = 32'b00000000000000010110110011100110;
assign LUT_3[5194] = 32'b00000000000000010010001111101101;
assign LUT_3[5195] = 32'b00000000000000011000111011001010;
assign LUT_3[5196] = 32'b00000000000000001101010101111111;
assign LUT_3[5197] = 32'b00000000000000010100000001011100;
assign LUT_3[5198] = 32'b00000000000000001111011101100011;
assign LUT_3[5199] = 32'b00000000000000010110001001000000;
assign LUT_3[5200] = 32'b00000000000000001110000010000110;
assign LUT_3[5201] = 32'b00000000000000010100101101100011;
assign LUT_3[5202] = 32'b00000000000000010000001001101010;
assign LUT_3[5203] = 32'b00000000000000010110110101000111;
assign LUT_3[5204] = 32'b00000000000000001011001111111100;
assign LUT_3[5205] = 32'b00000000000000010001111011011001;
assign LUT_3[5206] = 32'b00000000000000001101010111100000;
assign LUT_3[5207] = 32'b00000000000000010100000010111101;
assign LUT_3[5208] = 32'b00000000000000010011011011001100;
assign LUT_3[5209] = 32'b00000000000000011010000110101001;
assign LUT_3[5210] = 32'b00000000000000010101100010110000;
assign LUT_3[5211] = 32'b00000000000000011100001110001101;
assign LUT_3[5212] = 32'b00000000000000010000101001000010;
assign LUT_3[5213] = 32'b00000000000000010111010100011111;
assign LUT_3[5214] = 32'b00000000000000010010110000100110;
assign LUT_3[5215] = 32'b00000000000000011001011100000011;
assign LUT_3[5216] = 32'b00000000000000001011111101100011;
assign LUT_3[5217] = 32'b00000000000000010010101001000000;
assign LUT_3[5218] = 32'b00000000000000001110000101000111;
assign LUT_3[5219] = 32'b00000000000000010100110000100100;
assign LUT_3[5220] = 32'b00000000000000001001001011011001;
assign LUT_3[5221] = 32'b00000000000000001111110110110110;
assign LUT_3[5222] = 32'b00000000000000001011010010111101;
assign LUT_3[5223] = 32'b00000000000000010001111110011010;
assign LUT_3[5224] = 32'b00000000000000010001010110101001;
assign LUT_3[5225] = 32'b00000000000000011000000010000110;
assign LUT_3[5226] = 32'b00000000000000010011011110001101;
assign LUT_3[5227] = 32'b00000000000000011010001001101010;
assign LUT_3[5228] = 32'b00000000000000001110100100011111;
assign LUT_3[5229] = 32'b00000000000000010101001111111100;
assign LUT_3[5230] = 32'b00000000000000010000101100000011;
assign LUT_3[5231] = 32'b00000000000000010111010111100000;
assign LUT_3[5232] = 32'b00000000000000001111010000100110;
assign LUT_3[5233] = 32'b00000000000000010101111100000011;
assign LUT_3[5234] = 32'b00000000000000010001011000001010;
assign LUT_3[5235] = 32'b00000000000000011000000011100111;
assign LUT_3[5236] = 32'b00000000000000001100011110011100;
assign LUT_3[5237] = 32'b00000000000000010011001001111001;
assign LUT_3[5238] = 32'b00000000000000001110100110000000;
assign LUT_3[5239] = 32'b00000000000000010101010001011101;
assign LUT_3[5240] = 32'b00000000000000010100101001101100;
assign LUT_3[5241] = 32'b00000000000000011011010101001001;
assign LUT_3[5242] = 32'b00000000000000010110110001010000;
assign LUT_3[5243] = 32'b00000000000000011101011100101101;
assign LUT_3[5244] = 32'b00000000000000010001110111100010;
assign LUT_3[5245] = 32'b00000000000000011000100010111111;
assign LUT_3[5246] = 32'b00000000000000010011111111000110;
assign LUT_3[5247] = 32'b00000000000000011010101010100011;
assign LUT_3[5248] = 32'b00000000000000001101000001010110;
assign LUT_3[5249] = 32'b00000000000000010011101100110011;
assign LUT_3[5250] = 32'b00000000000000001111001000111010;
assign LUT_3[5251] = 32'b00000000000000010101110100010111;
assign LUT_3[5252] = 32'b00000000000000001010001111001100;
assign LUT_3[5253] = 32'b00000000000000010000111010101001;
assign LUT_3[5254] = 32'b00000000000000001100010110110000;
assign LUT_3[5255] = 32'b00000000000000010011000010001101;
assign LUT_3[5256] = 32'b00000000000000010010011010011100;
assign LUT_3[5257] = 32'b00000000000000011001000101111001;
assign LUT_3[5258] = 32'b00000000000000010100100010000000;
assign LUT_3[5259] = 32'b00000000000000011011001101011101;
assign LUT_3[5260] = 32'b00000000000000001111101000010010;
assign LUT_3[5261] = 32'b00000000000000010110010011101111;
assign LUT_3[5262] = 32'b00000000000000010001101111110110;
assign LUT_3[5263] = 32'b00000000000000011000011011010011;
assign LUT_3[5264] = 32'b00000000000000010000010100011001;
assign LUT_3[5265] = 32'b00000000000000010110111111110110;
assign LUT_3[5266] = 32'b00000000000000010010011011111101;
assign LUT_3[5267] = 32'b00000000000000011001000111011010;
assign LUT_3[5268] = 32'b00000000000000001101100010001111;
assign LUT_3[5269] = 32'b00000000000000010100001101101100;
assign LUT_3[5270] = 32'b00000000000000001111101001110011;
assign LUT_3[5271] = 32'b00000000000000010110010101010000;
assign LUT_3[5272] = 32'b00000000000000010101101101011111;
assign LUT_3[5273] = 32'b00000000000000011100011000111100;
assign LUT_3[5274] = 32'b00000000000000010111110101000011;
assign LUT_3[5275] = 32'b00000000000000011110100000100000;
assign LUT_3[5276] = 32'b00000000000000010010111011010101;
assign LUT_3[5277] = 32'b00000000000000011001100110110010;
assign LUT_3[5278] = 32'b00000000000000010101000010111001;
assign LUT_3[5279] = 32'b00000000000000011011101110010110;
assign LUT_3[5280] = 32'b00000000000000001110001111110110;
assign LUT_3[5281] = 32'b00000000000000010100111011010011;
assign LUT_3[5282] = 32'b00000000000000010000010111011010;
assign LUT_3[5283] = 32'b00000000000000010111000010110111;
assign LUT_3[5284] = 32'b00000000000000001011011101101100;
assign LUT_3[5285] = 32'b00000000000000010010001001001001;
assign LUT_3[5286] = 32'b00000000000000001101100101010000;
assign LUT_3[5287] = 32'b00000000000000010100010000101101;
assign LUT_3[5288] = 32'b00000000000000010011101000111100;
assign LUT_3[5289] = 32'b00000000000000011010010100011001;
assign LUT_3[5290] = 32'b00000000000000010101110000100000;
assign LUT_3[5291] = 32'b00000000000000011100011011111101;
assign LUT_3[5292] = 32'b00000000000000010000110110110010;
assign LUT_3[5293] = 32'b00000000000000010111100010001111;
assign LUT_3[5294] = 32'b00000000000000010010111110010110;
assign LUT_3[5295] = 32'b00000000000000011001101001110011;
assign LUT_3[5296] = 32'b00000000000000010001100010111001;
assign LUT_3[5297] = 32'b00000000000000011000001110010110;
assign LUT_3[5298] = 32'b00000000000000010011101010011101;
assign LUT_3[5299] = 32'b00000000000000011010010101111010;
assign LUT_3[5300] = 32'b00000000000000001110110000101111;
assign LUT_3[5301] = 32'b00000000000000010101011100001100;
assign LUT_3[5302] = 32'b00000000000000010000111000010011;
assign LUT_3[5303] = 32'b00000000000000010111100011110000;
assign LUT_3[5304] = 32'b00000000000000010110111011111111;
assign LUT_3[5305] = 32'b00000000000000011101100111011100;
assign LUT_3[5306] = 32'b00000000000000011001000011100011;
assign LUT_3[5307] = 32'b00000000000000011111101111000000;
assign LUT_3[5308] = 32'b00000000000000010100001001110101;
assign LUT_3[5309] = 32'b00000000000000011010110101010010;
assign LUT_3[5310] = 32'b00000000000000010110010001011001;
assign LUT_3[5311] = 32'b00000000000000011100111100110110;
assign LUT_3[5312] = 32'b00000000000000001100111010000001;
assign LUT_3[5313] = 32'b00000000000000010011100101011110;
assign LUT_3[5314] = 32'b00000000000000001111000001100101;
assign LUT_3[5315] = 32'b00000000000000010101101101000010;
assign LUT_3[5316] = 32'b00000000000000001010000111110111;
assign LUT_3[5317] = 32'b00000000000000010000110011010100;
assign LUT_3[5318] = 32'b00000000000000001100001111011011;
assign LUT_3[5319] = 32'b00000000000000010010111010111000;
assign LUT_3[5320] = 32'b00000000000000010010010011000111;
assign LUT_3[5321] = 32'b00000000000000011000111110100100;
assign LUT_3[5322] = 32'b00000000000000010100011010101011;
assign LUT_3[5323] = 32'b00000000000000011011000110001000;
assign LUT_3[5324] = 32'b00000000000000001111100000111101;
assign LUT_3[5325] = 32'b00000000000000010110001100011010;
assign LUT_3[5326] = 32'b00000000000000010001101000100001;
assign LUT_3[5327] = 32'b00000000000000011000010011111110;
assign LUT_3[5328] = 32'b00000000000000010000001101000100;
assign LUT_3[5329] = 32'b00000000000000010110111000100001;
assign LUT_3[5330] = 32'b00000000000000010010010100101000;
assign LUT_3[5331] = 32'b00000000000000011001000000000101;
assign LUT_3[5332] = 32'b00000000000000001101011010111010;
assign LUT_3[5333] = 32'b00000000000000010100000110010111;
assign LUT_3[5334] = 32'b00000000000000001111100010011110;
assign LUT_3[5335] = 32'b00000000000000010110001101111011;
assign LUT_3[5336] = 32'b00000000000000010101100110001010;
assign LUT_3[5337] = 32'b00000000000000011100010001100111;
assign LUT_3[5338] = 32'b00000000000000010111101101101110;
assign LUT_3[5339] = 32'b00000000000000011110011001001011;
assign LUT_3[5340] = 32'b00000000000000010010110100000000;
assign LUT_3[5341] = 32'b00000000000000011001011111011101;
assign LUT_3[5342] = 32'b00000000000000010100111011100100;
assign LUT_3[5343] = 32'b00000000000000011011100111000001;
assign LUT_3[5344] = 32'b00000000000000001110001000100001;
assign LUT_3[5345] = 32'b00000000000000010100110011111110;
assign LUT_3[5346] = 32'b00000000000000010000010000000101;
assign LUT_3[5347] = 32'b00000000000000010110111011100010;
assign LUT_3[5348] = 32'b00000000000000001011010110010111;
assign LUT_3[5349] = 32'b00000000000000010010000001110100;
assign LUT_3[5350] = 32'b00000000000000001101011101111011;
assign LUT_3[5351] = 32'b00000000000000010100001001011000;
assign LUT_3[5352] = 32'b00000000000000010011100001100111;
assign LUT_3[5353] = 32'b00000000000000011010001101000100;
assign LUT_3[5354] = 32'b00000000000000010101101001001011;
assign LUT_3[5355] = 32'b00000000000000011100010100101000;
assign LUT_3[5356] = 32'b00000000000000010000101111011101;
assign LUT_3[5357] = 32'b00000000000000010111011010111010;
assign LUT_3[5358] = 32'b00000000000000010010110111000001;
assign LUT_3[5359] = 32'b00000000000000011001100010011110;
assign LUT_3[5360] = 32'b00000000000000010001011011100100;
assign LUT_3[5361] = 32'b00000000000000011000000111000001;
assign LUT_3[5362] = 32'b00000000000000010011100011001000;
assign LUT_3[5363] = 32'b00000000000000011010001110100101;
assign LUT_3[5364] = 32'b00000000000000001110101001011010;
assign LUT_3[5365] = 32'b00000000000000010101010100110111;
assign LUT_3[5366] = 32'b00000000000000010000110000111110;
assign LUT_3[5367] = 32'b00000000000000010111011100011011;
assign LUT_3[5368] = 32'b00000000000000010110110100101010;
assign LUT_3[5369] = 32'b00000000000000011101100000000111;
assign LUT_3[5370] = 32'b00000000000000011000111100001110;
assign LUT_3[5371] = 32'b00000000000000011111100111101011;
assign LUT_3[5372] = 32'b00000000000000010100000010100000;
assign LUT_3[5373] = 32'b00000000000000011010101101111101;
assign LUT_3[5374] = 32'b00000000000000010110001010000100;
assign LUT_3[5375] = 32'b00000000000000011100110101100001;
assign LUT_3[5376] = 32'b00000000000000000111000101111001;
assign LUT_3[5377] = 32'b00000000000000001101110001010110;
assign LUT_3[5378] = 32'b00000000000000001001001101011101;
assign LUT_3[5379] = 32'b00000000000000001111111000111010;
assign LUT_3[5380] = 32'b00000000000000000100010011101111;
assign LUT_3[5381] = 32'b00000000000000001010111111001100;
assign LUT_3[5382] = 32'b00000000000000000110011011010011;
assign LUT_3[5383] = 32'b00000000000000001101000110110000;
assign LUT_3[5384] = 32'b00000000000000001100011110111111;
assign LUT_3[5385] = 32'b00000000000000010011001010011100;
assign LUT_3[5386] = 32'b00000000000000001110100110100011;
assign LUT_3[5387] = 32'b00000000000000010101010010000000;
assign LUT_3[5388] = 32'b00000000000000001001101100110101;
assign LUT_3[5389] = 32'b00000000000000010000011000010010;
assign LUT_3[5390] = 32'b00000000000000001011110100011001;
assign LUT_3[5391] = 32'b00000000000000010010011111110110;
assign LUT_3[5392] = 32'b00000000000000001010011000111100;
assign LUT_3[5393] = 32'b00000000000000010001000100011001;
assign LUT_3[5394] = 32'b00000000000000001100100000100000;
assign LUT_3[5395] = 32'b00000000000000010011001011111101;
assign LUT_3[5396] = 32'b00000000000000000111100110110010;
assign LUT_3[5397] = 32'b00000000000000001110010010001111;
assign LUT_3[5398] = 32'b00000000000000001001101110010110;
assign LUT_3[5399] = 32'b00000000000000010000011001110011;
assign LUT_3[5400] = 32'b00000000000000001111110010000010;
assign LUT_3[5401] = 32'b00000000000000010110011101011111;
assign LUT_3[5402] = 32'b00000000000000010001111001100110;
assign LUT_3[5403] = 32'b00000000000000011000100101000011;
assign LUT_3[5404] = 32'b00000000000000001100111111111000;
assign LUT_3[5405] = 32'b00000000000000010011101011010101;
assign LUT_3[5406] = 32'b00000000000000001111000111011100;
assign LUT_3[5407] = 32'b00000000000000010101110010111001;
assign LUT_3[5408] = 32'b00000000000000001000010100011001;
assign LUT_3[5409] = 32'b00000000000000001110111111110110;
assign LUT_3[5410] = 32'b00000000000000001010011011111101;
assign LUT_3[5411] = 32'b00000000000000010001000111011010;
assign LUT_3[5412] = 32'b00000000000000000101100010001111;
assign LUT_3[5413] = 32'b00000000000000001100001101101100;
assign LUT_3[5414] = 32'b00000000000000000111101001110011;
assign LUT_3[5415] = 32'b00000000000000001110010101010000;
assign LUT_3[5416] = 32'b00000000000000001101101101011111;
assign LUT_3[5417] = 32'b00000000000000010100011000111100;
assign LUT_3[5418] = 32'b00000000000000001111110101000011;
assign LUT_3[5419] = 32'b00000000000000010110100000100000;
assign LUT_3[5420] = 32'b00000000000000001010111011010101;
assign LUT_3[5421] = 32'b00000000000000010001100110110010;
assign LUT_3[5422] = 32'b00000000000000001101000010111001;
assign LUT_3[5423] = 32'b00000000000000010011101110010110;
assign LUT_3[5424] = 32'b00000000000000001011100111011100;
assign LUT_3[5425] = 32'b00000000000000010010010010111001;
assign LUT_3[5426] = 32'b00000000000000001101101111000000;
assign LUT_3[5427] = 32'b00000000000000010100011010011101;
assign LUT_3[5428] = 32'b00000000000000001000110101010010;
assign LUT_3[5429] = 32'b00000000000000001111100000101111;
assign LUT_3[5430] = 32'b00000000000000001010111100110110;
assign LUT_3[5431] = 32'b00000000000000010001101000010011;
assign LUT_3[5432] = 32'b00000000000000010001000000100010;
assign LUT_3[5433] = 32'b00000000000000010111101011111111;
assign LUT_3[5434] = 32'b00000000000000010011001000000110;
assign LUT_3[5435] = 32'b00000000000000011001110011100011;
assign LUT_3[5436] = 32'b00000000000000001110001110011000;
assign LUT_3[5437] = 32'b00000000000000010100111001110101;
assign LUT_3[5438] = 32'b00000000000000010000010101111100;
assign LUT_3[5439] = 32'b00000000000000010111000001011001;
assign LUT_3[5440] = 32'b00000000000000000110111110100100;
assign LUT_3[5441] = 32'b00000000000000001101101010000001;
assign LUT_3[5442] = 32'b00000000000000001001000110001000;
assign LUT_3[5443] = 32'b00000000000000001111110001100101;
assign LUT_3[5444] = 32'b00000000000000000100001100011010;
assign LUT_3[5445] = 32'b00000000000000001010110111110111;
assign LUT_3[5446] = 32'b00000000000000000110010011111110;
assign LUT_3[5447] = 32'b00000000000000001100111111011011;
assign LUT_3[5448] = 32'b00000000000000001100010111101010;
assign LUT_3[5449] = 32'b00000000000000010011000011000111;
assign LUT_3[5450] = 32'b00000000000000001110011111001110;
assign LUT_3[5451] = 32'b00000000000000010101001010101011;
assign LUT_3[5452] = 32'b00000000000000001001100101100000;
assign LUT_3[5453] = 32'b00000000000000010000010000111101;
assign LUT_3[5454] = 32'b00000000000000001011101101000100;
assign LUT_3[5455] = 32'b00000000000000010010011000100001;
assign LUT_3[5456] = 32'b00000000000000001010010001100111;
assign LUT_3[5457] = 32'b00000000000000010000111101000100;
assign LUT_3[5458] = 32'b00000000000000001100011001001011;
assign LUT_3[5459] = 32'b00000000000000010011000100101000;
assign LUT_3[5460] = 32'b00000000000000000111011111011101;
assign LUT_3[5461] = 32'b00000000000000001110001010111010;
assign LUT_3[5462] = 32'b00000000000000001001100111000001;
assign LUT_3[5463] = 32'b00000000000000010000010010011110;
assign LUT_3[5464] = 32'b00000000000000001111101010101101;
assign LUT_3[5465] = 32'b00000000000000010110010110001010;
assign LUT_3[5466] = 32'b00000000000000010001110010010001;
assign LUT_3[5467] = 32'b00000000000000011000011101101110;
assign LUT_3[5468] = 32'b00000000000000001100111000100011;
assign LUT_3[5469] = 32'b00000000000000010011100100000000;
assign LUT_3[5470] = 32'b00000000000000001111000000000111;
assign LUT_3[5471] = 32'b00000000000000010101101011100100;
assign LUT_3[5472] = 32'b00000000000000001000001101000100;
assign LUT_3[5473] = 32'b00000000000000001110111000100001;
assign LUT_3[5474] = 32'b00000000000000001010010100101000;
assign LUT_3[5475] = 32'b00000000000000010001000000000101;
assign LUT_3[5476] = 32'b00000000000000000101011010111010;
assign LUT_3[5477] = 32'b00000000000000001100000110010111;
assign LUT_3[5478] = 32'b00000000000000000111100010011110;
assign LUT_3[5479] = 32'b00000000000000001110001101111011;
assign LUT_3[5480] = 32'b00000000000000001101100110001010;
assign LUT_3[5481] = 32'b00000000000000010100010001100111;
assign LUT_3[5482] = 32'b00000000000000001111101101101110;
assign LUT_3[5483] = 32'b00000000000000010110011001001011;
assign LUT_3[5484] = 32'b00000000000000001010110100000000;
assign LUT_3[5485] = 32'b00000000000000010001011111011101;
assign LUT_3[5486] = 32'b00000000000000001100111011100100;
assign LUT_3[5487] = 32'b00000000000000010011100111000001;
assign LUT_3[5488] = 32'b00000000000000001011100000000111;
assign LUT_3[5489] = 32'b00000000000000010010001011100100;
assign LUT_3[5490] = 32'b00000000000000001101100111101011;
assign LUT_3[5491] = 32'b00000000000000010100010011001000;
assign LUT_3[5492] = 32'b00000000000000001000101101111101;
assign LUT_3[5493] = 32'b00000000000000001111011001011010;
assign LUT_3[5494] = 32'b00000000000000001010110101100001;
assign LUT_3[5495] = 32'b00000000000000010001100000111110;
assign LUT_3[5496] = 32'b00000000000000010000111001001101;
assign LUT_3[5497] = 32'b00000000000000010111100100101010;
assign LUT_3[5498] = 32'b00000000000000010011000000110001;
assign LUT_3[5499] = 32'b00000000000000011001101100001110;
assign LUT_3[5500] = 32'b00000000000000001110000111000011;
assign LUT_3[5501] = 32'b00000000000000010100110010100000;
assign LUT_3[5502] = 32'b00000000000000010000001110100111;
assign LUT_3[5503] = 32'b00000000000000010110111010000100;
assign LUT_3[5504] = 32'b00000000000000001001010000110111;
assign LUT_3[5505] = 32'b00000000000000001111111100010100;
assign LUT_3[5506] = 32'b00000000000000001011011000011011;
assign LUT_3[5507] = 32'b00000000000000010010000011111000;
assign LUT_3[5508] = 32'b00000000000000000110011110101101;
assign LUT_3[5509] = 32'b00000000000000001101001010001010;
assign LUT_3[5510] = 32'b00000000000000001000100110010001;
assign LUT_3[5511] = 32'b00000000000000001111010001101110;
assign LUT_3[5512] = 32'b00000000000000001110101001111101;
assign LUT_3[5513] = 32'b00000000000000010101010101011010;
assign LUT_3[5514] = 32'b00000000000000010000110001100001;
assign LUT_3[5515] = 32'b00000000000000010111011100111110;
assign LUT_3[5516] = 32'b00000000000000001011110111110011;
assign LUT_3[5517] = 32'b00000000000000010010100011010000;
assign LUT_3[5518] = 32'b00000000000000001101111111010111;
assign LUT_3[5519] = 32'b00000000000000010100101010110100;
assign LUT_3[5520] = 32'b00000000000000001100100011111010;
assign LUT_3[5521] = 32'b00000000000000010011001111010111;
assign LUT_3[5522] = 32'b00000000000000001110101011011110;
assign LUT_3[5523] = 32'b00000000000000010101010110111011;
assign LUT_3[5524] = 32'b00000000000000001001110001110000;
assign LUT_3[5525] = 32'b00000000000000010000011101001101;
assign LUT_3[5526] = 32'b00000000000000001011111001010100;
assign LUT_3[5527] = 32'b00000000000000010010100100110001;
assign LUT_3[5528] = 32'b00000000000000010001111101000000;
assign LUT_3[5529] = 32'b00000000000000011000101000011101;
assign LUT_3[5530] = 32'b00000000000000010100000100100100;
assign LUT_3[5531] = 32'b00000000000000011010110000000001;
assign LUT_3[5532] = 32'b00000000000000001111001010110110;
assign LUT_3[5533] = 32'b00000000000000010101110110010011;
assign LUT_3[5534] = 32'b00000000000000010001010010011010;
assign LUT_3[5535] = 32'b00000000000000010111111101110111;
assign LUT_3[5536] = 32'b00000000000000001010011111010111;
assign LUT_3[5537] = 32'b00000000000000010001001010110100;
assign LUT_3[5538] = 32'b00000000000000001100100110111011;
assign LUT_3[5539] = 32'b00000000000000010011010010011000;
assign LUT_3[5540] = 32'b00000000000000000111101101001101;
assign LUT_3[5541] = 32'b00000000000000001110011000101010;
assign LUT_3[5542] = 32'b00000000000000001001110100110001;
assign LUT_3[5543] = 32'b00000000000000010000100000001110;
assign LUT_3[5544] = 32'b00000000000000001111111000011101;
assign LUT_3[5545] = 32'b00000000000000010110100011111010;
assign LUT_3[5546] = 32'b00000000000000010010000000000001;
assign LUT_3[5547] = 32'b00000000000000011000101011011110;
assign LUT_3[5548] = 32'b00000000000000001101000110010011;
assign LUT_3[5549] = 32'b00000000000000010011110001110000;
assign LUT_3[5550] = 32'b00000000000000001111001101110111;
assign LUT_3[5551] = 32'b00000000000000010101111001010100;
assign LUT_3[5552] = 32'b00000000000000001101110010011010;
assign LUT_3[5553] = 32'b00000000000000010100011101110111;
assign LUT_3[5554] = 32'b00000000000000001111111001111110;
assign LUT_3[5555] = 32'b00000000000000010110100101011011;
assign LUT_3[5556] = 32'b00000000000000001011000000010000;
assign LUT_3[5557] = 32'b00000000000000010001101011101101;
assign LUT_3[5558] = 32'b00000000000000001101000111110100;
assign LUT_3[5559] = 32'b00000000000000010011110011010001;
assign LUT_3[5560] = 32'b00000000000000010011001011100000;
assign LUT_3[5561] = 32'b00000000000000011001110110111101;
assign LUT_3[5562] = 32'b00000000000000010101010011000100;
assign LUT_3[5563] = 32'b00000000000000011011111110100001;
assign LUT_3[5564] = 32'b00000000000000010000011001010110;
assign LUT_3[5565] = 32'b00000000000000010111000100110011;
assign LUT_3[5566] = 32'b00000000000000010010100000111010;
assign LUT_3[5567] = 32'b00000000000000011001001100010111;
assign LUT_3[5568] = 32'b00000000000000001001001001100010;
assign LUT_3[5569] = 32'b00000000000000001111110100111111;
assign LUT_3[5570] = 32'b00000000000000001011010001000110;
assign LUT_3[5571] = 32'b00000000000000010001111100100011;
assign LUT_3[5572] = 32'b00000000000000000110010111011000;
assign LUT_3[5573] = 32'b00000000000000001101000010110101;
assign LUT_3[5574] = 32'b00000000000000001000011110111100;
assign LUT_3[5575] = 32'b00000000000000001111001010011001;
assign LUT_3[5576] = 32'b00000000000000001110100010101000;
assign LUT_3[5577] = 32'b00000000000000010101001110000101;
assign LUT_3[5578] = 32'b00000000000000010000101010001100;
assign LUT_3[5579] = 32'b00000000000000010111010101101001;
assign LUT_3[5580] = 32'b00000000000000001011110000011110;
assign LUT_3[5581] = 32'b00000000000000010010011011111011;
assign LUT_3[5582] = 32'b00000000000000001101111000000010;
assign LUT_3[5583] = 32'b00000000000000010100100011011111;
assign LUT_3[5584] = 32'b00000000000000001100011100100101;
assign LUT_3[5585] = 32'b00000000000000010011001000000010;
assign LUT_3[5586] = 32'b00000000000000001110100100001001;
assign LUT_3[5587] = 32'b00000000000000010101001111100110;
assign LUT_3[5588] = 32'b00000000000000001001101010011011;
assign LUT_3[5589] = 32'b00000000000000010000010101111000;
assign LUT_3[5590] = 32'b00000000000000001011110001111111;
assign LUT_3[5591] = 32'b00000000000000010010011101011100;
assign LUT_3[5592] = 32'b00000000000000010001110101101011;
assign LUT_3[5593] = 32'b00000000000000011000100001001000;
assign LUT_3[5594] = 32'b00000000000000010011111101001111;
assign LUT_3[5595] = 32'b00000000000000011010101000101100;
assign LUT_3[5596] = 32'b00000000000000001111000011100001;
assign LUT_3[5597] = 32'b00000000000000010101101110111110;
assign LUT_3[5598] = 32'b00000000000000010001001011000101;
assign LUT_3[5599] = 32'b00000000000000010111110110100010;
assign LUT_3[5600] = 32'b00000000000000001010011000000010;
assign LUT_3[5601] = 32'b00000000000000010001000011011111;
assign LUT_3[5602] = 32'b00000000000000001100011111100110;
assign LUT_3[5603] = 32'b00000000000000010011001011000011;
assign LUT_3[5604] = 32'b00000000000000000111100101111000;
assign LUT_3[5605] = 32'b00000000000000001110010001010101;
assign LUT_3[5606] = 32'b00000000000000001001101101011100;
assign LUT_3[5607] = 32'b00000000000000010000011000111001;
assign LUT_3[5608] = 32'b00000000000000001111110001001000;
assign LUT_3[5609] = 32'b00000000000000010110011100100101;
assign LUT_3[5610] = 32'b00000000000000010001111000101100;
assign LUT_3[5611] = 32'b00000000000000011000100100001001;
assign LUT_3[5612] = 32'b00000000000000001100111110111110;
assign LUT_3[5613] = 32'b00000000000000010011101010011011;
assign LUT_3[5614] = 32'b00000000000000001111000110100010;
assign LUT_3[5615] = 32'b00000000000000010101110001111111;
assign LUT_3[5616] = 32'b00000000000000001101101011000101;
assign LUT_3[5617] = 32'b00000000000000010100010110100010;
assign LUT_3[5618] = 32'b00000000000000001111110010101001;
assign LUT_3[5619] = 32'b00000000000000010110011110000110;
assign LUT_3[5620] = 32'b00000000000000001010111000111011;
assign LUT_3[5621] = 32'b00000000000000010001100100011000;
assign LUT_3[5622] = 32'b00000000000000001101000000011111;
assign LUT_3[5623] = 32'b00000000000000010011101011111100;
assign LUT_3[5624] = 32'b00000000000000010011000100001011;
assign LUT_3[5625] = 32'b00000000000000011001101111101000;
assign LUT_3[5626] = 32'b00000000000000010101001011101111;
assign LUT_3[5627] = 32'b00000000000000011011110111001100;
assign LUT_3[5628] = 32'b00000000000000010000010010000001;
assign LUT_3[5629] = 32'b00000000000000010110111101011110;
assign LUT_3[5630] = 32'b00000000000000010010011001100101;
assign LUT_3[5631] = 32'b00000000000000011001000101000010;
assign LUT_3[5632] = 32'b00000000000000001110001011100100;
assign LUT_3[5633] = 32'b00000000000000010100110111000001;
assign LUT_3[5634] = 32'b00000000000000010000010011001000;
assign LUT_3[5635] = 32'b00000000000000010110111110100101;
assign LUT_3[5636] = 32'b00000000000000001011011001011010;
assign LUT_3[5637] = 32'b00000000000000010010000100110111;
assign LUT_3[5638] = 32'b00000000000000001101100000111110;
assign LUT_3[5639] = 32'b00000000000000010100001100011011;
assign LUT_3[5640] = 32'b00000000000000010011100100101010;
assign LUT_3[5641] = 32'b00000000000000011010010000000111;
assign LUT_3[5642] = 32'b00000000000000010101101100001110;
assign LUT_3[5643] = 32'b00000000000000011100010111101011;
assign LUT_3[5644] = 32'b00000000000000010000110010100000;
assign LUT_3[5645] = 32'b00000000000000010111011101111101;
assign LUT_3[5646] = 32'b00000000000000010010111010000100;
assign LUT_3[5647] = 32'b00000000000000011001100101100001;
assign LUT_3[5648] = 32'b00000000000000010001011110100111;
assign LUT_3[5649] = 32'b00000000000000011000001010000100;
assign LUT_3[5650] = 32'b00000000000000010011100110001011;
assign LUT_3[5651] = 32'b00000000000000011010010001101000;
assign LUT_3[5652] = 32'b00000000000000001110101100011101;
assign LUT_3[5653] = 32'b00000000000000010101010111111010;
assign LUT_3[5654] = 32'b00000000000000010000110100000001;
assign LUT_3[5655] = 32'b00000000000000010111011111011110;
assign LUT_3[5656] = 32'b00000000000000010110110111101101;
assign LUT_3[5657] = 32'b00000000000000011101100011001010;
assign LUT_3[5658] = 32'b00000000000000011000111111010001;
assign LUT_3[5659] = 32'b00000000000000011111101010101110;
assign LUT_3[5660] = 32'b00000000000000010100000101100011;
assign LUT_3[5661] = 32'b00000000000000011010110001000000;
assign LUT_3[5662] = 32'b00000000000000010110001101000111;
assign LUT_3[5663] = 32'b00000000000000011100111000100100;
assign LUT_3[5664] = 32'b00000000000000001111011010000100;
assign LUT_3[5665] = 32'b00000000000000010110000101100001;
assign LUT_3[5666] = 32'b00000000000000010001100001101000;
assign LUT_3[5667] = 32'b00000000000000011000001101000101;
assign LUT_3[5668] = 32'b00000000000000001100100111111010;
assign LUT_3[5669] = 32'b00000000000000010011010011010111;
assign LUT_3[5670] = 32'b00000000000000001110101111011110;
assign LUT_3[5671] = 32'b00000000000000010101011010111011;
assign LUT_3[5672] = 32'b00000000000000010100110011001010;
assign LUT_3[5673] = 32'b00000000000000011011011110100111;
assign LUT_3[5674] = 32'b00000000000000010110111010101110;
assign LUT_3[5675] = 32'b00000000000000011101100110001011;
assign LUT_3[5676] = 32'b00000000000000010010000001000000;
assign LUT_3[5677] = 32'b00000000000000011000101100011101;
assign LUT_3[5678] = 32'b00000000000000010100001000100100;
assign LUT_3[5679] = 32'b00000000000000011010110100000001;
assign LUT_3[5680] = 32'b00000000000000010010101101000111;
assign LUT_3[5681] = 32'b00000000000000011001011000100100;
assign LUT_3[5682] = 32'b00000000000000010100110100101011;
assign LUT_3[5683] = 32'b00000000000000011011100000001000;
assign LUT_3[5684] = 32'b00000000000000001111111010111101;
assign LUT_3[5685] = 32'b00000000000000010110100110011010;
assign LUT_3[5686] = 32'b00000000000000010010000010100001;
assign LUT_3[5687] = 32'b00000000000000011000101101111110;
assign LUT_3[5688] = 32'b00000000000000011000000110001101;
assign LUT_3[5689] = 32'b00000000000000011110110001101010;
assign LUT_3[5690] = 32'b00000000000000011010001101110001;
assign LUT_3[5691] = 32'b00000000000000100000111001001110;
assign LUT_3[5692] = 32'b00000000000000010101010100000011;
assign LUT_3[5693] = 32'b00000000000000011011111111100000;
assign LUT_3[5694] = 32'b00000000000000010111011011100111;
assign LUT_3[5695] = 32'b00000000000000011110000111000100;
assign LUT_3[5696] = 32'b00000000000000001110000100001111;
assign LUT_3[5697] = 32'b00000000000000010100101111101100;
assign LUT_3[5698] = 32'b00000000000000010000001011110011;
assign LUT_3[5699] = 32'b00000000000000010110110111010000;
assign LUT_3[5700] = 32'b00000000000000001011010010000101;
assign LUT_3[5701] = 32'b00000000000000010001111101100010;
assign LUT_3[5702] = 32'b00000000000000001101011001101001;
assign LUT_3[5703] = 32'b00000000000000010100000101000110;
assign LUT_3[5704] = 32'b00000000000000010011011101010101;
assign LUT_3[5705] = 32'b00000000000000011010001000110010;
assign LUT_3[5706] = 32'b00000000000000010101100100111001;
assign LUT_3[5707] = 32'b00000000000000011100010000010110;
assign LUT_3[5708] = 32'b00000000000000010000101011001011;
assign LUT_3[5709] = 32'b00000000000000010111010110101000;
assign LUT_3[5710] = 32'b00000000000000010010110010101111;
assign LUT_3[5711] = 32'b00000000000000011001011110001100;
assign LUT_3[5712] = 32'b00000000000000010001010111010010;
assign LUT_3[5713] = 32'b00000000000000011000000010101111;
assign LUT_3[5714] = 32'b00000000000000010011011110110110;
assign LUT_3[5715] = 32'b00000000000000011010001010010011;
assign LUT_3[5716] = 32'b00000000000000001110100101001000;
assign LUT_3[5717] = 32'b00000000000000010101010000100101;
assign LUT_3[5718] = 32'b00000000000000010000101100101100;
assign LUT_3[5719] = 32'b00000000000000010111011000001001;
assign LUT_3[5720] = 32'b00000000000000010110110000011000;
assign LUT_3[5721] = 32'b00000000000000011101011011110101;
assign LUT_3[5722] = 32'b00000000000000011000110111111100;
assign LUT_3[5723] = 32'b00000000000000011111100011011001;
assign LUT_3[5724] = 32'b00000000000000010011111110001110;
assign LUT_3[5725] = 32'b00000000000000011010101001101011;
assign LUT_3[5726] = 32'b00000000000000010110000101110010;
assign LUT_3[5727] = 32'b00000000000000011100110001001111;
assign LUT_3[5728] = 32'b00000000000000001111010010101111;
assign LUT_3[5729] = 32'b00000000000000010101111110001100;
assign LUT_3[5730] = 32'b00000000000000010001011010010011;
assign LUT_3[5731] = 32'b00000000000000011000000101110000;
assign LUT_3[5732] = 32'b00000000000000001100100000100101;
assign LUT_3[5733] = 32'b00000000000000010011001100000010;
assign LUT_3[5734] = 32'b00000000000000001110101000001001;
assign LUT_3[5735] = 32'b00000000000000010101010011100110;
assign LUT_3[5736] = 32'b00000000000000010100101011110101;
assign LUT_3[5737] = 32'b00000000000000011011010111010010;
assign LUT_3[5738] = 32'b00000000000000010110110011011001;
assign LUT_3[5739] = 32'b00000000000000011101011110110110;
assign LUT_3[5740] = 32'b00000000000000010001111001101011;
assign LUT_3[5741] = 32'b00000000000000011000100101001000;
assign LUT_3[5742] = 32'b00000000000000010100000001001111;
assign LUT_3[5743] = 32'b00000000000000011010101100101100;
assign LUT_3[5744] = 32'b00000000000000010010100101110010;
assign LUT_3[5745] = 32'b00000000000000011001010001001111;
assign LUT_3[5746] = 32'b00000000000000010100101101010110;
assign LUT_3[5747] = 32'b00000000000000011011011000110011;
assign LUT_3[5748] = 32'b00000000000000001111110011101000;
assign LUT_3[5749] = 32'b00000000000000010110011111000101;
assign LUT_3[5750] = 32'b00000000000000010001111011001100;
assign LUT_3[5751] = 32'b00000000000000011000100110101001;
assign LUT_3[5752] = 32'b00000000000000010111111110111000;
assign LUT_3[5753] = 32'b00000000000000011110101010010101;
assign LUT_3[5754] = 32'b00000000000000011010000110011100;
assign LUT_3[5755] = 32'b00000000000000100000110001111001;
assign LUT_3[5756] = 32'b00000000000000010101001100101110;
assign LUT_3[5757] = 32'b00000000000000011011111000001011;
assign LUT_3[5758] = 32'b00000000000000010111010100010010;
assign LUT_3[5759] = 32'b00000000000000011101111111101111;
assign LUT_3[5760] = 32'b00000000000000010000010110100010;
assign LUT_3[5761] = 32'b00000000000000010111000001111111;
assign LUT_3[5762] = 32'b00000000000000010010011110000110;
assign LUT_3[5763] = 32'b00000000000000011001001001100011;
assign LUT_3[5764] = 32'b00000000000000001101100100011000;
assign LUT_3[5765] = 32'b00000000000000010100001111110101;
assign LUT_3[5766] = 32'b00000000000000001111101011111100;
assign LUT_3[5767] = 32'b00000000000000010110010111011001;
assign LUT_3[5768] = 32'b00000000000000010101101111101000;
assign LUT_3[5769] = 32'b00000000000000011100011011000101;
assign LUT_3[5770] = 32'b00000000000000010111110111001100;
assign LUT_3[5771] = 32'b00000000000000011110100010101001;
assign LUT_3[5772] = 32'b00000000000000010010111101011110;
assign LUT_3[5773] = 32'b00000000000000011001101000111011;
assign LUT_3[5774] = 32'b00000000000000010101000101000010;
assign LUT_3[5775] = 32'b00000000000000011011110000011111;
assign LUT_3[5776] = 32'b00000000000000010011101001100101;
assign LUT_3[5777] = 32'b00000000000000011010010101000010;
assign LUT_3[5778] = 32'b00000000000000010101110001001001;
assign LUT_3[5779] = 32'b00000000000000011100011100100110;
assign LUT_3[5780] = 32'b00000000000000010000110111011011;
assign LUT_3[5781] = 32'b00000000000000010111100010111000;
assign LUT_3[5782] = 32'b00000000000000010010111110111111;
assign LUT_3[5783] = 32'b00000000000000011001101010011100;
assign LUT_3[5784] = 32'b00000000000000011001000010101011;
assign LUT_3[5785] = 32'b00000000000000011111101110001000;
assign LUT_3[5786] = 32'b00000000000000011011001010001111;
assign LUT_3[5787] = 32'b00000000000000100001110101101100;
assign LUT_3[5788] = 32'b00000000000000010110010000100001;
assign LUT_3[5789] = 32'b00000000000000011100111011111110;
assign LUT_3[5790] = 32'b00000000000000011000011000000101;
assign LUT_3[5791] = 32'b00000000000000011111000011100010;
assign LUT_3[5792] = 32'b00000000000000010001100101000010;
assign LUT_3[5793] = 32'b00000000000000011000010000011111;
assign LUT_3[5794] = 32'b00000000000000010011101100100110;
assign LUT_3[5795] = 32'b00000000000000011010011000000011;
assign LUT_3[5796] = 32'b00000000000000001110110010111000;
assign LUT_3[5797] = 32'b00000000000000010101011110010101;
assign LUT_3[5798] = 32'b00000000000000010000111010011100;
assign LUT_3[5799] = 32'b00000000000000010111100101111001;
assign LUT_3[5800] = 32'b00000000000000010110111110001000;
assign LUT_3[5801] = 32'b00000000000000011101101001100101;
assign LUT_3[5802] = 32'b00000000000000011001000101101100;
assign LUT_3[5803] = 32'b00000000000000011111110001001001;
assign LUT_3[5804] = 32'b00000000000000010100001011111110;
assign LUT_3[5805] = 32'b00000000000000011010110111011011;
assign LUT_3[5806] = 32'b00000000000000010110010011100010;
assign LUT_3[5807] = 32'b00000000000000011100111110111111;
assign LUT_3[5808] = 32'b00000000000000010100111000000101;
assign LUT_3[5809] = 32'b00000000000000011011100011100010;
assign LUT_3[5810] = 32'b00000000000000010110111111101001;
assign LUT_3[5811] = 32'b00000000000000011101101011000110;
assign LUT_3[5812] = 32'b00000000000000010010000101111011;
assign LUT_3[5813] = 32'b00000000000000011000110001011000;
assign LUT_3[5814] = 32'b00000000000000010100001101011111;
assign LUT_3[5815] = 32'b00000000000000011010111000111100;
assign LUT_3[5816] = 32'b00000000000000011010010001001011;
assign LUT_3[5817] = 32'b00000000000000100000111100101000;
assign LUT_3[5818] = 32'b00000000000000011100011000101111;
assign LUT_3[5819] = 32'b00000000000000100011000100001100;
assign LUT_3[5820] = 32'b00000000000000010111011111000001;
assign LUT_3[5821] = 32'b00000000000000011110001010011110;
assign LUT_3[5822] = 32'b00000000000000011001100110100101;
assign LUT_3[5823] = 32'b00000000000000100000010010000010;
assign LUT_3[5824] = 32'b00000000000000010000001111001101;
assign LUT_3[5825] = 32'b00000000000000010110111010101010;
assign LUT_3[5826] = 32'b00000000000000010010010110110001;
assign LUT_3[5827] = 32'b00000000000000011001000010001110;
assign LUT_3[5828] = 32'b00000000000000001101011101000011;
assign LUT_3[5829] = 32'b00000000000000010100001000100000;
assign LUT_3[5830] = 32'b00000000000000001111100100100111;
assign LUT_3[5831] = 32'b00000000000000010110010000000100;
assign LUT_3[5832] = 32'b00000000000000010101101000010011;
assign LUT_3[5833] = 32'b00000000000000011100010011110000;
assign LUT_3[5834] = 32'b00000000000000010111101111110111;
assign LUT_3[5835] = 32'b00000000000000011110011011010100;
assign LUT_3[5836] = 32'b00000000000000010010110110001001;
assign LUT_3[5837] = 32'b00000000000000011001100001100110;
assign LUT_3[5838] = 32'b00000000000000010100111101101101;
assign LUT_3[5839] = 32'b00000000000000011011101001001010;
assign LUT_3[5840] = 32'b00000000000000010011100010010000;
assign LUT_3[5841] = 32'b00000000000000011010001101101101;
assign LUT_3[5842] = 32'b00000000000000010101101001110100;
assign LUT_3[5843] = 32'b00000000000000011100010101010001;
assign LUT_3[5844] = 32'b00000000000000010000110000000110;
assign LUT_3[5845] = 32'b00000000000000010111011011100011;
assign LUT_3[5846] = 32'b00000000000000010010110111101010;
assign LUT_3[5847] = 32'b00000000000000011001100011000111;
assign LUT_3[5848] = 32'b00000000000000011000111011010110;
assign LUT_3[5849] = 32'b00000000000000011111100110110011;
assign LUT_3[5850] = 32'b00000000000000011011000010111010;
assign LUT_3[5851] = 32'b00000000000000100001101110010111;
assign LUT_3[5852] = 32'b00000000000000010110001001001100;
assign LUT_3[5853] = 32'b00000000000000011100110100101001;
assign LUT_3[5854] = 32'b00000000000000011000010000110000;
assign LUT_3[5855] = 32'b00000000000000011110111100001101;
assign LUT_3[5856] = 32'b00000000000000010001011101101101;
assign LUT_3[5857] = 32'b00000000000000011000001001001010;
assign LUT_3[5858] = 32'b00000000000000010011100101010001;
assign LUT_3[5859] = 32'b00000000000000011010010000101110;
assign LUT_3[5860] = 32'b00000000000000001110101011100011;
assign LUT_3[5861] = 32'b00000000000000010101010111000000;
assign LUT_3[5862] = 32'b00000000000000010000110011000111;
assign LUT_3[5863] = 32'b00000000000000010111011110100100;
assign LUT_3[5864] = 32'b00000000000000010110110110110011;
assign LUT_3[5865] = 32'b00000000000000011101100010010000;
assign LUT_3[5866] = 32'b00000000000000011000111110010111;
assign LUT_3[5867] = 32'b00000000000000011111101001110100;
assign LUT_3[5868] = 32'b00000000000000010100000100101001;
assign LUT_3[5869] = 32'b00000000000000011010110000000110;
assign LUT_3[5870] = 32'b00000000000000010110001100001101;
assign LUT_3[5871] = 32'b00000000000000011100110111101010;
assign LUT_3[5872] = 32'b00000000000000010100110000110000;
assign LUT_3[5873] = 32'b00000000000000011011011100001101;
assign LUT_3[5874] = 32'b00000000000000010110111000010100;
assign LUT_3[5875] = 32'b00000000000000011101100011110001;
assign LUT_3[5876] = 32'b00000000000000010001111110100110;
assign LUT_3[5877] = 32'b00000000000000011000101010000011;
assign LUT_3[5878] = 32'b00000000000000010100000110001010;
assign LUT_3[5879] = 32'b00000000000000011010110001100111;
assign LUT_3[5880] = 32'b00000000000000011010001001110110;
assign LUT_3[5881] = 32'b00000000000000100000110101010011;
assign LUT_3[5882] = 32'b00000000000000011100010001011010;
assign LUT_3[5883] = 32'b00000000000000100010111100110111;
assign LUT_3[5884] = 32'b00000000000000010111010111101100;
assign LUT_3[5885] = 32'b00000000000000011110000011001001;
assign LUT_3[5886] = 32'b00000000000000011001011111010000;
assign LUT_3[5887] = 32'b00000000000000100000001010101101;
assign LUT_3[5888] = 32'b00000000000000001010011011000101;
assign LUT_3[5889] = 32'b00000000000000010001000110100010;
assign LUT_3[5890] = 32'b00000000000000001100100010101001;
assign LUT_3[5891] = 32'b00000000000000010011001110000110;
assign LUT_3[5892] = 32'b00000000000000000111101000111011;
assign LUT_3[5893] = 32'b00000000000000001110010100011000;
assign LUT_3[5894] = 32'b00000000000000001001110000011111;
assign LUT_3[5895] = 32'b00000000000000010000011011111100;
assign LUT_3[5896] = 32'b00000000000000001111110100001011;
assign LUT_3[5897] = 32'b00000000000000010110011111101000;
assign LUT_3[5898] = 32'b00000000000000010001111011101111;
assign LUT_3[5899] = 32'b00000000000000011000100111001100;
assign LUT_3[5900] = 32'b00000000000000001101000010000001;
assign LUT_3[5901] = 32'b00000000000000010011101101011110;
assign LUT_3[5902] = 32'b00000000000000001111001001100101;
assign LUT_3[5903] = 32'b00000000000000010101110101000010;
assign LUT_3[5904] = 32'b00000000000000001101101110001000;
assign LUT_3[5905] = 32'b00000000000000010100011001100101;
assign LUT_3[5906] = 32'b00000000000000001111110101101100;
assign LUT_3[5907] = 32'b00000000000000010110100001001001;
assign LUT_3[5908] = 32'b00000000000000001010111011111110;
assign LUT_3[5909] = 32'b00000000000000010001100111011011;
assign LUT_3[5910] = 32'b00000000000000001101000011100010;
assign LUT_3[5911] = 32'b00000000000000010011101110111111;
assign LUT_3[5912] = 32'b00000000000000010011000111001110;
assign LUT_3[5913] = 32'b00000000000000011001110010101011;
assign LUT_3[5914] = 32'b00000000000000010101001110110010;
assign LUT_3[5915] = 32'b00000000000000011011111010001111;
assign LUT_3[5916] = 32'b00000000000000010000010101000100;
assign LUT_3[5917] = 32'b00000000000000010111000000100001;
assign LUT_3[5918] = 32'b00000000000000010010011100101000;
assign LUT_3[5919] = 32'b00000000000000011001001000000101;
assign LUT_3[5920] = 32'b00000000000000001011101001100101;
assign LUT_3[5921] = 32'b00000000000000010010010101000010;
assign LUT_3[5922] = 32'b00000000000000001101110001001001;
assign LUT_3[5923] = 32'b00000000000000010100011100100110;
assign LUT_3[5924] = 32'b00000000000000001000110111011011;
assign LUT_3[5925] = 32'b00000000000000001111100010111000;
assign LUT_3[5926] = 32'b00000000000000001010111110111111;
assign LUT_3[5927] = 32'b00000000000000010001101010011100;
assign LUT_3[5928] = 32'b00000000000000010001000010101011;
assign LUT_3[5929] = 32'b00000000000000010111101110001000;
assign LUT_3[5930] = 32'b00000000000000010011001010001111;
assign LUT_3[5931] = 32'b00000000000000011001110101101100;
assign LUT_3[5932] = 32'b00000000000000001110010000100001;
assign LUT_3[5933] = 32'b00000000000000010100111011111110;
assign LUT_3[5934] = 32'b00000000000000010000011000000101;
assign LUT_3[5935] = 32'b00000000000000010111000011100010;
assign LUT_3[5936] = 32'b00000000000000001110111100101000;
assign LUT_3[5937] = 32'b00000000000000010101101000000101;
assign LUT_3[5938] = 32'b00000000000000010001000100001100;
assign LUT_3[5939] = 32'b00000000000000010111101111101001;
assign LUT_3[5940] = 32'b00000000000000001100001010011110;
assign LUT_3[5941] = 32'b00000000000000010010110101111011;
assign LUT_3[5942] = 32'b00000000000000001110010010000010;
assign LUT_3[5943] = 32'b00000000000000010100111101011111;
assign LUT_3[5944] = 32'b00000000000000010100010101101110;
assign LUT_3[5945] = 32'b00000000000000011011000001001011;
assign LUT_3[5946] = 32'b00000000000000010110011101010010;
assign LUT_3[5947] = 32'b00000000000000011101001000101111;
assign LUT_3[5948] = 32'b00000000000000010001100011100100;
assign LUT_3[5949] = 32'b00000000000000011000001111000001;
assign LUT_3[5950] = 32'b00000000000000010011101011001000;
assign LUT_3[5951] = 32'b00000000000000011010010110100101;
assign LUT_3[5952] = 32'b00000000000000001010010011110000;
assign LUT_3[5953] = 32'b00000000000000010000111111001101;
assign LUT_3[5954] = 32'b00000000000000001100011011010100;
assign LUT_3[5955] = 32'b00000000000000010011000110110001;
assign LUT_3[5956] = 32'b00000000000000000111100001100110;
assign LUT_3[5957] = 32'b00000000000000001110001101000011;
assign LUT_3[5958] = 32'b00000000000000001001101001001010;
assign LUT_3[5959] = 32'b00000000000000010000010100100111;
assign LUT_3[5960] = 32'b00000000000000001111101100110110;
assign LUT_3[5961] = 32'b00000000000000010110011000010011;
assign LUT_3[5962] = 32'b00000000000000010001110100011010;
assign LUT_3[5963] = 32'b00000000000000011000011111110111;
assign LUT_3[5964] = 32'b00000000000000001100111010101100;
assign LUT_3[5965] = 32'b00000000000000010011100110001001;
assign LUT_3[5966] = 32'b00000000000000001111000010010000;
assign LUT_3[5967] = 32'b00000000000000010101101101101101;
assign LUT_3[5968] = 32'b00000000000000001101100110110011;
assign LUT_3[5969] = 32'b00000000000000010100010010010000;
assign LUT_3[5970] = 32'b00000000000000001111101110010111;
assign LUT_3[5971] = 32'b00000000000000010110011001110100;
assign LUT_3[5972] = 32'b00000000000000001010110100101001;
assign LUT_3[5973] = 32'b00000000000000010001100000000110;
assign LUT_3[5974] = 32'b00000000000000001100111100001101;
assign LUT_3[5975] = 32'b00000000000000010011100111101010;
assign LUT_3[5976] = 32'b00000000000000010010111111111001;
assign LUT_3[5977] = 32'b00000000000000011001101011010110;
assign LUT_3[5978] = 32'b00000000000000010101000111011101;
assign LUT_3[5979] = 32'b00000000000000011011110010111010;
assign LUT_3[5980] = 32'b00000000000000010000001101101111;
assign LUT_3[5981] = 32'b00000000000000010110111001001100;
assign LUT_3[5982] = 32'b00000000000000010010010101010011;
assign LUT_3[5983] = 32'b00000000000000011001000000110000;
assign LUT_3[5984] = 32'b00000000000000001011100010010000;
assign LUT_3[5985] = 32'b00000000000000010010001101101101;
assign LUT_3[5986] = 32'b00000000000000001101101001110100;
assign LUT_3[5987] = 32'b00000000000000010100010101010001;
assign LUT_3[5988] = 32'b00000000000000001000110000000110;
assign LUT_3[5989] = 32'b00000000000000001111011011100011;
assign LUT_3[5990] = 32'b00000000000000001010110111101010;
assign LUT_3[5991] = 32'b00000000000000010001100011000111;
assign LUT_3[5992] = 32'b00000000000000010000111011010110;
assign LUT_3[5993] = 32'b00000000000000010111100110110011;
assign LUT_3[5994] = 32'b00000000000000010011000010111010;
assign LUT_3[5995] = 32'b00000000000000011001101110010111;
assign LUT_3[5996] = 32'b00000000000000001110001001001100;
assign LUT_3[5997] = 32'b00000000000000010100110100101001;
assign LUT_3[5998] = 32'b00000000000000010000010000110000;
assign LUT_3[5999] = 32'b00000000000000010110111100001101;
assign LUT_3[6000] = 32'b00000000000000001110110101010011;
assign LUT_3[6001] = 32'b00000000000000010101100000110000;
assign LUT_3[6002] = 32'b00000000000000010000111100110111;
assign LUT_3[6003] = 32'b00000000000000010111101000010100;
assign LUT_3[6004] = 32'b00000000000000001100000011001001;
assign LUT_3[6005] = 32'b00000000000000010010101110100110;
assign LUT_3[6006] = 32'b00000000000000001110001010101101;
assign LUT_3[6007] = 32'b00000000000000010100110110001010;
assign LUT_3[6008] = 32'b00000000000000010100001110011001;
assign LUT_3[6009] = 32'b00000000000000011010111001110110;
assign LUT_3[6010] = 32'b00000000000000010110010101111101;
assign LUT_3[6011] = 32'b00000000000000011101000001011010;
assign LUT_3[6012] = 32'b00000000000000010001011100001111;
assign LUT_3[6013] = 32'b00000000000000011000000111101100;
assign LUT_3[6014] = 32'b00000000000000010011100011110011;
assign LUT_3[6015] = 32'b00000000000000011010001111010000;
assign LUT_3[6016] = 32'b00000000000000001100100110000011;
assign LUT_3[6017] = 32'b00000000000000010011010001100000;
assign LUT_3[6018] = 32'b00000000000000001110101101100111;
assign LUT_3[6019] = 32'b00000000000000010101011001000100;
assign LUT_3[6020] = 32'b00000000000000001001110011111001;
assign LUT_3[6021] = 32'b00000000000000010000011111010110;
assign LUT_3[6022] = 32'b00000000000000001011111011011101;
assign LUT_3[6023] = 32'b00000000000000010010100110111010;
assign LUT_3[6024] = 32'b00000000000000010001111111001001;
assign LUT_3[6025] = 32'b00000000000000011000101010100110;
assign LUT_3[6026] = 32'b00000000000000010100000110101101;
assign LUT_3[6027] = 32'b00000000000000011010110010001010;
assign LUT_3[6028] = 32'b00000000000000001111001100111111;
assign LUT_3[6029] = 32'b00000000000000010101111000011100;
assign LUT_3[6030] = 32'b00000000000000010001010100100011;
assign LUT_3[6031] = 32'b00000000000000011000000000000000;
assign LUT_3[6032] = 32'b00000000000000001111111001000110;
assign LUT_3[6033] = 32'b00000000000000010110100100100011;
assign LUT_3[6034] = 32'b00000000000000010010000000101010;
assign LUT_3[6035] = 32'b00000000000000011000101100000111;
assign LUT_3[6036] = 32'b00000000000000001101000110111100;
assign LUT_3[6037] = 32'b00000000000000010011110010011001;
assign LUT_3[6038] = 32'b00000000000000001111001110100000;
assign LUT_3[6039] = 32'b00000000000000010101111001111101;
assign LUT_3[6040] = 32'b00000000000000010101010010001100;
assign LUT_3[6041] = 32'b00000000000000011011111101101001;
assign LUT_3[6042] = 32'b00000000000000010111011001110000;
assign LUT_3[6043] = 32'b00000000000000011110000101001101;
assign LUT_3[6044] = 32'b00000000000000010010100000000010;
assign LUT_3[6045] = 32'b00000000000000011001001011011111;
assign LUT_3[6046] = 32'b00000000000000010100100111100110;
assign LUT_3[6047] = 32'b00000000000000011011010011000011;
assign LUT_3[6048] = 32'b00000000000000001101110100100011;
assign LUT_3[6049] = 32'b00000000000000010100100000000000;
assign LUT_3[6050] = 32'b00000000000000001111111100000111;
assign LUT_3[6051] = 32'b00000000000000010110100111100100;
assign LUT_3[6052] = 32'b00000000000000001011000010011001;
assign LUT_3[6053] = 32'b00000000000000010001101101110110;
assign LUT_3[6054] = 32'b00000000000000001101001001111101;
assign LUT_3[6055] = 32'b00000000000000010011110101011010;
assign LUT_3[6056] = 32'b00000000000000010011001101101001;
assign LUT_3[6057] = 32'b00000000000000011001111001000110;
assign LUT_3[6058] = 32'b00000000000000010101010101001101;
assign LUT_3[6059] = 32'b00000000000000011100000000101010;
assign LUT_3[6060] = 32'b00000000000000010000011011011111;
assign LUT_3[6061] = 32'b00000000000000010111000110111100;
assign LUT_3[6062] = 32'b00000000000000010010100011000011;
assign LUT_3[6063] = 32'b00000000000000011001001110100000;
assign LUT_3[6064] = 32'b00000000000000010001000111100110;
assign LUT_3[6065] = 32'b00000000000000010111110011000011;
assign LUT_3[6066] = 32'b00000000000000010011001111001010;
assign LUT_3[6067] = 32'b00000000000000011001111010100111;
assign LUT_3[6068] = 32'b00000000000000001110010101011100;
assign LUT_3[6069] = 32'b00000000000000010101000000111001;
assign LUT_3[6070] = 32'b00000000000000010000011101000000;
assign LUT_3[6071] = 32'b00000000000000010111001000011101;
assign LUT_3[6072] = 32'b00000000000000010110100000101100;
assign LUT_3[6073] = 32'b00000000000000011101001100001001;
assign LUT_3[6074] = 32'b00000000000000011000101000010000;
assign LUT_3[6075] = 32'b00000000000000011111010011101101;
assign LUT_3[6076] = 32'b00000000000000010011101110100010;
assign LUT_3[6077] = 32'b00000000000000011010011001111111;
assign LUT_3[6078] = 32'b00000000000000010101110110000110;
assign LUT_3[6079] = 32'b00000000000000011100100001100011;
assign LUT_3[6080] = 32'b00000000000000001100011110101110;
assign LUT_3[6081] = 32'b00000000000000010011001010001011;
assign LUT_3[6082] = 32'b00000000000000001110100110010010;
assign LUT_3[6083] = 32'b00000000000000010101010001101111;
assign LUT_3[6084] = 32'b00000000000000001001101100100100;
assign LUT_3[6085] = 32'b00000000000000010000011000000001;
assign LUT_3[6086] = 32'b00000000000000001011110100001000;
assign LUT_3[6087] = 32'b00000000000000010010011111100101;
assign LUT_3[6088] = 32'b00000000000000010001110111110100;
assign LUT_3[6089] = 32'b00000000000000011000100011010001;
assign LUT_3[6090] = 32'b00000000000000010011111111011000;
assign LUT_3[6091] = 32'b00000000000000011010101010110101;
assign LUT_3[6092] = 32'b00000000000000001111000101101010;
assign LUT_3[6093] = 32'b00000000000000010101110001000111;
assign LUT_3[6094] = 32'b00000000000000010001001101001110;
assign LUT_3[6095] = 32'b00000000000000010111111000101011;
assign LUT_3[6096] = 32'b00000000000000001111110001110001;
assign LUT_3[6097] = 32'b00000000000000010110011101001110;
assign LUT_3[6098] = 32'b00000000000000010001111001010101;
assign LUT_3[6099] = 32'b00000000000000011000100100110010;
assign LUT_3[6100] = 32'b00000000000000001100111111100111;
assign LUT_3[6101] = 32'b00000000000000010011101011000100;
assign LUT_3[6102] = 32'b00000000000000001111000111001011;
assign LUT_3[6103] = 32'b00000000000000010101110010101000;
assign LUT_3[6104] = 32'b00000000000000010101001010110111;
assign LUT_3[6105] = 32'b00000000000000011011110110010100;
assign LUT_3[6106] = 32'b00000000000000010111010010011011;
assign LUT_3[6107] = 32'b00000000000000011101111101111000;
assign LUT_3[6108] = 32'b00000000000000010010011000101101;
assign LUT_3[6109] = 32'b00000000000000011001000100001010;
assign LUT_3[6110] = 32'b00000000000000010100100000010001;
assign LUT_3[6111] = 32'b00000000000000011011001011101110;
assign LUT_3[6112] = 32'b00000000000000001101101101001110;
assign LUT_3[6113] = 32'b00000000000000010100011000101011;
assign LUT_3[6114] = 32'b00000000000000001111110100110010;
assign LUT_3[6115] = 32'b00000000000000010110100000001111;
assign LUT_3[6116] = 32'b00000000000000001010111011000100;
assign LUT_3[6117] = 32'b00000000000000010001100110100001;
assign LUT_3[6118] = 32'b00000000000000001101000010101000;
assign LUT_3[6119] = 32'b00000000000000010011101110000101;
assign LUT_3[6120] = 32'b00000000000000010011000110010100;
assign LUT_3[6121] = 32'b00000000000000011001110001110001;
assign LUT_3[6122] = 32'b00000000000000010101001101111000;
assign LUT_3[6123] = 32'b00000000000000011011111001010101;
assign LUT_3[6124] = 32'b00000000000000010000010100001010;
assign LUT_3[6125] = 32'b00000000000000010110111111100111;
assign LUT_3[6126] = 32'b00000000000000010010011011101110;
assign LUT_3[6127] = 32'b00000000000000011001000111001011;
assign LUT_3[6128] = 32'b00000000000000010001000000010001;
assign LUT_3[6129] = 32'b00000000000000010111101011101110;
assign LUT_3[6130] = 32'b00000000000000010011000111110101;
assign LUT_3[6131] = 32'b00000000000000011001110011010010;
assign LUT_3[6132] = 32'b00000000000000001110001110000111;
assign LUT_3[6133] = 32'b00000000000000010100111001100100;
assign LUT_3[6134] = 32'b00000000000000010000010101101011;
assign LUT_3[6135] = 32'b00000000000000010111000001001000;
assign LUT_3[6136] = 32'b00000000000000010110011001010111;
assign LUT_3[6137] = 32'b00000000000000011101000100110100;
assign LUT_3[6138] = 32'b00000000000000011000100000111011;
assign LUT_3[6139] = 32'b00000000000000011111001100011000;
assign LUT_3[6140] = 32'b00000000000000010011100111001101;
assign LUT_3[6141] = 32'b00000000000000011010010010101010;
assign LUT_3[6142] = 32'b00000000000000010101101110110001;
assign LUT_3[6143] = 32'b00000000000000011100011010001110;
assign LUT_3[6144] = 32'b00000000000000000110000111101001;
assign LUT_3[6145] = 32'b00000000000000001100110011000110;
assign LUT_3[6146] = 32'b00000000000000001000001111001101;
assign LUT_3[6147] = 32'b00000000000000001110111010101010;
assign LUT_3[6148] = 32'b00000000000000000011010101011111;
assign LUT_3[6149] = 32'b00000000000000001010000000111100;
assign LUT_3[6150] = 32'b00000000000000000101011101000011;
assign LUT_3[6151] = 32'b00000000000000001100001000100000;
assign LUT_3[6152] = 32'b00000000000000001011100000101111;
assign LUT_3[6153] = 32'b00000000000000010010001100001100;
assign LUT_3[6154] = 32'b00000000000000001101101000010011;
assign LUT_3[6155] = 32'b00000000000000010100010011110000;
assign LUT_3[6156] = 32'b00000000000000001000101110100101;
assign LUT_3[6157] = 32'b00000000000000001111011010000010;
assign LUT_3[6158] = 32'b00000000000000001010110110001001;
assign LUT_3[6159] = 32'b00000000000000010001100001100110;
assign LUT_3[6160] = 32'b00000000000000001001011010101100;
assign LUT_3[6161] = 32'b00000000000000010000000110001001;
assign LUT_3[6162] = 32'b00000000000000001011100010010000;
assign LUT_3[6163] = 32'b00000000000000010010001101101101;
assign LUT_3[6164] = 32'b00000000000000000110101000100010;
assign LUT_3[6165] = 32'b00000000000000001101010011111111;
assign LUT_3[6166] = 32'b00000000000000001000110000000110;
assign LUT_3[6167] = 32'b00000000000000001111011011100011;
assign LUT_3[6168] = 32'b00000000000000001110110011110010;
assign LUT_3[6169] = 32'b00000000000000010101011111001111;
assign LUT_3[6170] = 32'b00000000000000010000111011010110;
assign LUT_3[6171] = 32'b00000000000000010111100110110011;
assign LUT_3[6172] = 32'b00000000000000001100000001101000;
assign LUT_3[6173] = 32'b00000000000000010010101101000101;
assign LUT_3[6174] = 32'b00000000000000001110001001001100;
assign LUT_3[6175] = 32'b00000000000000010100110100101001;
assign LUT_3[6176] = 32'b00000000000000000111010110001001;
assign LUT_3[6177] = 32'b00000000000000001110000001100110;
assign LUT_3[6178] = 32'b00000000000000001001011101101101;
assign LUT_3[6179] = 32'b00000000000000010000001001001010;
assign LUT_3[6180] = 32'b00000000000000000100100011111111;
assign LUT_3[6181] = 32'b00000000000000001011001111011100;
assign LUT_3[6182] = 32'b00000000000000000110101011100011;
assign LUT_3[6183] = 32'b00000000000000001101010111000000;
assign LUT_3[6184] = 32'b00000000000000001100101111001111;
assign LUT_3[6185] = 32'b00000000000000010011011010101100;
assign LUT_3[6186] = 32'b00000000000000001110110110110011;
assign LUT_3[6187] = 32'b00000000000000010101100010010000;
assign LUT_3[6188] = 32'b00000000000000001001111101000101;
assign LUT_3[6189] = 32'b00000000000000010000101000100010;
assign LUT_3[6190] = 32'b00000000000000001100000100101001;
assign LUT_3[6191] = 32'b00000000000000010010110000000110;
assign LUT_3[6192] = 32'b00000000000000001010101001001100;
assign LUT_3[6193] = 32'b00000000000000010001010100101001;
assign LUT_3[6194] = 32'b00000000000000001100110000110000;
assign LUT_3[6195] = 32'b00000000000000010011011100001101;
assign LUT_3[6196] = 32'b00000000000000000111110111000010;
assign LUT_3[6197] = 32'b00000000000000001110100010011111;
assign LUT_3[6198] = 32'b00000000000000001001111110100110;
assign LUT_3[6199] = 32'b00000000000000010000101010000011;
assign LUT_3[6200] = 32'b00000000000000010000000010010010;
assign LUT_3[6201] = 32'b00000000000000010110101101101111;
assign LUT_3[6202] = 32'b00000000000000010010001001110110;
assign LUT_3[6203] = 32'b00000000000000011000110101010011;
assign LUT_3[6204] = 32'b00000000000000001101010000001000;
assign LUT_3[6205] = 32'b00000000000000010011111011100101;
assign LUT_3[6206] = 32'b00000000000000001111010111101100;
assign LUT_3[6207] = 32'b00000000000000010110000011001001;
assign LUT_3[6208] = 32'b00000000000000000110000000010100;
assign LUT_3[6209] = 32'b00000000000000001100101011110001;
assign LUT_3[6210] = 32'b00000000000000001000000111111000;
assign LUT_3[6211] = 32'b00000000000000001110110011010101;
assign LUT_3[6212] = 32'b00000000000000000011001110001010;
assign LUT_3[6213] = 32'b00000000000000001001111001100111;
assign LUT_3[6214] = 32'b00000000000000000101010101101110;
assign LUT_3[6215] = 32'b00000000000000001100000001001011;
assign LUT_3[6216] = 32'b00000000000000001011011001011010;
assign LUT_3[6217] = 32'b00000000000000010010000100110111;
assign LUT_3[6218] = 32'b00000000000000001101100000111110;
assign LUT_3[6219] = 32'b00000000000000010100001100011011;
assign LUT_3[6220] = 32'b00000000000000001000100111010000;
assign LUT_3[6221] = 32'b00000000000000001111010010101101;
assign LUT_3[6222] = 32'b00000000000000001010101110110100;
assign LUT_3[6223] = 32'b00000000000000010001011010010001;
assign LUT_3[6224] = 32'b00000000000000001001010011010111;
assign LUT_3[6225] = 32'b00000000000000001111111110110100;
assign LUT_3[6226] = 32'b00000000000000001011011010111011;
assign LUT_3[6227] = 32'b00000000000000010010000110011000;
assign LUT_3[6228] = 32'b00000000000000000110100001001101;
assign LUT_3[6229] = 32'b00000000000000001101001100101010;
assign LUT_3[6230] = 32'b00000000000000001000101000110001;
assign LUT_3[6231] = 32'b00000000000000001111010100001110;
assign LUT_3[6232] = 32'b00000000000000001110101100011101;
assign LUT_3[6233] = 32'b00000000000000010101010111111010;
assign LUT_3[6234] = 32'b00000000000000010000110100000001;
assign LUT_3[6235] = 32'b00000000000000010111011111011110;
assign LUT_3[6236] = 32'b00000000000000001011111010010011;
assign LUT_3[6237] = 32'b00000000000000010010100101110000;
assign LUT_3[6238] = 32'b00000000000000001110000001110111;
assign LUT_3[6239] = 32'b00000000000000010100101101010100;
assign LUT_3[6240] = 32'b00000000000000000111001110110100;
assign LUT_3[6241] = 32'b00000000000000001101111010010001;
assign LUT_3[6242] = 32'b00000000000000001001010110011000;
assign LUT_3[6243] = 32'b00000000000000010000000001110101;
assign LUT_3[6244] = 32'b00000000000000000100011100101010;
assign LUT_3[6245] = 32'b00000000000000001011001000000111;
assign LUT_3[6246] = 32'b00000000000000000110100100001110;
assign LUT_3[6247] = 32'b00000000000000001101001111101011;
assign LUT_3[6248] = 32'b00000000000000001100100111111010;
assign LUT_3[6249] = 32'b00000000000000010011010011010111;
assign LUT_3[6250] = 32'b00000000000000001110101111011110;
assign LUT_3[6251] = 32'b00000000000000010101011010111011;
assign LUT_3[6252] = 32'b00000000000000001001110101110000;
assign LUT_3[6253] = 32'b00000000000000010000100001001101;
assign LUT_3[6254] = 32'b00000000000000001011111101010100;
assign LUT_3[6255] = 32'b00000000000000010010101000110001;
assign LUT_3[6256] = 32'b00000000000000001010100001110111;
assign LUT_3[6257] = 32'b00000000000000010001001101010100;
assign LUT_3[6258] = 32'b00000000000000001100101001011011;
assign LUT_3[6259] = 32'b00000000000000010011010100111000;
assign LUT_3[6260] = 32'b00000000000000000111101111101101;
assign LUT_3[6261] = 32'b00000000000000001110011011001010;
assign LUT_3[6262] = 32'b00000000000000001001110111010001;
assign LUT_3[6263] = 32'b00000000000000010000100010101110;
assign LUT_3[6264] = 32'b00000000000000001111111010111101;
assign LUT_3[6265] = 32'b00000000000000010110100110011010;
assign LUT_3[6266] = 32'b00000000000000010010000010100001;
assign LUT_3[6267] = 32'b00000000000000011000101101111110;
assign LUT_3[6268] = 32'b00000000000000001101001000110011;
assign LUT_3[6269] = 32'b00000000000000010011110100010000;
assign LUT_3[6270] = 32'b00000000000000001111010000010111;
assign LUT_3[6271] = 32'b00000000000000010101111011110100;
assign LUT_3[6272] = 32'b00000000000000001000010010100111;
assign LUT_3[6273] = 32'b00000000000000001110111110000100;
assign LUT_3[6274] = 32'b00000000000000001010011010001011;
assign LUT_3[6275] = 32'b00000000000000010001000101101000;
assign LUT_3[6276] = 32'b00000000000000000101100000011101;
assign LUT_3[6277] = 32'b00000000000000001100001011111010;
assign LUT_3[6278] = 32'b00000000000000000111101000000001;
assign LUT_3[6279] = 32'b00000000000000001110010011011110;
assign LUT_3[6280] = 32'b00000000000000001101101011101101;
assign LUT_3[6281] = 32'b00000000000000010100010111001010;
assign LUT_3[6282] = 32'b00000000000000001111110011010001;
assign LUT_3[6283] = 32'b00000000000000010110011110101110;
assign LUT_3[6284] = 32'b00000000000000001010111001100011;
assign LUT_3[6285] = 32'b00000000000000010001100101000000;
assign LUT_3[6286] = 32'b00000000000000001101000001000111;
assign LUT_3[6287] = 32'b00000000000000010011101100100100;
assign LUT_3[6288] = 32'b00000000000000001011100101101010;
assign LUT_3[6289] = 32'b00000000000000010010010001000111;
assign LUT_3[6290] = 32'b00000000000000001101101101001110;
assign LUT_3[6291] = 32'b00000000000000010100011000101011;
assign LUT_3[6292] = 32'b00000000000000001000110011100000;
assign LUT_3[6293] = 32'b00000000000000001111011110111101;
assign LUT_3[6294] = 32'b00000000000000001010111011000100;
assign LUT_3[6295] = 32'b00000000000000010001100110100001;
assign LUT_3[6296] = 32'b00000000000000010000111110110000;
assign LUT_3[6297] = 32'b00000000000000010111101010001101;
assign LUT_3[6298] = 32'b00000000000000010011000110010100;
assign LUT_3[6299] = 32'b00000000000000011001110001110001;
assign LUT_3[6300] = 32'b00000000000000001110001100100110;
assign LUT_3[6301] = 32'b00000000000000010100111000000011;
assign LUT_3[6302] = 32'b00000000000000010000010100001010;
assign LUT_3[6303] = 32'b00000000000000010110111111100111;
assign LUT_3[6304] = 32'b00000000000000001001100001000111;
assign LUT_3[6305] = 32'b00000000000000010000001100100100;
assign LUT_3[6306] = 32'b00000000000000001011101000101011;
assign LUT_3[6307] = 32'b00000000000000010010010100001000;
assign LUT_3[6308] = 32'b00000000000000000110101110111101;
assign LUT_3[6309] = 32'b00000000000000001101011010011010;
assign LUT_3[6310] = 32'b00000000000000001000110110100001;
assign LUT_3[6311] = 32'b00000000000000001111100001111110;
assign LUT_3[6312] = 32'b00000000000000001110111010001101;
assign LUT_3[6313] = 32'b00000000000000010101100101101010;
assign LUT_3[6314] = 32'b00000000000000010001000001110001;
assign LUT_3[6315] = 32'b00000000000000010111101101001110;
assign LUT_3[6316] = 32'b00000000000000001100001000000011;
assign LUT_3[6317] = 32'b00000000000000010010110011100000;
assign LUT_3[6318] = 32'b00000000000000001110001111100111;
assign LUT_3[6319] = 32'b00000000000000010100111011000100;
assign LUT_3[6320] = 32'b00000000000000001100110100001010;
assign LUT_3[6321] = 32'b00000000000000010011011111100111;
assign LUT_3[6322] = 32'b00000000000000001110111011101110;
assign LUT_3[6323] = 32'b00000000000000010101100111001011;
assign LUT_3[6324] = 32'b00000000000000001010000010000000;
assign LUT_3[6325] = 32'b00000000000000010000101101011101;
assign LUT_3[6326] = 32'b00000000000000001100001001100100;
assign LUT_3[6327] = 32'b00000000000000010010110101000001;
assign LUT_3[6328] = 32'b00000000000000010010001101010000;
assign LUT_3[6329] = 32'b00000000000000011000111000101101;
assign LUT_3[6330] = 32'b00000000000000010100010100110100;
assign LUT_3[6331] = 32'b00000000000000011011000000010001;
assign LUT_3[6332] = 32'b00000000000000001111011011000110;
assign LUT_3[6333] = 32'b00000000000000010110000110100011;
assign LUT_3[6334] = 32'b00000000000000010001100010101010;
assign LUT_3[6335] = 32'b00000000000000011000001110000111;
assign LUT_3[6336] = 32'b00000000000000001000001011010010;
assign LUT_3[6337] = 32'b00000000000000001110110110101111;
assign LUT_3[6338] = 32'b00000000000000001010010010110110;
assign LUT_3[6339] = 32'b00000000000000010000111110010011;
assign LUT_3[6340] = 32'b00000000000000000101011001001000;
assign LUT_3[6341] = 32'b00000000000000001100000100100101;
assign LUT_3[6342] = 32'b00000000000000000111100000101100;
assign LUT_3[6343] = 32'b00000000000000001110001100001001;
assign LUT_3[6344] = 32'b00000000000000001101100100011000;
assign LUT_3[6345] = 32'b00000000000000010100001111110101;
assign LUT_3[6346] = 32'b00000000000000001111101011111100;
assign LUT_3[6347] = 32'b00000000000000010110010111011001;
assign LUT_3[6348] = 32'b00000000000000001010110010001110;
assign LUT_3[6349] = 32'b00000000000000010001011101101011;
assign LUT_3[6350] = 32'b00000000000000001100111001110010;
assign LUT_3[6351] = 32'b00000000000000010011100101001111;
assign LUT_3[6352] = 32'b00000000000000001011011110010101;
assign LUT_3[6353] = 32'b00000000000000010010001001110010;
assign LUT_3[6354] = 32'b00000000000000001101100101111001;
assign LUT_3[6355] = 32'b00000000000000010100010001010110;
assign LUT_3[6356] = 32'b00000000000000001000101100001011;
assign LUT_3[6357] = 32'b00000000000000001111010111101000;
assign LUT_3[6358] = 32'b00000000000000001010110011101111;
assign LUT_3[6359] = 32'b00000000000000010001011111001100;
assign LUT_3[6360] = 32'b00000000000000010000110111011011;
assign LUT_3[6361] = 32'b00000000000000010111100010111000;
assign LUT_3[6362] = 32'b00000000000000010010111110111111;
assign LUT_3[6363] = 32'b00000000000000011001101010011100;
assign LUT_3[6364] = 32'b00000000000000001110000101010001;
assign LUT_3[6365] = 32'b00000000000000010100110000101110;
assign LUT_3[6366] = 32'b00000000000000010000001100110101;
assign LUT_3[6367] = 32'b00000000000000010110111000010010;
assign LUT_3[6368] = 32'b00000000000000001001011001110010;
assign LUT_3[6369] = 32'b00000000000000010000000101001111;
assign LUT_3[6370] = 32'b00000000000000001011100001010110;
assign LUT_3[6371] = 32'b00000000000000010010001100110011;
assign LUT_3[6372] = 32'b00000000000000000110100111101000;
assign LUT_3[6373] = 32'b00000000000000001101010011000101;
assign LUT_3[6374] = 32'b00000000000000001000101111001100;
assign LUT_3[6375] = 32'b00000000000000001111011010101001;
assign LUT_3[6376] = 32'b00000000000000001110110010111000;
assign LUT_3[6377] = 32'b00000000000000010101011110010101;
assign LUT_3[6378] = 32'b00000000000000010000111010011100;
assign LUT_3[6379] = 32'b00000000000000010111100101111001;
assign LUT_3[6380] = 32'b00000000000000001100000000101110;
assign LUT_3[6381] = 32'b00000000000000010010101100001011;
assign LUT_3[6382] = 32'b00000000000000001110001000010010;
assign LUT_3[6383] = 32'b00000000000000010100110011101111;
assign LUT_3[6384] = 32'b00000000000000001100101100110101;
assign LUT_3[6385] = 32'b00000000000000010011011000010010;
assign LUT_3[6386] = 32'b00000000000000001110110100011001;
assign LUT_3[6387] = 32'b00000000000000010101011111110110;
assign LUT_3[6388] = 32'b00000000000000001001111010101011;
assign LUT_3[6389] = 32'b00000000000000010000100110001000;
assign LUT_3[6390] = 32'b00000000000000001100000010001111;
assign LUT_3[6391] = 32'b00000000000000010010101101101100;
assign LUT_3[6392] = 32'b00000000000000010010000101111011;
assign LUT_3[6393] = 32'b00000000000000011000110001011000;
assign LUT_3[6394] = 32'b00000000000000010100001101011111;
assign LUT_3[6395] = 32'b00000000000000011010111000111100;
assign LUT_3[6396] = 32'b00000000000000001111010011110001;
assign LUT_3[6397] = 32'b00000000000000010101111111001110;
assign LUT_3[6398] = 32'b00000000000000010001011011010101;
assign LUT_3[6399] = 32'b00000000000000011000000110110010;
assign LUT_3[6400] = 32'b00000000000000000010010111001010;
assign LUT_3[6401] = 32'b00000000000000001001000010100111;
assign LUT_3[6402] = 32'b00000000000000000100011110101110;
assign LUT_3[6403] = 32'b00000000000000001011001010001011;
assign LUT_3[6404] = 32'b11111111111111111111100101000000;
assign LUT_3[6405] = 32'b00000000000000000110010000011101;
assign LUT_3[6406] = 32'b00000000000000000001101100100100;
assign LUT_3[6407] = 32'b00000000000000001000011000000001;
assign LUT_3[6408] = 32'b00000000000000000111110000010000;
assign LUT_3[6409] = 32'b00000000000000001110011011101101;
assign LUT_3[6410] = 32'b00000000000000001001110111110100;
assign LUT_3[6411] = 32'b00000000000000010000100011010001;
assign LUT_3[6412] = 32'b00000000000000000100111110000110;
assign LUT_3[6413] = 32'b00000000000000001011101001100011;
assign LUT_3[6414] = 32'b00000000000000000111000101101010;
assign LUT_3[6415] = 32'b00000000000000001101110001000111;
assign LUT_3[6416] = 32'b00000000000000000101101010001101;
assign LUT_3[6417] = 32'b00000000000000001100010101101010;
assign LUT_3[6418] = 32'b00000000000000000111110001110001;
assign LUT_3[6419] = 32'b00000000000000001110011101001110;
assign LUT_3[6420] = 32'b00000000000000000010111000000011;
assign LUT_3[6421] = 32'b00000000000000001001100011100000;
assign LUT_3[6422] = 32'b00000000000000000100111111100111;
assign LUT_3[6423] = 32'b00000000000000001011101011000100;
assign LUT_3[6424] = 32'b00000000000000001011000011010011;
assign LUT_3[6425] = 32'b00000000000000010001101110110000;
assign LUT_3[6426] = 32'b00000000000000001101001010110111;
assign LUT_3[6427] = 32'b00000000000000010011110110010100;
assign LUT_3[6428] = 32'b00000000000000001000010001001001;
assign LUT_3[6429] = 32'b00000000000000001110111100100110;
assign LUT_3[6430] = 32'b00000000000000001010011000101101;
assign LUT_3[6431] = 32'b00000000000000010001000100001010;
assign LUT_3[6432] = 32'b00000000000000000011100101101010;
assign LUT_3[6433] = 32'b00000000000000001010010001000111;
assign LUT_3[6434] = 32'b00000000000000000101101101001110;
assign LUT_3[6435] = 32'b00000000000000001100011000101011;
assign LUT_3[6436] = 32'b00000000000000000000110011100000;
assign LUT_3[6437] = 32'b00000000000000000111011110111101;
assign LUT_3[6438] = 32'b00000000000000000010111011000100;
assign LUT_3[6439] = 32'b00000000000000001001100110100001;
assign LUT_3[6440] = 32'b00000000000000001000111110110000;
assign LUT_3[6441] = 32'b00000000000000001111101010001101;
assign LUT_3[6442] = 32'b00000000000000001011000110010100;
assign LUT_3[6443] = 32'b00000000000000010001110001110001;
assign LUT_3[6444] = 32'b00000000000000000110001100100110;
assign LUT_3[6445] = 32'b00000000000000001100111000000011;
assign LUT_3[6446] = 32'b00000000000000001000010100001010;
assign LUT_3[6447] = 32'b00000000000000001110111111100111;
assign LUT_3[6448] = 32'b00000000000000000110111000101101;
assign LUT_3[6449] = 32'b00000000000000001101100100001010;
assign LUT_3[6450] = 32'b00000000000000001001000000010001;
assign LUT_3[6451] = 32'b00000000000000001111101011101110;
assign LUT_3[6452] = 32'b00000000000000000100000110100011;
assign LUT_3[6453] = 32'b00000000000000001010110010000000;
assign LUT_3[6454] = 32'b00000000000000000110001110000111;
assign LUT_3[6455] = 32'b00000000000000001100111001100100;
assign LUT_3[6456] = 32'b00000000000000001100010001110011;
assign LUT_3[6457] = 32'b00000000000000010010111101010000;
assign LUT_3[6458] = 32'b00000000000000001110011001010111;
assign LUT_3[6459] = 32'b00000000000000010101000100110100;
assign LUT_3[6460] = 32'b00000000000000001001011111101001;
assign LUT_3[6461] = 32'b00000000000000010000001011000110;
assign LUT_3[6462] = 32'b00000000000000001011100111001101;
assign LUT_3[6463] = 32'b00000000000000010010010010101010;
assign LUT_3[6464] = 32'b00000000000000000010001111110101;
assign LUT_3[6465] = 32'b00000000000000001000111011010010;
assign LUT_3[6466] = 32'b00000000000000000100010111011001;
assign LUT_3[6467] = 32'b00000000000000001011000010110110;
assign LUT_3[6468] = 32'b11111111111111111111011101101011;
assign LUT_3[6469] = 32'b00000000000000000110001001001000;
assign LUT_3[6470] = 32'b00000000000000000001100101001111;
assign LUT_3[6471] = 32'b00000000000000001000010000101100;
assign LUT_3[6472] = 32'b00000000000000000111101000111011;
assign LUT_3[6473] = 32'b00000000000000001110010100011000;
assign LUT_3[6474] = 32'b00000000000000001001110000011111;
assign LUT_3[6475] = 32'b00000000000000010000011011111100;
assign LUT_3[6476] = 32'b00000000000000000100110110110001;
assign LUT_3[6477] = 32'b00000000000000001011100010001110;
assign LUT_3[6478] = 32'b00000000000000000110111110010101;
assign LUT_3[6479] = 32'b00000000000000001101101001110010;
assign LUT_3[6480] = 32'b00000000000000000101100010111000;
assign LUT_3[6481] = 32'b00000000000000001100001110010101;
assign LUT_3[6482] = 32'b00000000000000000111101010011100;
assign LUT_3[6483] = 32'b00000000000000001110010101111001;
assign LUT_3[6484] = 32'b00000000000000000010110000101110;
assign LUT_3[6485] = 32'b00000000000000001001011100001011;
assign LUT_3[6486] = 32'b00000000000000000100111000010010;
assign LUT_3[6487] = 32'b00000000000000001011100011101111;
assign LUT_3[6488] = 32'b00000000000000001010111011111110;
assign LUT_3[6489] = 32'b00000000000000010001100111011011;
assign LUT_3[6490] = 32'b00000000000000001101000011100010;
assign LUT_3[6491] = 32'b00000000000000010011101110111111;
assign LUT_3[6492] = 32'b00000000000000001000001001110100;
assign LUT_3[6493] = 32'b00000000000000001110110101010001;
assign LUT_3[6494] = 32'b00000000000000001010010001011000;
assign LUT_3[6495] = 32'b00000000000000010000111100110101;
assign LUT_3[6496] = 32'b00000000000000000011011110010101;
assign LUT_3[6497] = 32'b00000000000000001010001001110010;
assign LUT_3[6498] = 32'b00000000000000000101100101111001;
assign LUT_3[6499] = 32'b00000000000000001100010001010110;
assign LUT_3[6500] = 32'b00000000000000000000101100001011;
assign LUT_3[6501] = 32'b00000000000000000111010111101000;
assign LUT_3[6502] = 32'b00000000000000000010110011101111;
assign LUT_3[6503] = 32'b00000000000000001001011111001100;
assign LUT_3[6504] = 32'b00000000000000001000110111011011;
assign LUT_3[6505] = 32'b00000000000000001111100010111000;
assign LUT_3[6506] = 32'b00000000000000001010111110111111;
assign LUT_3[6507] = 32'b00000000000000010001101010011100;
assign LUT_3[6508] = 32'b00000000000000000110000101010001;
assign LUT_3[6509] = 32'b00000000000000001100110000101110;
assign LUT_3[6510] = 32'b00000000000000001000001100110101;
assign LUT_3[6511] = 32'b00000000000000001110111000010010;
assign LUT_3[6512] = 32'b00000000000000000110110001011000;
assign LUT_3[6513] = 32'b00000000000000001101011100110101;
assign LUT_3[6514] = 32'b00000000000000001000111000111100;
assign LUT_3[6515] = 32'b00000000000000001111100100011001;
assign LUT_3[6516] = 32'b00000000000000000011111111001110;
assign LUT_3[6517] = 32'b00000000000000001010101010101011;
assign LUT_3[6518] = 32'b00000000000000000110000110110010;
assign LUT_3[6519] = 32'b00000000000000001100110010001111;
assign LUT_3[6520] = 32'b00000000000000001100001010011110;
assign LUT_3[6521] = 32'b00000000000000010010110101111011;
assign LUT_3[6522] = 32'b00000000000000001110010010000010;
assign LUT_3[6523] = 32'b00000000000000010100111101011111;
assign LUT_3[6524] = 32'b00000000000000001001011000010100;
assign LUT_3[6525] = 32'b00000000000000010000000011110001;
assign LUT_3[6526] = 32'b00000000000000001011011111111000;
assign LUT_3[6527] = 32'b00000000000000010010001011010101;
assign LUT_3[6528] = 32'b00000000000000000100100010001000;
assign LUT_3[6529] = 32'b00000000000000001011001101100101;
assign LUT_3[6530] = 32'b00000000000000000110101001101100;
assign LUT_3[6531] = 32'b00000000000000001101010101001001;
assign LUT_3[6532] = 32'b00000000000000000001101111111110;
assign LUT_3[6533] = 32'b00000000000000001000011011011011;
assign LUT_3[6534] = 32'b00000000000000000011110111100010;
assign LUT_3[6535] = 32'b00000000000000001010100010111111;
assign LUT_3[6536] = 32'b00000000000000001001111011001110;
assign LUT_3[6537] = 32'b00000000000000010000100110101011;
assign LUT_3[6538] = 32'b00000000000000001100000010110010;
assign LUT_3[6539] = 32'b00000000000000010010101110001111;
assign LUT_3[6540] = 32'b00000000000000000111001001000100;
assign LUT_3[6541] = 32'b00000000000000001101110100100001;
assign LUT_3[6542] = 32'b00000000000000001001010000101000;
assign LUT_3[6543] = 32'b00000000000000001111111100000101;
assign LUT_3[6544] = 32'b00000000000000000111110101001011;
assign LUT_3[6545] = 32'b00000000000000001110100000101000;
assign LUT_3[6546] = 32'b00000000000000001001111100101111;
assign LUT_3[6547] = 32'b00000000000000010000101000001100;
assign LUT_3[6548] = 32'b00000000000000000101000011000001;
assign LUT_3[6549] = 32'b00000000000000001011101110011110;
assign LUT_3[6550] = 32'b00000000000000000111001010100101;
assign LUT_3[6551] = 32'b00000000000000001101110110000010;
assign LUT_3[6552] = 32'b00000000000000001101001110010001;
assign LUT_3[6553] = 32'b00000000000000010011111001101110;
assign LUT_3[6554] = 32'b00000000000000001111010101110101;
assign LUT_3[6555] = 32'b00000000000000010110000001010010;
assign LUT_3[6556] = 32'b00000000000000001010011100000111;
assign LUT_3[6557] = 32'b00000000000000010001000111100100;
assign LUT_3[6558] = 32'b00000000000000001100100011101011;
assign LUT_3[6559] = 32'b00000000000000010011001111001000;
assign LUT_3[6560] = 32'b00000000000000000101110000101000;
assign LUT_3[6561] = 32'b00000000000000001100011100000101;
assign LUT_3[6562] = 32'b00000000000000000111111000001100;
assign LUT_3[6563] = 32'b00000000000000001110100011101001;
assign LUT_3[6564] = 32'b00000000000000000010111110011110;
assign LUT_3[6565] = 32'b00000000000000001001101001111011;
assign LUT_3[6566] = 32'b00000000000000000101000110000010;
assign LUT_3[6567] = 32'b00000000000000001011110001011111;
assign LUT_3[6568] = 32'b00000000000000001011001001101110;
assign LUT_3[6569] = 32'b00000000000000010001110101001011;
assign LUT_3[6570] = 32'b00000000000000001101010001010010;
assign LUT_3[6571] = 32'b00000000000000010011111100101111;
assign LUT_3[6572] = 32'b00000000000000001000010111100100;
assign LUT_3[6573] = 32'b00000000000000001111000011000001;
assign LUT_3[6574] = 32'b00000000000000001010011111001000;
assign LUT_3[6575] = 32'b00000000000000010001001010100101;
assign LUT_3[6576] = 32'b00000000000000001001000011101011;
assign LUT_3[6577] = 32'b00000000000000001111101111001000;
assign LUT_3[6578] = 32'b00000000000000001011001011001111;
assign LUT_3[6579] = 32'b00000000000000010001110110101100;
assign LUT_3[6580] = 32'b00000000000000000110010001100001;
assign LUT_3[6581] = 32'b00000000000000001100111100111110;
assign LUT_3[6582] = 32'b00000000000000001000011001000101;
assign LUT_3[6583] = 32'b00000000000000001111000100100010;
assign LUT_3[6584] = 32'b00000000000000001110011100110001;
assign LUT_3[6585] = 32'b00000000000000010101001000001110;
assign LUT_3[6586] = 32'b00000000000000010000100100010101;
assign LUT_3[6587] = 32'b00000000000000010111001111110010;
assign LUT_3[6588] = 32'b00000000000000001011101010100111;
assign LUT_3[6589] = 32'b00000000000000010010010110000100;
assign LUT_3[6590] = 32'b00000000000000001101110010001011;
assign LUT_3[6591] = 32'b00000000000000010100011101101000;
assign LUT_3[6592] = 32'b00000000000000000100011010110011;
assign LUT_3[6593] = 32'b00000000000000001011000110010000;
assign LUT_3[6594] = 32'b00000000000000000110100010010111;
assign LUT_3[6595] = 32'b00000000000000001101001101110100;
assign LUT_3[6596] = 32'b00000000000000000001101000101001;
assign LUT_3[6597] = 32'b00000000000000001000010100000110;
assign LUT_3[6598] = 32'b00000000000000000011110000001101;
assign LUT_3[6599] = 32'b00000000000000001010011011101010;
assign LUT_3[6600] = 32'b00000000000000001001110011111001;
assign LUT_3[6601] = 32'b00000000000000010000011111010110;
assign LUT_3[6602] = 32'b00000000000000001011111011011101;
assign LUT_3[6603] = 32'b00000000000000010010100110111010;
assign LUT_3[6604] = 32'b00000000000000000111000001101111;
assign LUT_3[6605] = 32'b00000000000000001101101101001100;
assign LUT_3[6606] = 32'b00000000000000001001001001010011;
assign LUT_3[6607] = 32'b00000000000000001111110100110000;
assign LUT_3[6608] = 32'b00000000000000000111101101110110;
assign LUT_3[6609] = 32'b00000000000000001110011001010011;
assign LUT_3[6610] = 32'b00000000000000001001110101011010;
assign LUT_3[6611] = 32'b00000000000000010000100000110111;
assign LUT_3[6612] = 32'b00000000000000000100111011101100;
assign LUT_3[6613] = 32'b00000000000000001011100111001001;
assign LUT_3[6614] = 32'b00000000000000000111000011010000;
assign LUT_3[6615] = 32'b00000000000000001101101110101101;
assign LUT_3[6616] = 32'b00000000000000001101000110111100;
assign LUT_3[6617] = 32'b00000000000000010011110010011001;
assign LUT_3[6618] = 32'b00000000000000001111001110100000;
assign LUT_3[6619] = 32'b00000000000000010101111001111101;
assign LUT_3[6620] = 32'b00000000000000001010010100110010;
assign LUT_3[6621] = 32'b00000000000000010001000000001111;
assign LUT_3[6622] = 32'b00000000000000001100011100010110;
assign LUT_3[6623] = 32'b00000000000000010011000111110011;
assign LUT_3[6624] = 32'b00000000000000000101101001010011;
assign LUT_3[6625] = 32'b00000000000000001100010100110000;
assign LUT_3[6626] = 32'b00000000000000000111110000110111;
assign LUT_3[6627] = 32'b00000000000000001110011100010100;
assign LUT_3[6628] = 32'b00000000000000000010110111001001;
assign LUT_3[6629] = 32'b00000000000000001001100010100110;
assign LUT_3[6630] = 32'b00000000000000000100111110101101;
assign LUT_3[6631] = 32'b00000000000000001011101010001010;
assign LUT_3[6632] = 32'b00000000000000001011000010011001;
assign LUT_3[6633] = 32'b00000000000000010001101101110110;
assign LUT_3[6634] = 32'b00000000000000001101001001111101;
assign LUT_3[6635] = 32'b00000000000000010011110101011010;
assign LUT_3[6636] = 32'b00000000000000001000010000001111;
assign LUT_3[6637] = 32'b00000000000000001110111011101100;
assign LUT_3[6638] = 32'b00000000000000001010010111110011;
assign LUT_3[6639] = 32'b00000000000000010001000011010000;
assign LUT_3[6640] = 32'b00000000000000001000111100010110;
assign LUT_3[6641] = 32'b00000000000000001111100111110011;
assign LUT_3[6642] = 32'b00000000000000001011000011111010;
assign LUT_3[6643] = 32'b00000000000000010001101111010111;
assign LUT_3[6644] = 32'b00000000000000000110001010001100;
assign LUT_3[6645] = 32'b00000000000000001100110101101001;
assign LUT_3[6646] = 32'b00000000000000001000010001110000;
assign LUT_3[6647] = 32'b00000000000000001110111101001101;
assign LUT_3[6648] = 32'b00000000000000001110010101011100;
assign LUT_3[6649] = 32'b00000000000000010101000000111001;
assign LUT_3[6650] = 32'b00000000000000010000011101000000;
assign LUT_3[6651] = 32'b00000000000000010111001000011101;
assign LUT_3[6652] = 32'b00000000000000001011100011010010;
assign LUT_3[6653] = 32'b00000000000000010010001110101111;
assign LUT_3[6654] = 32'b00000000000000001101101010110110;
assign LUT_3[6655] = 32'b00000000000000010100010110010011;
assign LUT_3[6656] = 32'b00000000000000001001011100110101;
assign LUT_3[6657] = 32'b00000000000000010000001000010010;
assign LUT_3[6658] = 32'b00000000000000001011100100011001;
assign LUT_3[6659] = 32'b00000000000000010010001111110110;
assign LUT_3[6660] = 32'b00000000000000000110101010101011;
assign LUT_3[6661] = 32'b00000000000000001101010110001000;
assign LUT_3[6662] = 32'b00000000000000001000110010001111;
assign LUT_3[6663] = 32'b00000000000000001111011101101100;
assign LUT_3[6664] = 32'b00000000000000001110110101111011;
assign LUT_3[6665] = 32'b00000000000000010101100001011000;
assign LUT_3[6666] = 32'b00000000000000010000111101011111;
assign LUT_3[6667] = 32'b00000000000000010111101000111100;
assign LUT_3[6668] = 32'b00000000000000001100000011110001;
assign LUT_3[6669] = 32'b00000000000000010010101111001110;
assign LUT_3[6670] = 32'b00000000000000001110001011010101;
assign LUT_3[6671] = 32'b00000000000000010100110110110010;
assign LUT_3[6672] = 32'b00000000000000001100101111111000;
assign LUT_3[6673] = 32'b00000000000000010011011011010101;
assign LUT_3[6674] = 32'b00000000000000001110110111011100;
assign LUT_3[6675] = 32'b00000000000000010101100010111001;
assign LUT_3[6676] = 32'b00000000000000001001111101101110;
assign LUT_3[6677] = 32'b00000000000000010000101001001011;
assign LUT_3[6678] = 32'b00000000000000001100000101010010;
assign LUT_3[6679] = 32'b00000000000000010010110000101111;
assign LUT_3[6680] = 32'b00000000000000010010001000111110;
assign LUT_3[6681] = 32'b00000000000000011000110100011011;
assign LUT_3[6682] = 32'b00000000000000010100010000100010;
assign LUT_3[6683] = 32'b00000000000000011010111011111111;
assign LUT_3[6684] = 32'b00000000000000001111010110110100;
assign LUT_3[6685] = 32'b00000000000000010110000010010001;
assign LUT_3[6686] = 32'b00000000000000010001011110011000;
assign LUT_3[6687] = 32'b00000000000000011000001001110101;
assign LUT_3[6688] = 32'b00000000000000001010101011010101;
assign LUT_3[6689] = 32'b00000000000000010001010110110010;
assign LUT_3[6690] = 32'b00000000000000001100110010111001;
assign LUT_3[6691] = 32'b00000000000000010011011110010110;
assign LUT_3[6692] = 32'b00000000000000000111111001001011;
assign LUT_3[6693] = 32'b00000000000000001110100100101000;
assign LUT_3[6694] = 32'b00000000000000001010000000101111;
assign LUT_3[6695] = 32'b00000000000000010000101100001100;
assign LUT_3[6696] = 32'b00000000000000010000000100011011;
assign LUT_3[6697] = 32'b00000000000000010110101111111000;
assign LUT_3[6698] = 32'b00000000000000010010001011111111;
assign LUT_3[6699] = 32'b00000000000000011000110111011100;
assign LUT_3[6700] = 32'b00000000000000001101010010010001;
assign LUT_3[6701] = 32'b00000000000000010011111101101110;
assign LUT_3[6702] = 32'b00000000000000001111011001110101;
assign LUT_3[6703] = 32'b00000000000000010110000101010010;
assign LUT_3[6704] = 32'b00000000000000001101111110011000;
assign LUT_3[6705] = 32'b00000000000000010100101001110101;
assign LUT_3[6706] = 32'b00000000000000010000000101111100;
assign LUT_3[6707] = 32'b00000000000000010110110001011001;
assign LUT_3[6708] = 32'b00000000000000001011001100001110;
assign LUT_3[6709] = 32'b00000000000000010001110111101011;
assign LUT_3[6710] = 32'b00000000000000001101010011110010;
assign LUT_3[6711] = 32'b00000000000000010011111111001111;
assign LUT_3[6712] = 32'b00000000000000010011010111011110;
assign LUT_3[6713] = 32'b00000000000000011010000010111011;
assign LUT_3[6714] = 32'b00000000000000010101011111000010;
assign LUT_3[6715] = 32'b00000000000000011100001010011111;
assign LUT_3[6716] = 32'b00000000000000010000100101010100;
assign LUT_3[6717] = 32'b00000000000000010111010000110001;
assign LUT_3[6718] = 32'b00000000000000010010101100111000;
assign LUT_3[6719] = 32'b00000000000000011001011000010101;
assign LUT_3[6720] = 32'b00000000000000001001010101100000;
assign LUT_3[6721] = 32'b00000000000000010000000000111101;
assign LUT_3[6722] = 32'b00000000000000001011011101000100;
assign LUT_3[6723] = 32'b00000000000000010010001000100001;
assign LUT_3[6724] = 32'b00000000000000000110100011010110;
assign LUT_3[6725] = 32'b00000000000000001101001110110011;
assign LUT_3[6726] = 32'b00000000000000001000101010111010;
assign LUT_3[6727] = 32'b00000000000000001111010110010111;
assign LUT_3[6728] = 32'b00000000000000001110101110100110;
assign LUT_3[6729] = 32'b00000000000000010101011010000011;
assign LUT_3[6730] = 32'b00000000000000010000110110001010;
assign LUT_3[6731] = 32'b00000000000000010111100001100111;
assign LUT_3[6732] = 32'b00000000000000001011111100011100;
assign LUT_3[6733] = 32'b00000000000000010010100111111001;
assign LUT_3[6734] = 32'b00000000000000001110000100000000;
assign LUT_3[6735] = 32'b00000000000000010100101111011101;
assign LUT_3[6736] = 32'b00000000000000001100101000100011;
assign LUT_3[6737] = 32'b00000000000000010011010100000000;
assign LUT_3[6738] = 32'b00000000000000001110110000000111;
assign LUT_3[6739] = 32'b00000000000000010101011011100100;
assign LUT_3[6740] = 32'b00000000000000001001110110011001;
assign LUT_3[6741] = 32'b00000000000000010000100001110110;
assign LUT_3[6742] = 32'b00000000000000001011111101111101;
assign LUT_3[6743] = 32'b00000000000000010010101001011010;
assign LUT_3[6744] = 32'b00000000000000010010000001101001;
assign LUT_3[6745] = 32'b00000000000000011000101101000110;
assign LUT_3[6746] = 32'b00000000000000010100001001001101;
assign LUT_3[6747] = 32'b00000000000000011010110100101010;
assign LUT_3[6748] = 32'b00000000000000001111001111011111;
assign LUT_3[6749] = 32'b00000000000000010101111010111100;
assign LUT_3[6750] = 32'b00000000000000010001010111000011;
assign LUT_3[6751] = 32'b00000000000000011000000010100000;
assign LUT_3[6752] = 32'b00000000000000001010100100000000;
assign LUT_3[6753] = 32'b00000000000000010001001111011101;
assign LUT_3[6754] = 32'b00000000000000001100101011100100;
assign LUT_3[6755] = 32'b00000000000000010011010111000001;
assign LUT_3[6756] = 32'b00000000000000000111110001110110;
assign LUT_3[6757] = 32'b00000000000000001110011101010011;
assign LUT_3[6758] = 32'b00000000000000001001111001011010;
assign LUT_3[6759] = 32'b00000000000000010000100100110111;
assign LUT_3[6760] = 32'b00000000000000001111111101000110;
assign LUT_3[6761] = 32'b00000000000000010110101000100011;
assign LUT_3[6762] = 32'b00000000000000010010000100101010;
assign LUT_3[6763] = 32'b00000000000000011000110000000111;
assign LUT_3[6764] = 32'b00000000000000001101001010111100;
assign LUT_3[6765] = 32'b00000000000000010011110110011001;
assign LUT_3[6766] = 32'b00000000000000001111010010100000;
assign LUT_3[6767] = 32'b00000000000000010101111101111101;
assign LUT_3[6768] = 32'b00000000000000001101110111000011;
assign LUT_3[6769] = 32'b00000000000000010100100010100000;
assign LUT_3[6770] = 32'b00000000000000001111111110100111;
assign LUT_3[6771] = 32'b00000000000000010110101010000100;
assign LUT_3[6772] = 32'b00000000000000001011000100111001;
assign LUT_3[6773] = 32'b00000000000000010001110000010110;
assign LUT_3[6774] = 32'b00000000000000001101001100011101;
assign LUT_3[6775] = 32'b00000000000000010011110111111010;
assign LUT_3[6776] = 32'b00000000000000010011010000001001;
assign LUT_3[6777] = 32'b00000000000000011001111011100110;
assign LUT_3[6778] = 32'b00000000000000010101010111101101;
assign LUT_3[6779] = 32'b00000000000000011100000011001010;
assign LUT_3[6780] = 32'b00000000000000010000011101111111;
assign LUT_3[6781] = 32'b00000000000000010111001001011100;
assign LUT_3[6782] = 32'b00000000000000010010100101100011;
assign LUT_3[6783] = 32'b00000000000000011001010001000000;
assign LUT_3[6784] = 32'b00000000000000001011100111110011;
assign LUT_3[6785] = 32'b00000000000000010010010011010000;
assign LUT_3[6786] = 32'b00000000000000001101101111010111;
assign LUT_3[6787] = 32'b00000000000000010100011010110100;
assign LUT_3[6788] = 32'b00000000000000001000110101101001;
assign LUT_3[6789] = 32'b00000000000000001111100001000110;
assign LUT_3[6790] = 32'b00000000000000001010111101001101;
assign LUT_3[6791] = 32'b00000000000000010001101000101010;
assign LUT_3[6792] = 32'b00000000000000010001000000111001;
assign LUT_3[6793] = 32'b00000000000000010111101100010110;
assign LUT_3[6794] = 32'b00000000000000010011001000011101;
assign LUT_3[6795] = 32'b00000000000000011001110011111010;
assign LUT_3[6796] = 32'b00000000000000001110001110101111;
assign LUT_3[6797] = 32'b00000000000000010100111010001100;
assign LUT_3[6798] = 32'b00000000000000010000010110010011;
assign LUT_3[6799] = 32'b00000000000000010111000001110000;
assign LUT_3[6800] = 32'b00000000000000001110111010110110;
assign LUT_3[6801] = 32'b00000000000000010101100110010011;
assign LUT_3[6802] = 32'b00000000000000010001000010011010;
assign LUT_3[6803] = 32'b00000000000000010111101101110111;
assign LUT_3[6804] = 32'b00000000000000001100001000101100;
assign LUT_3[6805] = 32'b00000000000000010010110100001001;
assign LUT_3[6806] = 32'b00000000000000001110010000010000;
assign LUT_3[6807] = 32'b00000000000000010100111011101101;
assign LUT_3[6808] = 32'b00000000000000010100010011111100;
assign LUT_3[6809] = 32'b00000000000000011010111111011001;
assign LUT_3[6810] = 32'b00000000000000010110011011100000;
assign LUT_3[6811] = 32'b00000000000000011101000110111101;
assign LUT_3[6812] = 32'b00000000000000010001100001110010;
assign LUT_3[6813] = 32'b00000000000000011000001101001111;
assign LUT_3[6814] = 32'b00000000000000010011101001010110;
assign LUT_3[6815] = 32'b00000000000000011010010100110011;
assign LUT_3[6816] = 32'b00000000000000001100110110010011;
assign LUT_3[6817] = 32'b00000000000000010011100001110000;
assign LUT_3[6818] = 32'b00000000000000001110111101110111;
assign LUT_3[6819] = 32'b00000000000000010101101001010100;
assign LUT_3[6820] = 32'b00000000000000001010000100001001;
assign LUT_3[6821] = 32'b00000000000000010000101111100110;
assign LUT_3[6822] = 32'b00000000000000001100001011101101;
assign LUT_3[6823] = 32'b00000000000000010010110111001010;
assign LUT_3[6824] = 32'b00000000000000010010001111011001;
assign LUT_3[6825] = 32'b00000000000000011000111010110110;
assign LUT_3[6826] = 32'b00000000000000010100010110111101;
assign LUT_3[6827] = 32'b00000000000000011011000010011010;
assign LUT_3[6828] = 32'b00000000000000001111011101001111;
assign LUT_3[6829] = 32'b00000000000000010110001000101100;
assign LUT_3[6830] = 32'b00000000000000010001100100110011;
assign LUT_3[6831] = 32'b00000000000000011000010000010000;
assign LUT_3[6832] = 32'b00000000000000010000001001010110;
assign LUT_3[6833] = 32'b00000000000000010110110100110011;
assign LUT_3[6834] = 32'b00000000000000010010010000111010;
assign LUT_3[6835] = 32'b00000000000000011000111100010111;
assign LUT_3[6836] = 32'b00000000000000001101010111001100;
assign LUT_3[6837] = 32'b00000000000000010100000010101001;
assign LUT_3[6838] = 32'b00000000000000001111011110110000;
assign LUT_3[6839] = 32'b00000000000000010110001010001101;
assign LUT_3[6840] = 32'b00000000000000010101100010011100;
assign LUT_3[6841] = 32'b00000000000000011100001101111001;
assign LUT_3[6842] = 32'b00000000000000010111101010000000;
assign LUT_3[6843] = 32'b00000000000000011110010101011101;
assign LUT_3[6844] = 32'b00000000000000010010110000010010;
assign LUT_3[6845] = 32'b00000000000000011001011011101111;
assign LUT_3[6846] = 32'b00000000000000010100110111110110;
assign LUT_3[6847] = 32'b00000000000000011011100011010011;
assign LUT_3[6848] = 32'b00000000000000001011100000011110;
assign LUT_3[6849] = 32'b00000000000000010010001011111011;
assign LUT_3[6850] = 32'b00000000000000001101101000000010;
assign LUT_3[6851] = 32'b00000000000000010100010011011111;
assign LUT_3[6852] = 32'b00000000000000001000101110010100;
assign LUT_3[6853] = 32'b00000000000000001111011001110001;
assign LUT_3[6854] = 32'b00000000000000001010110101111000;
assign LUT_3[6855] = 32'b00000000000000010001100001010101;
assign LUT_3[6856] = 32'b00000000000000010000111001100100;
assign LUT_3[6857] = 32'b00000000000000010111100101000001;
assign LUT_3[6858] = 32'b00000000000000010011000001001000;
assign LUT_3[6859] = 32'b00000000000000011001101100100101;
assign LUT_3[6860] = 32'b00000000000000001110000111011010;
assign LUT_3[6861] = 32'b00000000000000010100110010110111;
assign LUT_3[6862] = 32'b00000000000000010000001110111110;
assign LUT_3[6863] = 32'b00000000000000010110111010011011;
assign LUT_3[6864] = 32'b00000000000000001110110011100001;
assign LUT_3[6865] = 32'b00000000000000010101011110111110;
assign LUT_3[6866] = 32'b00000000000000010000111011000101;
assign LUT_3[6867] = 32'b00000000000000010111100110100010;
assign LUT_3[6868] = 32'b00000000000000001100000001010111;
assign LUT_3[6869] = 32'b00000000000000010010101100110100;
assign LUT_3[6870] = 32'b00000000000000001110001000111011;
assign LUT_3[6871] = 32'b00000000000000010100110100011000;
assign LUT_3[6872] = 32'b00000000000000010100001100100111;
assign LUT_3[6873] = 32'b00000000000000011010111000000100;
assign LUT_3[6874] = 32'b00000000000000010110010100001011;
assign LUT_3[6875] = 32'b00000000000000011100111111101000;
assign LUT_3[6876] = 32'b00000000000000010001011010011101;
assign LUT_3[6877] = 32'b00000000000000011000000101111010;
assign LUT_3[6878] = 32'b00000000000000010011100010000001;
assign LUT_3[6879] = 32'b00000000000000011010001101011110;
assign LUT_3[6880] = 32'b00000000000000001100101110111110;
assign LUT_3[6881] = 32'b00000000000000010011011010011011;
assign LUT_3[6882] = 32'b00000000000000001110110110100010;
assign LUT_3[6883] = 32'b00000000000000010101100001111111;
assign LUT_3[6884] = 32'b00000000000000001001111100110100;
assign LUT_3[6885] = 32'b00000000000000010000101000010001;
assign LUT_3[6886] = 32'b00000000000000001100000100011000;
assign LUT_3[6887] = 32'b00000000000000010010101111110101;
assign LUT_3[6888] = 32'b00000000000000010010001000000100;
assign LUT_3[6889] = 32'b00000000000000011000110011100001;
assign LUT_3[6890] = 32'b00000000000000010100001111101000;
assign LUT_3[6891] = 32'b00000000000000011010111011000101;
assign LUT_3[6892] = 32'b00000000000000001111010101111010;
assign LUT_3[6893] = 32'b00000000000000010110000001010111;
assign LUT_3[6894] = 32'b00000000000000010001011101011110;
assign LUT_3[6895] = 32'b00000000000000011000001000111011;
assign LUT_3[6896] = 32'b00000000000000010000000010000001;
assign LUT_3[6897] = 32'b00000000000000010110101101011110;
assign LUT_3[6898] = 32'b00000000000000010010001001100101;
assign LUT_3[6899] = 32'b00000000000000011000110101000010;
assign LUT_3[6900] = 32'b00000000000000001101001111110111;
assign LUT_3[6901] = 32'b00000000000000010011111011010100;
assign LUT_3[6902] = 32'b00000000000000001111010111011011;
assign LUT_3[6903] = 32'b00000000000000010110000010111000;
assign LUT_3[6904] = 32'b00000000000000010101011011000111;
assign LUT_3[6905] = 32'b00000000000000011100000110100100;
assign LUT_3[6906] = 32'b00000000000000010111100010101011;
assign LUT_3[6907] = 32'b00000000000000011110001110001000;
assign LUT_3[6908] = 32'b00000000000000010010101000111101;
assign LUT_3[6909] = 32'b00000000000000011001010100011010;
assign LUT_3[6910] = 32'b00000000000000010100110000100001;
assign LUT_3[6911] = 32'b00000000000000011011011011111110;
assign LUT_3[6912] = 32'b00000000000000000101101100010110;
assign LUT_3[6913] = 32'b00000000000000001100010111110011;
assign LUT_3[6914] = 32'b00000000000000000111110011111010;
assign LUT_3[6915] = 32'b00000000000000001110011111010111;
assign LUT_3[6916] = 32'b00000000000000000010111010001100;
assign LUT_3[6917] = 32'b00000000000000001001100101101001;
assign LUT_3[6918] = 32'b00000000000000000101000001110000;
assign LUT_3[6919] = 32'b00000000000000001011101101001101;
assign LUT_3[6920] = 32'b00000000000000001011000101011100;
assign LUT_3[6921] = 32'b00000000000000010001110000111001;
assign LUT_3[6922] = 32'b00000000000000001101001101000000;
assign LUT_3[6923] = 32'b00000000000000010011111000011101;
assign LUT_3[6924] = 32'b00000000000000001000010011010010;
assign LUT_3[6925] = 32'b00000000000000001110111110101111;
assign LUT_3[6926] = 32'b00000000000000001010011010110110;
assign LUT_3[6927] = 32'b00000000000000010001000110010011;
assign LUT_3[6928] = 32'b00000000000000001000111111011001;
assign LUT_3[6929] = 32'b00000000000000001111101010110110;
assign LUT_3[6930] = 32'b00000000000000001011000110111101;
assign LUT_3[6931] = 32'b00000000000000010001110010011010;
assign LUT_3[6932] = 32'b00000000000000000110001101001111;
assign LUT_3[6933] = 32'b00000000000000001100111000101100;
assign LUT_3[6934] = 32'b00000000000000001000010100110011;
assign LUT_3[6935] = 32'b00000000000000001111000000010000;
assign LUT_3[6936] = 32'b00000000000000001110011000011111;
assign LUT_3[6937] = 32'b00000000000000010101000011111100;
assign LUT_3[6938] = 32'b00000000000000010000100000000011;
assign LUT_3[6939] = 32'b00000000000000010111001011100000;
assign LUT_3[6940] = 32'b00000000000000001011100110010101;
assign LUT_3[6941] = 32'b00000000000000010010010001110010;
assign LUT_3[6942] = 32'b00000000000000001101101101111001;
assign LUT_3[6943] = 32'b00000000000000010100011001010110;
assign LUT_3[6944] = 32'b00000000000000000110111010110110;
assign LUT_3[6945] = 32'b00000000000000001101100110010011;
assign LUT_3[6946] = 32'b00000000000000001001000010011010;
assign LUT_3[6947] = 32'b00000000000000001111101101110111;
assign LUT_3[6948] = 32'b00000000000000000100001000101100;
assign LUT_3[6949] = 32'b00000000000000001010110100001001;
assign LUT_3[6950] = 32'b00000000000000000110010000010000;
assign LUT_3[6951] = 32'b00000000000000001100111011101101;
assign LUT_3[6952] = 32'b00000000000000001100010011111100;
assign LUT_3[6953] = 32'b00000000000000010010111111011001;
assign LUT_3[6954] = 32'b00000000000000001110011011100000;
assign LUT_3[6955] = 32'b00000000000000010101000110111101;
assign LUT_3[6956] = 32'b00000000000000001001100001110010;
assign LUT_3[6957] = 32'b00000000000000010000001101001111;
assign LUT_3[6958] = 32'b00000000000000001011101001010110;
assign LUT_3[6959] = 32'b00000000000000010010010100110011;
assign LUT_3[6960] = 32'b00000000000000001010001101111001;
assign LUT_3[6961] = 32'b00000000000000010000111001010110;
assign LUT_3[6962] = 32'b00000000000000001100010101011101;
assign LUT_3[6963] = 32'b00000000000000010011000000111010;
assign LUT_3[6964] = 32'b00000000000000000111011011101111;
assign LUT_3[6965] = 32'b00000000000000001110000111001100;
assign LUT_3[6966] = 32'b00000000000000001001100011010011;
assign LUT_3[6967] = 32'b00000000000000010000001110110000;
assign LUT_3[6968] = 32'b00000000000000001111100110111111;
assign LUT_3[6969] = 32'b00000000000000010110010010011100;
assign LUT_3[6970] = 32'b00000000000000010001101110100011;
assign LUT_3[6971] = 32'b00000000000000011000011010000000;
assign LUT_3[6972] = 32'b00000000000000001100110100110101;
assign LUT_3[6973] = 32'b00000000000000010011100000010010;
assign LUT_3[6974] = 32'b00000000000000001110111100011001;
assign LUT_3[6975] = 32'b00000000000000010101100111110110;
assign LUT_3[6976] = 32'b00000000000000000101100101000001;
assign LUT_3[6977] = 32'b00000000000000001100010000011110;
assign LUT_3[6978] = 32'b00000000000000000111101100100101;
assign LUT_3[6979] = 32'b00000000000000001110011000000010;
assign LUT_3[6980] = 32'b00000000000000000010110010110111;
assign LUT_3[6981] = 32'b00000000000000001001011110010100;
assign LUT_3[6982] = 32'b00000000000000000100111010011011;
assign LUT_3[6983] = 32'b00000000000000001011100101111000;
assign LUT_3[6984] = 32'b00000000000000001010111110000111;
assign LUT_3[6985] = 32'b00000000000000010001101001100100;
assign LUT_3[6986] = 32'b00000000000000001101000101101011;
assign LUT_3[6987] = 32'b00000000000000010011110001001000;
assign LUT_3[6988] = 32'b00000000000000001000001011111101;
assign LUT_3[6989] = 32'b00000000000000001110110111011010;
assign LUT_3[6990] = 32'b00000000000000001010010011100001;
assign LUT_3[6991] = 32'b00000000000000010000111110111110;
assign LUT_3[6992] = 32'b00000000000000001000111000000100;
assign LUT_3[6993] = 32'b00000000000000001111100011100001;
assign LUT_3[6994] = 32'b00000000000000001010111111101000;
assign LUT_3[6995] = 32'b00000000000000010001101011000101;
assign LUT_3[6996] = 32'b00000000000000000110000101111010;
assign LUT_3[6997] = 32'b00000000000000001100110001010111;
assign LUT_3[6998] = 32'b00000000000000001000001101011110;
assign LUT_3[6999] = 32'b00000000000000001110111000111011;
assign LUT_3[7000] = 32'b00000000000000001110010001001010;
assign LUT_3[7001] = 32'b00000000000000010100111100100111;
assign LUT_3[7002] = 32'b00000000000000010000011000101110;
assign LUT_3[7003] = 32'b00000000000000010111000100001011;
assign LUT_3[7004] = 32'b00000000000000001011011111000000;
assign LUT_3[7005] = 32'b00000000000000010010001010011101;
assign LUT_3[7006] = 32'b00000000000000001101100110100100;
assign LUT_3[7007] = 32'b00000000000000010100010010000001;
assign LUT_3[7008] = 32'b00000000000000000110110011100001;
assign LUT_3[7009] = 32'b00000000000000001101011110111110;
assign LUT_3[7010] = 32'b00000000000000001000111011000101;
assign LUT_3[7011] = 32'b00000000000000001111100110100010;
assign LUT_3[7012] = 32'b00000000000000000100000001010111;
assign LUT_3[7013] = 32'b00000000000000001010101100110100;
assign LUT_3[7014] = 32'b00000000000000000110001000111011;
assign LUT_3[7015] = 32'b00000000000000001100110100011000;
assign LUT_3[7016] = 32'b00000000000000001100001100100111;
assign LUT_3[7017] = 32'b00000000000000010010111000000100;
assign LUT_3[7018] = 32'b00000000000000001110010100001011;
assign LUT_3[7019] = 32'b00000000000000010100111111101000;
assign LUT_3[7020] = 32'b00000000000000001001011010011101;
assign LUT_3[7021] = 32'b00000000000000010000000101111010;
assign LUT_3[7022] = 32'b00000000000000001011100010000001;
assign LUT_3[7023] = 32'b00000000000000010010001101011110;
assign LUT_3[7024] = 32'b00000000000000001010000110100100;
assign LUT_3[7025] = 32'b00000000000000010000110010000001;
assign LUT_3[7026] = 32'b00000000000000001100001110001000;
assign LUT_3[7027] = 32'b00000000000000010010111001100101;
assign LUT_3[7028] = 32'b00000000000000000111010100011010;
assign LUT_3[7029] = 32'b00000000000000001101111111110111;
assign LUT_3[7030] = 32'b00000000000000001001011011111110;
assign LUT_3[7031] = 32'b00000000000000010000000111011011;
assign LUT_3[7032] = 32'b00000000000000001111011111101010;
assign LUT_3[7033] = 32'b00000000000000010110001011000111;
assign LUT_3[7034] = 32'b00000000000000010001100111001110;
assign LUT_3[7035] = 32'b00000000000000011000010010101011;
assign LUT_3[7036] = 32'b00000000000000001100101101100000;
assign LUT_3[7037] = 32'b00000000000000010011011000111101;
assign LUT_3[7038] = 32'b00000000000000001110110101000100;
assign LUT_3[7039] = 32'b00000000000000010101100000100001;
assign LUT_3[7040] = 32'b00000000000000000111110111010100;
assign LUT_3[7041] = 32'b00000000000000001110100010110001;
assign LUT_3[7042] = 32'b00000000000000001001111110111000;
assign LUT_3[7043] = 32'b00000000000000010000101010010101;
assign LUT_3[7044] = 32'b00000000000000000101000101001010;
assign LUT_3[7045] = 32'b00000000000000001011110000100111;
assign LUT_3[7046] = 32'b00000000000000000111001100101110;
assign LUT_3[7047] = 32'b00000000000000001101111000001011;
assign LUT_3[7048] = 32'b00000000000000001101010000011010;
assign LUT_3[7049] = 32'b00000000000000010011111011110111;
assign LUT_3[7050] = 32'b00000000000000001111010111111110;
assign LUT_3[7051] = 32'b00000000000000010110000011011011;
assign LUT_3[7052] = 32'b00000000000000001010011110010000;
assign LUT_3[7053] = 32'b00000000000000010001001001101101;
assign LUT_3[7054] = 32'b00000000000000001100100101110100;
assign LUT_3[7055] = 32'b00000000000000010011010001010001;
assign LUT_3[7056] = 32'b00000000000000001011001010010111;
assign LUT_3[7057] = 32'b00000000000000010001110101110100;
assign LUT_3[7058] = 32'b00000000000000001101010001111011;
assign LUT_3[7059] = 32'b00000000000000010011111101011000;
assign LUT_3[7060] = 32'b00000000000000001000011000001101;
assign LUT_3[7061] = 32'b00000000000000001111000011101010;
assign LUT_3[7062] = 32'b00000000000000001010011111110001;
assign LUT_3[7063] = 32'b00000000000000010001001011001110;
assign LUT_3[7064] = 32'b00000000000000010000100011011101;
assign LUT_3[7065] = 32'b00000000000000010111001110111010;
assign LUT_3[7066] = 32'b00000000000000010010101011000001;
assign LUT_3[7067] = 32'b00000000000000011001010110011110;
assign LUT_3[7068] = 32'b00000000000000001101110001010011;
assign LUT_3[7069] = 32'b00000000000000010100011100110000;
assign LUT_3[7070] = 32'b00000000000000001111111000110111;
assign LUT_3[7071] = 32'b00000000000000010110100100010100;
assign LUT_3[7072] = 32'b00000000000000001001000101110100;
assign LUT_3[7073] = 32'b00000000000000001111110001010001;
assign LUT_3[7074] = 32'b00000000000000001011001101011000;
assign LUT_3[7075] = 32'b00000000000000010001111000110101;
assign LUT_3[7076] = 32'b00000000000000000110010011101010;
assign LUT_3[7077] = 32'b00000000000000001100111111000111;
assign LUT_3[7078] = 32'b00000000000000001000011011001110;
assign LUT_3[7079] = 32'b00000000000000001111000110101011;
assign LUT_3[7080] = 32'b00000000000000001110011110111010;
assign LUT_3[7081] = 32'b00000000000000010101001010010111;
assign LUT_3[7082] = 32'b00000000000000010000100110011110;
assign LUT_3[7083] = 32'b00000000000000010111010001111011;
assign LUT_3[7084] = 32'b00000000000000001011101100110000;
assign LUT_3[7085] = 32'b00000000000000010010011000001101;
assign LUT_3[7086] = 32'b00000000000000001101110100010100;
assign LUT_3[7087] = 32'b00000000000000010100011111110001;
assign LUT_3[7088] = 32'b00000000000000001100011000110111;
assign LUT_3[7089] = 32'b00000000000000010011000100010100;
assign LUT_3[7090] = 32'b00000000000000001110100000011011;
assign LUT_3[7091] = 32'b00000000000000010101001011111000;
assign LUT_3[7092] = 32'b00000000000000001001100110101101;
assign LUT_3[7093] = 32'b00000000000000010000010010001010;
assign LUT_3[7094] = 32'b00000000000000001011101110010001;
assign LUT_3[7095] = 32'b00000000000000010010011001101110;
assign LUT_3[7096] = 32'b00000000000000010001110001111101;
assign LUT_3[7097] = 32'b00000000000000011000011101011010;
assign LUT_3[7098] = 32'b00000000000000010011111001100001;
assign LUT_3[7099] = 32'b00000000000000011010100100111110;
assign LUT_3[7100] = 32'b00000000000000001110111111110011;
assign LUT_3[7101] = 32'b00000000000000010101101011010000;
assign LUT_3[7102] = 32'b00000000000000010001000111010111;
assign LUT_3[7103] = 32'b00000000000000010111110010110100;
assign LUT_3[7104] = 32'b00000000000000000111101111111111;
assign LUT_3[7105] = 32'b00000000000000001110011011011100;
assign LUT_3[7106] = 32'b00000000000000001001110111100011;
assign LUT_3[7107] = 32'b00000000000000010000100011000000;
assign LUT_3[7108] = 32'b00000000000000000100111101110101;
assign LUT_3[7109] = 32'b00000000000000001011101001010010;
assign LUT_3[7110] = 32'b00000000000000000111000101011001;
assign LUT_3[7111] = 32'b00000000000000001101110000110110;
assign LUT_3[7112] = 32'b00000000000000001101001001000101;
assign LUT_3[7113] = 32'b00000000000000010011110100100010;
assign LUT_3[7114] = 32'b00000000000000001111010000101001;
assign LUT_3[7115] = 32'b00000000000000010101111100000110;
assign LUT_3[7116] = 32'b00000000000000001010010110111011;
assign LUT_3[7117] = 32'b00000000000000010001000010011000;
assign LUT_3[7118] = 32'b00000000000000001100011110011111;
assign LUT_3[7119] = 32'b00000000000000010011001001111100;
assign LUT_3[7120] = 32'b00000000000000001011000011000010;
assign LUT_3[7121] = 32'b00000000000000010001101110011111;
assign LUT_3[7122] = 32'b00000000000000001101001010100110;
assign LUT_3[7123] = 32'b00000000000000010011110110000011;
assign LUT_3[7124] = 32'b00000000000000001000010000111000;
assign LUT_3[7125] = 32'b00000000000000001110111100010101;
assign LUT_3[7126] = 32'b00000000000000001010011000011100;
assign LUT_3[7127] = 32'b00000000000000010001000011111001;
assign LUT_3[7128] = 32'b00000000000000010000011100001000;
assign LUT_3[7129] = 32'b00000000000000010111000111100101;
assign LUT_3[7130] = 32'b00000000000000010010100011101100;
assign LUT_3[7131] = 32'b00000000000000011001001111001001;
assign LUT_3[7132] = 32'b00000000000000001101101001111110;
assign LUT_3[7133] = 32'b00000000000000010100010101011011;
assign LUT_3[7134] = 32'b00000000000000001111110001100010;
assign LUT_3[7135] = 32'b00000000000000010110011100111111;
assign LUT_3[7136] = 32'b00000000000000001000111110011111;
assign LUT_3[7137] = 32'b00000000000000001111101001111100;
assign LUT_3[7138] = 32'b00000000000000001011000110000011;
assign LUT_3[7139] = 32'b00000000000000010001110001100000;
assign LUT_3[7140] = 32'b00000000000000000110001100010101;
assign LUT_3[7141] = 32'b00000000000000001100110111110010;
assign LUT_3[7142] = 32'b00000000000000001000010011111001;
assign LUT_3[7143] = 32'b00000000000000001110111111010110;
assign LUT_3[7144] = 32'b00000000000000001110010111100101;
assign LUT_3[7145] = 32'b00000000000000010101000011000010;
assign LUT_3[7146] = 32'b00000000000000010000011111001001;
assign LUT_3[7147] = 32'b00000000000000010111001010100110;
assign LUT_3[7148] = 32'b00000000000000001011100101011011;
assign LUT_3[7149] = 32'b00000000000000010010010000111000;
assign LUT_3[7150] = 32'b00000000000000001101101100111111;
assign LUT_3[7151] = 32'b00000000000000010100011000011100;
assign LUT_3[7152] = 32'b00000000000000001100010001100010;
assign LUT_3[7153] = 32'b00000000000000010010111100111111;
assign LUT_3[7154] = 32'b00000000000000001110011001000110;
assign LUT_3[7155] = 32'b00000000000000010101000100100011;
assign LUT_3[7156] = 32'b00000000000000001001011111011000;
assign LUT_3[7157] = 32'b00000000000000010000001010110101;
assign LUT_3[7158] = 32'b00000000000000001011100110111100;
assign LUT_3[7159] = 32'b00000000000000010010010010011001;
assign LUT_3[7160] = 32'b00000000000000010001101010101000;
assign LUT_3[7161] = 32'b00000000000000011000010110000101;
assign LUT_3[7162] = 32'b00000000000000010011110010001100;
assign LUT_3[7163] = 32'b00000000000000011010011101101001;
assign LUT_3[7164] = 32'b00000000000000001110111000011110;
assign LUT_3[7165] = 32'b00000000000000010101100011111011;
assign LUT_3[7166] = 32'b00000000000000010001000000000010;
assign LUT_3[7167] = 32'b00000000000000010111101011011111;
assign LUT_3[7168] = 32'b00000000000000001100101100100110;
assign LUT_3[7169] = 32'b00000000000000010011011000000011;
assign LUT_3[7170] = 32'b00000000000000001110110100001010;
assign LUT_3[7171] = 32'b00000000000000010101011111100111;
assign LUT_3[7172] = 32'b00000000000000001001111010011100;
assign LUT_3[7173] = 32'b00000000000000010000100101111001;
assign LUT_3[7174] = 32'b00000000000000001100000010000000;
assign LUT_3[7175] = 32'b00000000000000010010101101011101;
assign LUT_3[7176] = 32'b00000000000000010010000101101100;
assign LUT_3[7177] = 32'b00000000000000011000110001001001;
assign LUT_3[7178] = 32'b00000000000000010100001101010000;
assign LUT_3[7179] = 32'b00000000000000011010111000101101;
assign LUT_3[7180] = 32'b00000000000000001111010011100010;
assign LUT_3[7181] = 32'b00000000000000010101111110111111;
assign LUT_3[7182] = 32'b00000000000000010001011011000110;
assign LUT_3[7183] = 32'b00000000000000011000000110100011;
assign LUT_3[7184] = 32'b00000000000000001111111111101001;
assign LUT_3[7185] = 32'b00000000000000010110101011000110;
assign LUT_3[7186] = 32'b00000000000000010010000111001101;
assign LUT_3[7187] = 32'b00000000000000011000110010101010;
assign LUT_3[7188] = 32'b00000000000000001101001101011111;
assign LUT_3[7189] = 32'b00000000000000010011111000111100;
assign LUT_3[7190] = 32'b00000000000000001111010101000011;
assign LUT_3[7191] = 32'b00000000000000010110000000100000;
assign LUT_3[7192] = 32'b00000000000000010101011000101111;
assign LUT_3[7193] = 32'b00000000000000011100000100001100;
assign LUT_3[7194] = 32'b00000000000000010111100000010011;
assign LUT_3[7195] = 32'b00000000000000011110001011110000;
assign LUT_3[7196] = 32'b00000000000000010010100110100101;
assign LUT_3[7197] = 32'b00000000000000011001010010000010;
assign LUT_3[7198] = 32'b00000000000000010100101110001001;
assign LUT_3[7199] = 32'b00000000000000011011011001100110;
assign LUT_3[7200] = 32'b00000000000000001101111011000110;
assign LUT_3[7201] = 32'b00000000000000010100100110100011;
assign LUT_3[7202] = 32'b00000000000000010000000010101010;
assign LUT_3[7203] = 32'b00000000000000010110101110000111;
assign LUT_3[7204] = 32'b00000000000000001011001000111100;
assign LUT_3[7205] = 32'b00000000000000010001110100011001;
assign LUT_3[7206] = 32'b00000000000000001101010000100000;
assign LUT_3[7207] = 32'b00000000000000010011111011111101;
assign LUT_3[7208] = 32'b00000000000000010011010100001100;
assign LUT_3[7209] = 32'b00000000000000011001111111101001;
assign LUT_3[7210] = 32'b00000000000000010101011011110000;
assign LUT_3[7211] = 32'b00000000000000011100000111001101;
assign LUT_3[7212] = 32'b00000000000000010000100010000010;
assign LUT_3[7213] = 32'b00000000000000010111001101011111;
assign LUT_3[7214] = 32'b00000000000000010010101001100110;
assign LUT_3[7215] = 32'b00000000000000011001010101000011;
assign LUT_3[7216] = 32'b00000000000000010001001110001001;
assign LUT_3[7217] = 32'b00000000000000010111111001100110;
assign LUT_3[7218] = 32'b00000000000000010011010101101101;
assign LUT_3[7219] = 32'b00000000000000011010000001001010;
assign LUT_3[7220] = 32'b00000000000000001110011011111111;
assign LUT_3[7221] = 32'b00000000000000010101000111011100;
assign LUT_3[7222] = 32'b00000000000000010000100011100011;
assign LUT_3[7223] = 32'b00000000000000010111001111000000;
assign LUT_3[7224] = 32'b00000000000000010110100111001111;
assign LUT_3[7225] = 32'b00000000000000011101010010101100;
assign LUT_3[7226] = 32'b00000000000000011000101110110011;
assign LUT_3[7227] = 32'b00000000000000011111011010010000;
assign LUT_3[7228] = 32'b00000000000000010011110101000101;
assign LUT_3[7229] = 32'b00000000000000011010100000100010;
assign LUT_3[7230] = 32'b00000000000000010101111100101001;
assign LUT_3[7231] = 32'b00000000000000011100101000000110;
assign LUT_3[7232] = 32'b00000000000000001100100101010001;
assign LUT_3[7233] = 32'b00000000000000010011010000101110;
assign LUT_3[7234] = 32'b00000000000000001110101100110101;
assign LUT_3[7235] = 32'b00000000000000010101011000010010;
assign LUT_3[7236] = 32'b00000000000000001001110011000111;
assign LUT_3[7237] = 32'b00000000000000010000011110100100;
assign LUT_3[7238] = 32'b00000000000000001011111010101011;
assign LUT_3[7239] = 32'b00000000000000010010100110001000;
assign LUT_3[7240] = 32'b00000000000000010001111110010111;
assign LUT_3[7241] = 32'b00000000000000011000101001110100;
assign LUT_3[7242] = 32'b00000000000000010100000101111011;
assign LUT_3[7243] = 32'b00000000000000011010110001011000;
assign LUT_3[7244] = 32'b00000000000000001111001100001101;
assign LUT_3[7245] = 32'b00000000000000010101110111101010;
assign LUT_3[7246] = 32'b00000000000000010001010011110001;
assign LUT_3[7247] = 32'b00000000000000010111111111001110;
assign LUT_3[7248] = 32'b00000000000000001111111000010100;
assign LUT_3[7249] = 32'b00000000000000010110100011110001;
assign LUT_3[7250] = 32'b00000000000000010001111111111000;
assign LUT_3[7251] = 32'b00000000000000011000101011010101;
assign LUT_3[7252] = 32'b00000000000000001101000110001010;
assign LUT_3[7253] = 32'b00000000000000010011110001100111;
assign LUT_3[7254] = 32'b00000000000000001111001101101110;
assign LUT_3[7255] = 32'b00000000000000010101111001001011;
assign LUT_3[7256] = 32'b00000000000000010101010001011010;
assign LUT_3[7257] = 32'b00000000000000011011111100110111;
assign LUT_3[7258] = 32'b00000000000000010111011000111110;
assign LUT_3[7259] = 32'b00000000000000011110000100011011;
assign LUT_3[7260] = 32'b00000000000000010010011111010000;
assign LUT_3[7261] = 32'b00000000000000011001001010101101;
assign LUT_3[7262] = 32'b00000000000000010100100110110100;
assign LUT_3[7263] = 32'b00000000000000011011010010010001;
assign LUT_3[7264] = 32'b00000000000000001101110011110001;
assign LUT_3[7265] = 32'b00000000000000010100011111001110;
assign LUT_3[7266] = 32'b00000000000000001111111011010101;
assign LUT_3[7267] = 32'b00000000000000010110100110110010;
assign LUT_3[7268] = 32'b00000000000000001011000001100111;
assign LUT_3[7269] = 32'b00000000000000010001101101000100;
assign LUT_3[7270] = 32'b00000000000000001101001001001011;
assign LUT_3[7271] = 32'b00000000000000010011110100101000;
assign LUT_3[7272] = 32'b00000000000000010011001100110111;
assign LUT_3[7273] = 32'b00000000000000011001111000010100;
assign LUT_3[7274] = 32'b00000000000000010101010100011011;
assign LUT_3[7275] = 32'b00000000000000011011111111111000;
assign LUT_3[7276] = 32'b00000000000000010000011010101101;
assign LUT_3[7277] = 32'b00000000000000010111000110001010;
assign LUT_3[7278] = 32'b00000000000000010010100010010001;
assign LUT_3[7279] = 32'b00000000000000011001001101101110;
assign LUT_3[7280] = 32'b00000000000000010001000110110100;
assign LUT_3[7281] = 32'b00000000000000010111110010010001;
assign LUT_3[7282] = 32'b00000000000000010011001110011000;
assign LUT_3[7283] = 32'b00000000000000011001111001110101;
assign LUT_3[7284] = 32'b00000000000000001110010100101010;
assign LUT_3[7285] = 32'b00000000000000010101000000000111;
assign LUT_3[7286] = 32'b00000000000000010000011100001110;
assign LUT_3[7287] = 32'b00000000000000010111000111101011;
assign LUT_3[7288] = 32'b00000000000000010110011111111010;
assign LUT_3[7289] = 32'b00000000000000011101001011010111;
assign LUT_3[7290] = 32'b00000000000000011000100111011110;
assign LUT_3[7291] = 32'b00000000000000011111010010111011;
assign LUT_3[7292] = 32'b00000000000000010011101101110000;
assign LUT_3[7293] = 32'b00000000000000011010011001001101;
assign LUT_3[7294] = 32'b00000000000000010101110101010100;
assign LUT_3[7295] = 32'b00000000000000011100100000110001;
assign LUT_3[7296] = 32'b00000000000000001110110111100100;
assign LUT_3[7297] = 32'b00000000000000010101100011000001;
assign LUT_3[7298] = 32'b00000000000000010000111111001000;
assign LUT_3[7299] = 32'b00000000000000010111101010100101;
assign LUT_3[7300] = 32'b00000000000000001100000101011010;
assign LUT_3[7301] = 32'b00000000000000010010110000110111;
assign LUT_3[7302] = 32'b00000000000000001110001100111110;
assign LUT_3[7303] = 32'b00000000000000010100111000011011;
assign LUT_3[7304] = 32'b00000000000000010100010000101010;
assign LUT_3[7305] = 32'b00000000000000011010111100000111;
assign LUT_3[7306] = 32'b00000000000000010110011000001110;
assign LUT_3[7307] = 32'b00000000000000011101000011101011;
assign LUT_3[7308] = 32'b00000000000000010001011110100000;
assign LUT_3[7309] = 32'b00000000000000011000001001111101;
assign LUT_3[7310] = 32'b00000000000000010011100110000100;
assign LUT_3[7311] = 32'b00000000000000011010010001100001;
assign LUT_3[7312] = 32'b00000000000000010010001010100111;
assign LUT_3[7313] = 32'b00000000000000011000110110000100;
assign LUT_3[7314] = 32'b00000000000000010100010010001011;
assign LUT_3[7315] = 32'b00000000000000011010111101101000;
assign LUT_3[7316] = 32'b00000000000000001111011000011101;
assign LUT_3[7317] = 32'b00000000000000010110000011111010;
assign LUT_3[7318] = 32'b00000000000000010001100000000001;
assign LUT_3[7319] = 32'b00000000000000011000001011011110;
assign LUT_3[7320] = 32'b00000000000000010111100011101101;
assign LUT_3[7321] = 32'b00000000000000011110001111001010;
assign LUT_3[7322] = 32'b00000000000000011001101011010001;
assign LUT_3[7323] = 32'b00000000000000100000010110101110;
assign LUT_3[7324] = 32'b00000000000000010100110001100011;
assign LUT_3[7325] = 32'b00000000000000011011011101000000;
assign LUT_3[7326] = 32'b00000000000000010110111001000111;
assign LUT_3[7327] = 32'b00000000000000011101100100100100;
assign LUT_3[7328] = 32'b00000000000000010000000110000100;
assign LUT_3[7329] = 32'b00000000000000010110110001100001;
assign LUT_3[7330] = 32'b00000000000000010010001101101000;
assign LUT_3[7331] = 32'b00000000000000011000111001000101;
assign LUT_3[7332] = 32'b00000000000000001101010011111010;
assign LUT_3[7333] = 32'b00000000000000010011111111010111;
assign LUT_3[7334] = 32'b00000000000000001111011011011110;
assign LUT_3[7335] = 32'b00000000000000010110000110111011;
assign LUT_3[7336] = 32'b00000000000000010101011111001010;
assign LUT_3[7337] = 32'b00000000000000011100001010100111;
assign LUT_3[7338] = 32'b00000000000000010111100110101110;
assign LUT_3[7339] = 32'b00000000000000011110010010001011;
assign LUT_3[7340] = 32'b00000000000000010010101101000000;
assign LUT_3[7341] = 32'b00000000000000011001011000011101;
assign LUT_3[7342] = 32'b00000000000000010100110100100100;
assign LUT_3[7343] = 32'b00000000000000011011100000000001;
assign LUT_3[7344] = 32'b00000000000000010011011001000111;
assign LUT_3[7345] = 32'b00000000000000011010000100100100;
assign LUT_3[7346] = 32'b00000000000000010101100000101011;
assign LUT_3[7347] = 32'b00000000000000011100001100001000;
assign LUT_3[7348] = 32'b00000000000000010000100110111101;
assign LUT_3[7349] = 32'b00000000000000010111010010011010;
assign LUT_3[7350] = 32'b00000000000000010010101110100001;
assign LUT_3[7351] = 32'b00000000000000011001011001111110;
assign LUT_3[7352] = 32'b00000000000000011000110010001101;
assign LUT_3[7353] = 32'b00000000000000011111011101101010;
assign LUT_3[7354] = 32'b00000000000000011010111001110001;
assign LUT_3[7355] = 32'b00000000000000100001100101001110;
assign LUT_3[7356] = 32'b00000000000000010110000000000011;
assign LUT_3[7357] = 32'b00000000000000011100101011100000;
assign LUT_3[7358] = 32'b00000000000000011000000111100111;
assign LUT_3[7359] = 32'b00000000000000011110110011000100;
assign LUT_3[7360] = 32'b00000000000000001110110000001111;
assign LUT_3[7361] = 32'b00000000000000010101011011101100;
assign LUT_3[7362] = 32'b00000000000000010000110111110011;
assign LUT_3[7363] = 32'b00000000000000010111100011010000;
assign LUT_3[7364] = 32'b00000000000000001011111110000101;
assign LUT_3[7365] = 32'b00000000000000010010101001100010;
assign LUT_3[7366] = 32'b00000000000000001110000101101001;
assign LUT_3[7367] = 32'b00000000000000010100110001000110;
assign LUT_3[7368] = 32'b00000000000000010100001001010101;
assign LUT_3[7369] = 32'b00000000000000011010110100110010;
assign LUT_3[7370] = 32'b00000000000000010110010000111001;
assign LUT_3[7371] = 32'b00000000000000011100111100010110;
assign LUT_3[7372] = 32'b00000000000000010001010111001011;
assign LUT_3[7373] = 32'b00000000000000011000000010101000;
assign LUT_3[7374] = 32'b00000000000000010011011110101111;
assign LUT_3[7375] = 32'b00000000000000011010001010001100;
assign LUT_3[7376] = 32'b00000000000000010010000011010010;
assign LUT_3[7377] = 32'b00000000000000011000101110101111;
assign LUT_3[7378] = 32'b00000000000000010100001010110110;
assign LUT_3[7379] = 32'b00000000000000011010110110010011;
assign LUT_3[7380] = 32'b00000000000000001111010001001000;
assign LUT_3[7381] = 32'b00000000000000010101111100100101;
assign LUT_3[7382] = 32'b00000000000000010001011000101100;
assign LUT_3[7383] = 32'b00000000000000011000000100001001;
assign LUT_3[7384] = 32'b00000000000000010111011100011000;
assign LUT_3[7385] = 32'b00000000000000011110000111110101;
assign LUT_3[7386] = 32'b00000000000000011001100011111100;
assign LUT_3[7387] = 32'b00000000000000100000001111011001;
assign LUT_3[7388] = 32'b00000000000000010100101010001110;
assign LUT_3[7389] = 32'b00000000000000011011010101101011;
assign LUT_3[7390] = 32'b00000000000000010110110001110010;
assign LUT_3[7391] = 32'b00000000000000011101011101001111;
assign LUT_3[7392] = 32'b00000000000000001111111110101111;
assign LUT_3[7393] = 32'b00000000000000010110101010001100;
assign LUT_3[7394] = 32'b00000000000000010010000110010011;
assign LUT_3[7395] = 32'b00000000000000011000110001110000;
assign LUT_3[7396] = 32'b00000000000000001101001100100101;
assign LUT_3[7397] = 32'b00000000000000010011111000000010;
assign LUT_3[7398] = 32'b00000000000000001111010100001001;
assign LUT_3[7399] = 32'b00000000000000010101111111100110;
assign LUT_3[7400] = 32'b00000000000000010101010111110101;
assign LUT_3[7401] = 32'b00000000000000011100000011010010;
assign LUT_3[7402] = 32'b00000000000000010111011111011001;
assign LUT_3[7403] = 32'b00000000000000011110001010110110;
assign LUT_3[7404] = 32'b00000000000000010010100101101011;
assign LUT_3[7405] = 32'b00000000000000011001010001001000;
assign LUT_3[7406] = 32'b00000000000000010100101101001111;
assign LUT_3[7407] = 32'b00000000000000011011011000101100;
assign LUT_3[7408] = 32'b00000000000000010011010001110010;
assign LUT_3[7409] = 32'b00000000000000011001111101001111;
assign LUT_3[7410] = 32'b00000000000000010101011001010110;
assign LUT_3[7411] = 32'b00000000000000011100000100110011;
assign LUT_3[7412] = 32'b00000000000000010000011111101000;
assign LUT_3[7413] = 32'b00000000000000010111001011000101;
assign LUT_3[7414] = 32'b00000000000000010010100111001100;
assign LUT_3[7415] = 32'b00000000000000011001010010101001;
assign LUT_3[7416] = 32'b00000000000000011000101010111000;
assign LUT_3[7417] = 32'b00000000000000011111010110010101;
assign LUT_3[7418] = 32'b00000000000000011010110010011100;
assign LUT_3[7419] = 32'b00000000000000100001011101111001;
assign LUT_3[7420] = 32'b00000000000000010101111000101110;
assign LUT_3[7421] = 32'b00000000000000011100100100001011;
assign LUT_3[7422] = 32'b00000000000000011000000000010010;
assign LUT_3[7423] = 32'b00000000000000011110101011101111;
assign LUT_3[7424] = 32'b00000000000000001000111100000111;
assign LUT_3[7425] = 32'b00000000000000001111100111100100;
assign LUT_3[7426] = 32'b00000000000000001011000011101011;
assign LUT_3[7427] = 32'b00000000000000010001101111001000;
assign LUT_3[7428] = 32'b00000000000000000110001001111101;
assign LUT_3[7429] = 32'b00000000000000001100110101011010;
assign LUT_3[7430] = 32'b00000000000000001000010001100001;
assign LUT_3[7431] = 32'b00000000000000001110111100111110;
assign LUT_3[7432] = 32'b00000000000000001110010101001101;
assign LUT_3[7433] = 32'b00000000000000010101000000101010;
assign LUT_3[7434] = 32'b00000000000000010000011100110001;
assign LUT_3[7435] = 32'b00000000000000010111001000001110;
assign LUT_3[7436] = 32'b00000000000000001011100011000011;
assign LUT_3[7437] = 32'b00000000000000010010001110100000;
assign LUT_3[7438] = 32'b00000000000000001101101010100111;
assign LUT_3[7439] = 32'b00000000000000010100010110000100;
assign LUT_3[7440] = 32'b00000000000000001100001111001010;
assign LUT_3[7441] = 32'b00000000000000010010111010100111;
assign LUT_3[7442] = 32'b00000000000000001110010110101110;
assign LUT_3[7443] = 32'b00000000000000010101000010001011;
assign LUT_3[7444] = 32'b00000000000000001001011101000000;
assign LUT_3[7445] = 32'b00000000000000010000001000011101;
assign LUT_3[7446] = 32'b00000000000000001011100100100100;
assign LUT_3[7447] = 32'b00000000000000010010010000000001;
assign LUT_3[7448] = 32'b00000000000000010001101000010000;
assign LUT_3[7449] = 32'b00000000000000011000010011101101;
assign LUT_3[7450] = 32'b00000000000000010011101111110100;
assign LUT_3[7451] = 32'b00000000000000011010011011010001;
assign LUT_3[7452] = 32'b00000000000000001110110110000110;
assign LUT_3[7453] = 32'b00000000000000010101100001100011;
assign LUT_3[7454] = 32'b00000000000000010000111101101010;
assign LUT_3[7455] = 32'b00000000000000010111101001000111;
assign LUT_3[7456] = 32'b00000000000000001010001010100111;
assign LUT_3[7457] = 32'b00000000000000010000110110000100;
assign LUT_3[7458] = 32'b00000000000000001100010010001011;
assign LUT_3[7459] = 32'b00000000000000010010111101101000;
assign LUT_3[7460] = 32'b00000000000000000111011000011101;
assign LUT_3[7461] = 32'b00000000000000001110000011111010;
assign LUT_3[7462] = 32'b00000000000000001001100000000001;
assign LUT_3[7463] = 32'b00000000000000010000001011011110;
assign LUT_3[7464] = 32'b00000000000000001111100011101101;
assign LUT_3[7465] = 32'b00000000000000010110001111001010;
assign LUT_3[7466] = 32'b00000000000000010001101011010001;
assign LUT_3[7467] = 32'b00000000000000011000010110101110;
assign LUT_3[7468] = 32'b00000000000000001100110001100011;
assign LUT_3[7469] = 32'b00000000000000010011011101000000;
assign LUT_3[7470] = 32'b00000000000000001110111001000111;
assign LUT_3[7471] = 32'b00000000000000010101100100100100;
assign LUT_3[7472] = 32'b00000000000000001101011101101010;
assign LUT_3[7473] = 32'b00000000000000010100001001000111;
assign LUT_3[7474] = 32'b00000000000000001111100101001110;
assign LUT_3[7475] = 32'b00000000000000010110010000101011;
assign LUT_3[7476] = 32'b00000000000000001010101011100000;
assign LUT_3[7477] = 32'b00000000000000010001010110111101;
assign LUT_3[7478] = 32'b00000000000000001100110011000100;
assign LUT_3[7479] = 32'b00000000000000010011011110100001;
assign LUT_3[7480] = 32'b00000000000000010010110110110000;
assign LUT_3[7481] = 32'b00000000000000011001100010001101;
assign LUT_3[7482] = 32'b00000000000000010100111110010100;
assign LUT_3[7483] = 32'b00000000000000011011101001110001;
assign LUT_3[7484] = 32'b00000000000000010000000100100110;
assign LUT_3[7485] = 32'b00000000000000010110110000000011;
assign LUT_3[7486] = 32'b00000000000000010010001100001010;
assign LUT_3[7487] = 32'b00000000000000011000110111100111;
assign LUT_3[7488] = 32'b00000000000000001000110100110010;
assign LUT_3[7489] = 32'b00000000000000001111100000001111;
assign LUT_3[7490] = 32'b00000000000000001010111100010110;
assign LUT_3[7491] = 32'b00000000000000010001100111110011;
assign LUT_3[7492] = 32'b00000000000000000110000010101000;
assign LUT_3[7493] = 32'b00000000000000001100101110000101;
assign LUT_3[7494] = 32'b00000000000000001000001010001100;
assign LUT_3[7495] = 32'b00000000000000001110110101101001;
assign LUT_3[7496] = 32'b00000000000000001110001101111000;
assign LUT_3[7497] = 32'b00000000000000010100111001010101;
assign LUT_3[7498] = 32'b00000000000000010000010101011100;
assign LUT_3[7499] = 32'b00000000000000010111000000111001;
assign LUT_3[7500] = 32'b00000000000000001011011011101110;
assign LUT_3[7501] = 32'b00000000000000010010000111001011;
assign LUT_3[7502] = 32'b00000000000000001101100011010010;
assign LUT_3[7503] = 32'b00000000000000010100001110101111;
assign LUT_3[7504] = 32'b00000000000000001100000111110101;
assign LUT_3[7505] = 32'b00000000000000010010110011010010;
assign LUT_3[7506] = 32'b00000000000000001110001111011001;
assign LUT_3[7507] = 32'b00000000000000010100111010110110;
assign LUT_3[7508] = 32'b00000000000000001001010101101011;
assign LUT_3[7509] = 32'b00000000000000010000000001001000;
assign LUT_3[7510] = 32'b00000000000000001011011101001111;
assign LUT_3[7511] = 32'b00000000000000010010001000101100;
assign LUT_3[7512] = 32'b00000000000000010001100000111011;
assign LUT_3[7513] = 32'b00000000000000011000001100011000;
assign LUT_3[7514] = 32'b00000000000000010011101000011111;
assign LUT_3[7515] = 32'b00000000000000011010010011111100;
assign LUT_3[7516] = 32'b00000000000000001110101110110001;
assign LUT_3[7517] = 32'b00000000000000010101011010001110;
assign LUT_3[7518] = 32'b00000000000000010000110110010101;
assign LUT_3[7519] = 32'b00000000000000010111100001110010;
assign LUT_3[7520] = 32'b00000000000000001010000011010010;
assign LUT_3[7521] = 32'b00000000000000010000101110101111;
assign LUT_3[7522] = 32'b00000000000000001100001010110110;
assign LUT_3[7523] = 32'b00000000000000010010110110010011;
assign LUT_3[7524] = 32'b00000000000000000111010001001000;
assign LUT_3[7525] = 32'b00000000000000001101111100100101;
assign LUT_3[7526] = 32'b00000000000000001001011000101100;
assign LUT_3[7527] = 32'b00000000000000010000000100001001;
assign LUT_3[7528] = 32'b00000000000000001111011100011000;
assign LUT_3[7529] = 32'b00000000000000010110000111110101;
assign LUT_3[7530] = 32'b00000000000000010001100011111100;
assign LUT_3[7531] = 32'b00000000000000011000001111011001;
assign LUT_3[7532] = 32'b00000000000000001100101010001110;
assign LUT_3[7533] = 32'b00000000000000010011010101101011;
assign LUT_3[7534] = 32'b00000000000000001110110001110010;
assign LUT_3[7535] = 32'b00000000000000010101011101001111;
assign LUT_3[7536] = 32'b00000000000000001101010110010101;
assign LUT_3[7537] = 32'b00000000000000010100000001110010;
assign LUT_3[7538] = 32'b00000000000000001111011101111001;
assign LUT_3[7539] = 32'b00000000000000010110001001010110;
assign LUT_3[7540] = 32'b00000000000000001010100100001011;
assign LUT_3[7541] = 32'b00000000000000010001001111101000;
assign LUT_3[7542] = 32'b00000000000000001100101011101111;
assign LUT_3[7543] = 32'b00000000000000010011010111001100;
assign LUT_3[7544] = 32'b00000000000000010010101111011011;
assign LUT_3[7545] = 32'b00000000000000011001011010111000;
assign LUT_3[7546] = 32'b00000000000000010100110110111111;
assign LUT_3[7547] = 32'b00000000000000011011100010011100;
assign LUT_3[7548] = 32'b00000000000000001111111101010001;
assign LUT_3[7549] = 32'b00000000000000010110101000101110;
assign LUT_3[7550] = 32'b00000000000000010010000100110101;
assign LUT_3[7551] = 32'b00000000000000011000110000010010;
assign LUT_3[7552] = 32'b00000000000000001011000111000101;
assign LUT_3[7553] = 32'b00000000000000010001110010100010;
assign LUT_3[7554] = 32'b00000000000000001101001110101001;
assign LUT_3[7555] = 32'b00000000000000010011111010000110;
assign LUT_3[7556] = 32'b00000000000000001000010100111011;
assign LUT_3[7557] = 32'b00000000000000001111000000011000;
assign LUT_3[7558] = 32'b00000000000000001010011100011111;
assign LUT_3[7559] = 32'b00000000000000010001000111111100;
assign LUT_3[7560] = 32'b00000000000000010000100000001011;
assign LUT_3[7561] = 32'b00000000000000010111001011101000;
assign LUT_3[7562] = 32'b00000000000000010010100111101111;
assign LUT_3[7563] = 32'b00000000000000011001010011001100;
assign LUT_3[7564] = 32'b00000000000000001101101110000001;
assign LUT_3[7565] = 32'b00000000000000010100011001011110;
assign LUT_3[7566] = 32'b00000000000000001111110101100101;
assign LUT_3[7567] = 32'b00000000000000010110100001000010;
assign LUT_3[7568] = 32'b00000000000000001110011010001000;
assign LUT_3[7569] = 32'b00000000000000010101000101100101;
assign LUT_3[7570] = 32'b00000000000000010000100001101100;
assign LUT_3[7571] = 32'b00000000000000010111001101001001;
assign LUT_3[7572] = 32'b00000000000000001011100111111110;
assign LUT_3[7573] = 32'b00000000000000010010010011011011;
assign LUT_3[7574] = 32'b00000000000000001101101111100010;
assign LUT_3[7575] = 32'b00000000000000010100011010111111;
assign LUT_3[7576] = 32'b00000000000000010011110011001110;
assign LUT_3[7577] = 32'b00000000000000011010011110101011;
assign LUT_3[7578] = 32'b00000000000000010101111010110010;
assign LUT_3[7579] = 32'b00000000000000011100100110001111;
assign LUT_3[7580] = 32'b00000000000000010001000001000100;
assign LUT_3[7581] = 32'b00000000000000010111101100100001;
assign LUT_3[7582] = 32'b00000000000000010011001000101000;
assign LUT_3[7583] = 32'b00000000000000011001110100000101;
assign LUT_3[7584] = 32'b00000000000000001100010101100101;
assign LUT_3[7585] = 32'b00000000000000010011000001000010;
assign LUT_3[7586] = 32'b00000000000000001110011101001001;
assign LUT_3[7587] = 32'b00000000000000010101001000100110;
assign LUT_3[7588] = 32'b00000000000000001001100011011011;
assign LUT_3[7589] = 32'b00000000000000010000001110111000;
assign LUT_3[7590] = 32'b00000000000000001011101010111111;
assign LUT_3[7591] = 32'b00000000000000010010010110011100;
assign LUT_3[7592] = 32'b00000000000000010001101110101011;
assign LUT_3[7593] = 32'b00000000000000011000011010001000;
assign LUT_3[7594] = 32'b00000000000000010011110110001111;
assign LUT_3[7595] = 32'b00000000000000011010100001101100;
assign LUT_3[7596] = 32'b00000000000000001110111100100001;
assign LUT_3[7597] = 32'b00000000000000010101100111111110;
assign LUT_3[7598] = 32'b00000000000000010001000100000101;
assign LUT_3[7599] = 32'b00000000000000010111101111100010;
assign LUT_3[7600] = 32'b00000000000000001111101000101000;
assign LUT_3[7601] = 32'b00000000000000010110010100000101;
assign LUT_3[7602] = 32'b00000000000000010001110000001100;
assign LUT_3[7603] = 32'b00000000000000011000011011101001;
assign LUT_3[7604] = 32'b00000000000000001100110110011110;
assign LUT_3[7605] = 32'b00000000000000010011100001111011;
assign LUT_3[7606] = 32'b00000000000000001110111110000010;
assign LUT_3[7607] = 32'b00000000000000010101101001011111;
assign LUT_3[7608] = 32'b00000000000000010101000001101110;
assign LUT_3[7609] = 32'b00000000000000011011101101001011;
assign LUT_3[7610] = 32'b00000000000000010111001001010010;
assign LUT_3[7611] = 32'b00000000000000011101110100101111;
assign LUT_3[7612] = 32'b00000000000000010010001111100100;
assign LUT_3[7613] = 32'b00000000000000011000111011000001;
assign LUT_3[7614] = 32'b00000000000000010100010111001000;
assign LUT_3[7615] = 32'b00000000000000011011000010100101;
assign LUT_3[7616] = 32'b00000000000000001010111111110000;
assign LUT_3[7617] = 32'b00000000000000010001101011001101;
assign LUT_3[7618] = 32'b00000000000000001101000111010100;
assign LUT_3[7619] = 32'b00000000000000010011110010110001;
assign LUT_3[7620] = 32'b00000000000000001000001101100110;
assign LUT_3[7621] = 32'b00000000000000001110111001000011;
assign LUT_3[7622] = 32'b00000000000000001010010101001010;
assign LUT_3[7623] = 32'b00000000000000010001000000100111;
assign LUT_3[7624] = 32'b00000000000000010000011000110110;
assign LUT_3[7625] = 32'b00000000000000010111000100010011;
assign LUT_3[7626] = 32'b00000000000000010010100000011010;
assign LUT_3[7627] = 32'b00000000000000011001001011110111;
assign LUT_3[7628] = 32'b00000000000000001101100110101100;
assign LUT_3[7629] = 32'b00000000000000010100010010001001;
assign LUT_3[7630] = 32'b00000000000000001111101110010000;
assign LUT_3[7631] = 32'b00000000000000010110011001101101;
assign LUT_3[7632] = 32'b00000000000000001110010010110011;
assign LUT_3[7633] = 32'b00000000000000010100111110010000;
assign LUT_3[7634] = 32'b00000000000000010000011010010111;
assign LUT_3[7635] = 32'b00000000000000010111000101110100;
assign LUT_3[7636] = 32'b00000000000000001011100000101001;
assign LUT_3[7637] = 32'b00000000000000010010001100000110;
assign LUT_3[7638] = 32'b00000000000000001101101000001101;
assign LUT_3[7639] = 32'b00000000000000010100010011101010;
assign LUT_3[7640] = 32'b00000000000000010011101011111001;
assign LUT_3[7641] = 32'b00000000000000011010010111010110;
assign LUT_3[7642] = 32'b00000000000000010101110011011101;
assign LUT_3[7643] = 32'b00000000000000011100011110111010;
assign LUT_3[7644] = 32'b00000000000000010000111001101111;
assign LUT_3[7645] = 32'b00000000000000010111100101001100;
assign LUT_3[7646] = 32'b00000000000000010011000001010011;
assign LUT_3[7647] = 32'b00000000000000011001101100110000;
assign LUT_3[7648] = 32'b00000000000000001100001110010000;
assign LUT_3[7649] = 32'b00000000000000010010111001101101;
assign LUT_3[7650] = 32'b00000000000000001110010101110100;
assign LUT_3[7651] = 32'b00000000000000010101000001010001;
assign LUT_3[7652] = 32'b00000000000000001001011100000110;
assign LUT_3[7653] = 32'b00000000000000010000000111100011;
assign LUT_3[7654] = 32'b00000000000000001011100011101010;
assign LUT_3[7655] = 32'b00000000000000010010001111000111;
assign LUT_3[7656] = 32'b00000000000000010001100111010110;
assign LUT_3[7657] = 32'b00000000000000011000010010110011;
assign LUT_3[7658] = 32'b00000000000000010011101110111010;
assign LUT_3[7659] = 32'b00000000000000011010011010010111;
assign LUT_3[7660] = 32'b00000000000000001110110101001100;
assign LUT_3[7661] = 32'b00000000000000010101100000101001;
assign LUT_3[7662] = 32'b00000000000000010000111100110000;
assign LUT_3[7663] = 32'b00000000000000010111101000001101;
assign LUT_3[7664] = 32'b00000000000000001111100001010011;
assign LUT_3[7665] = 32'b00000000000000010110001100110000;
assign LUT_3[7666] = 32'b00000000000000010001101000110111;
assign LUT_3[7667] = 32'b00000000000000011000010100010100;
assign LUT_3[7668] = 32'b00000000000000001100101111001001;
assign LUT_3[7669] = 32'b00000000000000010011011010100110;
assign LUT_3[7670] = 32'b00000000000000001110110110101101;
assign LUT_3[7671] = 32'b00000000000000010101100010001010;
assign LUT_3[7672] = 32'b00000000000000010100111010011001;
assign LUT_3[7673] = 32'b00000000000000011011100101110110;
assign LUT_3[7674] = 32'b00000000000000010111000001111101;
assign LUT_3[7675] = 32'b00000000000000011101101101011010;
assign LUT_3[7676] = 32'b00000000000000010010001000001111;
assign LUT_3[7677] = 32'b00000000000000011000110011101100;
assign LUT_3[7678] = 32'b00000000000000010100001111110011;
assign LUT_3[7679] = 32'b00000000000000011010111011010000;
assign LUT_3[7680] = 32'b00000000000000010000000001110010;
assign LUT_3[7681] = 32'b00000000000000010110101101001111;
assign LUT_3[7682] = 32'b00000000000000010010001001010110;
assign LUT_3[7683] = 32'b00000000000000011000110100110011;
assign LUT_3[7684] = 32'b00000000000000001101001111101000;
assign LUT_3[7685] = 32'b00000000000000010011111011000101;
assign LUT_3[7686] = 32'b00000000000000001111010111001100;
assign LUT_3[7687] = 32'b00000000000000010110000010101001;
assign LUT_3[7688] = 32'b00000000000000010101011010111000;
assign LUT_3[7689] = 32'b00000000000000011100000110010101;
assign LUT_3[7690] = 32'b00000000000000010111100010011100;
assign LUT_3[7691] = 32'b00000000000000011110001101111001;
assign LUT_3[7692] = 32'b00000000000000010010101000101110;
assign LUT_3[7693] = 32'b00000000000000011001010100001011;
assign LUT_3[7694] = 32'b00000000000000010100110000010010;
assign LUT_3[7695] = 32'b00000000000000011011011011101111;
assign LUT_3[7696] = 32'b00000000000000010011010100110101;
assign LUT_3[7697] = 32'b00000000000000011010000000010010;
assign LUT_3[7698] = 32'b00000000000000010101011100011001;
assign LUT_3[7699] = 32'b00000000000000011100000111110110;
assign LUT_3[7700] = 32'b00000000000000010000100010101011;
assign LUT_3[7701] = 32'b00000000000000010111001110001000;
assign LUT_3[7702] = 32'b00000000000000010010101010001111;
assign LUT_3[7703] = 32'b00000000000000011001010101101100;
assign LUT_3[7704] = 32'b00000000000000011000101101111011;
assign LUT_3[7705] = 32'b00000000000000011111011001011000;
assign LUT_3[7706] = 32'b00000000000000011010110101011111;
assign LUT_3[7707] = 32'b00000000000000100001100000111100;
assign LUT_3[7708] = 32'b00000000000000010101111011110001;
assign LUT_3[7709] = 32'b00000000000000011100100111001110;
assign LUT_3[7710] = 32'b00000000000000011000000011010101;
assign LUT_3[7711] = 32'b00000000000000011110101110110010;
assign LUT_3[7712] = 32'b00000000000000010001010000010010;
assign LUT_3[7713] = 32'b00000000000000010111111011101111;
assign LUT_3[7714] = 32'b00000000000000010011010111110110;
assign LUT_3[7715] = 32'b00000000000000011010000011010011;
assign LUT_3[7716] = 32'b00000000000000001110011110001000;
assign LUT_3[7717] = 32'b00000000000000010101001001100101;
assign LUT_3[7718] = 32'b00000000000000010000100101101100;
assign LUT_3[7719] = 32'b00000000000000010111010001001001;
assign LUT_3[7720] = 32'b00000000000000010110101001011000;
assign LUT_3[7721] = 32'b00000000000000011101010100110101;
assign LUT_3[7722] = 32'b00000000000000011000110000111100;
assign LUT_3[7723] = 32'b00000000000000011111011100011001;
assign LUT_3[7724] = 32'b00000000000000010011110111001110;
assign LUT_3[7725] = 32'b00000000000000011010100010101011;
assign LUT_3[7726] = 32'b00000000000000010101111110110010;
assign LUT_3[7727] = 32'b00000000000000011100101010001111;
assign LUT_3[7728] = 32'b00000000000000010100100011010101;
assign LUT_3[7729] = 32'b00000000000000011011001110110010;
assign LUT_3[7730] = 32'b00000000000000010110101010111001;
assign LUT_3[7731] = 32'b00000000000000011101010110010110;
assign LUT_3[7732] = 32'b00000000000000010001110001001011;
assign LUT_3[7733] = 32'b00000000000000011000011100101000;
assign LUT_3[7734] = 32'b00000000000000010011111000101111;
assign LUT_3[7735] = 32'b00000000000000011010100100001100;
assign LUT_3[7736] = 32'b00000000000000011001111100011011;
assign LUT_3[7737] = 32'b00000000000000100000100111111000;
assign LUT_3[7738] = 32'b00000000000000011100000011111111;
assign LUT_3[7739] = 32'b00000000000000100010101111011100;
assign LUT_3[7740] = 32'b00000000000000010111001010010001;
assign LUT_3[7741] = 32'b00000000000000011101110101101110;
assign LUT_3[7742] = 32'b00000000000000011001010001110101;
assign LUT_3[7743] = 32'b00000000000000011111111101010010;
assign LUT_3[7744] = 32'b00000000000000001111111010011101;
assign LUT_3[7745] = 32'b00000000000000010110100101111010;
assign LUT_3[7746] = 32'b00000000000000010010000010000001;
assign LUT_3[7747] = 32'b00000000000000011000101101011110;
assign LUT_3[7748] = 32'b00000000000000001101001000010011;
assign LUT_3[7749] = 32'b00000000000000010011110011110000;
assign LUT_3[7750] = 32'b00000000000000001111001111110111;
assign LUT_3[7751] = 32'b00000000000000010101111011010100;
assign LUT_3[7752] = 32'b00000000000000010101010011100011;
assign LUT_3[7753] = 32'b00000000000000011011111111000000;
assign LUT_3[7754] = 32'b00000000000000010111011011000111;
assign LUT_3[7755] = 32'b00000000000000011110000110100100;
assign LUT_3[7756] = 32'b00000000000000010010100001011001;
assign LUT_3[7757] = 32'b00000000000000011001001100110110;
assign LUT_3[7758] = 32'b00000000000000010100101000111101;
assign LUT_3[7759] = 32'b00000000000000011011010100011010;
assign LUT_3[7760] = 32'b00000000000000010011001101100000;
assign LUT_3[7761] = 32'b00000000000000011001111000111101;
assign LUT_3[7762] = 32'b00000000000000010101010101000100;
assign LUT_3[7763] = 32'b00000000000000011100000000100001;
assign LUT_3[7764] = 32'b00000000000000010000011011010110;
assign LUT_3[7765] = 32'b00000000000000010111000110110011;
assign LUT_3[7766] = 32'b00000000000000010010100010111010;
assign LUT_3[7767] = 32'b00000000000000011001001110010111;
assign LUT_3[7768] = 32'b00000000000000011000100110100110;
assign LUT_3[7769] = 32'b00000000000000011111010010000011;
assign LUT_3[7770] = 32'b00000000000000011010101110001010;
assign LUT_3[7771] = 32'b00000000000000100001011001100111;
assign LUT_3[7772] = 32'b00000000000000010101110100011100;
assign LUT_3[7773] = 32'b00000000000000011100011111111001;
assign LUT_3[7774] = 32'b00000000000000010111111100000000;
assign LUT_3[7775] = 32'b00000000000000011110100111011101;
assign LUT_3[7776] = 32'b00000000000000010001001000111101;
assign LUT_3[7777] = 32'b00000000000000010111110100011010;
assign LUT_3[7778] = 32'b00000000000000010011010000100001;
assign LUT_3[7779] = 32'b00000000000000011001111011111110;
assign LUT_3[7780] = 32'b00000000000000001110010110110011;
assign LUT_3[7781] = 32'b00000000000000010101000010010000;
assign LUT_3[7782] = 32'b00000000000000010000011110010111;
assign LUT_3[7783] = 32'b00000000000000010111001001110100;
assign LUT_3[7784] = 32'b00000000000000010110100010000011;
assign LUT_3[7785] = 32'b00000000000000011101001101100000;
assign LUT_3[7786] = 32'b00000000000000011000101001100111;
assign LUT_3[7787] = 32'b00000000000000011111010101000100;
assign LUT_3[7788] = 32'b00000000000000010011101111111001;
assign LUT_3[7789] = 32'b00000000000000011010011011010110;
assign LUT_3[7790] = 32'b00000000000000010101110111011101;
assign LUT_3[7791] = 32'b00000000000000011100100010111010;
assign LUT_3[7792] = 32'b00000000000000010100011100000000;
assign LUT_3[7793] = 32'b00000000000000011011000111011101;
assign LUT_3[7794] = 32'b00000000000000010110100011100100;
assign LUT_3[7795] = 32'b00000000000000011101001111000001;
assign LUT_3[7796] = 32'b00000000000000010001101001110110;
assign LUT_3[7797] = 32'b00000000000000011000010101010011;
assign LUT_3[7798] = 32'b00000000000000010011110001011010;
assign LUT_3[7799] = 32'b00000000000000011010011100110111;
assign LUT_3[7800] = 32'b00000000000000011001110101000110;
assign LUT_3[7801] = 32'b00000000000000100000100000100011;
assign LUT_3[7802] = 32'b00000000000000011011111100101010;
assign LUT_3[7803] = 32'b00000000000000100010101000000111;
assign LUT_3[7804] = 32'b00000000000000010111000010111100;
assign LUT_3[7805] = 32'b00000000000000011101101110011001;
assign LUT_3[7806] = 32'b00000000000000011001001010100000;
assign LUT_3[7807] = 32'b00000000000000011111110101111101;
assign LUT_3[7808] = 32'b00000000000000010010001100110000;
assign LUT_3[7809] = 32'b00000000000000011000111000001101;
assign LUT_3[7810] = 32'b00000000000000010100010100010100;
assign LUT_3[7811] = 32'b00000000000000011010111111110001;
assign LUT_3[7812] = 32'b00000000000000001111011010100110;
assign LUT_3[7813] = 32'b00000000000000010110000110000011;
assign LUT_3[7814] = 32'b00000000000000010001100010001010;
assign LUT_3[7815] = 32'b00000000000000011000001101100111;
assign LUT_3[7816] = 32'b00000000000000010111100101110110;
assign LUT_3[7817] = 32'b00000000000000011110010001010011;
assign LUT_3[7818] = 32'b00000000000000011001101101011010;
assign LUT_3[7819] = 32'b00000000000000100000011000110111;
assign LUT_3[7820] = 32'b00000000000000010100110011101100;
assign LUT_3[7821] = 32'b00000000000000011011011111001001;
assign LUT_3[7822] = 32'b00000000000000010110111011010000;
assign LUT_3[7823] = 32'b00000000000000011101100110101101;
assign LUT_3[7824] = 32'b00000000000000010101011111110011;
assign LUT_3[7825] = 32'b00000000000000011100001011010000;
assign LUT_3[7826] = 32'b00000000000000010111100111010111;
assign LUT_3[7827] = 32'b00000000000000011110010010110100;
assign LUT_3[7828] = 32'b00000000000000010010101101101001;
assign LUT_3[7829] = 32'b00000000000000011001011001000110;
assign LUT_3[7830] = 32'b00000000000000010100110101001101;
assign LUT_3[7831] = 32'b00000000000000011011100000101010;
assign LUT_3[7832] = 32'b00000000000000011010111000111001;
assign LUT_3[7833] = 32'b00000000000000100001100100010110;
assign LUT_3[7834] = 32'b00000000000000011101000000011101;
assign LUT_3[7835] = 32'b00000000000000100011101011111010;
assign LUT_3[7836] = 32'b00000000000000011000000110101111;
assign LUT_3[7837] = 32'b00000000000000011110110010001100;
assign LUT_3[7838] = 32'b00000000000000011010001110010011;
assign LUT_3[7839] = 32'b00000000000000100000111001110000;
assign LUT_3[7840] = 32'b00000000000000010011011011010000;
assign LUT_3[7841] = 32'b00000000000000011010000110101101;
assign LUT_3[7842] = 32'b00000000000000010101100010110100;
assign LUT_3[7843] = 32'b00000000000000011100001110010001;
assign LUT_3[7844] = 32'b00000000000000010000101001000110;
assign LUT_3[7845] = 32'b00000000000000010111010100100011;
assign LUT_3[7846] = 32'b00000000000000010010110000101010;
assign LUT_3[7847] = 32'b00000000000000011001011100000111;
assign LUT_3[7848] = 32'b00000000000000011000110100010110;
assign LUT_3[7849] = 32'b00000000000000011111011111110011;
assign LUT_3[7850] = 32'b00000000000000011010111011111010;
assign LUT_3[7851] = 32'b00000000000000100001100111010111;
assign LUT_3[7852] = 32'b00000000000000010110000010001100;
assign LUT_3[7853] = 32'b00000000000000011100101101101001;
assign LUT_3[7854] = 32'b00000000000000011000001001110000;
assign LUT_3[7855] = 32'b00000000000000011110110101001101;
assign LUT_3[7856] = 32'b00000000000000010110101110010011;
assign LUT_3[7857] = 32'b00000000000000011101011001110000;
assign LUT_3[7858] = 32'b00000000000000011000110101110111;
assign LUT_3[7859] = 32'b00000000000000011111100001010100;
assign LUT_3[7860] = 32'b00000000000000010011111100001001;
assign LUT_3[7861] = 32'b00000000000000011010100111100110;
assign LUT_3[7862] = 32'b00000000000000010110000011101101;
assign LUT_3[7863] = 32'b00000000000000011100101111001010;
assign LUT_3[7864] = 32'b00000000000000011100000111011001;
assign LUT_3[7865] = 32'b00000000000000100010110010110110;
assign LUT_3[7866] = 32'b00000000000000011110001110111101;
assign LUT_3[7867] = 32'b00000000000000100100111010011010;
assign LUT_3[7868] = 32'b00000000000000011001010101001111;
assign LUT_3[7869] = 32'b00000000000000100000000000101100;
assign LUT_3[7870] = 32'b00000000000000011011011100110011;
assign LUT_3[7871] = 32'b00000000000000100010001000010000;
assign LUT_3[7872] = 32'b00000000000000010010000101011011;
assign LUT_3[7873] = 32'b00000000000000011000110000111000;
assign LUT_3[7874] = 32'b00000000000000010100001100111111;
assign LUT_3[7875] = 32'b00000000000000011010111000011100;
assign LUT_3[7876] = 32'b00000000000000001111010011010001;
assign LUT_3[7877] = 32'b00000000000000010101111110101110;
assign LUT_3[7878] = 32'b00000000000000010001011010110101;
assign LUT_3[7879] = 32'b00000000000000011000000110010010;
assign LUT_3[7880] = 32'b00000000000000010111011110100001;
assign LUT_3[7881] = 32'b00000000000000011110001001111110;
assign LUT_3[7882] = 32'b00000000000000011001100110000101;
assign LUT_3[7883] = 32'b00000000000000100000010001100010;
assign LUT_3[7884] = 32'b00000000000000010100101100010111;
assign LUT_3[7885] = 32'b00000000000000011011010111110100;
assign LUT_3[7886] = 32'b00000000000000010110110011111011;
assign LUT_3[7887] = 32'b00000000000000011101011111011000;
assign LUT_3[7888] = 32'b00000000000000010101011000011110;
assign LUT_3[7889] = 32'b00000000000000011100000011111011;
assign LUT_3[7890] = 32'b00000000000000010111100000000010;
assign LUT_3[7891] = 32'b00000000000000011110001011011111;
assign LUT_3[7892] = 32'b00000000000000010010100110010100;
assign LUT_3[7893] = 32'b00000000000000011001010001110001;
assign LUT_3[7894] = 32'b00000000000000010100101101111000;
assign LUT_3[7895] = 32'b00000000000000011011011001010101;
assign LUT_3[7896] = 32'b00000000000000011010110001100100;
assign LUT_3[7897] = 32'b00000000000000100001011101000001;
assign LUT_3[7898] = 32'b00000000000000011100111001001000;
assign LUT_3[7899] = 32'b00000000000000100011100100100101;
assign LUT_3[7900] = 32'b00000000000000010111111111011010;
assign LUT_3[7901] = 32'b00000000000000011110101010110111;
assign LUT_3[7902] = 32'b00000000000000011010000110111110;
assign LUT_3[7903] = 32'b00000000000000100000110010011011;
assign LUT_3[7904] = 32'b00000000000000010011010011111011;
assign LUT_3[7905] = 32'b00000000000000011001111111011000;
assign LUT_3[7906] = 32'b00000000000000010101011011011111;
assign LUT_3[7907] = 32'b00000000000000011100000110111100;
assign LUT_3[7908] = 32'b00000000000000010000100001110001;
assign LUT_3[7909] = 32'b00000000000000010111001101001110;
assign LUT_3[7910] = 32'b00000000000000010010101001010101;
assign LUT_3[7911] = 32'b00000000000000011001010100110010;
assign LUT_3[7912] = 32'b00000000000000011000101101000001;
assign LUT_3[7913] = 32'b00000000000000011111011000011110;
assign LUT_3[7914] = 32'b00000000000000011010110100100101;
assign LUT_3[7915] = 32'b00000000000000100001100000000010;
assign LUT_3[7916] = 32'b00000000000000010101111010110111;
assign LUT_3[7917] = 32'b00000000000000011100100110010100;
assign LUT_3[7918] = 32'b00000000000000011000000010011011;
assign LUT_3[7919] = 32'b00000000000000011110101101111000;
assign LUT_3[7920] = 32'b00000000000000010110100110111110;
assign LUT_3[7921] = 32'b00000000000000011101010010011011;
assign LUT_3[7922] = 32'b00000000000000011000101110100010;
assign LUT_3[7923] = 32'b00000000000000011111011001111111;
assign LUT_3[7924] = 32'b00000000000000010011110100110100;
assign LUT_3[7925] = 32'b00000000000000011010100000010001;
assign LUT_3[7926] = 32'b00000000000000010101111100011000;
assign LUT_3[7927] = 32'b00000000000000011100100111110101;
assign LUT_3[7928] = 32'b00000000000000011100000000000100;
assign LUT_3[7929] = 32'b00000000000000100010101011100001;
assign LUT_3[7930] = 32'b00000000000000011110000111101000;
assign LUT_3[7931] = 32'b00000000000000100100110011000101;
assign LUT_3[7932] = 32'b00000000000000011001001101111010;
assign LUT_3[7933] = 32'b00000000000000011111111001010111;
assign LUT_3[7934] = 32'b00000000000000011011010101011110;
assign LUT_3[7935] = 32'b00000000000000100010000000111011;
assign LUT_3[7936] = 32'b00000000000000001100010001010011;
assign LUT_3[7937] = 32'b00000000000000010010111100110000;
assign LUT_3[7938] = 32'b00000000000000001110011000110111;
assign LUT_3[7939] = 32'b00000000000000010101000100010100;
assign LUT_3[7940] = 32'b00000000000000001001011111001001;
assign LUT_3[7941] = 32'b00000000000000010000001010100110;
assign LUT_3[7942] = 32'b00000000000000001011100110101101;
assign LUT_3[7943] = 32'b00000000000000010010010010001010;
assign LUT_3[7944] = 32'b00000000000000010001101010011001;
assign LUT_3[7945] = 32'b00000000000000011000010101110110;
assign LUT_3[7946] = 32'b00000000000000010011110001111101;
assign LUT_3[7947] = 32'b00000000000000011010011101011010;
assign LUT_3[7948] = 32'b00000000000000001110111000001111;
assign LUT_3[7949] = 32'b00000000000000010101100011101100;
assign LUT_3[7950] = 32'b00000000000000010000111111110011;
assign LUT_3[7951] = 32'b00000000000000010111101011010000;
assign LUT_3[7952] = 32'b00000000000000001111100100010110;
assign LUT_3[7953] = 32'b00000000000000010110001111110011;
assign LUT_3[7954] = 32'b00000000000000010001101011111010;
assign LUT_3[7955] = 32'b00000000000000011000010111010111;
assign LUT_3[7956] = 32'b00000000000000001100110010001100;
assign LUT_3[7957] = 32'b00000000000000010011011101101001;
assign LUT_3[7958] = 32'b00000000000000001110111001110000;
assign LUT_3[7959] = 32'b00000000000000010101100101001101;
assign LUT_3[7960] = 32'b00000000000000010100111101011100;
assign LUT_3[7961] = 32'b00000000000000011011101000111001;
assign LUT_3[7962] = 32'b00000000000000010111000101000000;
assign LUT_3[7963] = 32'b00000000000000011101110000011101;
assign LUT_3[7964] = 32'b00000000000000010010001011010010;
assign LUT_3[7965] = 32'b00000000000000011000110110101111;
assign LUT_3[7966] = 32'b00000000000000010100010010110110;
assign LUT_3[7967] = 32'b00000000000000011010111110010011;
assign LUT_3[7968] = 32'b00000000000000001101011111110011;
assign LUT_3[7969] = 32'b00000000000000010100001011010000;
assign LUT_3[7970] = 32'b00000000000000001111100111010111;
assign LUT_3[7971] = 32'b00000000000000010110010010110100;
assign LUT_3[7972] = 32'b00000000000000001010101101101001;
assign LUT_3[7973] = 32'b00000000000000010001011001000110;
assign LUT_3[7974] = 32'b00000000000000001100110101001101;
assign LUT_3[7975] = 32'b00000000000000010011100000101010;
assign LUT_3[7976] = 32'b00000000000000010010111000111001;
assign LUT_3[7977] = 32'b00000000000000011001100100010110;
assign LUT_3[7978] = 32'b00000000000000010101000000011101;
assign LUT_3[7979] = 32'b00000000000000011011101011111010;
assign LUT_3[7980] = 32'b00000000000000010000000110101111;
assign LUT_3[7981] = 32'b00000000000000010110110010001100;
assign LUT_3[7982] = 32'b00000000000000010010001110010011;
assign LUT_3[7983] = 32'b00000000000000011000111001110000;
assign LUT_3[7984] = 32'b00000000000000010000110010110110;
assign LUT_3[7985] = 32'b00000000000000010111011110010011;
assign LUT_3[7986] = 32'b00000000000000010010111010011010;
assign LUT_3[7987] = 32'b00000000000000011001100101110111;
assign LUT_3[7988] = 32'b00000000000000001110000000101100;
assign LUT_3[7989] = 32'b00000000000000010100101100001001;
assign LUT_3[7990] = 32'b00000000000000010000001000010000;
assign LUT_3[7991] = 32'b00000000000000010110110011101101;
assign LUT_3[7992] = 32'b00000000000000010110001011111100;
assign LUT_3[7993] = 32'b00000000000000011100110111011001;
assign LUT_3[7994] = 32'b00000000000000011000010011100000;
assign LUT_3[7995] = 32'b00000000000000011110111110111101;
assign LUT_3[7996] = 32'b00000000000000010011011001110010;
assign LUT_3[7997] = 32'b00000000000000011010000101001111;
assign LUT_3[7998] = 32'b00000000000000010101100001010110;
assign LUT_3[7999] = 32'b00000000000000011100001100110011;
assign LUT_3[8000] = 32'b00000000000000001100001001111110;
assign LUT_3[8001] = 32'b00000000000000010010110101011011;
assign LUT_3[8002] = 32'b00000000000000001110010001100010;
assign LUT_3[8003] = 32'b00000000000000010100111100111111;
assign LUT_3[8004] = 32'b00000000000000001001010111110100;
assign LUT_3[8005] = 32'b00000000000000010000000011010001;
assign LUT_3[8006] = 32'b00000000000000001011011111011000;
assign LUT_3[8007] = 32'b00000000000000010010001010110101;
assign LUT_3[8008] = 32'b00000000000000010001100011000100;
assign LUT_3[8009] = 32'b00000000000000011000001110100001;
assign LUT_3[8010] = 32'b00000000000000010011101010101000;
assign LUT_3[8011] = 32'b00000000000000011010010110000101;
assign LUT_3[8012] = 32'b00000000000000001110110000111010;
assign LUT_3[8013] = 32'b00000000000000010101011100010111;
assign LUT_3[8014] = 32'b00000000000000010000111000011110;
assign LUT_3[8015] = 32'b00000000000000010111100011111011;
assign LUT_3[8016] = 32'b00000000000000001111011101000001;
assign LUT_3[8017] = 32'b00000000000000010110001000011110;
assign LUT_3[8018] = 32'b00000000000000010001100100100101;
assign LUT_3[8019] = 32'b00000000000000011000010000000010;
assign LUT_3[8020] = 32'b00000000000000001100101010110111;
assign LUT_3[8021] = 32'b00000000000000010011010110010100;
assign LUT_3[8022] = 32'b00000000000000001110110010011011;
assign LUT_3[8023] = 32'b00000000000000010101011101111000;
assign LUT_3[8024] = 32'b00000000000000010100110110000111;
assign LUT_3[8025] = 32'b00000000000000011011100001100100;
assign LUT_3[8026] = 32'b00000000000000010110111101101011;
assign LUT_3[8027] = 32'b00000000000000011101101001001000;
assign LUT_3[8028] = 32'b00000000000000010010000011111101;
assign LUT_3[8029] = 32'b00000000000000011000101111011010;
assign LUT_3[8030] = 32'b00000000000000010100001011100001;
assign LUT_3[8031] = 32'b00000000000000011010110110111110;
assign LUT_3[8032] = 32'b00000000000000001101011000011110;
assign LUT_3[8033] = 32'b00000000000000010100000011111011;
assign LUT_3[8034] = 32'b00000000000000001111100000000010;
assign LUT_3[8035] = 32'b00000000000000010110001011011111;
assign LUT_3[8036] = 32'b00000000000000001010100110010100;
assign LUT_3[8037] = 32'b00000000000000010001010001110001;
assign LUT_3[8038] = 32'b00000000000000001100101101111000;
assign LUT_3[8039] = 32'b00000000000000010011011001010101;
assign LUT_3[8040] = 32'b00000000000000010010110001100100;
assign LUT_3[8041] = 32'b00000000000000011001011101000001;
assign LUT_3[8042] = 32'b00000000000000010100111001001000;
assign LUT_3[8043] = 32'b00000000000000011011100100100101;
assign LUT_3[8044] = 32'b00000000000000001111111111011010;
assign LUT_3[8045] = 32'b00000000000000010110101010110111;
assign LUT_3[8046] = 32'b00000000000000010010000110111110;
assign LUT_3[8047] = 32'b00000000000000011000110010011011;
assign LUT_3[8048] = 32'b00000000000000010000101011100001;
assign LUT_3[8049] = 32'b00000000000000010111010110111110;
assign LUT_3[8050] = 32'b00000000000000010010110011000101;
assign LUT_3[8051] = 32'b00000000000000011001011110100010;
assign LUT_3[8052] = 32'b00000000000000001101111001010111;
assign LUT_3[8053] = 32'b00000000000000010100100100110100;
assign LUT_3[8054] = 32'b00000000000000010000000000111011;
assign LUT_3[8055] = 32'b00000000000000010110101100011000;
assign LUT_3[8056] = 32'b00000000000000010110000100100111;
assign LUT_3[8057] = 32'b00000000000000011100110000000100;
assign LUT_3[8058] = 32'b00000000000000011000001100001011;
assign LUT_3[8059] = 32'b00000000000000011110110111101000;
assign LUT_3[8060] = 32'b00000000000000010011010010011101;
assign LUT_3[8061] = 32'b00000000000000011001111101111010;
assign LUT_3[8062] = 32'b00000000000000010101011010000001;
assign LUT_3[8063] = 32'b00000000000000011100000101011110;
assign LUT_3[8064] = 32'b00000000000000001110011100010001;
assign LUT_3[8065] = 32'b00000000000000010101000111101110;
assign LUT_3[8066] = 32'b00000000000000010000100011110101;
assign LUT_3[8067] = 32'b00000000000000010111001111010010;
assign LUT_3[8068] = 32'b00000000000000001011101010000111;
assign LUT_3[8069] = 32'b00000000000000010010010101100100;
assign LUT_3[8070] = 32'b00000000000000001101110001101011;
assign LUT_3[8071] = 32'b00000000000000010100011101001000;
assign LUT_3[8072] = 32'b00000000000000010011110101010111;
assign LUT_3[8073] = 32'b00000000000000011010100000110100;
assign LUT_3[8074] = 32'b00000000000000010101111100111011;
assign LUT_3[8075] = 32'b00000000000000011100101000011000;
assign LUT_3[8076] = 32'b00000000000000010001000011001101;
assign LUT_3[8077] = 32'b00000000000000010111101110101010;
assign LUT_3[8078] = 32'b00000000000000010011001010110001;
assign LUT_3[8079] = 32'b00000000000000011001110110001110;
assign LUT_3[8080] = 32'b00000000000000010001101111010100;
assign LUT_3[8081] = 32'b00000000000000011000011010110001;
assign LUT_3[8082] = 32'b00000000000000010011110110111000;
assign LUT_3[8083] = 32'b00000000000000011010100010010101;
assign LUT_3[8084] = 32'b00000000000000001110111101001010;
assign LUT_3[8085] = 32'b00000000000000010101101000100111;
assign LUT_3[8086] = 32'b00000000000000010001000100101110;
assign LUT_3[8087] = 32'b00000000000000010111110000001011;
assign LUT_3[8088] = 32'b00000000000000010111001000011010;
assign LUT_3[8089] = 32'b00000000000000011101110011110111;
assign LUT_3[8090] = 32'b00000000000000011001001111111110;
assign LUT_3[8091] = 32'b00000000000000011111111011011011;
assign LUT_3[8092] = 32'b00000000000000010100010110010000;
assign LUT_3[8093] = 32'b00000000000000011011000001101101;
assign LUT_3[8094] = 32'b00000000000000010110011101110100;
assign LUT_3[8095] = 32'b00000000000000011101001001010001;
assign LUT_3[8096] = 32'b00000000000000001111101010110001;
assign LUT_3[8097] = 32'b00000000000000010110010110001110;
assign LUT_3[8098] = 32'b00000000000000010001110010010101;
assign LUT_3[8099] = 32'b00000000000000011000011101110010;
assign LUT_3[8100] = 32'b00000000000000001100111000100111;
assign LUT_3[8101] = 32'b00000000000000010011100100000100;
assign LUT_3[8102] = 32'b00000000000000001111000000001011;
assign LUT_3[8103] = 32'b00000000000000010101101011101000;
assign LUT_3[8104] = 32'b00000000000000010101000011110111;
assign LUT_3[8105] = 32'b00000000000000011011101111010100;
assign LUT_3[8106] = 32'b00000000000000010111001011011011;
assign LUT_3[8107] = 32'b00000000000000011101110110111000;
assign LUT_3[8108] = 32'b00000000000000010010010001101101;
assign LUT_3[8109] = 32'b00000000000000011000111101001010;
assign LUT_3[8110] = 32'b00000000000000010100011001010001;
assign LUT_3[8111] = 32'b00000000000000011011000100101110;
assign LUT_3[8112] = 32'b00000000000000010010111101110100;
assign LUT_3[8113] = 32'b00000000000000011001101001010001;
assign LUT_3[8114] = 32'b00000000000000010101000101011000;
assign LUT_3[8115] = 32'b00000000000000011011110000110101;
assign LUT_3[8116] = 32'b00000000000000010000001011101010;
assign LUT_3[8117] = 32'b00000000000000010110110111000111;
assign LUT_3[8118] = 32'b00000000000000010010010011001110;
assign LUT_3[8119] = 32'b00000000000000011000111110101011;
assign LUT_3[8120] = 32'b00000000000000011000010110111010;
assign LUT_3[8121] = 32'b00000000000000011111000010010111;
assign LUT_3[8122] = 32'b00000000000000011010011110011110;
assign LUT_3[8123] = 32'b00000000000000100001001001111011;
assign LUT_3[8124] = 32'b00000000000000010101100100110000;
assign LUT_3[8125] = 32'b00000000000000011100010000001101;
assign LUT_3[8126] = 32'b00000000000000010111101100010100;
assign LUT_3[8127] = 32'b00000000000000011110010111110001;
assign LUT_3[8128] = 32'b00000000000000001110010100111100;
assign LUT_3[8129] = 32'b00000000000000010101000000011001;
assign LUT_3[8130] = 32'b00000000000000010000011100100000;
assign LUT_3[8131] = 32'b00000000000000010111000111111101;
assign LUT_3[8132] = 32'b00000000000000001011100010110010;
assign LUT_3[8133] = 32'b00000000000000010010001110001111;
assign LUT_3[8134] = 32'b00000000000000001101101010010110;
assign LUT_3[8135] = 32'b00000000000000010100010101110011;
assign LUT_3[8136] = 32'b00000000000000010011101110000010;
assign LUT_3[8137] = 32'b00000000000000011010011001011111;
assign LUT_3[8138] = 32'b00000000000000010101110101100110;
assign LUT_3[8139] = 32'b00000000000000011100100001000011;
assign LUT_3[8140] = 32'b00000000000000010000111011111000;
assign LUT_3[8141] = 32'b00000000000000010111100111010101;
assign LUT_3[8142] = 32'b00000000000000010011000011011100;
assign LUT_3[8143] = 32'b00000000000000011001101110111001;
assign LUT_3[8144] = 32'b00000000000000010001100111111111;
assign LUT_3[8145] = 32'b00000000000000011000010011011100;
assign LUT_3[8146] = 32'b00000000000000010011101111100011;
assign LUT_3[8147] = 32'b00000000000000011010011011000000;
assign LUT_3[8148] = 32'b00000000000000001110110101110101;
assign LUT_3[8149] = 32'b00000000000000010101100001010010;
assign LUT_3[8150] = 32'b00000000000000010000111101011001;
assign LUT_3[8151] = 32'b00000000000000010111101000110110;
assign LUT_3[8152] = 32'b00000000000000010111000001000101;
assign LUT_3[8153] = 32'b00000000000000011101101100100010;
assign LUT_3[8154] = 32'b00000000000000011001001000101001;
assign LUT_3[8155] = 32'b00000000000000011111110100000110;
assign LUT_3[8156] = 32'b00000000000000010100001110111011;
assign LUT_3[8157] = 32'b00000000000000011010111010011000;
assign LUT_3[8158] = 32'b00000000000000010110010110011111;
assign LUT_3[8159] = 32'b00000000000000011101000001111100;
assign LUT_3[8160] = 32'b00000000000000001111100011011100;
assign LUT_3[8161] = 32'b00000000000000010110001110111001;
assign LUT_3[8162] = 32'b00000000000000010001101011000000;
assign LUT_3[8163] = 32'b00000000000000011000010110011101;
assign LUT_3[8164] = 32'b00000000000000001100110001010010;
assign LUT_3[8165] = 32'b00000000000000010011011100101111;
assign LUT_3[8166] = 32'b00000000000000001110111000110110;
assign LUT_3[8167] = 32'b00000000000000010101100100010011;
assign LUT_3[8168] = 32'b00000000000000010100111100100010;
assign LUT_3[8169] = 32'b00000000000000011011100111111111;
assign LUT_3[8170] = 32'b00000000000000010111000100000110;
assign LUT_3[8171] = 32'b00000000000000011101101111100011;
assign LUT_3[8172] = 32'b00000000000000010010001010011000;
assign LUT_3[8173] = 32'b00000000000000011000110101110101;
assign LUT_3[8174] = 32'b00000000000000010100010001111100;
assign LUT_3[8175] = 32'b00000000000000011010111101011001;
assign LUT_3[8176] = 32'b00000000000000010010110110011111;
assign LUT_3[8177] = 32'b00000000000000011001100001111100;
assign LUT_3[8178] = 32'b00000000000000010100111110000011;
assign LUT_3[8179] = 32'b00000000000000011011101001100000;
assign LUT_3[8180] = 32'b00000000000000010000000100010101;
assign LUT_3[8181] = 32'b00000000000000010110101111110010;
assign LUT_3[8182] = 32'b00000000000000010010001011111001;
assign LUT_3[8183] = 32'b00000000000000011000110111010110;
assign LUT_3[8184] = 32'b00000000000000011000001111100101;
assign LUT_3[8185] = 32'b00000000000000011110111011000010;
assign LUT_3[8186] = 32'b00000000000000011010010111001001;
assign LUT_3[8187] = 32'b00000000000000100001000010100110;
assign LUT_3[8188] = 32'b00000000000000010101011101011011;
assign LUT_3[8189] = 32'b00000000000000011100001000111000;
assign LUT_3[8190] = 32'b00000000000000010111100100111111;
assign LUT_3[8191] = 32'b00000000000000011110010000011100;
assign LUT_3[8192] = 32'b00000000000000000110010101011011;
assign LUT_3[8193] = 32'b00000000000000001101000000111000;
assign LUT_3[8194] = 32'b00000000000000001000011100111111;
assign LUT_3[8195] = 32'b00000000000000001111001000011100;
assign LUT_3[8196] = 32'b00000000000000000011100011010001;
assign LUT_3[8197] = 32'b00000000000000001010001110101110;
assign LUT_3[8198] = 32'b00000000000000000101101010110101;
assign LUT_3[8199] = 32'b00000000000000001100010110010010;
assign LUT_3[8200] = 32'b00000000000000001011101110100001;
assign LUT_3[8201] = 32'b00000000000000010010011001111110;
assign LUT_3[8202] = 32'b00000000000000001101110110000101;
assign LUT_3[8203] = 32'b00000000000000010100100001100010;
assign LUT_3[8204] = 32'b00000000000000001000111100010111;
assign LUT_3[8205] = 32'b00000000000000001111100111110100;
assign LUT_3[8206] = 32'b00000000000000001011000011111011;
assign LUT_3[8207] = 32'b00000000000000010001101111011000;
assign LUT_3[8208] = 32'b00000000000000001001101000011110;
assign LUT_3[8209] = 32'b00000000000000010000010011111011;
assign LUT_3[8210] = 32'b00000000000000001011110000000010;
assign LUT_3[8211] = 32'b00000000000000010010011011011111;
assign LUT_3[8212] = 32'b00000000000000000110110110010100;
assign LUT_3[8213] = 32'b00000000000000001101100001110001;
assign LUT_3[8214] = 32'b00000000000000001000111101111000;
assign LUT_3[8215] = 32'b00000000000000001111101001010101;
assign LUT_3[8216] = 32'b00000000000000001111000001100100;
assign LUT_3[8217] = 32'b00000000000000010101101101000001;
assign LUT_3[8218] = 32'b00000000000000010001001001001000;
assign LUT_3[8219] = 32'b00000000000000010111110100100101;
assign LUT_3[8220] = 32'b00000000000000001100001111011010;
assign LUT_3[8221] = 32'b00000000000000010010111010110111;
assign LUT_3[8222] = 32'b00000000000000001110010110111110;
assign LUT_3[8223] = 32'b00000000000000010101000010011011;
assign LUT_3[8224] = 32'b00000000000000000111100011111011;
assign LUT_3[8225] = 32'b00000000000000001110001111011000;
assign LUT_3[8226] = 32'b00000000000000001001101011011111;
assign LUT_3[8227] = 32'b00000000000000010000010110111100;
assign LUT_3[8228] = 32'b00000000000000000100110001110001;
assign LUT_3[8229] = 32'b00000000000000001011011101001110;
assign LUT_3[8230] = 32'b00000000000000000110111001010101;
assign LUT_3[8231] = 32'b00000000000000001101100100110010;
assign LUT_3[8232] = 32'b00000000000000001100111101000001;
assign LUT_3[8233] = 32'b00000000000000010011101000011110;
assign LUT_3[8234] = 32'b00000000000000001111000100100101;
assign LUT_3[8235] = 32'b00000000000000010101110000000010;
assign LUT_3[8236] = 32'b00000000000000001010001010110111;
assign LUT_3[8237] = 32'b00000000000000010000110110010100;
assign LUT_3[8238] = 32'b00000000000000001100010010011011;
assign LUT_3[8239] = 32'b00000000000000010010111101111000;
assign LUT_3[8240] = 32'b00000000000000001010110110111110;
assign LUT_3[8241] = 32'b00000000000000010001100010011011;
assign LUT_3[8242] = 32'b00000000000000001100111110100010;
assign LUT_3[8243] = 32'b00000000000000010011101001111111;
assign LUT_3[8244] = 32'b00000000000000001000000100110100;
assign LUT_3[8245] = 32'b00000000000000001110110000010001;
assign LUT_3[8246] = 32'b00000000000000001010001100011000;
assign LUT_3[8247] = 32'b00000000000000010000110111110101;
assign LUT_3[8248] = 32'b00000000000000010000010000000100;
assign LUT_3[8249] = 32'b00000000000000010110111011100001;
assign LUT_3[8250] = 32'b00000000000000010010010111101000;
assign LUT_3[8251] = 32'b00000000000000011001000011000101;
assign LUT_3[8252] = 32'b00000000000000001101011101111010;
assign LUT_3[8253] = 32'b00000000000000010100001001010111;
assign LUT_3[8254] = 32'b00000000000000001111100101011110;
assign LUT_3[8255] = 32'b00000000000000010110010000111011;
assign LUT_3[8256] = 32'b00000000000000000110001110000110;
assign LUT_3[8257] = 32'b00000000000000001100111001100011;
assign LUT_3[8258] = 32'b00000000000000001000010101101010;
assign LUT_3[8259] = 32'b00000000000000001111000001000111;
assign LUT_3[8260] = 32'b00000000000000000011011011111100;
assign LUT_3[8261] = 32'b00000000000000001010000111011001;
assign LUT_3[8262] = 32'b00000000000000000101100011100000;
assign LUT_3[8263] = 32'b00000000000000001100001110111101;
assign LUT_3[8264] = 32'b00000000000000001011100111001100;
assign LUT_3[8265] = 32'b00000000000000010010010010101001;
assign LUT_3[8266] = 32'b00000000000000001101101110110000;
assign LUT_3[8267] = 32'b00000000000000010100011010001101;
assign LUT_3[8268] = 32'b00000000000000001000110101000010;
assign LUT_3[8269] = 32'b00000000000000001111100000011111;
assign LUT_3[8270] = 32'b00000000000000001010111100100110;
assign LUT_3[8271] = 32'b00000000000000010001101000000011;
assign LUT_3[8272] = 32'b00000000000000001001100001001001;
assign LUT_3[8273] = 32'b00000000000000010000001100100110;
assign LUT_3[8274] = 32'b00000000000000001011101000101101;
assign LUT_3[8275] = 32'b00000000000000010010010100001010;
assign LUT_3[8276] = 32'b00000000000000000110101110111111;
assign LUT_3[8277] = 32'b00000000000000001101011010011100;
assign LUT_3[8278] = 32'b00000000000000001000110110100011;
assign LUT_3[8279] = 32'b00000000000000001111100010000000;
assign LUT_3[8280] = 32'b00000000000000001110111010001111;
assign LUT_3[8281] = 32'b00000000000000010101100101101100;
assign LUT_3[8282] = 32'b00000000000000010001000001110011;
assign LUT_3[8283] = 32'b00000000000000010111101101010000;
assign LUT_3[8284] = 32'b00000000000000001100001000000101;
assign LUT_3[8285] = 32'b00000000000000010010110011100010;
assign LUT_3[8286] = 32'b00000000000000001110001111101001;
assign LUT_3[8287] = 32'b00000000000000010100111011000110;
assign LUT_3[8288] = 32'b00000000000000000111011100100110;
assign LUT_3[8289] = 32'b00000000000000001110001000000011;
assign LUT_3[8290] = 32'b00000000000000001001100100001010;
assign LUT_3[8291] = 32'b00000000000000010000001111100111;
assign LUT_3[8292] = 32'b00000000000000000100101010011100;
assign LUT_3[8293] = 32'b00000000000000001011010101111001;
assign LUT_3[8294] = 32'b00000000000000000110110010000000;
assign LUT_3[8295] = 32'b00000000000000001101011101011101;
assign LUT_3[8296] = 32'b00000000000000001100110101101100;
assign LUT_3[8297] = 32'b00000000000000010011100001001001;
assign LUT_3[8298] = 32'b00000000000000001110111101010000;
assign LUT_3[8299] = 32'b00000000000000010101101000101101;
assign LUT_3[8300] = 32'b00000000000000001010000011100010;
assign LUT_3[8301] = 32'b00000000000000010000101110111111;
assign LUT_3[8302] = 32'b00000000000000001100001011000110;
assign LUT_3[8303] = 32'b00000000000000010010110110100011;
assign LUT_3[8304] = 32'b00000000000000001010101111101001;
assign LUT_3[8305] = 32'b00000000000000010001011011000110;
assign LUT_3[8306] = 32'b00000000000000001100110111001101;
assign LUT_3[8307] = 32'b00000000000000010011100010101010;
assign LUT_3[8308] = 32'b00000000000000000111111101011111;
assign LUT_3[8309] = 32'b00000000000000001110101000111100;
assign LUT_3[8310] = 32'b00000000000000001010000101000011;
assign LUT_3[8311] = 32'b00000000000000010000110000100000;
assign LUT_3[8312] = 32'b00000000000000010000001000101111;
assign LUT_3[8313] = 32'b00000000000000010110110100001100;
assign LUT_3[8314] = 32'b00000000000000010010010000010011;
assign LUT_3[8315] = 32'b00000000000000011000111011110000;
assign LUT_3[8316] = 32'b00000000000000001101010110100101;
assign LUT_3[8317] = 32'b00000000000000010100000010000010;
assign LUT_3[8318] = 32'b00000000000000001111011110001001;
assign LUT_3[8319] = 32'b00000000000000010110001001100110;
assign LUT_3[8320] = 32'b00000000000000001000100000011001;
assign LUT_3[8321] = 32'b00000000000000001111001011110110;
assign LUT_3[8322] = 32'b00000000000000001010100111111101;
assign LUT_3[8323] = 32'b00000000000000010001010011011010;
assign LUT_3[8324] = 32'b00000000000000000101101110001111;
assign LUT_3[8325] = 32'b00000000000000001100011001101100;
assign LUT_3[8326] = 32'b00000000000000000111110101110011;
assign LUT_3[8327] = 32'b00000000000000001110100001010000;
assign LUT_3[8328] = 32'b00000000000000001101111001011111;
assign LUT_3[8329] = 32'b00000000000000010100100100111100;
assign LUT_3[8330] = 32'b00000000000000010000000001000011;
assign LUT_3[8331] = 32'b00000000000000010110101100100000;
assign LUT_3[8332] = 32'b00000000000000001011000111010101;
assign LUT_3[8333] = 32'b00000000000000010001110010110010;
assign LUT_3[8334] = 32'b00000000000000001101001110111001;
assign LUT_3[8335] = 32'b00000000000000010011111010010110;
assign LUT_3[8336] = 32'b00000000000000001011110011011100;
assign LUT_3[8337] = 32'b00000000000000010010011110111001;
assign LUT_3[8338] = 32'b00000000000000001101111011000000;
assign LUT_3[8339] = 32'b00000000000000010100100110011101;
assign LUT_3[8340] = 32'b00000000000000001001000001010010;
assign LUT_3[8341] = 32'b00000000000000001111101100101111;
assign LUT_3[8342] = 32'b00000000000000001011001000110110;
assign LUT_3[8343] = 32'b00000000000000010001110100010011;
assign LUT_3[8344] = 32'b00000000000000010001001100100010;
assign LUT_3[8345] = 32'b00000000000000010111110111111111;
assign LUT_3[8346] = 32'b00000000000000010011010100000110;
assign LUT_3[8347] = 32'b00000000000000011001111111100011;
assign LUT_3[8348] = 32'b00000000000000001110011010011000;
assign LUT_3[8349] = 32'b00000000000000010101000101110101;
assign LUT_3[8350] = 32'b00000000000000010000100001111100;
assign LUT_3[8351] = 32'b00000000000000010111001101011001;
assign LUT_3[8352] = 32'b00000000000000001001101110111001;
assign LUT_3[8353] = 32'b00000000000000010000011010010110;
assign LUT_3[8354] = 32'b00000000000000001011110110011101;
assign LUT_3[8355] = 32'b00000000000000010010100001111010;
assign LUT_3[8356] = 32'b00000000000000000110111100101111;
assign LUT_3[8357] = 32'b00000000000000001101101000001100;
assign LUT_3[8358] = 32'b00000000000000001001000100010011;
assign LUT_3[8359] = 32'b00000000000000001111101111110000;
assign LUT_3[8360] = 32'b00000000000000001111000111111111;
assign LUT_3[8361] = 32'b00000000000000010101110011011100;
assign LUT_3[8362] = 32'b00000000000000010001001111100011;
assign LUT_3[8363] = 32'b00000000000000010111111011000000;
assign LUT_3[8364] = 32'b00000000000000001100010101110101;
assign LUT_3[8365] = 32'b00000000000000010011000001010010;
assign LUT_3[8366] = 32'b00000000000000001110011101011001;
assign LUT_3[8367] = 32'b00000000000000010101001000110110;
assign LUT_3[8368] = 32'b00000000000000001101000001111100;
assign LUT_3[8369] = 32'b00000000000000010011101101011001;
assign LUT_3[8370] = 32'b00000000000000001111001001100000;
assign LUT_3[8371] = 32'b00000000000000010101110100111101;
assign LUT_3[8372] = 32'b00000000000000001010001111110010;
assign LUT_3[8373] = 32'b00000000000000010000111011001111;
assign LUT_3[8374] = 32'b00000000000000001100010111010110;
assign LUT_3[8375] = 32'b00000000000000010011000010110011;
assign LUT_3[8376] = 32'b00000000000000010010011011000010;
assign LUT_3[8377] = 32'b00000000000000011001000110011111;
assign LUT_3[8378] = 32'b00000000000000010100100010100110;
assign LUT_3[8379] = 32'b00000000000000011011001110000011;
assign LUT_3[8380] = 32'b00000000000000001111101000111000;
assign LUT_3[8381] = 32'b00000000000000010110010100010101;
assign LUT_3[8382] = 32'b00000000000000010001110000011100;
assign LUT_3[8383] = 32'b00000000000000011000011011111001;
assign LUT_3[8384] = 32'b00000000000000001000011001000100;
assign LUT_3[8385] = 32'b00000000000000001111000100100001;
assign LUT_3[8386] = 32'b00000000000000001010100000101000;
assign LUT_3[8387] = 32'b00000000000000010001001100000101;
assign LUT_3[8388] = 32'b00000000000000000101100110111010;
assign LUT_3[8389] = 32'b00000000000000001100010010010111;
assign LUT_3[8390] = 32'b00000000000000000111101110011110;
assign LUT_3[8391] = 32'b00000000000000001110011001111011;
assign LUT_3[8392] = 32'b00000000000000001101110010001010;
assign LUT_3[8393] = 32'b00000000000000010100011101100111;
assign LUT_3[8394] = 32'b00000000000000001111111001101110;
assign LUT_3[8395] = 32'b00000000000000010110100101001011;
assign LUT_3[8396] = 32'b00000000000000001011000000000000;
assign LUT_3[8397] = 32'b00000000000000010001101011011101;
assign LUT_3[8398] = 32'b00000000000000001101000111100100;
assign LUT_3[8399] = 32'b00000000000000010011110011000001;
assign LUT_3[8400] = 32'b00000000000000001011101100000111;
assign LUT_3[8401] = 32'b00000000000000010010010111100100;
assign LUT_3[8402] = 32'b00000000000000001101110011101011;
assign LUT_3[8403] = 32'b00000000000000010100011111001000;
assign LUT_3[8404] = 32'b00000000000000001000111001111101;
assign LUT_3[8405] = 32'b00000000000000001111100101011010;
assign LUT_3[8406] = 32'b00000000000000001011000001100001;
assign LUT_3[8407] = 32'b00000000000000010001101100111110;
assign LUT_3[8408] = 32'b00000000000000010001000101001101;
assign LUT_3[8409] = 32'b00000000000000010111110000101010;
assign LUT_3[8410] = 32'b00000000000000010011001100110001;
assign LUT_3[8411] = 32'b00000000000000011001111000001110;
assign LUT_3[8412] = 32'b00000000000000001110010011000011;
assign LUT_3[8413] = 32'b00000000000000010100111110100000;
assign LUT_3[8414] = 32'b00000000000000010000011010100111;
assign LUT_3[8415] = 32'b00000000000000010111000110000100;
assign LUT_3[8416] = 32'b00000000000000001001100111100100;
assign LUT_3[8417] = 32'b00000000000000010000010011000001;
assign LUT_3[8418] = 32'b00000000000000001011101111001000;
assign LUT_3[8419] = 32'b00000000000000010010011010100101;
assign LUT_3[8420] = 32'b00000000000000000110110101011010;
assign LUT_3[8421] = 32'b00000000000000001101100000110111;
assign LUT_3[8422] = 32'b00000000000000001000111100111110;
assign LUT_3[8423] = 32'b00000000000000001111101000011011;
assign LUT_3[8424] = 32'b00000000000000001111000000101010;
assign LUT_3[8425] = 32'b00000000000000010101101100000111;
assign LUT_3[8426] = 32'b00000000000000010001001000001110;
assign LUT_3[8427] = 32'b00000000000000010111110011101011;
assign LUT_3[8428] = 32'b00000000000000001100001110100000;
assign LUT_3[8429] = 32'b00000000000000010010111001111101;
assign LUT_3[8430] = 32'b00000000000000001110010110000100;
assign LUT_3[8431] = 32'b00000000000000010101000001100001;
assign LUT_3[8432] = 32'b00000000000000001100111010100111;
assign LUT_3[8433] = 32'b00000000000000010011100110000100;
assign LUT_3[8434] = 32'b00000000000000001111000010001011;
assign LUT_3[8435] = 32'b00000000000000010101101101101000;
assign LUT_3[8436] = 32'b00000000000000001010001000011101;
assign LUT_3[8437] = 32'b00000000000000010000110011111010;
assign LUT_3[8438] = 32'b00000000000000001100010000000001;
assign LUT_3[8439] = 32'b00000000000000010010111011011110;
assign LUT_3[8440] = 32'b00000000000000010010010011101101;
assign LUT_3[8441] = 32'b00000000000000011000111111001010;
assign LUT_3[8442] = 32'b00000000000000010100011011010001;
assign LUT_3[8443] = 32'b00000000000000011011000110101110;
assign LUT_3[8444] = 32'b00000000000000001111100001100011;
assign LUT_3[8445] = 32'b00000000000000010110001101000000;
assign LUT_3[8446] = 32'b00000000000000010001101001000111;
assign LUT_3[8447] = 32'b00000000000000011000010100100100;
assign LUT_3[8448] = 32'b00000000000000000010100100111100;
assign LUT_3[8449] = 32'b00000000000000001001010000011001;
assign LUT_3[8450] = 32'b00000000000000000100101100100000;
assign LUT_3[8451] = 32'b00000000000000001011010111111101;
assign LUT_3[8452] = 32'b11111111111111111111110010110010;
assign LUT_3[8453] = 32'b00000000000000000110011110001111;
assign LUT_3[8454] = 32'b00000000000000000001111010010110;
assign LUT_3[8455] = 32'b00000000000000001000100101110011;
assign LUT_3[8456] = 32'b00000000000000000111111110000010;
assign LUT_3[8457] = 32'b00000000000000001110101001011111;
assign LUT_3[8458] = 32'b00000000000000001010000101100110;
assign LUT_3[8459] = 32'b00000000000000010000110001000011;
assign LUT_3[8460] = 32'b00000000000000000101001011111000;
assign LUT_3[8461] = 32'b00000000000000001011110111010101;
assign LUT_3[8462] = 32'b00000000000000000111010011011100;
assign LUT_3[8463] = 32'b00000000000000001101111110111001;
assign LUT_3[8464] = 32'b00000000000000000101110111111111;
assign LUT_3[8465] = 32'b00000000000000001100100011011100;
assign LUT_3[8466] = 32'b00000000000000000111111111100011;
assign LUT_3[8467] = 32'b00000000000000001110101011000000;
assign LUT_3[8468] = 32'b00000000000000000011000101110101;
assign LUT_3[8469] = 32'b00000000000000001001110001010010;
assign LUT_3[8470] = 32'b00000000000000000101001101011001;
assign LUT_3[8471] = 32'b00000000000000001011111000110110;
assign LUT_3[8472] = 32'b00000000000000001011010001000101;
assign LUT_3[8473] = 32'b00000000000000010001111100100010;
assign LUT_3[8474] = 32'b00000000000000001101011000101001;
assign LUT_3[8475] = 32'b00000000000000010100000100000110;
assign LUT_3[8476] = 32'b00000000000000001000011110111011;
assign LUT_3[8477] = 32'b00000000000000001111001010011000;
assign LUT_3[8478] = 32'b00000000000000001010100110011111;
assign LUT_3[8479] = 32'b00000000000000010001010001111100;
assign LUT_3[8480] = 32'b00000000000000000011110011011100;
assign LUT_3[8481] = 32'b00000000000000001010011110111001;
assign LUT_3[8482] = 32'b00000000000000000101111011000000;
assign LUT_3[8483] = 32'b00000000000000001100100110011101;
assign LUT_3[8484] = 32'b00000000000000000001000001010010;
assign LUT_3[8485] = 32'b00000000000000000111101100101111;
assign LUT_3[8486] = 32'b00000000000000000011001000110110;
assign LUT_3[8487] = 32'b00000000000000001001110100010011;
assign LUT_3[8488] = 32'b00000000000000001001001100100010;
assign LUT_3[8489] = 32'b00000000000000001111110111111111;
assign LUT_3[8490] = 32'b00000000000000001011010100000110;
assign LUT_3[8491] = 32'b00000000000000010001111111100011;
assign LUT_3[8492] = 32'b00000000000000000110011010011000;
assign LUT_3[8493] = 32'b00000000000000001101000101110101;
assign LUT_3[8494] = 32'b00000000000000001000100001111100;
assign LUT_3[8495] = 32'b00000000000000001111001101011001;
assign LUT_3[8496] = 32'b00000000000000000111000110011111;
assign LUT_3[8497] = 32'b00000000000000001101110001111100;
assign LUT_3[8498] = 32'b00000000000000001001001110000011;
assign LUT_3[8499] = 32'b00000000000000001111111001100000;
assign LUT_3[8500] = 32'b00000000000000000100010100010101;
assign LUT_3[8501] = 32'b00000000000000001010111111110010;
assign LUT_3[8502] = 32'b00000000000000000110011011111001;
assign LUT_3[8503] = 32'b00000000000000001101000111010110;
assign LUT_3[8504] = 32'b00000000000000001100011111100101;
assign LUT_3[8505] = 32'b00000000000000010011001011000010;
assign LUT_3[8506] = 32'b00000000000000001110100111001001;
assign LUT_3[8507] = 32'b00000000000000010101010010100110;
assign LUT_3[8508] = 32'b00000000000000001001101101011011;
assign LUT_3[8509] = 32'b00000000000000010000011000111000;
assign LUT_3[8510] = 32'b00000000000000001011110100111111;
assign LUT_3[8511] = 32'b00000000000000010010100000011100;
assign LUT_3[8512] = 32'b00000000000000000010011101100111;
assign LUT_3[8513] = 32'b00000000000000001001001001000100;
assign LUT_3[8514] = 32'b00000000000000000100100101001011;
assign LUT_3[8515] = 32'b00000000000000001011010000101000;
assign LUT_3[8516] = 32'b11111111111111111111101011011101;
assign LUT_3[8517] = 32'b00000000000000000110010110111010;
assign LUT_3[8518] = 32'b00000000000000000001110011000001;
assign LUT_3[8519] = 32'b00000000000000001000011110011110;
assign LUT_3[8520] = 32'b00000000000000000111110110101101;
assign LUT_3[8521] = 32'b00000000000000001110100010001010;
assign LUT_3[8522] = 32'b00000000000000001001111110010001;
assign LUT_3[8523] = 32'b00000000000000010000101001101110;
assign LUT_3[8524] = 32'b00000000000000000101000100100011;
assign LUT_3[8525] = 32'b00000000000000001011110000000000;
assign LUT_3[8526] = 32'b00000000000000000111001100000111;
assign LUT_3[8527] = 32'b00000000000000001101110111100100;
assign LUT_3[8528] = 32'b00000000000000000101110000101010;
assign LUT_3[8529] = 32'b00000000000000001100011100000111;
assign LUT_3[8530] = 32'b00000000000000000111111000001110;
assign LUT_3[8531] = 32'b00000000000000001110100011101011;
assign LUT_3[8532] = 32'b00000000000000000010111110100000;
assign LUT_3[8533] = 32'b00000000000000001001101001111101;
assign LUT_3[8534] = 32'b00000000000000000101000110000100;
assign LUT_3[8535] = 32'b00000000000000001011110001100001;
assign LUT_3[8536] = 32'b00000000000000001011001001110000;
assign LUT_3[8537] = 32'b00000000000000010001110101001101;
assign LUT_3[8538] = 32'b00000000000000001101010001010100;
assign LUT_3[8539] = 32'b00000000000000010011111100110001;
assign LUT_3[8540] = 32'b00000000000000001000010111100110;
assign LUT_3[8541] = 32'b00000000000000001111000011000011;
assign LUT_3[8542] = 32'b00000000000000001010011111001010;
assign LUT_3[8543] = 32'b00000000000000010001001010100111;
assign LUT_3[8544] = 32'b00000000000000000011101100000111;
assign LUT_3[8545] = 32'b00000000000000001010010111100100;
assign LUT_3[8546] = 32'b00000000000000000101110011101011;
assign LUT_3[8547] = 32'b00000000000000001100011111001000;
assign LUT_3[8548] = 32'b00000000000000000000111001111101;
assign LUT_3[8549] = 32'b00000000000000000111100101011010;
assign LUT_3[8550] = 32'b00000000000000000011000001100001;
assign LUT_3[8551] = 32'b00000000000000001001101100111110;
assign LUT_3[8552] = 32'b00000000000000001001000101001101;
assign LUT_3[8553] = 32'b00000000000000001111110000101010;
assign LUT_3[8554] = 32'b00000000000000001011001100110001;
assign LUT_3[8555] = 32'b00000000000000010001111000001110;
assign LUT_3[8556] = 32'b00000000000000000110010011000011;
assign LUT_3[8557] = 32'b00000000000000001100111110100000;
assign LUT_3[8558] = 32'b00000000000000001000011010100111;
assign LUT_3[8559] = 32'b00000000000000001111000110000100;
assign LUT_3[8560] = 32'b00000000000000000110111111001010;
assign LUT_3[8561] = 32'b00000000000000001101101010100111;
assign LUT_3[8562] = 32'b00000000000000001001000110101110;
assign LUT_3[8563] = 32'b00000000000000001111110010001011;
assign LUT_3[8564] = 32'b00000000000000000100001101000000;
assign LUT_3[8565] = 32'b00000000000000001010111000011101;
assign LUT_3[8566] = 32'b00000000000000000110010100100100;
assign LUT_3[8567] = 32'b00000000000000001101000000000001;
assign LUT_3[8568] = 32'b00000000000000001100011000010000;
assign LUT_3[8569] = 32'b00000000000000010011000011101101;
assign LUT_3[8570] = 32'b00000000000000001110011111110100;
assign LUT_3[8571] = 32'b00000000000000010101001011010001;
assign LUT_3[8572] = 32'b00000000000000001001100110000110;
assign LUT_3[8573] = 32'b00000000000000010000010001100011;
assign LUT_3[8574] = 32'b00000000000000001011101101101010;
assign LUT_3[8575] = 32'b00000000000000010010011001000111;
assign LUT_3[8576] = 32'b00000000000000000100101111111010;
assign LUT_3[8577] = 32'b00000000000000001011011011010111;
assign LUT_3[8578] = 32'b00000000000000000110110111011110;
assign LUT_3[8579] = 32'b00000000000000001101100010111011;
assign LUT_3[8580] = 32'b00000000000000000001111101110000;
assign LUT_3[8581] = 32'b00000000000000001000101001001101;
assign LUT_3[8582] = 32'b00000000000000000100000101010100;
assign LUT_3[8583] = 32'b00000000000000001010110000110001;
assign LUT_3[8584] = 32'b00000000000000001010001001000000;
assign LUT_3[8585] = 32'b00000000000000010000110100011101;
assign LUT_3[8586] = 32'b00000000000000001100010000100100;
assign LUT_3[8587] = 32'b00000000000000010010111100000001;
assign LUT_3[8588] = 32'b00000000000000000111010110110110;
assign LUT_3[8589] = 32'b00000000000000001110000010010011;
assign LUT_3[8590] = 32'b00000000000000001001011110011010;
assign LUT_3[8591] = 32'b00000000000000010000001001110111;
assign LUT_3[8592] = 32'b00000000000000001000000010111101;
assign LUT_3[8593] = 32'b00000000000000001110101110011010;
assign LUT_3[8594] = 32'b00000000000000001010001010100001;
assign LUT_3[8595] = 32'b00000000000000010000110101111110;
assign LUT_3[8596] = 32'b00000000000000000101010000110011;
assign LUT_3[8597] = 32'b00000000000000001011111100010000;
assign LUT_3[8598] = 32'b00000000000000000111011000010111;
assign LUT_3[8599] = 32'b00000000000000001110000011110100;
assign LUT_3[8600] = 32'b00000000000000001101011100000011;
assign LUT_3[8601] = 32'b00000000000000010100000111100000;
assign LUT_3[8602] = 32'b00000000000000001111100011100111;
assign LUT_3[8603] = 32'b00000000000000010110001111000100;
assign LUT_3[8604] = 32'b00000000000000001010101001111001;
assign LUT_3[8605] = 32'b00000000000000010001010101010110;
assign LUT_3[8606] = 32'b00000000000000001100110001011101;
assign LUT_3[8607] = 32'b00000000000000010011011100111010;
assign LUT_3[8608] = 32'b00000000000000000101111110011010;
assign LUT_3[8609] = 32'b00000000000000001100101001110111;
assign LUT_3[8610] = 32'b00000000000000001000000101111110;
assign LUT_3[8611] = 32'b00000000000000001110110001011011;
assign LUT_3[8612] = 32'b00000000000000000011001100010000;
assign LUT_3[8613] = 32'b00000000000000001001110111101101;
assign LUT_3[8614] = 32'b00000000000000000101010011110100;
assign LUT_3[8615] = 32'b00000000000000001011111111010001;
assign LUT_3[8616] = 32'b00000000000000001011010111100000;
assign LUT_3[8617] = 32'b00000000000000010010000010111101;
assign LUT_3[8618] = 32'b00000000000000001101011111000100;
assign LUT_3[8619] = 32'b00000000000000010100001010100001;
assign LUT_3[8620] = 32'b00000000000000001000100101010110;
assign LUT_3[8621] = 32'b00000000000000001111010000110011;
assign LUT_3[8622] = 32'b00000000000000001010101100111010;
assign LUT_3[8623] = 32'b00000000000000010001011000010111;
assign LUT_3[8624] = 32'b00000000000000001001010001011101;
assign LUT_3[8625] = 32'b00000000000000001111111100111010;
assign LUT_3[8626] = 32'b00000000000000001011011001000001;
assign LUT_3[8627] = 32'b00000000000000010010000100011110;
assign LUT_3[8628] = 32'b00000000000000000110011111010011;
assign LUT_3[8629] = 32'b00000000000000001101001010110000;
assign LUT_3[8630] = 32'b00000000000000001000100110110111;
assign LUT_3[8631] = 32'b00000000000000001111010010010100;
assign LUT_3[8632] = 32'b00000000000000001110101010100011;
assign LUT_3[8633] = 32'b00000000000000010101010110000000;
assign LUT_3[8634] = 32'b00000000000000010000110010000111;
assign LUT_3[8635] = 32'b00000000000000010111011101100100;
assign LUT_3[8636] = 32'b00000000000000001011111000011001;
assign LUT_3[8637] = 32'b00000000000000010010100011110110;
assign LUT_3[8638] = 32'b00000000000000001101111111111101;
assign LUT_3[8639] = 32'b00000000000000010100101011011010;
assign LUT_3[8640] = 32'b00000000000000000100101000100101;
assign LUT_3[8641] = 32'b00000000000000001011010100000010;
assign LUT_3[8642] = 32'b00000000000000000110110000001001;
assign LUT_3[8643] = 32'b00000000000000001101011011100110;
assign LUT_3[8644] = 32'b00000000000000000001110110011011;
assign LUT_3[8645] = 32'b00000000000000001000100001111000;
assign LUT_3[8646] = 32'b00000000000000000011111101111111;
assign LUT_3[8647] = 32'b00000000000000001010101001011100;
assign LUT_3[8648] = 32'b00000000000000001010000001101011;
assign LUT_3[8649] = 32'b00000000000000010000101101001000;
assign LUT_3[8650] = 32'b00000000000000001100001001001111;
assign LUT_3[8651] = 32'b00000000000000010010110100101100;
assign LUT_3[8652] = 32'b00000000000000000111001111100001;
assign LUT_3[8653] = 32'b00000000000000001101111010111110;
assign LUT_3[8654] = 32'b00000000000000001001010111000101;
assign LUT_3[8655] = 32'b00000000000000010000000010100010;
assign LUT_3[8656] = 32'b00000000000000000111111011101000;
assign LUT_3[8657] = 32'b00000000000000001110100111000101;
assign LUT_3[8658] = 32'b00000000000000001010000011001100;
assign LUT_3[8659] = 32'b00000000000000010000101110101001;
assign LUT_3[8660] = 32'b00000000000000000101001001011110;
assign LUT_3[8661] = 32'b00000000000000001011110100111011;
assign LUT_3[8662] = 32'b00000000000000000111010001000010;
assign LUT_3[8663] = 32'b00000000000000001101111100011111;
assign LUT_3[8664] = 32'b00000000000000001101010100101110;
assign LUT_3[8665] = 32'b00000000000000010100000000001011;
assign LUT_3[8666] = 32'b00000000000000001111011100010010;
assign LUT_3[8667] = 32'b00000000000000010110000111101111;
assign LUT_3[8668] = 32'b00000000000000001010100010100100;
assign LUT_3[8669] = 32'b00000000000000010001001110000001;
assign LUT_3[8670] = 32'b00000000000000001100101010001000;
assign LUT_3[8671] = 32'b00000000000000010011010101100101;
assign LUT_3[8672] = 32'b00000000000000000101110111000101;
assign LUT_3[8673] = 32'b00000000000000001100100010100010;
assign LUT_3[8674] = 32'b00000000000000000111111110101001;
assign LUT_3[8675] = 32'b00000000000000001110101010000110;
assign LUT_3[8676] = 32'b00000000000000000011000100111011;
assign LUT_3[8677] = 32'b00000000000000001001110000011000;
assign LUT_3[8678] = 32'b00000000000000000101001100011111;
assign LUT_3[8679] = 32'b00000000000000001011110111111100;
assign LUT_3[8680] = 32'b00000000000000001011010000001011;
assign LUT_3[8681] = 32'b00000000000000010001111011101000;
assign LUT_3[8682] = 32'b00000000000000001101010111101111;
assign LUT_3[8683] = 32'b00000000000000010100000011001100;
assign LUT_3[8684] = 32'b00000000000000001000011110000001;
assign LUT_3[8685] = 32'b00000000000000001111001001011110;
assign LUT_3[8686] = 32'b00000000000000001010100101100101;
assign LUT_3[8687] = 32'b00000000000000010001010001000010;
assign LUT_3[8688] = 32'b00000000000000001001001010001000;
assign LUT_3[8689] = 32'b00000000000000001111110101100101;
assign LUT_3[8690] = 32'b00000000000000001011010001101100;
assign LUT_3[8691] = 32'b00000000000000010001111101001001;
assign LUT_3[8692] = 32'b00000000000000000110010111111110;
assign LUT_3[8693] = 32'b00000000000000001101000011011011;
assign LUT_3[8694] = 32'b00000000000000001000011111100010;
assign LUT_3[8695] = 32'b00000000000000001111001010111111;
assign LUT_3[8696] = 32'b00000000000000001110100011001110;
assign LUT_3[8697] = 32'b00000000000000010101001110101011;
assign LUT_3[8698] = 32'b00000000000000010000101010110010;
assign LUT_3[8699] = 32'b00000000000000010111010110001111;
assign LUT_3[8700] = 32'b00000000000000001011110001000100;
assign LUT_3[8701] = 32'b00000000000000010010011100100001;
assign LUT_3[8702] = 32'b00000000000000001101111000101000;
assign LUT_3[8703] = 32'b00000000000000010100100100000101;
assign LUT_3[8704] = 32'b00000000000000001001101010100111;
assign LUT_3[8705] = 32'b00000000000000010000010110000100;
assign LUT_3[8706] = 32'b00000000000000001011110010001011;
assign LUT_3[8707] = 32'b00000000000000010010011101101000;
assign LUT_3[8708] = 32'b00000000000000000110111000011101;
assign LUT_3[8709] = 32'b00000000000000001101100011111010;
assign LUT_3[8710] = 32'b00000000000000001001000000000001;
assign LUT_3[8711] = 32'b00000000000000001111101011011110;
assign LUT_3[8712] = 32'b00000000000000001111000011101101;
assign LUT_3[8713] = 32'b00000000000000010101101111001010;
assign LUT_3[8714] = 32'b00000000000000010001001011010001;
assign LUT_3[8715] = 32'b00000000000000010111110110101110;
assign LUT_3[8716] = 32'b00000000000000001100010001100011;
assign LUT_3[8717] = 32'b00000000000000010010111101000000;
assign LUT_3[8718] = 32'b00000000000000001110011001000111;
assign LUT_3[8719] = 32'b00000000000000010101000100100100;
assign LUT_3[8720] = 32'b00000000000000001100111101101010;
assign LUT_3[8721] = 32'b00000000000000010011101001000111;
assign LUT_3[8722] = 32'b00000000000000001111000101001110;
assign LUT_3[8723] = 32'b00000000000000010101110000101011;
assign LUT_3[8724] = 32'b00000000000000001010001011100000;
assign LUT_3[8725] = 32'b00000000000000010000110110111101;
assign LUT_3[8726] = 32'b00000000000000001100010011000100;
assign LUT_3[8727] = 32'b00000000000000010010111110100001;
assign LUT_3[8728] = 32'b00000000000000010010010110110000;
assign LUT_3[8729] = 32'b00000000000000011001000010001101;
assign LUT_3[8730] = 32'b00000000000000010100011110010100;
assign LUT_3[8731] = 32'b00000000000000011011001001110001;
assign LUT_3[8732] = 32'b00000000000000001111100100100110;
assign LUT_3[8733] = 32'b00000000000000010110010000000011;
assign LUT_3[8734] = 32'b00000000000000010001101100001010;
assign LUT_3[8735] = 32'b00000000000000011000010111100111;
assign LUT_3[8736] = 32'b00000000000000001010111001000111;
assign LUT_3[8737] = 32'b00000000000000010001100100100100;
assign LUT_3[8738] = 32'b00000000000000001101000000101011;
assign LUT_3[8739] = 32'b00000000000000010011101100001000;
assign LUT_3[8740] = 32'b00000000000000001000000110111101;
assign LUT_3[8741] = 32'b00000000000000001110110010011010;
assign LUT_3[8742] = 32'b00000000000000001010001110100001;
assign LUT_3[8743] = 32'b00000000000000010000111001111110;
assign LUT_3[8744] = 32'b00000000000000010000010010001101;
assign LUT_3[8745] = 32'b00000000000000010110111101101010;
assign LUT_3[8746] = 32'b00000000000000010010011001110001;
assign LUT_3[8747] = 32'b00000000000000011001000101001110;
assign LUT_3[8748] = 32'b00000000000000001101100000000011;
assign LUT_3[8749] = 32'b00000000000000010100001011100000;
assign LUT_3[8750] = 32'b00000000000000001111100111100111;
assign LUT_3[8751] = 32'b00000000000000010110010011000100;
assign LUT_3[8752] = 32'b00000000000000001110001100001010;
assign LUT_3[8753] = 32'b00000000000000010100110111100111;
assign LUT_3[8754] = 32'b00000000000000010000010011101110;
assign LUT_3[8755] = 32'b00000000000000010110111111001011;
assign LUT_3[8756] = 32'b00000000000000001011011010000000;
assign LUT_3[8757] = 32'b00000000000000010010000101011101;
assign LUT_3[8758] = 32'b00000000000000001101100001100100;
assign LUT_3[8759] = 32'b00000000000000010100001101000001;
assign LUT_3[8760] = 32'b00000000000000010011100101010000;
assign LUT_3[8761] = 32'b00000000000000011010010000101101;
assign LUT_3[8762] = 32'b00000000000000010101101100110100;
assign LUT_3[8763] = 32'b00000000000000011100011000010001;
assign LUT_3[8764] = 32'b00000000000000010000110011000110;
assign LUT_3[8765] = 32'b00000000000000010111011110100011;
assign LUT_3[8766] = 32'b00000000000000010010111010101010;
assign LUT_3[8767] = 32'b00000000000000011001100110000111;
assign LUT_3[8768] = 32'b00000000000000001001100011010010;
assign LUT_3[8769] = 32'b00000000000000010000001110101111;
assign LUT_3[8770] = 32'b00000000000000001011101010110110;
assign LUT_3[8771] = 32'b00000000000000010010010110010011;
assign LUT_3[8772] = 32'b00000000000000000110110001001000;
assign LUT_3[8773] = 32'b00000000000000001101011100100101;
assign LUT_3[8774] = 32'b00000000000000001000111000101100;
assign LUT_3[8775] = 32'b00000000000000001111100100001001;
assign LUT_3[8776] = 32'b00000000000000001110111100011000;
assign LUT_3[8777] = 32'b00000000000000010101100111110101;
assign LUT_3[8778] = 32'b00000000000000010001000011111100;
assign LUT_3[8779] = 32'b00000000000000010111101111011001;
assign LUT_3[8780] = 32'b00000000000000001100001010001110;
assign LUT_3[8781] = 32'b00000000000000010010110101101011;
assign LUT_3[8782] = 32'b00000000000000001110010001110010;
assign LUT_3[8783] = 32'b00000000000000010100111101001111;
assign LUT_3[8784] = 32'b00000000000000001100110110010101;
assign LUT_3[8785] = 32'b00000000000000010011100001110010;
assign LUT_3[8786] = 32'b00000000000000001110111101111001;
assign LUT_3[8787] = 32'b00000000000000010101101001010110;
assign LUT_3[8788] = 32'b00000000000000001010000100001011;
assign LUT_3[8789] = 32'b00000000000000010000101111101000;
assign LUT_3[8790] = 32'b00000000000000001100001011101111;
assign LUT_3[8791] = 32'b00000000000000010010110111001100;
assign LUT_3[8792] = 32'b00000000000000010010001111011011;
assign LUT_3[8793] = 32'b00000000000000011000111010111000;
assign LUT_3[8794] = 32'b00000000000000010100010110111111;
assign LUT_3[8795] = 32'b00000000000000011011000010011100;
assign LUT_3[8796] = 32'b00000000000000001111011101010001;
assign LUT_3[8797] = 32'b00000000000000010110001000101110;
assign LUT_3[8798] = 32'b00000000000000010001100100110101;
assign LUT_3[8799] = 32'b00000000000000011000010000010010;
assign LUT_3[8800] = 32'b00000000000000001010110001110010;
assign LUT_3[8801] = 32'b00000000000000010001011101001111;
assign LUT_3[8802] = 32'b00000000000000001100111001010110;
assign LUT_3[8803] = 32'b00000000000000010011100100110011;
assign LUT_3[8804] = 32'b00000000000000000111111111101000;
assign LUT_3[8805] = 32'b00000000000000001110101011000101;
assign LUT_3[8806] = 32'b00000000000000001010000111001100;
assign LUT_3[8807] = 32'b00000000000000010000110010101001;
assign LUT_3[8808] = 32'b00000000000000010000001010111000;
assign LUT_3[8809] = 32'b00000000000000010110110110010101;
assign LUT_3[8810] = 32'b00000000000000010010010010011100;
assign LUT_3[8811] = 32'b00000000000000011000111101111001;
assign LUT_3[8812] = 32'b00000000000000001101011000101110;
assign LUT_3[8813] = 32'b00000000000000010100000100001011;
assign LUT_3[8814] = 32'b00000000000000001111100000010010;
assign LUT_3[8815] = 32'b00000000000000010110001011101111;
assign LUT_3[8816] = 32'b00000000000000001110000100110101;
assign LUT_3[8817] = 32'b00000000000000010100110000010010;
assign LUT_3[8818] = 32'b00000000000000010000001100011001;
assign LUT_3[8819] = 32'b00000000000000010110110111110110;
assign LUT_3[8820] = 32'b00000000000000001011010010101011;
assign LUT_3[8821] = 32'b00000000000000010001111110001000;
assign LUT_3[8822] = 32'b00000000000000001101011010001111;
assign LUT_3[8823] = 32'b00000000000000010100000101101100;
assign LUT_3[8824] = 32'b00000000000000010011011101111011;
assign LUT_3[8825] = 32'b00000000000000011010001001011000;
assign LUT_3[8826] = 32'b00000000000000010101100101011111;
assign LUT_3[8827] = 32'b00000000000000011100010000111100;
assign LUT_3[8828] = 32'b00000000000000010000101011110001;
assign LUT_3[8829] = 32'b00000000000000010111010111001110;
assign LUT_3[8830] = 32'b00000000000000010010110011010101;
assign LUT_3[8831] = 32'b00000000000000011001011110110010;
assign LUT_3[8832] = 32'b00000000000000001011110101100101;
assign LUT_3[8833] = 32'b00000000000000010010100001000010;
assign LUT_3[8834] = 32'b00000000000000001101111101001001;
assign LUT_3[8835] = 32'b00000000000000010100101000100110;
assign LUT_3[8836] = 32'b00000000000000001001000011011011;
assign LUT_3[8837] = 32'b00000000000000001111101110111000;
assign LUT_3[8838] = 32'b00000000000000001011001010111111;
assign LUT_3[8839] = 32'b00000000000000010001110110011100;
assign LUT_3[8840] = 32'b00000000000000010001001110101011;
assign LUT_3[8841] = 32'b00000000000000010111111010001000;
assign LUT_3[8842] = 32'b00000000000000010011010110001111;
assign LUT_3[8843] = 32'b00000000000000011010000001101100;
assign LUT_3[8844] = 32'b00000000000000001110011100100001;
assign LUT_3[8845] = 32'b00000000000000010101000111111110;
assign LUT_3[8846] = 32'b00000000000000010000100100000101;
assign LUT_3[8847] = 32'b00000000000000010111001111100010;
assign LUT_3[8848] = 32'b00000000000000001111001000101000;
assign LUT_3[8849] = 32'b00000000000000010101110100000101;
assign LUT_3[8850] = 32'b00000000000000010001010000001100;
assign LUT_3[8851] = 32'b00000000000000010111111011101001;
assign LUT_3[8852] = 32'b00000000000000001100010110011110;
assign LUT_3[8853] = 32'b00000000000000010011000001111011;
assign LUT_3[8854] = 32'b00000000000000001110011110000010;
assign LUT_3[8855] = 32'b00000000000000010101001001011111;
assign LUT_3[8856] = 32'b00000000000000010100100001101110;
assign LUT_3[8857] = 32'b00000000000000011011001101001011;
assign LUT_3[8858] = 32'b00000000000000010110101001010010;
assign LUT_3[8859] = 32'b00000000000000011101010100101111;
assign LUT_3[8860] = 32'b00000000000000010001101111100100;
assign LUT_3[8861] = 32'b00000000000000011000011011000001;
assign LUT_3[8862] = 32'b00000000000000010011110111001000;
assign LUT_3[8863] = 32'b00000000000000011010100010100101;
assign LUT_3[8864] = 32'b00000000000000001101000100000101;
assign LUT_3[8865] = 32'b00000000000000010011101111100010;
assign LUT_3[8866] = 32'b00000000000000001111001011101001;
assign LUT_3[8867] = 32'b00000000000000010101110111000110;
assign LUT_3[8868] = 32'b00000000000000001010010001111011;
assign LUT_3[8869] = 32'b00000000000000010000111101011000;
assign LUT_3[8870] = 32'b00000000000000001100011001011111;
assign LUT_3[8871] = 32'b00000000000000010011000100111100;
assign LUT_3[8872] = 32'b00000000000000010010011101001011;
assign LUT_3[8873] = 32'b00000000000000011001001000101000;
assign LUT_3[8874] = 32'b00000000000000010100100100101111;
assign LUT_3[8875] = 32'b00000000000000011011010000001100;
assign LUT_3[8876] = 32'b00000000000000001111101011000001;
assign LUT_3[8877] = 32'b00000000000000010110010110011110;
assign LUT_3[8878] = 32'b00000000000000010001110010100101;
assign LUT_3[8879] = 32'b00000000000000011000011110000010;
assign LUT_3[8880] = 32'b00000000000000010000010111001000;
assign LUT_3[8881] = 32'b00000000000000010111000010100101;
assign LUT_3[8882] = 32'b00000000000000010010011110101100;
assign LUT_3[8883] = 32'b00000000000000011001001010001001;
assign LUT_3[8884] = 32'b00000000000000001101100100111110;
assign LUT_3[8885] = 32'b00000000000000010100010000011011;
assign LUT_3[8886] = 32'b00000000000000001111101100100010;
assign LUT_3[8887] = 32'b00000000000000010110010111111111;
assign LUT_3[8888] = 32'b00000000000000010101110000001110;
assign LUT_3[8889] = 32'b00000000000000011100011011101011;
assign LUT_3[8890] = 32'b00000000000000010111110111110010;
assign LUT_3[8891] = 32'b00000000000000011110100011001111;
assign LUT_3[8892] = 32'b00000000000000010010111110000100;
assign LUT_3[8893] = 32'b00000000000000011001101001100001;
assign LUT_3[8894] = 32'b00000000000000010101000101101000;
assign LUT_3[8895] = 32'b00000000000000011011110001000101;
assign LUT_3[8896] = 32'b00000000000000001011101110010000;
assign LUT_3[8897] = 32'b00000000000000010010011001101101;
assign LUT_3[8898] = 32'b00000000000000001101110101110100;
assign LUT_3[8899] = 32'b00000000000000010100100001010001;
assign LUT_3[8900] = 32'b00000000000000001000111100000110;
assign LUT_3[8901] = 32'b00000000000000001111100111100011;
assign LUT_3[8902] = 32'b00000000000000001011000011101010;
assign LUT_3[8903] = 32'b00000000000000010001101111000111;
assign LUT_3[8904] = 32'b00000000000000010001000111010110;
assign LUT_3[8905] = 32'b00000000000000010111110010110011;
assign LUT_3[8906] = 32'b00000000000000010011001110111010;
assign LUT_3[8907] = 32'b00000000000000011001111010010111;
assign LUT_3[8908] = 32'b00000000000000001110010101001100;
assign LUT_3[8909] = 32'b00000000000000010101000000101001;
assign LUT_3[8910] = 32'b00000000000000010000011100110000;
assign LUT_3[8911] = 32'b00000000000000010111001000001101;
assign LUT_3[8912] = 32'b00000000000000001111000001010011;
assign LUT_3[8913] = 32'b00000000000000010101101100110000;
assign LUT_3[8914] = 32'b00000000000000010001001000110111;
assign LUT_3[8915] = 32'b00000000000000010111110100010100;
assign LUT_3[8916] = 32'b00000000000000001100001111001001;
assign LUT_3[8917] = 32'b00000000000000010010111010100110;
assign LUT_3[8918] = 32'b00000000000000001110010110101101;
assign LUT_3[8919] = 32'b00000000000000010101000010001010;
assign LUT_3[8920] = 32'b00000000000000010100011010011001;
assign LUT_3[8921] = 32'b00000000000000011011000101110110;
assign LUT_3[8922] = 32'b00000000000000010110100001111101;
assign LUT_3[8923] = 32'b00000000000000011101001101011010;
assign LUT_3[8924] = 32'b00000000000000010001101000001111;
assign LUT_3[8925] = 32'b00000000000000011000010011101100;
assign LUT_3[8926] = 32'b00000000000000010011101111110011;
assign LUT_3[8927] = 32'b00000000000000011010011011010000;
assign LUT_3[8928] = 32'b00000000000000001100111100110000;
assign LUT_3[8929] = 32'b00000000000000010011101000001101;
assign LUT_3[8930] = 32'b00000000000000001111000100010100;
assign LUT_3[8931] = 32'b00000000000000010101101111110001;
assign LUT_3[8932] = 32'b00000000000000001010001010100110;
assign LUT_3[8933] = 32'b00000000000000010000110110000011;
assign LUT_3[8934] = 32'b00000000000000001100010010001010;
assign LUT_3[8935] = 32'b00000000000000010010111101100111;
assign LUT_3[8936] = 32'b00000000000000010010010101110110;
assign LUT_3[8937] = 32'b00000000000000011001000001010011;
assign LUT_3[8938] = 32'b00000000000000010100011101011010;
assign LUT_3[8939] = 32'b00000000000000011011001000110111;
assign LUT_3[8940] = 32'b00000000000000001111100011101100;
assign LUT_3[8941] = 32'b00000000000000010110001111001001;
assign LUT_3[8942] = 32'b00000000000000010001101011010000;
assign LUT_3[8943] = 32'b00000000000000011000010110101101;
assign LUT_3[8944] = 32'b00000000000000010000001111110011;
assign LUT_3[8945] = 32'b00000000000000010110111011010000;
assign LUT_3[8946] = 32'b00000000000000010010010111010111;
assign LUT_3[8947] = 32'b00000000000000011001000010110100;
assign LUT_3[8948] = 32'b00000000000000001101011101101001;
assign LUT_3[8949] = 32'b00000000000000010100001001000110;
assign LUT_3[8950] = 32'b00000000000000001111100101001101;
assign LUT_3[8951] = 32'b00000000000000010110010000101010;
assign LUT_3[8952] = 32'b00000000000000010101101000111001;
assign LUT_3[8953] = 32'b00000000000000011100010100010110;
assign LUT_3[8954] = 32'b00000000000000010111110000011101;
assign LUT_3[8955] = 32'b00000000000000011110011011111010;
assign LUT_3[8956] = 32'b00000000000000010010110110101111;
assign LUT_3[8957] = 32'b00000000000000011001100010001100;
assign LUT_3[8958] = 32'b00000000000000010100111110010011;
assign LUT_3[8959] = 32'b00000000000000011011101001110000;
assign LUT_3[8960] = 32'b00000000000000000101111010001000;
assign LUT_3[8961] = 32'b00000000000000001100100101100101;
assign LUT_3[8962] = 32'b00000000000000001000000001101100;
assign LUT_3[8963] = 32'b00000000000000001110101101001001;
assign LUT_3[8964] = 32'b00000000000000000011000111111110;
assign LUT_3[8965] = 32'b00000000000000001001110011011011;
assign LUT_3[8966] = 32'b00000000000000000101001111100010;
assign LUT_3[8967] = 32'b00000000000000001011111010111111;
assign LUT_3[8968] = 32'b00000000000000001011010011001110;
assign LUT_3[8969] = 32'b00000000000000010001111110101011;
assign LUT_3[8970] = 32'b00000000000000001101011010110010;
assign LUT_3[8971] = 32'b00000000000000010100000110001111;
assign LUT_3[8972] = 32'b00000000000000001000100001000100;
assign LUT_3[8973] = 32'b00000000000000001111001100100001;
assign LUT_3[8974] = 32'b00000000000000001010101000101000;
assign LUT_3[8975] = 32'b00000000000000010001010100000101;
assign LUT_3[8976] = 32'b00000000000000001001001101001011;
assign LUT_3[8977] = 32'b00000000000000001111111000101000;
assign LUT_3[8978] = 32'b00000000000000001011010100101111;
assign LUT_3[8979] = 32'b00000000000000010010000000001100;
assign LUT_3[8980] = 32'b00000000000000000110011011000001;
assign LUT_3[8981] = 32'b00000000000000001101000110011110;
assign LUT_3[8982] = 32'b00000000000000001000100010100101;
assign LUT_3[8983] = 32'b00000000000000001111001110000010;
assign LUT_3[8984] = 32'b00000000000000001110100110010001;
assign LUT_3[8985] = 32'b00000000000000010101010001101110;
assign LUT_3[8986] = 32'b00000000000000010000101101110101;
assign LUT_3[8987] = 32'b00000000000000010111011001010010;
assign LUT_3[8988] = 32'b00000000000000001011110100000111;
assign LUT_3[8989] = 32'b00000000000000010010011111100100;
assign LUT_3[8990] = 32'b00000000000000001101111011101011;
assign LUT_3[8991] = 32'b00000000000000010100100111001000;
assign LUT_3[8992] = 32'b00000000000000000111001000101000;
assign LUT_3[8993] = 32'b00000000000000001101110100000101;
assign LUT_3[8994] = 32'b00000000000000001001010000001100;
assign LUT_3[8995] = 32'b00000000000000001111111011101001;
assign LUT_3[8996] = 32'b00000000000000000100010110011110;
assign LUT_3[8997] = 32'b00000000000000001011000001111011;
assign LUT_3[8998] = 32'b00000000000000000110011110000010;
assign LUT_3[8999] = 32'b00000000000000001101001001011111;
assign LUT_3[9000] = 32'b00000000000000001100100001101110;
assign LUT_3[9001] = 32'b00000000000000010011001101001011;
assign LUT_3[9002] = 32'b00000000000000001110101001010010;
assign LUT_3[9003] = 32'b00000000000000010101010100101111;
assign LUT_3[9004] = 32'b00000000000000001001101111100100;
assign LUT_3[9005] = 32'b00000000000000010000011011000001;
assign LUT_3[9006] = 32'b00000000000000001011110111001000;
assign LUT_3[9007] = 32'b00000000000000010010100010100101;
assign LUT_3[9008] = 32'b00000000000000001010011011101011;
assign LUT_3[9009] = 32'b00000000000000010001000111001000;
assign LUT_3[9010] = 32'b00000000000000001100100011001111;
assign LUT_3[9011] = 32'b00000000000000010011001110101100;
assign LUT_3[9012] = 32'b00000000000000000111101001100001;
assign LUT_3[9013] = 32'b00000000000000001110010100111110;
assign LUT_3[9014] = 32'b00000000000000001001110001000101;
assign LUT_3[9015] = 32'b00000000000000010000011100100010;
assign LUT_3[9016] = 32'b00000000000000001111110100110001;
assign LUT_3[9017] = 32'b00000000000000010110100000001110;
assign LUT_3[9018] = 32'b00000000000000010001111100010101;
assign LUT_3[9019] = 32'b00000000000000011000100111110010;
assign LUT_3[9020] = 32'b00000000000000001101000010100111;
assign LUT_3[9021] = 32'b00000000000000010011101110000100;
assign LUT_3[9022] = 32'b00000000000000001111001010001011;
assign LUT_3[9023] = 32'b00000000000000010101110101101000;
assign LUT_3[9024] = 32'b00000000000000000101110010110011;
assign LUT_3[9025] = 32'b00000000000000001100011110010000;
assign LUT_3[9026] = 32'b00000000000000000111111010010111;
assign LUT_3[9027] = 32'b00000000000000001110100101110100;
assign LUT_3[9028] = 32'b00000000000000000011000000101001;
assign LUT_3[9029] = 32'b00000000000000001001101100000110;
assign LUT_3[9030] = 32'b00000000000000000101001000001101;
assign LUT_3[9031] = 32'b00000000000000001011110011101010;
assign LUT_3[9032] = 32'b00000000000000001011001011111001;
assign LUT_3[9033] = 32'b00000000000000010001110111010110;
assign LUT_3[9034] = 32'b00000000000000001101010011011101;
assign LUT_3[9035] = 32'b00000000000000010011111110111010;
assign LUT_3[9036] = 32'b00000000000000001000011001101111;
assign LUT_3[9037] = 32'b00000000000000001111000101001100;
assign LUT_3[9038] = 32'b00000000000000001010100001010011;
assign LUT_3[9039] = 32'b00000000000000010001001100110000;
assign LUT_3[9040] = 32'b00000000000000001001000101110110;
assign LUT_3[9041] = 32'b00000000000000001111110001010011;
assign LUT_3[9042] = 32'b00000000000000001011001101011010;
assign LUT_3[9043] = 32'b00000000000000010001111000110111;
assign LUT_3[9044] = 32'b00000000000000000110010011101100;
assign LUT_3[9045] = 32'b00000000000000001100111111001001;
assign LUT_3[9046] = 32'b00000000000000001000011011010000;
assign LUT_3[9047] = 32'b00000000000000001111000110101101;
assign LUT_3[9048] = 32'b00000000000000001110011110111100;
assign LUT_3[9049] = 32'b00000000000000010101001010011001;
assign LUT_3[9050] = 32'b00000000000000010000100110100000;
assign LUT_3[9051] = 32'b00000000000000010111010001111101;
assign LUT_3[9052] = 32'b00000000000000001011101100110010;
assign LUT_3[9053] = 32'b00000000000000010010011000001111;
assign LUT_3[9054] = 32'b00000000000000001101110100010110;
assign LUT_3[9055] = 32'b00000000000000010100011111110011;
assign LUT_3[9056] = 32'b00000000000000000111000001010011;
assign LUT_3[9057] = 32'b00000000000000001101101100110000;
assign LUT_3[9058] = 32'b00000000000000001001001000110111;
assign LUT_3[9059] = 32'b00000000000000001111110100010100;
assign LUT_3[9060] = 32'b00000000000000000100001111001001;
assign LUT_3[9061] = 32'b00000000000000001010111010100110;
assign LUT_3[9062] = 32'b00000000000000000110010110101101;
assign LUT_3[9063] = 32'b00000000000000001101000010001010;
assign LUT_3[9064] = 32'b00000000000000001100011010011001;
assign LUT_3[9065] = 32'b00000000000000010011000101110110;
assign LUT_3[9066] = 32'b00000000000000001110100001111101;
assign LUT_3[9067] = 32'b00000000000000010101001101011010;
assign LUT_3[9068] = 32'b00000000000000001001101000001111;
assign LUT_3[9069] = 32'b00000000000000010000010011101100;
assign LUT_3[9070] = 32'b00000000000000001011101111110011;
assign LUT_3[9071] = 32'b00000000000000010010011011010000;
assign LUT_3[9072] = 32'b00000000000000001010010100010110;
assign LUT_3[9073] = 32'b00000000000000010000111111110011;
assign LUT_3[9074] = 32'b00000000000000001100011011111010;
assign LUT_3[9075] = 32'b00000000000000010011000111010111;
assign LUT_3[9076] = 32'b00000000000000000111100010001100;
assign LUT_3[9077] = 32'b00000000000000001110001101101001;
assign LUT_3[9078] = 32'b00000000000000001001101001110000;
assign LUT_3[9079] = 32'b00000000000000010000010101001101;
assign LUT_3[9080] = 32'b00000000000000001111101101011100;
assign LUT_3[9081] = 32'b00000000000000010110011000111001;
assign LUT_3[9082] = 32'b00000000000000010001110101000000;
assign LUT_3[9083] = 32'b00000000000000011000100000011101;
assign LUT_3[9084] = 32'b00000000000000001100111011010010;
assign LUT_3[9085] = 32'b00000000000000010011100110101111;
assign LUT_3[9086] = 32'b00000000000000001111000010110110;
assign LUT_3[9087] = 32'b00000000000000010101101110010011;
assign LUT_3[9088] = 32'b00000000000000001000000101000110;
assign LUT_3[9089] = 32'b00000000000000001110110000100011;
assign LUT_3[9090] = 32'b00000000000000001010001100101010;
assign LUT_3[9091] = 32'b00000000000000010000111000000111;
assign LUT_3[9092] = 32'b00000000000000000101010010111100;
assign LUT_3[9093] = 32'b00000000000000001011111110011001;
assign LUT_3[9094] = 32'b00000000000000000111011010100000;
assign LUT_3[9095] = 32'b00000000000000001110000101111101;
assign LUT_3[9096] = 32'b00000000000000001101011110001100;
assign LUT_3[9097] = 32'b00000000000000010100001001101001;
assign LUT_3[9098] = 32'b00000000000000001111100101110000;
assign LUT_3[9099] = 32'b00000000000000010110010001001101;
assign LUT_3[9100] = 32'b00000000000000001010101100000010;
assign LUT_3[9101] = 32'b00000000000000010001010111011111;
assign LUT_3[9102] = 32'b00000000000000001100110011100110;
assign LUT_3[9103] = 32'b00000000000000010011011111000011;
assign LUT_3[9104] = 32'b00000000000000001011011000001001;
assign LUT_3[9105] = 32'b00000000000000010010000011100110;
assign LUT_3[9106] = 32'b00000000000000001101011111101101;
assign LUT_3[9107] = 32'b00000000000000010100001011001010;
assign LUT_3[9108] = 32'b00000000000000001000100101111111;
assign LUT_3[9109] = 32'b00000000000000001111010001011100;
assign LUT_3[9110] = 32'b00000000000000001010101101100011;
assign LUT_3[9111] = 32'b00000000000000010001011001000000;
assign LUT_3[9112] = 32'b00000000000000010000110001001111;
assign LUT_3[9113] = 32'b00000000000000010111011100101100;
assign LUT_3[9114] = 32'b00000000000000010010111000110011;
assign LUT_3[9115] = 32'b00000000000000011001100100010000;
assign LUT_3[9116] = 32'b00000000000000001101111111000101;
assign LUT_3[9117] = 32'b00000000000000010100101010100010;
assign LUT_3[9118] = 32'b00000000000000010000000110101001;
assign LUT_3[9119] = 32'b00000000000000010110110010000110;
assign LUT_3[9120] = 32'b00000000000000001001010011100110;
assign LUT_3[9121] = 32'b00000000000000001111111111000011;
assign LUT_3[9122] = 32'b00000000000000001011011011001010;
assign LUT_3[9123] = 32'b00000000000000010010000110100111;
assign LUT_3[9124] = 32'b00000000000000000110100001011100;
assign LUT_3[9125] = 32'b00000000000000001101001100111001;
assign LUT_3[9126] = 32'b00000000000000001000101001000000;
assign LUT_3[9127] = 32'b00000000000000001111010100011101;
assign LUT_3[9128] = 32'b00000000000000001110101100101100;
assign LUT_3[9129] = 32'b00000000000000010101011000001001;
assign LUT_3[9130] = 32'b00000000000000010000110100010000;
assign LUT_3[9131] = 32'b00000000000000010111011111101101;
assign LUT_3[9132] = 32'b00000000000000001011111010100010;
assign LUT_3[9133] = 32'b00000000000000010010100101111111;
assign LUT_3[9134] = 32'b00000000000000001110000010000110;
assign LUT_3[9135] = 32'b00000000000000010100101101100011;
assign LUT_3[9136] = 32'b00000000000000001100100110101001;
assign LUT_3[9137] = 32'b00000000000000010011010010000110;
assign LUT_3[9138] = 32'b00000000000000001110101110001101;
assign LUT_3[9139] = 32'b00000000000000010101011001101010;
assign LUT_3[9140] = 32'b00000000000000001001110100011111;
assign LUT_3[9141] = 32'b00000000000000010000011111111100;
assign LUT_3[9142] = 32'b00000000000000001011111100000011;
assign LUT_3[9143] = 32'b00000000000000010010100111100000;
assign LUT_3[9144] = 32'b00000000000000010001111111101111;
assign LUT_3[9145] = 32'b00000000000000011000101011001100;
assign LUT_3[9146] = 32'b00000000000000010100000111010011;
assign LUT_3[9147] = 32'b00000000000000011010110010110000;
assign LUT_3[9148] = 32'b00000000000000001111001101100101;
assign LUT_3[9149] = 32'b00000000000000010101111001000010;
assign LUT_3[9150] = 32'b00000000000000010001010101001001;
assign LUT_3[9151] = 32'b00000000000000011000000000100110;
assign LUT_3[9152] = 32'b00000000000000000111111101110001;
assign LUT_3[9153] = 32'b00000000000000001110101001001110;
assign LUT_3[9154] = 32'b00000000000000001010000101010101;
assign LUT_3[9155] = 32'b00000000000000010000110000110010;
assign LUT_3[9156] = 32'b00000000000000000101001011100111;
assign LUT_3[9157] = 32'b00000000000000001011110111000100;
assign LUT_3[9158] = 32'b00000000000000000111010011001011;
assign LUT_3[9159] = 32'b00000000000000001101111110101000;
assign LUT_3[9160] = 32'b00000000000000001101010110110111;
assign LUT_3[9161] = 32'b00000000000000010100000010010100;
assign LUT_3[9162] = 32'b00000000000000001111011110011011;
assign LUT_3[9163] = 32'b00000000000000010110001001111000;
assign LUT_3[9164] = 32'b00000000000000001010100100101101;
assign LUT_3[9165] = 32'b00000000000000010001010000001010;
assign LUT_3[9166] = 32'b00000000000000001100101100010001;
assign LUT_3[9167] = 32'b00000000000000010011010111101110;
assign LUT_3[9168] = 32'b00000000000000001011010000110100;
assign LUT_3[9169] = 32'b00000000000000010001111100010001;
assign LUT_3[9170] = 32'b00000000000000001101011000011000;
assign LUT_3[9171] = 32'b00000000000000010100000011110101;
assign LUT_3[9172] = 32'b00000000000000001000011110101010;
assign LUT_3[9173] = 32'b00000000000000001111001010000111;
assign LUT_3[9174] = 32'b00000000000000001010100110001110;
assign LUT_3[9175] = 32'b00000000000000010001010001101011;
assign LUT_3[9176] = 32'b00000000000000010000101001111010;
assign LUT_3[9177] = 32'b00000000000000010111010101010111;
assign LUT_3[9178] = 32'b00000000000000010010110001011110;
assign LUT_3[9179] = 32'b00000000000000011001011100111011;
assign LUT_3[9180] = 32'b00000000000000001101110111110000;
assign LUT_3[9181] = 32'b00000000000000010100100011001101;
assign LUT_3[9182] = 32'b00000000000000001111111111010100;
assign LUT_3[9183] = 32'b00000000000000010110101010110001;
assign LUT_3[9184] = 32'b00000000000000001001001100010001;
assign LUT_3[9185] = 32'b00000000000000001111110111101110;
assign LUT_3[9186] = 32'b00000000000000001011010011110101;
assign LUT_3[9187] = 32'b00000000000000010001111111010010;
assign LUT_3[9188] = 32'b00000000000000000110011010000111;
assign LUT_3[9189] = 32'b00000000000000001101000101100100;
assign LUT_3[9190] = 32'b00000000000000001000100001101011;
assign LUT_3[9191] = 32'b00000000000000001111001101001000;
assign LUT_3[9192] = 32'b00000000000000001110100101010111;
assign LUT_3[9193] = 32'b00000000000000010101010000110100;
assign LUT_3[9194] = 32'b00000000000000010000101100111011;
assign LUT_3[9195] = 32'b00000000000000010111011000011000;
assign LUT_3[9196] = 32'b00000000000000001011110011001101;
assign LUT_3[9197] = 32'b00000000000000010010011110101010;
assign LUT_3[9198] = 32'b00000000000000001101111010110001;
assign LUT_3[9199] = 32'b00000000000000010100100110001110;
assign LUT_3[9200] = 32'b00000000000000001100011111010100;
assign LUT_3[9201] = 32'b00000000000000010011001010110001;
assign LUT_3[9202] = 32'b00000000000000001110100110111000;
assign LUT_3[9203] = 32'b00000000000000010101010010010101;
assign LUT_3[9204] = 32'b00000000000000001001101101001010;
assign LUT_3[9205] = 32'b00000000000000010000011000100111;
assign LUT_3[9206] = 32'b00000000000000001011110100101110;
assign LUT_3[9207] = 32'b00000000000000010010100000001011;
assign LUT_3[9208] = 32'b00000000000000010001111000011010;
assign LUT_3[9209] = 32'b00000000000000011000100011110111;
assign LUT_3[9210] = 32'b00000000000000010011111111111110;
assign LUT_3[9211] = 32'b00000000000000011010101011011011;
assign LUT_3[9212] = 32'b00000000000000001111000110010000;
assign LUT_3[9213] = 32'b00000000000000010101110001101101;
assign LUT_3[9214] = 32'b00000000000000010001001101110100;
assign LUT_3[9215] = 32'b00000000000000010111111001010001;
assign LUT_3[9216] = 32'b00000000000000001100111010011000;
assign LUT_3[9217] = 32'b00000000000000010011100101110101;
assign LUT_3[9218] = 32'b00000000000000001111000001111100;
assign LUT_3[9219] = 32'b00000000000000010101101101011001;
assign LUT_3[9220] = 32'b00000000000000001010001000001110;
assign LUT_3[9221] = 32'b00000000000000010000110011101011;
assign LUT_3[9222] = 32'b00000000000000001100001111110010;
assign LUT_3[9223] = 32'b00000000000000010010111011001111;
assign LUT_3[9224] = 32'b00000000000000010010010011011110;
assign LUT_3[9225] = 32'b00000000000000011000111110111011;
assign LUT_3[9226] = 32'b00000000000000010100011011000010;
assign LUT_3[9227] = 32'b00000000000000011011000110011111;
assign LUT_3[9228] = 32'b00000000000000001111100001010100;
assign LUT_3[9229] = 32'b00000000000000010110001100110001;
assign LUT_3[9230] = 32'b00000000000000010001101000111000;
assign LUT_3[9231] = 32'b00000000000000011000010100010101;
assign LUT_3[9232] = 32'b00000000000000010000001101011011;
assign LUT_3[9233] = 32'b00000000000000010110111000111000;
assign LUT_3[9234] = 32'b00000000000000010010010100111111;
assign LUT_3[9235] = 32'b00000000000000011001000000011100;
assign LUT_3[9236] = 32'b00000000000000001101011011010001;
assign LUT_3[9237] = 32'b00000000000000010100000110101110;
assign LUT_3[9238] = 32'b00000000000000001111100010110101;
assign LUT_3[9239] = 32'b00000000000000010110001110010010;
assign LUT_3[9240] = 32'b00000000000000010101100110100001;
assign LUT_3[9241] = 32'b00000000000000011100010001111110;
assign LUT_3[9242] = 32'b00000000000000010111101110000101;
assign LUT_3[9243] = 32'b00000000000000011110011001100010;
assign LUT_3[9244] = 32'b00000000000000010010110100010111;
assign LUT_3[9245] = 32'b00000000000000011001011111110100;
assign LUT_3[9246] = 32'b00000000000000010100111011111011;
assign LUT_3[9247] = 32'b00000000000000011011100111011000;
assign LUT_3[9248] = 32'b00000000000000001110001000111000;
assign LUT_3[9249] = 32'b00000000000000010100110100010101;
assign LUT_3[9250] = 32'b00000000000000010000010000011100;
assign LUT_3[9251] = 32'b00000000000000010110111011111001;
assign LUT_3[9252] = 32'b00000000000000001011010110101110;
assign LUT_3[9253] = 32'b00000000000000010010000010001011;
assign LUT_3[9254] = 32'b00000000000000001101011110010010;
assign LUT_3[9255] = 32'b00000000000000010100001001101111;
assign LUT_3[9256] = 32'b00000000000000010011100001111110;
assign LUT_3[9257] = 32'b00000000000000011010001101011011;
assign LUT_3[9258] = 32'b00000000000000010101101001100010;
assign LUT_3[9259] = 32'b00000000000000011100010100111111;
assign LUT_3[9260] = 32'b00000000000000010000101111110100;
assign LUT_3[9261] = 32'b00000000000000010111011011010001;
assign LUT_3[9262] = 32'b00000000000000010010110111011000;
assign LUT_3[9263] = 32'b00000000000000011001100010110101;
assign LUT_3[9264] = 32'b00000000000000010001011011111011;
assign LUT_3[9265] = 32'b00000000000000011000000111011000;
assign LUT_3[9266] = 32'b00000000000000010011100011011111;
assign LUT_3[9267] = 32'b00000000000000011010001110111100;
assign LUT_3[9268] = 32'b00000000000000001110101001110001;
assign LUT_3[9269] = 32'b00000000000000010101010101001110;
assign LUT_3[9270] = 32'b00000000000000010000110001010101;
assign LUT_3[9271] = 32'b00000000000000010111011100110010;
assign LUT_3[9272] = 32'b00000000000000010110110101000001;
assign LUT_3[9273] = 32'b00000000000000011101100000011110;
assign LUT_3[9274] = 32'b00000000000000011000111100100101;
assign LUT_3[9275] = 32'b00000000000000011111101000000010;
assign LUT_3[9276] = 32'b00000000000000010100000010110111;
assign LUT_3[9277] = 32'b00000000000000011010101110010100;
assign LUT_3[9278] = 32'b00000000000000010110001010011011;
assign LUT_3[9279] = 32'b00000000000000011100110101111000;
assign LUT_3[9280] = 32'b00000000000000001100110011000011;
assign LUT_3[9281] = 32'b00000000000000010011011110100000;
assign LUT_3[9282] = 32'b00000000000000001110111010100111;
assign LUT_3[9283] = 32'b00000000000000010101100110000100;
assign LUT_3[9284] = 32'b00000000000000001010000000111001;
assign LUT_3[9285] = 32'b00000000000000010000101100010110;
assign LUT_3[9286] = 32'b00000000000000001100001000011101;
assign LUT_3[9287] = 32'b00000000000000010010110011111010;
assign LUT_3[9288] = 32'b00000000000000010010001100001001;
assign LUT_3[9289] = 32'b00000000000000011000110111100110;
assign LUT_3[9290] = 32'b00000000000000010100010011101101;
assign LUT_3[9291] = 32'b00000000000000011010111111001010;
assign LUT_3[9292] = 32'b00000000000000001111011001111111;
assign LUT_3[9293] = 32'b00000000000000010110000101011100;
assign LUT_3[9294] = 32'b00000000000000010001100001100011;
assign LUT_3[9295] = 32'b00000000000000011000001101000000;
assign LUT_3[9296] = 32'b00000000000000010000000110000110;
assign LUT_3[9297] = 32'b00000000000000010110110001100011;
assign LUT_3[9298] = 32'b00000000000000010010001101101010;
assign LUT_3[9299] = 32'b00000000000000011000111001000111;
assign LUT_3[9300] = 32'b00000000000000001101010011111100;
assign LUT_3[9301] = 32'b00000000000000010011111111011001;
assign LUT_3[9302] = 32'b00000000000000001111011011100000;
assign LUT_3[9303] = 32'b00000000000000010110000110111101;
assign LUT_3[9304] = 32'b00000000000000010101011111001100;
assign LUT_3[9305] = 32'b00000000000000011100001010101001;
assign LUT_3[9306] = 32'b00000000000000010111100110110000;
assign LUT_3[9307] = 32'b00000000000000011110010010001101;
assign LUT_3[9308] = 32'b00000000000000010010101101000010;
assign LUT_3[9309] = 32'b00000000000000011001011000011111;
assign LUT_3[9310] = 32'b00000000000000010100110100100110;
assign LUT_3[9311] = 32'b00000000000000011011100000000011;
assign LUT_3[9312] = 32'b00000000000000001110000001100011;
assign LUT_3[9313] = 32'b00000000000000010100101101000000;
assign LUT_3[9314] = 32'b00000000000000010000001001000111;
assign LUT_3[9315] = 32'b00000000000000010110110100100100;
assign LUT_3[9316] = 32'b00000000000000001011001111011001;
assign LUT_3[9317] = 32'b00000000000000010001111010110110;
assign LUT_3[9318] = 32'b00000000000000001101010110111101;
assign LUT_3[9319] = 32'b00000000000000010100000010011010;
assign LUT_3[9320] = 32'b00000000000000010011011010101001;
assign LUT_3[9321] = 32'b00000000000000011010000110000110;
assign LUT_3[9322] = 32'b00000000000000010101100010001101;
assign LUT_3[9323] = 32'b00000000000000011100001101101010;
assign LUT_3[9324] = 32'b00000000000000010000101000011111;
assign LUT_3[9325] = 32'b00000000000000010111010011111100;
assign LUT_3[9326] = 32'b00000000000000010010110000000011;
assign LUT_3[9327] = 32'b00000000000000011001011011100000;
assign LUT_3[9328] = 32'b00000000000000010001010100100110;
assign LUT_3[9329] = 32'b00000000000000011000000000000011;
assign LUT_3[9330] = 32'b00000000000000010011011100001010;
assign LUT_3[9331] = 32'b00000000000000011010000111100111;
assign LUT_3[9332] = 32'b00000000000000001110100010011100;
assign LUT_3[9333] = 32'b00000000000000010101001101111001;
assign LUT_3[9334] = 32'b00000000000000010000101010000000;
assign LUT_3[9335] = 32'b00000000000000010111010101011101;
assign LUT_3[9336] = 32'b00000000000000010110101101101100;
assign LUT_3[9337] = 32'b00000000000000011101011001001001;
assign LUT_3[9338] = 32'b00000000000000011000110101010000;
assign LUT_3[9339] = 32'b00000000000000011111100000101101;
assign LUT_3[9340] = 32'b00000000000000010011111011100010;
assign LUT_3[9341] = 32'b00000000000000011010100110111111;
assign LUT_3[9342] = 32'b00000000000000010110000011000110;
assign LUT_3[9343] = 32'b00000000000000011100101110100011;
assign LUT_3[9344] = 32'b00000000000000001111000101010110;
assign LUT_3[9345] = 32'b00000000000000010101110000110011;
assign LUT_3[9346] = 32'b00000000000000010001001100111010;
assign LUT_3[9347] = 32'b00000000000000010111111000010111;
assign LUT_3[9348] = 32'b00000000000000001100010011001100;
assign LUT_3[9349] = 32'b00000000000000010010111110101001;
assign LUT_3[9350] = 32'b00000000000000001110011010110000;
assign LUT_3[9351] = 32'b00000000000000010101000110001101;
assign LUT_3[9352] = 32'b00000000000000010100011110011100;
assign LUT_3[9353] = 32'b00000000000000011011001001111001;
assign LUT_3[9354] = 32'b00000000000000010110100110000000;
assign LUT_3[9355] = 32'b00000000000000011101010001011101;
assign LUT_3[9356] = 32'b00000000000000010001101100010010;
assign LUT_3[9357] = 32'b00000000000000011000010111101111;
assign LUT_3[9358] = 32'b00000000000000010011110011110110;
assign LUT_3[9359] = 32'b00000000000000011010011111010011;
assign LUT_3[9360] = 32'b00000000000000010010011000011001;
assign LUT_3[9361] = 32'b00000000000000011001000011110110;
assign LUT_3[9362] = 32'b00000000000000010100011111111101;
assign LUT_3[9363] = 32'b00000000000000011011001011011010;
assign LUT_3[9364] = 32'b00000000000000001111100110001111;
assign LUT_3[9365] = 32'b00000000000000010110010001101100;
assign LUT_3[9366] = 32'b00000000000000010001101101110011;
assign LUT_3[9367] = 32'b00000000000000011000011001010000;
assign LUT_3[9368] = 32'b00000000000000010111110001011111;
assign LUT_3[9369] = 32'b00000000000000011110011100111100;
assign LUT_3[9370] = 32'b00000000000000011001111001000011;
assign LUT_3[9371] = 32'b00000000000000100000100100100000;
assign LUT_3[9372] = 32'b00000000000000010100111111010101;
assign LUT_3[9373] = 32'b00000000000000011011101010110010;
assign LUT_3[9374] = 32'b00000000000000010111000110111001;
assign LUT_3[9375] = 32'b00000000000000011101110010010110;
assign LUT_3[9376] = 32'b00000000000000010000010011110110;
assign LUT_3[9377] = 32'b00000000000000010110111111010011;
assign LUT_3[9378] = 32'b00000000000000010010011011011010;
assign LUT_3[9379] = 32'b00000000000000011001000110110111;
assign LUT_3[9380] = 32'b00000000000000001101100001101100;
assign LUT_3[9381] = 32'b00000000000000010100001101001001;
assign LUT_3[9382] = 32'b00000000000000001111101001010000;
assign LUT_3[9383] = 32'b00000000000000010110010100101101;
assign LUT_3[9384] = 32'b00000000000000010101101100111100;
assign LUT_3[9385] = 32'b00000000000000011100011000011001;
assign LUT_3[9386] = 32'b00000000000000010111110100100000;
assign LUT_3[9387] = 32'b00000000000000011110011111111101;
assign LUT_3[9388] = 32'b00000000000000010010111010110010;
assign LUT_3[9389] = 32'b00000000000000011001100110001111;
assign LUT_3[9390] = 32'b00000000000000010101000010010110;
assign LUT_3[9391] = 32'b00000000000000011011101101110011;
assign LUT_3[9392] = 32'b00000000000000010011100110111001;
assign LUT_3[9393] = 32'b00000000000000011010010010010110;
assign LUT_3[9394] = 32'b00000000000000010101101110011101;
assign LUT_3[9395] = 32'b00000000000000011100011001111010;
assign LUT_3[9396] = 32'b00000000000000010000110100101111;
assign LUT_3[9397] = 32'b00000000000000010111100000001100;
assign LUT_3[9398] = 32'b00000000000000010010111100010011;
assign LUT_3[9399] = 32'b00000000000000011001100111110000;
assign LUT_3[9400] = 32'b00000000000000011000111111111111;
assign LUT_3[9401] = 32'b00000000000000011111101011011100;
assign LUT_3[9402] = 32'b00000000000000011011000111100011;
assign LUT_3[9403] = 32'b00000000000000100001110011000000;
assign LUT_3[9404] = 32'b00000000000000010110001101110101;
assign LUT_3[9405] = 32'b00000000000000011100111001010010;
assign LUT_3[9406] = 32'b00000000000000011000010101011001;
assign LUT_3[9407] = 32'b00000000000000011111000000110110;
assign LUT_3[9408] = 32'b00000000000000001110111110000001;
assign LUT_3[9409] = 32'b00000000000000010101101001011110;
assign LUT_3[9410] = 32'b00000000000000010001000101100101;
assign LUT_3[9411] = 32'b00000000000000010111110001000010;
assign LUT_3[9412] = 32'b00000000000000001100001011110111;
assign LUT_3[9413] = 32'b00000000000000010010110111010100;
assign LUT_3[9414] = 32'b00000000000000001110010011011011;
assign LUT_3[9415] = 32'b00000000000000010100111110111000;
assign LUT_3[9416] = 32'b00000000000000010100010111000111;
assign LUT_3[9417] = 32'b00000000000000011011000010100100;
assign LUT_3[9418] = 32'b00000000000000010110011110101011;
assign LUT_3[9419] = 32'b00000000000000011101001010001000;
assign LUT_3[9420] = 32'b00000000000000010001100100111101;
assign LUT_3[9421] = 32'b00000000000000011000010000011010;
assign LUT_3[9422] = 32'b00000000000000010011101100100001;
assign LUT_3[9423] = 32'b00000000000000011010010111111110;
assign LUT_3[9424] = 32'b00000000000000010010010001000100;
assign LUT_3[9425] = 32'b00000000000000011000111100100001;
assign LUT_3[9426] = 32'b00000000000000010100011000101000;
assign LUT_3[9427] = 32'b00000000000000011011000100000101;
assign LUT_3[9428] = 32'b00000000000000001111011110111010;
assign LUT_3[9429] = 32'b00000000000000010110001010010111;
assign LUT_3[9430] = 32'b00000000000000010001100110011110;
assign LUT_3[9431] = 32'b00000000000000011000010001111011;
assign LUT_3[9432] = 32'b00000000000000010111101010001010;
assign LUT_3[9433] = 32'b00000000000000011110010101100111;
assign LUT_3[9434] = 32'b00000000000000011001110001101110;
assign LUT_3[9435] = 32'b00000000000000100000011101001011;
assign LUT_3[9436] = 32'b00000000000000010100111000000000;
assign LUT_3[9437] = 32'b00000000000000011011100011011101;
assign LUT_3[9438] = 32'b00000000000000010110111111100100;
assign LUT_3[9439] = 32'b00000000000000011101101011000001;
assign LUT_3[9440] = 32'b00000000000000010000001100100001;
assign LUT_3[9441] = 32'b00000000000000010110110111111110;
assign LUT_3[9442] = 32'b00000000000000010010010100000101;
assign LUT_3[9443] = 32'b00000000000000011000111111100010;
assign LUT_3[9444] = 32'b00000000000000001101011010010111;
assign LUT_3[9445] = 32'b00000000000000010100000101110100;
assign LUT_3[9446] = 32'b00000000000000001111100001111011;
assign LUT_3[9447] = 32'b00000000000000010110001101011000;
assign LUT_3[9448] = 32'b00000000000000010101100101100111;
assign LUT_3[9449] = 32'b00000000000000011100010001000100;
assign LUT_3[9450] = 32'b00000000000000010111101101001011;
assign LUT_3[9451] = 32'b00000000000000011110011000101000;
assign LUT_3[9452] = 32'b00000000000000010010110011011101;
assign LUT_3[9453] = 32'b00000000000000011001011110111010;
assign LUT_3[9454] = 32'b00000000000000010100111011000001;
assign LUT_3[9455] = 32'b00000000000000011011100110011110;
assign LUT_3[9456] = 32'b00000000000000010011011111100100;
assign LUT_3[9457] = 32'b00000000000000011010001011000001;
assign LUT_3[9458] = 32'b00000000000000010101100111001000;
assign LUT_3[9459] = 32'b00000000000000011100010010100101;
assign LUT_3[9460] = 32'b00000000000000010000101101011010;
assign LUT_3[9461] = 32'b00000000000000010111011000110111;
assign LUT_3[9462] = 32'b00000000000000010010110100111110;
assign LUT_3[9463] = 32'b00000000000000011001100000011011;
assign LUT_3[9464] = 32'b00000000000000011000111000101010;
assign LUT_3[9465] = 32'b00000000000000011111100100000111;
assign LUT_3[9466] = 32'b00000000000000011011000000001110;
assign LUT_3[9467] = 32'b00000000000000100001101011101011;
assign LUT_3[9468] = 32'b00000000000000010110000110100000;
assign LUT_3[9469] = 32'b00000000000000011100110001111101;
assign LUT_3[9470] = 32'b00000000000000011000001110000100;
assign LUT_3[9471] = 32'b00000000000000011110111001100001;
assign LUT_3[9472] = 32'b00000000000000001001001001111001;
assign LUT_3[9473] = 32'b00000000000000001111110101010110;
assign LUT_3[9474] = 32'b00000000000000001011010001011101;
assign LUT_3[9475] = 32'b00000000000000010001111100111010;
assign LUT_3[9476] = 32'b00000000000000000110010111101111;
assign LUT_3[9477] = 32'b00000000000000001101000011001100;
assign LUT_3[9478] = 32'b00000000000000001000011111010011;
assign LUT_3[9479] = 32'b00000000000000001111001010110000;
assign LUT_3[9480] = 32'b00000000000000001110100010111111;
assign LUT_3[9481] = 32'b00000000000000010101001110011100;
assign LUT_3[9482] = 32'b00000000000000010000101010100011;
assign LUT_3[9483] = 32'b00000000000000010111010110000000;
assign LUT_3[9484] = 32'b00000000000000001011110000110101;
assign LUT_3[9485] = 32'b00000000000000010010011100010010;
assign LUT_3[9486] = 32'b00000000000000001101111000011001;
assign LUT_3[9487] = 32'b00000000000000010100100011110110;
assign LUT_3[9488] = 32'b00000000000000001100011100111100;
assign LUT_3[9489] = 32'b00000000000000010011001000011001;
assign LUT_3[9490] = 32'b00000000000000001110100100100000;
assign LUT_3[9491] = 32'b00000000000000010101001111111101;
assign LUT_3[9492] = 32'b00000000000000001001101010110010;
assign LUT_3[9493] = 32'b00000000000000010000010110001111;
assign LUT_3[9494] = 32'b00000000000000001011110010010110;
assign LUT_3[9495] = 32'b00000000000000010010011101110011;
assign LUT_3[9496] = 32'b00000000000000010001110110000010;
assign LUT_3[9497] = 32'b00000000000000011000100001011111;
assign LUT_3[9498] = 32'b00000000000000010011111101100110;
assign LUT_3[9499] = 32'b00000000000000011010101001000011;
assign LUT_3[9500] = 32'b00000000000000001111000011111000;
assign LUT_3[9501] = 32'b00000000000000010101101111010101;
assign LUT_3[9502] = 32'b00000000000000010001001011011100;
assign LUT_3[9503] = 32'b00000000000000010111110110111001;
assign LUT_3[9504] = 32'b00000000000000001010011000011001;
assign LUT_3[9505] = 32'b00000000000000010001000011110110;
assign LUT_3[9506] = 32'b00000000000000001100011111111101;
assign LUT_3[9507] = 32'b00000000000000010011001011011010;
assign LUT_3[9508] = 32'b00000000000000000111100110001111;
assign LUT_3[9509] = 32'b00000000000000001110010001101100;
assign LUT_3[9510] = 32'b00000000000000001001101101110011;
assign LUT_3[9511] = 32'b00000000000000010000011001010000;
assign LUT_3[9512] = 32'b00000000000000001111110001011111;
assign LUT_3[9513] = 32'b00000000000000010110011100111100;
assign LUT_3[9514] = 32'b00000000000000010001111001000011;
assign LUT_3[9515] = 32'b00000000000000011000100100100000;
assign LUT_3[9516] = 32'b00000000000000001100111111010101;
assign LUT_3[9517] = 32'b00000000000000010011101010110010;
assign LUT_3[9518] = 32'b00000000000000001111000110111001;
assign LUT_3[9519] = 32'b00000000000000010101110010010110;
assign LUT_3[9520] = 32'b00000000000000001101101011011100;
assign LUT_3[9521] = 32'b00000000000000010100010110111001;
assign LUT_3[9522] = 32'b00000000000000001111110011000000;
assign LUT_3[9523] = 32'b00000000000000010110011110011101;
assign LUT_3[9524] = 32'b00000000000000001010111001010010;
assign LUT_3[9525] = 32'b00000000000000010001100100101111;
assign LUT_3[9526] = 32'b00000000000000001101000000110110;
assign LUT_3[9527] = 32'b00000000000000010011101100010011;
assign LUT_3[9528] = 32'b00000000000000010011000100100010;
assign LUT_3[9529] = 32'b00000000000000011001101111111111;
assign LUT_3[9530] = 32'b00000000000000010101001100000110;
assign LUT_3[9531] = 32'b00000000000000011011110111100011;
assign LUT_3[9532] = 32'b00000000000000010000010010011000;
assign LUT_3[9533] = 32'b00000000000000010110111101110101;
assign LUT_3[9534] = 32'b00000000000000010010011001111100;
assign LUT_3[9535] = 32'b00000000000000011001000101011001;
assign LUT_3[9536] = 32'b00000000000000001001000010100100;
assign LUT_3[9537] = 32'b00000000000000001111101110000001;
assign LUT_3[9538] = 32'b00000000000000001011001010001000;
assign LUT_3[9539] = 32'b00000000000000010001110101100101;
assign LUT_3[9540] = 32'b00000000000000000110010000011010;
assign LUT_3[9541] = 32'b00000000000000001100111011110111;
assign LUT_3[9542] = 32'b00000000000000001000010111111110;
assign LUT_3[9543] = 32'b00000000000000001111000011011011;
assign LUT_3[9544] = 32'b00000000000000001110011011101010;
assign LUT_3[9545] = 32'b00000000000000010101000111000111;
assign LUT_3[9546] = 32'b00000000000000010000100011001110;
assign LUT_3[9547] = 32'b00000000000000010111001110101011;
assign LUT_3[9548] = 32'b00000000000000001011101001100000;
assign LUT_3[9549] = 32'b00000000000000010010010100111101;
assign LUT_3[9550] = 32'b00000000000000001101110001000100;
assign LUT_3[9551] = 32'b00000000000000010100011100100001;
assign LUT_3[9552] = 32'b00000000000000001100010101100111;
assign LUT_3[9553] = 32'b00000000000000010011000001000100;
assign LUT_3[9554] = 32'b00000000000000001110011101001011;
assign LUT_3[9555] = 32'b00000000000000010101001000101000;
assign LUT_3[9556] = 32'b00000000000000001001100011011101;
assign LUT_3[9557] = 32'b00000000000000010000001110111010;
assign LUT_3[9558] = 32'b00000000000000001011101011000001;
assign LUT_3[9559] = 32'b00000000000000010010010110011110;
assign LUT_3[9560] = 32'b00000000000000010001101110101101;
assign LUT_3[9561] = 32'b00000000000000011000011010001010;
assign LUT_3[9562] = 32'b00000000000000010011110110010001;
assign LUT_3[9563] = 32'b00000000000000011010100001101110;
assign LUT_3[9564] = 32'b00000000000000001110111100100011;
assign LUT_3[9565] = 32'b00000000000000010101101000000000;
assign LUT_3[9566] = 32'b00000000000000010001000100000111;
assign LUT_3[9567] = 32'b00000000000000010111101111100100;
assign LUT_3[9568] = 32'b00000000000000001010010001000100;
assign LUT_3[9569] = 32'b00000000000000010000111100100001;
assign LUT_3[9570] = 32'b00000000000000001100011000101000;
assign LUT_3[9571] = 32'b00000000000000010011000100000101;
assign LUT_3[9572] = 32'b00000000000000000111011110111010;
assign LUT_3[9573] = 32'b00000000000000001110001010010111;
assign LUT_3[9574] = 32'b00000000000000001001100110011110;
assign LUT_3[9575] = 32'b00000000000000010000010001111011;
assign LUT_3[9576] = 32'b00000000000000001111101010001010;
assign LUT_3[9577] = 32'b00000000000000010110010101100111;
assign LUT_3[9578] = 32'b00000000000000010001110001101110;
assign LUT_3[9579] = 32'b00000000000000011000011101001011;
assign LUT_3[9580] = 32'b00000000000000001100111000000000;
assign LUT_3[9581] = 32'b00000000000000010011100011011101;
assign LUT_3[9582] = 32'b00000000000000001110111111100100;
assign LUT_3[9583] = 32'b00000000000000010101101011000001;
assign LUT_3[9584] = 32'b00000000000000001101100100000111;
assign LUT_3[9585] = 32'b00000000000000010100001111100100;
assign LUT_3[9586] = 32'b00000000000000001111101011101011;
assign LUT_3[9587] = 32'b00000000000000010110010111001000;
assign LUT_3[9588] = 32'b00000000000000001010110001111101;
assign LUT_3[9589] = 32'b00000000000000010001011101011010;
assign LUT_3[9590] = 32'b00000000000000001100111001100001;
assign LUT_3[9591] = 32'b00000000000000010011100100111110;
assign LUT_3[9592] = 32'b00000000000000010010111101001101;
assign LUT_3[9593] = 32'b00000000000000011001101000101010;
assign LUT_3[9594] = 32'b00000000000000010101000100110001;
assign LUT_3[9595] = 32'b00000000000000011011110000001110;
assign LUT_3[9596] = 32'b00000000000000010000001011000011;
assign LUT_3[9597] = 32'b00000000000000010110110110100000;
assign LUT_3[9598] = 32'b00000000000000010010010010100111;
assign LUT_3[9599] = 32'b00000000000000011000111110000100;
assign LUT_3[9600] = 32'b00000000000000001011010100110111;
assign LUT_3[9601] = 32'b00000000000000010010000000010100;
assign LUT_3[9602] = 32'b00000000000000001101011100011011;
assign LUT_3[9603] = 32'b00000000000000010100000111111000;
assign LUT_3[9604] = 32'b00000000000000001000100010101101;
assign LUT_3[9605] = 32'b00000000000000001111001110001010;
assign LUT_3[9606] = 32'b00000000000000001010101010010001;
assign LUT_3[9607] = 32'b00000000000000010001010101101110;
assign LUT_3[9608] = 32'b00000000000000010000101101111101;
assign LUT_3[9609] = 32'b00000000000000010111011001011010;
assign LUT_3[9610] = 32'b00000000000000010010110101100001;
assign LUT_3[9611] = 32'b00000000000000011001100000111110;
assign LUT_3[9612] = 32'b00000000000000001101111011110011;
assign LUT_3[9613] = 32'b00000000000000010100100111010000;
assign LUT_3[9614] = 32'b00000000000000010000000011010111;
assign LUT_3[9615] = 32'b00000000000000010110101110110100;
assign LUT_3[9616] = 32'b00000000000000001110100111111010;
assign LUT_3[9617] = 32'b00000000000000010101010011010111;
assign LUT_3[9618] = 32'b00000000000000010000101111011110;
assign LUT_3[9619] = 32'b00000000000000010111011010111011;
assign LUT_3[9620] = 32'b00000000000000001011110101110000;
assign LUT_3[9621] = 32'b00000000000000010010100001001101;
assign LUT_3[9622] = 32'b00000000000000001101111101010100;
assign LUT_3[9623] = 32'b00000000000000010100101000110001;
assign LUT_3[9624] = 32'b00000000000000010100000001000000;
assign LUT_3[9625] = 32'b00000000000000011010101100011101;
assign LUT_3[9626] = 32'b00000000000000010110001000100100;
assign LUT_3[9627] = 32'b00000000000000011100110100000001;
assign LUT_3[9628] = 32'b00000000000000010001001110110110;
assign LUT_3[9629] = 32'b00000000000000010111111010010011;
assign LUT_3[9630] = 32'b00000000000000010011010110011010;
assign LUT_3[9631] = 32'b00000000000000011010000001110111;
assign LUT_3[9632] = 32'b00000000000000001100100011010111;
assign LUT_3[9633] = 32'b00000000000000010011001110110100;
assign LUT_3[9634] = 32'b00000000000000001110101010111011;
assign LUT_3[9635] = 32'b00000000000000010101010110011000;
assign LUT_3[9636] = 32'b00000000000000001001110001001101;
assign LUT_3[9637] = 32'b00000000000000010000011100101010;
assign LUT_3[9638] = 32'b00000000000000001011111000110001;
assign LUT_3[9639] = 32'b00000000000000010010100100001110;
assign LUT_3[9640] = 32'b00000000000000010001111100011101;
assign LUT_3[9641] = 32'b00000000000000011000100111111010;
assign LUT_3[9642] = 32'b00000000000000010100000100000001;
assign LUT_3[9643] = 32'b00000000000000011010101111011110;
assign LUT_3[9644] = 32'b00000000000000001111001010010011;
assign LUT_3[9645] = 32'b00000000000000010101110101110000;
assign LUT_3[9646] = 32'b00000000000000010001010001110111;
assign LUT_3[9647] = 32'b00000000000000010111111101010100;
assign LUT_3[9648] = 32'b00000000000000001111110110011010;
assign LUT_3[9649] = 32'b00000000000000010110100001110111;
assign LUT_3[9650] = 32'b00000000000000010001111101111110;
assign LUT_3[9651] = 32'b00000000000000011000101001011011;
assign LUT_3[9652] = 32'b00000000000000001101000100010000;
assign LUT_3[9653] = 32'b00000000000000010011101111101101;
assign LUT_3[9654] = 32'b00000000000000001111001011110100;
assign LUT_3[9655] = 32'b00000000000000010101110111010001;
assign LUT_3[9656] = 32'b00000000000000010101001111100000;
assign LUT_3[9657] = 32'b00000000000000011011111010111101;
assign LUT_3[9658] = 32'b00000000000000010111010111000100;
assign LUT_3[9659] = 32'b00000000000000011110000010100001;
assign LUT_3[9660] = 32'b00000000000000010010011101010110;
assign LUT_3[9661] = 32'b00000000000000011001001000110011;
assign LUT_3[9662] = 32'b00000000000000010100100100111010;
assign LUT_3[9663] = 32'b00000000000000011011010000010111;
assign LUT_3[9664] = 32'b00000000000000001011001101100010;
assign LUT_3[9665] = 32'b00000000000000010001111000111111;
assign LUT_3[9666] = 32'b00000000000000001101010101000110;
assign LUT_3[9667] = 32'b00000000000000010100000000100011;
assign LUT_3[9668] = 32'b00000000000000001000011011011000;
assign LUT_3[9669] = 32'b00000000000000001111000110110101;
assign LUT_3[9670] = 32'b00000000000000001010100010111100;
assign LUT_3[9671] = 32'b00000000000000010001001110011001;
assign LUT_3[9672] = 32'b00000000000000010000100110101000;
assign LUT_3[9673] = 32'b00000000000000010111010010000101;
assign LUT_3[9674] = 32'b00000000000000010010101110001100;
assign LUT_3[9675] = 32'b00000000000000011001011001101001;
assign LUT_3[9676] = 32'b00000000000000001101110100011110;
assign LUT_3[9677] = 32'b00000000000000010100011111111011;
assign LUT_3[9678] = 32'b00000000000000001111111100000010;
assign LUT_3[9679] = 32'b00000000000000010110100111011111;
assign LUT_3[9680] = 32'b00000000000000001110100000100101;
assign LUT_3[9681] = 32'b00000000000000010101001100000010;
assign LUT_3[9682] = 32'b00000000000000010000101000001001;
assign LUT_3[9683] = 32'b00000000000000010111010011100110;
assign LUT_3[9684] = 32'b00000000000000001011101110011011;
assign LUT_3[9685] = 32'b00000000000000010010011001111000;
assign LUT_3[9686] = 32'b00000000000000001101110101111111;
assign LUT_3[9687] = 32'b00000000000000010100100001011100;
assign LUT_3[9688] = 32'b00000000000000010011111001101011;
assign LUT_3[9689] = 32'b00000000000000011010100101001000;
assign LUT_3[9690] = 32'b00000000000000010110000001001111;
assign LUT_3[9691] = 32'b00000000000000011100101100101100;
assign LUT_3[9692] = 32'b00000000000000010001000111100001;
assign LUT_3[9693] = 32'b00000000000000010111110010111110;
assign LUT_3[9694] = 32'b00000000000000010011001111000101;
assign LUT_3[9695] = 32'b00000000000000011001111010100010;
assign LUT_3[9696] = 32'b00000000000000001100011100000010;
assign LUT_3[9697] = 32'b00000000000000010011000111011111;
assign LUT_3[9698] = 32'b00000000000000001110100011100110;
assign LUT_3[9699] = 32'b00000000000000010101001111000011;
assign LUT_3[9700] = 32'b00000000000000001001101001111000;
assign LUT_3[9701] = 32'b00000000000000010000010101010101;
assign LUT_3[9702] = 32'b00000000000000001011110001011100;
assign LUT_3[9703] = 32'b00000000000000010010011100111001;
assign LUT_3[9704] = 32'b00000000000000010001110101001000;
assign LUT_3[9705] = 32'b00000000000000011000100000100101;
assign LUT_3[9706] = 32'b00000000000000010011111100101100;
assign LUT_3[9707] = 32'b00000000000000011010101000001001;
assign LUT_3[9708] = 32'b00000000000000001111000010111110;
assign LUT_3[9709] = 32'b00000000000000010101101110011011;
assign LUT_3[9710] = 32'b00000000000000010001001010100010;
assign LUT_3[9711] = 32'b00000000000000010111110101111111;
assign LUT_3[9712] = 32'b00000000000000001111101111000101;
assign LUT_3[9713] = 32'b00000000000000010110011010100010;
assign LUT_3[9714] = 32'b00000000000000010001110110101001;
assign LUT_3[9715] = 32'b00000000000000011000100010000110;
assign LUT_3[9716] = 32'b00000000000000001100111100111011;
assign LUT_3[9717] = 32'b00000000000000010011101000011000;
assign LUT_3[9718] = 32'b00000000000000001111000100011111;
assign LUT_3[9719] = 32'b00000000000000010101101111111100;
assign LUT_3[9720] = 32'b00000000000000010101001000001011;
assign LUT_3[9721] = 32'b00000000000000011011110011101000;
assign LUT_3[9722] = 32'b00000000000000010111001111101111;
assign LUT_3[9723] = 32'b00000000000000011101111011001100;
assign LUT_3[9724] = 32'b00000000000000010010010110000001;
assign LUT_3[9725] = 32'b00000000000000011001000001011110;
assign LUT_3[9726] = 32'b00000000000000010100011101100101;
assign LUT_3[9727] = 32'b00000000000000011011001001000010;
assign LUT_3[9728] = 32'b00000000000000010000001111100100;
assign LUT_3[9729] = 32'b00000000000000010110111011000001;
assign LUT_3[9730] = 32'b00000000000000010010010111001000;
assign LUT_3[9731] = 32'b00000000000000011001000010100101;
assign LUT_3[9732] = 32'b00000000000000001101011101011010;
assign LUT_3[9733] = 32'b00000000000000010100001000110111;
assign LUT_3[9734] = 32'b00000000000000001111100100111110;
assign LUT_3[9735] = 32'b00000000000000010110010000011011;
assign LUT_3[9736] = 32'b00000000000000010101101000101010;
assign LUT_3[9737] = 32'b00000000000000011100010100000111;
assign LUT_3[9738] = 32'b00000000000000010111110000001110;
assign LUT_3[9739] = 32'b00000000000000011110011011101011;
assign LUT_3[9740] = 32'b00000000000000010010110110100000;
assign LUT_3[9741] = 32'b00000000000000011001100001111101;
assign LUT_3[9742] = 32'b00000000000000010100111110000100;
assign LUT_3[9743] = 32'b00000000000000011011101001100001;
assign LUT_3[9744] = 32'b00000000000000010011100010100111;
assign LUT_3[9745] = 32'b00000000000000011010001110000100;
assign LUT_3[9746] = 32'b00000000000000010101101010001011;
assign LUT_3[9747] = 32'b00000000000000011100010101101000;
assign LUT_3[9748] = 32'b00000000000000010000110000011101;
assign LUT_3[9749] = 32'b00000000000000010111011011111010;
assign LUT_3[9750] = 32'b00000000000000010010111000000001;
assign LUT_3[9751] = 32'b00000000000000011001100011011110;
assign LUT_3[9752] = 32'b00000000000000011000111011101101;
assign LUT_3[9753] = 32'b00000000000000011111100111001010;
assign LUT_3[9754] = 32'b00000000000000011011000011010001;
assign LUT_3[9755] = 32'b00000000000000100001101110101110;
assign LUT_3[9756] = 32'b00000000000000010110001001100011;
assign LUT_3[9757] = 32'b00000000000000011100110101000000;
assign LUT_3[9758] = 32'b00000000000000011000010001000111;
assign LUT_3[9759] = 32'b00000000000000011110111100100100;
assign LUT_3[9760] = 32'b00000000000000010001011110000100;
assign LUT_3[9761] = 32'b00000000000000011000001001100001;
assign LUT_3[9762] = 32'b00000000000000010011100101101000;
assign LUT_3[9763] = 32'b00000000000000011010010001000101;
assign LUT_3[9764] = 32'b00000000000000001110101011111010;
assign LUT_3[9765] = 32'b00000000000000010101010111010111;
assign LUT_3[9766] = 32'b00000000000000010000110011011110;
assign LUT_3[9767] = 32'b00000000000000010111011110111011;
assign LUT_3[9768] = 32'b00000000000000010110110111001010;
assign LUT_3[9769] = 32'b00000000000000011101100010100111;
assign LUT_3[9770] = 32'b00000000000000011000111110101110;
assign LUT_3[9771] = 32'b00000000000000011111101010001011;
assign LUT_3[9772] = 32'b00000000000000010100000101000000;
assign LUT_3[9773] = 32'b00000000000000011010110000011101;
assign LUT_3[9774] = 32'b00000000000000010110001100100100;
assign LUT_3[9775] = 32'b00000000000000011100111000000001;
assign LUT_3[9776] = 32'b00000000000000010100110001000111;
assign LUT_3[9777] = 32'b00000000000000011011011100100100;
assign LUT_3[9778] = 32'b00000000000000010110111000101011;
assign LUT_3[9779] = 32'b00000000000000011101100100001000;
assign LUT_3[9780] = 32'b00000000000000010001111110111101;
assign LUT_3[9781] = 32'b00000000000000011000101010011010;
assign LUT_3[9782] = 32'b00000000000000010100000110100001;
assign LUT_3[9783] = 32'b00000000000000011010110001111110;
assign LUT_3[9784] = 32'b00000000000000011010001010001101;
assign LUT_3[9785] = 32'b00000000000000100000110101101010;
assign LUT_3[9786] = 32'b00000000000000011100010001110001;
assign LUT_3[9787] = 32'b00000000000000100010111101001110;
assign LUT_3[9788] = 32'b00000000000000010111011000000011;
assign LUT_3[9789] = 32'b00000000000000011110000011100000;
assign LUT_3[9790] = 32'b00000000000000011001011111100111;
assign LUT_3[9791] = 32'b00000000000000100000001011000100;
assign LUT_3[9792] = 32'b00000000000000010000001000001111;
assign LUT_3[9793] = 32'b00000000000000010110110011101100;
assign LUT_3[9794] = 32'b00000000000000010010001111110011;
assign LUT_3[9795] = 32'b00000000000000011000111011010000;
assign LUT_3[9796] = 32'b00000000000000001101010110000101;
assign LUT_3[9797] = 32'b00000000000000010100000001100010;
assign LUT_3[9798] = 32'b00000000000000001111011101101001;
assign LUT_3[9799] = 32'b00000000000000010110001001000110;
assign LUT_3[9800] = 32'b00000000000000010101100001010101;
assign LUT_3[9801] = 32'b00000000000000011100001100110010;
assign LUT_3[9802] = 32'b00000000000000010111101000111001;
assign LUT_3[9803] = 32'b00000000000000011110010100010110;
assign LUT_3[9804] = 32'b00000000000000010010101111001011;
assign LUT_3[9805] = 32'b00000000000000011001011010101000;
assign LUT_3[9806] = 32'b00000000000000010100110110101111;
assign LUT_3[9807] = 32'b00000000000000011011100010001100;
assign LUT_3[9808] = 32'b00000000000000010011011011010010;
assign LUT_3[9809] = 32'b00000000000000011010000110101111;
assign LUT_3[9810] = 32'b00000000000000010101100010110110;
assign LUT_3[9811] = 32'b00000000000000011100001110010011;
assign LUT_3[9812] = 32'b00000000000000010000101001001000;
assign LUT_3[9813] = 32'b00000000000000010111010100100101;
assign LUT_3[9814] = 32'b00000000000000010010110000101100;
assign LUT_3[9815] = 32'b00000000000000011001011100001001;
assign LUT_3[9816] = 32'b00000000000000011000110100011000;
assign LUT_3[9817] = 32'b00000000000000011111011111110101;
assign LUT_3[9818] = 32'b00000000000000011010111011111100;
assign LUT_3[9819] = 32'b00000000000000100001100111011001;
assign LUT_3[9820] = 32'b00000000000000010110000010001110;
assign LUT_3[9821] = 32'b00000000000000011100101101101011;
assign LUT_3[9822] = 32'b00000000000000011000001001110010;
assign LUT_3[9823] = 32'b00000000000000011110110101001111;
assign LUT_3[9824] = 32'b00000000000000010001010110101111;
assign LUT_3[9825] = 32'b00000000000000011000000010001100;
assign LUT_3[9826] = 32'b00000000000000010011011110010011;
assign LUT_3[9827] = 32'b00000000000000011010001001110000;
assign LUT_3[9828] = 32'b00000000000000001110100100100101;
assign LUT_3[9829] = 32'b00000000000000010101010000000010;
assign LUT_3[9830] = 32'b00000000000000010000101100001001;
assign LUT_3[9831] = 32'b00000000000000010111010111100110;
assign LUT_3[9832] = 32'b00000000000000010110101111110101;
assign LUT_3[9833] = 32'b00000000000000011101011011010010;
assign LUT_3[9834] = 32'b00000000000000011000110111011001;
assign LUT_3[9835] = 32'b00000000000000011111100010110110;
assign LUT_3[9836] = 32'b00000000000000010011111101101011;
assign LUT_3[9837] = 32'b00000000000000011010101001001000;
assign LUT_3[9838] = 32'b00000000000000010110000101001111;
assign LUT_3[9839] = 32'b00000000000000011100110000101100;
assign LUT_3[9840] = 32'b00000000000000010100101001110010;
assign LUT_3[9841] = 32'b00000000000000011011010101001111;
assign LUT_3[9842] = 32'b00000000000000010110110001010110;
assign LUT_3[9843] = 32'b00000000000000011101011100110011;
assign LUT_3[9844] = 32'b00000000000000010001110111101000;
assign LUT_3[9845] = 32'b00000000000000011000100011000101;
assign LUT_3[9846] = 32'b00000000000000010011111111001100;
assign LUT_3[9847] = 32'b00000000000000011010101010101001;
assign LUT_3[9848] = 32'b00000000000000011010000010111000;
assign LUT_3[9849] = 32'b00000000000000100000101110010101;
assign LUT_3[9850] = 32'b00000000000000011100001010011100;
assign LUT_3[9851] = 32'b00000000000000100010110101111001;
assign LUT_3[9852] = 32'b00000000000000010111010000101110;
assign LUT_3[9853] = 32'b00000000000000011101111100001011;
assign LUT_3[9854] = 32'b00000000000000011001011000010010;
assign LUT_3[9855] = 32'b00000000000000100000000011101111;
assign LUT_3[9856] = 32'b00000000000000010010011010100010;
assign LUT_3[9857] = 32'b00000000000000011001000101111111;
assign LUT_3[9858] = 32'b00000000000000010100100010000110;
assign LUT_3[9859] = 32'b00000000000000011011001101100011;
assign LUT_3[9860] = 32'b00000000000000001111101000011000;
assign LUT_3[9861] = 32'b00000000000000010110010011110101;
assign LUT_3[9862] = 32'b00000000000000010001101111111100;
assign LUT_3[9863] = 32'b00000000000000011000011011011001;
assign LUT_3[9864] = 32'b00000000000000010111110011101000;
assign LUT_3[9865] = 32'b00000000000000011110011111000101;
assign LUT_3[9866] = 32'b00000000000000011001111011001100;
assign LUT_3[9867] = 32'b00000000000000100000100110101001;
assign LUT_3[9868] = 32'b00000000000000010101000001011110;
assign LUT_3[9869] = 32'b00000000000000011011101100111011;
assign LUT_3[9870] = 32'b00000000000000010111001001000010;
assign LUT_3[9871] = 32'b00000000000000011101110100011111;
assign LUT_3[9872] = 32'b00000000000000010101101101100101;
assign LUT_3[9873] = 32'b00000000000000011100011001000010;
assign LUT_3[9874] = 32'b00000000000000010111110101001001;
assign LUT_3[9875] = 32'b00000000000000011110100000100110;
assign LUT_3[9876] = 32'b00000000000000010010111011011011;
assign LUT_3[9877] = 32'b00000000000000011001100110111000;
assign LUT_3[9878] = 32'b00000000000000010101000010111111;
assign LUT_3[9879] = 32'b00000000000000011011101110011100;
assign LUT_3[9880] = 32'b00000000000000011011000110101011;
assign LUT_3[9881] = 32'b00000000000000100001110010001000;
assign LUT_3[9882] = 32'b00000000000000011101001110001111;
assign LUT_3[9883] = 32'b00000000000000100011111001101100;
assign LUT_3[9884] = 32'b00000000000000011000010100100001;
assign LUT_3[9885] = 32'b00000000000000011110111111111110;
assign LUT_3[9886] = 32'b00000000000000011010011100000101;
assign LUT_3[9887] = 32'b00000000000000100001000111100010;
assign LUT_3[9888] = 32'b00000000000000010011101001000010;
assign LUT_3[9889] = 32'b00000000000000011010010100011111;
assign LUT_3[9890] = 32'b00000000000000010101110000100110;
assign LUT_3[9891] = 32'b00000000000000011100011100000011;
assign LUT_3[9892] = 32'b00000000000000010000110110111000;
assign LUT_3[9893] = 32'b00000000000000010111100010010101;
assign LUT_3[9894] = 32'b00000000000000010010111110011100;
assign LUT_3[9895] = 32'b00000000000000011001101001111001;
assign LUT_3[9896] = 32'b00000000000000011001000010001000;
assign LUT_3[9897] = 32'b00000000000000011111101101100101;
assign LUT_3[9898] = 32'b00000000000000011011001001101100;
assign LUT_3[9899] = 32'b00000000000000100001110101001001;
assign LUT_3[9900] = 32'b00000000000000010110001111111110;
assign LUT_3[9901] = 32'b00000000000000011100111011011011;
assign LUT_3[9902] = 32'b00000000000000011000010111100010;
assign LUT_3[9903] = 32'b00000000000000011111000010111111;
assign LUT_3[9904] = 32'b00000000000000010110111100000101;
assign LUT_3[9905] = 32'b00000000000000011101100111100010;
assign LUT_3[9906] = 32'b00000000000000011001000011101001;
assign LUT_3[9907] = 32'b00000000000000011111101111000110;
assign LUT_3[9908] = 32'b00000000000000010100001001111011;
assign LUT_3[9909] = 32'b00000000000000011010110101011000;
assign LUT_3[9910] = 32'b00000000000000010110010001011111;
assign LUT_3[9911] = 32'b00000000000000011100111100111100;
assign LUT_3[9912] = 32'b00000000000000011100010101001011;
assign LUT_3[9913] = 32'b00000000000000100011000000101000;
assign LUT_3[9914] = 32'b00000000000000011110011100101111;
assign LUT_3[9915] = 32'b00000000000000100101001000001100;
assign LUT_3[9916] = 32'b00000000000000011001100011000001;
assign LUT_3[9917] = 32'b00000000000000100000001110011110;
assign LUT_3[9918] = 32'b00000000000000011011101010100101;
assign LUT_3[9919] = 32'b00000000000000100010010110000010;
assign LUT_3[9920] = 32'b00000000000000010010010011001101;
assign LUT_3[9921] = 32'b00000000000000011000111110101010;
assign LUT_3[9922] = 32'b00000000000000010100011010110001;
assign LUT_3[9923] = 32'b00000000000000011011000110001110;
assign LUT_3[9924] = 32'b00000000000000001111100001000011;
assign LUT_3[9925] = 32'b00000000000000010110001100100000;
assign LUT_3[9926] = 32'b00000000000000010001101000100111;
assign LUT_3[9927] = 32'b00000000000000011000010100000100;
assign LUT_3[9928] = 32'b00000000000000010111101100010011;
assign LUT_3[9929] = 32'b00000000000000011110010111110000;
assign LUT_3[9930] = 32'b00000000000000011001110011110111;
assign LUT_3[9931] = 32'b00000000000000100000011111010100;
assign LUT_3[9932] = 32'b00000000000000010100111010001001;
assign LUT_3[9933] = 32'b00000000000000011011100101100110;
assign LUT_3[9934] = 32'b00000000000000010111000001101101;
assign LUT_3[9935] = 32'b00000000000000011101101101001010;
assign LUT_3[9936] = 32'b00000000000000010101100110010000;
assign LUT_3[9937] = 32'b00000000000000011100010001101101;
assign LUT_3[9938] = 32'b00000000000000010111101101110100;
assign LUT_3[9939] = 32'b00000000000000011110011001010001;
assign LUT_3[9940] = 32'b00000000000000010010110100000110;
assign LUT_3[9941] = 32'b00000000000000011001011111100011;
assign LUT_3[9942] = 32'b00000000000000010100111011101010;
assign LUT_3[9943] = 32'b00000000000000011011100111000111;
assign LUT_3[9944] = 32'b00000000000000011010111111010110;
assign LUT_3[9945] = 32'b00000000000000100001101010110011;
assign LUT_3[9946] = 32'b00000000000000011101000110111010;
assign LUT_3[9947] = 32'b00000000000000100011110010010111;
assign LUT_3[9948] = 32'b00000000000000011000001101001100;
assign LUT_3[9949] = 32'b00000000000000011110111000101001;
assign LUT_3[9950] = 32'b00000000000000011010010100110000;
assign LUT_3[9951] = 32'b00000000000000100001000000001101;
assign LUT_3[9952] = 32'b00000000000000010011100001101101;
assign LUT_3[9953] = 32'b00000000000000011010001101001010;
assign LUT_3[9954] = 32'b00000000000000010101101001010001;
assign LUT_3[9955] = 32'b00000000000000011100010100101110;
assign LUT_3[9956] = 32'b00000000000000010000101111100011;
assign LUT_3[9957] = 32'b00000000000000010111011011000000;
assign LUT_3[9958] = 32'b00000000000000010010110111000111;
assign LUT_3[9959] = 32'b00000000000000011001100010100100;
assign LUT_3[9960] = 32'b00000000000000011000111010110011;
assign LUT_3[9961] = 32'b00000000000000011111100110010000;
assign LUT_3[9962] = 32'b00000000000000011011000010010111;
assign LUT_3[9963] = 32'b00000000000000100001101101110100;
assign LUT_3[9964] = 32'b00000000000000010110001000101001;
assign LUT_3[9965] = 32'b00000000000000011100110100000110;
assign LUT_3[9966] = 32'b00000000000000011000010000001101;
assign LUT_3[9967] = 32'b00000000000000011110111011101010;
assign LUT_3[9968] = 32'b00000000000000010110110100110000;
assign LUT_3[9969] = 32'b00000000000000011101100000001101;
assign LUT_3[9970] = 32'b00000000000000011000111100010100;
assign LUT_3[9971] = 32'b00000000000000011111100111110001;
assign LUT_3[9972] = 32'b00000000000000010100000010100110;
assign LUT_3[9973] = 32'b00000000000000011010101110000011;
assign LUT_3[9974] = 32'b00000000000000010110001010001010;
assign LUT_3[9975] = 32'b00000000000000011100110101100111;
assign LUT_3[9976] = 32'b00000000000000011100001101110110;
assign LUT_3[9977] = 32'b00000000000000100010111001010011;
assign LUT_3[9978] = 32'b00000000000000011110010101011010;
assign LUT_3[9979] = 32'b00000000000000100101000000110111;
assign LUT_3[9980] = 32'b00000000000000011001011011101100;
assign LUT_3[9981] = 32'b00000000000000100000000111001001;
assign LUT_3[9982] = 32'b00000000000000011011100011010000;
assign LUT_3[9983] = 32'b00000000000000100010001110101101;
assign LUT_3[9984] = 32'b00000000000000001100011111000101;
assign LUT_3[9985] = 32'b00000000000000010011001010100010;
assign LUT_3[9986] = 32'b00000000000000001110100110101001;
assign LUT_3[9987] = 32'b00000000000000010101010010000110;
assign LUT_3[9988] = 32'b00000000000000001001101100111011;
assign LUT_3[9989] = 32'b00000000000000010000011000011000;
assign LUT_3[9990] = 32'b00000000000000001011110100011111;
assign LUT_3[9991] = 32'b00000000000000010010011111111100;
assign LUT_3[9992] = 32'b00000000000000010001111000001011;
assign LUT_3[9993] = 32'b00000000000000011000100011101000;
assign LUT_3[9994] = 32'b00000000000000010011111111101111;
assign LUT_3[9995] = 32'b00000000000000011010101011001100;
assign LUT_3[9996] = 32'b00000000000000001111000110000001;
assign LUT_3[9997] = 32'b00000000000000010101110001011110;
assign LUT_3[9998] = 32'b00000000000000010001001101100101;
assign LUT_3[9999] = 32'b00000000000000010111111001000010;
assign LUT_3[10000] = 32'b00000000000000001111110010001000;
assign LUT_3[10001] = 32'b00000000000000010110011101100101;
assign LUT_3[10002] = 32'b00000000000000010001111001101100;
assign LUT_3[10003] = 32'b00000000000000011000100101001001;
assign LUT_3[10004] = 32'b00000000000000001100111111111110;
assign LUT_3[10005] = 32'b00000000000000010011101011011011;
assign LUT_3[10006] = 32'b00000000000000001111000111100010;
assign LUT_3[10007] = 32'b00000000000000010101110010111111;
assign LUT_3[10008] = 32'b00000000000000010101001011001110;
assign LUT_3[10009] = 32'b00000000000000011011110110101011;
assign LUT_3[10010] = 32'b00000000000000010111010010110010;
assign LUT_3[10011] = 32'b00000000000000011101111110001111;
assign LUT_3[10012] = 32'b00000000000000010010011001000100;
assign LUT_3[10013] = 32'b00000000000000011001000100100001;
assign LUT_3[10014] = 32'b00000000000000010100100000101000;
assign LUT_3[10015] = 32'b00000000000000011011001100000101;
assign LUT_3[10016] = 32'b00000000000000001101101101100101;
assign LUT_3[10017] = 32'b00000000000000010100011001000010;
assign LUT_3[10018] = 32'b00000000000000001111110101001001;
assign LUT_3[10019] = 32'b00000000000000010110100000100110;
assign LUT_3[10020] = 32'b00000000000000001010111011011011;
assign LUT_3[10021] = 32'b00000000000000010001100110111000;
assign LUT_3[10022] = 32'b00000000000000001101000010111111;
assign LUT_3[10023] = 32'b00000000000000010011101110011100;
assign LUT_3[10024] = 32'b00000000000000010011000110101011;
assign LUT_3[10025] = 32'b00000000000000011001110010001000;
assign LUT_3[10026] = 32'b00000000000000010101001110001111;
assign LUT_3[10027] = 32'b00000000000000011011111001101100;
assign LUT_3[10028] = 32'b00000000000000010000010100100001;
assign LUT_3[10029] = 32'b00000000000000010110111111111110;
assign LUT_3[10030] = 32'b00000000000000010010011100000101;
assign LUT_3[10031] = 32'b00000000000000011001000111100010;
assign LUT_3[10032] = 32'b00000000000000010001000000101000;
assign LUT_3[10033] = 32'b00000000000000010111101100000101;
assign LUT_3[10034] = 32'b00000000000000010011001000001100;
assign LUT_3[10035] = 32'b00000000000000011001110011101001;
assign LUT_3[10036] = 32'b00000000000000001110001110011110;
assign LUT_3[10037] = 32'b00000000000000010100111001111011;
assign LUT_3[10038] = 32'b00000000000000010000010110000010;
assign LUT_3[10039] = 32'b00000000000000010111000001011111;
assign LUT_3[10040] = 32'b00000000000000010110011001101110;
assign LUT_3[10041] = 32'b00000000000000011101000101001011;
assign LUT_3[10042] = 32'b00000000000000011000100001010010;
assign LUT_3[10043] = 32'b00000000000000011111001100101111;
assign LUT_3[10044] = 32'b00000000000000010011100111100100;
assign LUT_3[10045] = 32'b00000000000000011010010011000001;
assign LUT_3[10046] = 32'b00000000000000010101101111001000;
assign LUT_3[10047] = 32'b00000000000000011100011010100101;
assign LUT_3[10048] = 32'b00000000000000001100010111110000;
assign LUT_3[10049] = 32'b00000000000000010011000011001101;
assign LUT_3[10050] = 32'b00000000000000001110011111010100;
assign LUT_3[10051] = 32'b00000000000000010101001010110001;
assign LUT_3[10052] = 32'b00000000000000001001100101100110;
assign LUT_3[10053] = 32'b00000000000000010000010001000011;
assign LUT_3[10054] = 32'b00000000000000001011101101001010;
assign LUT_3[10055] = 32'b00000000000000010010011000100111;
assign LUT_3[10056] = 32'b00000000000000010001110000110110;
assign LUT_3[10057] = 32'b00000000000000011000011100010011;
assign LUT_3[10058] = 32'b00000000000000010011111000011010;
assign LUT_3[10059] = 32'b00000000000000011010100011110111;
assign LUT_3[10060] = 32'b00000000000000001110111110101100;
assign LUT_3[10061] = 32'b00000000000000010101101010001001;
assign LUT_3[10062] = 32'b00000000000000010001000110010000;
assign LUT_3[10063] = 32'b00000000000000010111110001101101;
assign LUT_3[10064] = 32'b00000000000000001111101010110011;
assign LUT_3[10065] = 32'b00000000000000010110010110010000;
assign LUT_3[10066] = 32'b00000000000000010001110010010111;
assign LUT_3[10067] = 32'b00000000000000011000011101110100;
assign LUT_3[10068] = 32'b00000000000000001100111000101001;
assign LUT_3[10069] = 32'b00000000000000010011100100000110;
assign LUT_3[10070] = 32'b00000000000000001111000000001101;
assign LUT_3[10071] = 32'b00000000000000010101101011101010;
assign LUT_3[10072] = 32'b00000000000000010101000011111001;
assign LUT_3[10073] = 32'b00000000000000011011101111010110;
assign LUT_3[10074] = 32'b00000000000000010111001011011101;
assign LUT_3[10075] = 32'b00000000000000011101110110111010;
assign LUT_3[10076] = 32'b00000000000000010010010001101111;
assign LUT_3[10077] = 32'b00000000000000011000111101001100;
assign LUT_3[10078] = 32'b00000000000000010100011001010011;
assign LUT_3[10079] = 32'b00000000000000011011000100110000;
assign LUT_3[10080] = 32'b00000000000000001101100110010000;
assign LUT_3[10081] = 32'b00000000000000010100010001101101;
assign LUT_3[10082] = 32'b00000000000000001111101101110100;
assign LUT_3[10083] = 32'b00000000000000010110011001010001;
assign LUT_3[10084] = 32'b00000000000000001010110100000110;
assign LUT_3[10085] = 32'b00000000000000010001011111100011;
assign LUT_3[10086] = 32'b00000000000000001100111011101010;
assign LUT_3[10087] = 32'b00000000000000010011100111000111;
assign LUT_3[10088] = 32'b00000000000000010010111111010110;
assign LUT_3[10089] = 32'b00000000000000011001101010110011;
assign LUT_3[10090] = 32'b00000000000000010101000110111010;
assign LUT_3[10091] = 32'b00000000000000011011110010010111;
assign LUT_3[10092] = 32'b00000000000000010000001101001100;
assign LUT_3[10093] = 32'b00000000000000010110111000101001;
assign LUT_3[10094] = 32'b00000000000000010010010100110000;
assign LUT_3[10095] = 32'b00000000000000011001000000001101;
assign LUT_3[10096] = 32'b00000000000000010000111001010011;
assign LUT_3[10097] = 32'b00000000000000010111100100110000;
assign LUT_3[10098] = 32'b00000000000000010011000000110111;
assign LUT_3[10099] = 32'b00000000000000011001101100010100;
assign LUT_3[10100] = 32'b00000000000000001110000111001001;
assign LUT_3[10101] = 32'b00000000000000010100110010100110;
assign LUT_3[10102] = 32'b00000000000000010000001110101101;
assign LUT_3[10103] = 32'b00000000000000010110111010001010;
assign LUT_3[10104] = 32'b00000000000000010110010010011001;
assign LUT_3[10105] = 32'b00000000000000011100111101110110;
assign LUT_3[10106] = 32'b00000000000000011000011001111101;
assign LUT_3[10107] = 32'b00000000000000011111000101011010;
assign LUT_3[10108] = 32'b00000000000000010011100000001111;
assign LUT_3[10109] = 32'b00000000000000011010001011101100;
assign LUT_3[10110] = 32'b00000000000000010101100111110011;
assign LUT_3[10111] = 32'b00000000000000011100010011010000;
assign LUT_3[10112] = 32'b00000000000000001110101010000011;
assign LUT_3[10113] = 32'b00000000000000010101010101100000;
assign LUT_3[10114] = 32'b00000000000000010000110001100111;
assign LUT_3[10115] = 32'b00000000000000010111011101000100;
assign LUT_3[10116] = 32'b00000000000000001011110111111001;
assign LUT_3[10117] = 32'b00000000000000010010100011010110;
assign LUT_3[10118] = 32'b00000000000000001101111111011101;
assign LUT_3[10119] = 32'b00000000000000010100101010111010;
assign LUT_3[10120] = 32'b00000000000000010100000011001001;
assign LUT_3[10121] = 32'b00000000000000011010101110100110;
assign LUT_3[10122] = 32'b00000000000000010110001010101101;
assign LUT_3[10123] = 32'b00000000000000011100110110001010;
assign LUT_3[10124] = 32'b00000000000000010001010000111111;
assign LUT_3[10125] = 32'b00000000000000010111111100011100;
assign LUT_3[10126] = 32'b00000000000000010011011000100011;
assign LUT_3[10127] = 32'b00000000000000011010000100000000;
assign LUT_3[10128] = 32'b00000000000000010001111101000110;
assign LUT_3[10129] = 32'b00000000000000011000101000100011;
assign LUT_3[10130] = 32'b00000000000000010100000100101010;
assign LUT_3[10131] = 32'b00000000000000011010110000000111;
assign LUT_3[10132] = 32'b00000000000000001111001010111100;
assign LUT_3[10133] = 32'b00000000000000010101110110011001;
assign LUT_3[10134] = 32'b00000000000000010001010010100000;
assign LUT_3[10135] = 32'b00000000000000010111111101111101;
assign LUT_3[10136] = 32'b00000000000000010111010110001100;
assign LUT_3[10137] = 32'b00000000000000011110000001101001;
assign LUT_3[10138] = 32'b00000000000000011001011101110000;
assign LUT_3[10139] = 32'b00000000000000100000001001001101;
assign LUT_3[10140] = 32'b00000000000000010100100100000010;
assign LUT_3[10141] = 32'b00000000000000011011001111011111;
assign LUT_3[10142] = 32'b00000000000000010110101011100110;
assign LUT_3[10143] = 32'b00000000000000011101010111000011;
assign LUT_3[10144] = 32'b00000000000000001111111000100011;
assign LUT_3[10145] = 32'b00000000000000010110100100000000;
assign LUT_3[10146] = 32'b00000000000000010010000000000111;
assign LUT_3[10147] = 32'b00000000000000011000101011100100;
assign LUT_3[10148] = 32'b00000000000000001101000110011001;
assign LUT_3[10149] = 32'b00000000000000010011110001110110;
assign LUT_3[10150] = 32'b00000000000000001111001101111101;
assign LUT_3[10151] = 32'b00000000000000010101111001011010;
assign LUT_3[10152] = 32'b00000000000000010101010001101001;
assign LUT_3[10153] = 32'b00000000000000011011111101000110;
assign LUT_3[10154] = 32'b00000000000000010111011001001101;
assign LUT_3[10155] = 32'b00000000000000011110000100101010;
assign LUT_3[10156] = 32'b00000000000000010010011111011111;
assign LUT_3[10157] = 32'b00000000000000011001001010111100;
assign LUT_3[10158] = 32'b00000000000000010100100111000011;
assign LUT_3[10159] = 32'b00000000000000011011010010100000;
assign LUT_3[10160] = 32'b00000000000000010011001011100110;
assign LUT_3[10161] = 32'b00000000000000011001110111000011;
assign LUT_3[10162] = 32'b00000000000000010101010011001010;
assign LUT_3[10163] = 32'b00000000000000011011111110100111;
assign LUT_3[10164] = 32'b00000000000000010000011001011100;
assign LUT_3[10165] = 32'b00000000000000010111000100111001;
assign LUT_3[10166] = 32'b00000000000000010010100001000000;
assign LUT_3[10167] = 32'b00000000000000011001001100011101;
assign LUT_3[10168] = 32'b00000000000000011000100100101100;
assign LUT_3[10169] = 32'b00000000000000011111010000001001;
assign LUT_3[10170] = 32'b00000000000000011010101100010000;
assign LUT_3[10171] = 32'b00000000000000100001010111101101;
assign LUT_3[10172] = 32'b00000000000000010101110010100010;
assign LUT_3[10173] = 32'b00000000000000011100011101111111;
assign LUT_3[10174] = 32'b00000000000000010111111010000110;
assign LUT_3[10175] = 32'b00000000000000011110100101100011;
assign LUT_3[10176] = 32'b00000000000000001110100010101110;
assign LUT_3[10177] = 32'b00000000000000010101001110001011;
assign LUT_3[10178] = 32'b00000000000000010000101010010010;
assign LUT_3[10179] = 32'b00000000000000010111010101101111;
assign LUT_3[10180] = 32'b00000000000000001011110000100100;
assign LUT_3[10181] = 32'b00000000000000010010011100000001;
assign LUT_3[10182] = 32'b00000000000000001101111000001000;
assign LUT_3[10183] = 32'b00000000000000010100100011100101;
assign LUT_3[10184] = 32'b00000000000000010011111011110100;
assign LUT_3[10185] = 32'b00000000000000011010100111010001;
assign LUT_3[10186] = 32'b00000000000000010110000011011000;
assign LUT_3[10187] = 32'b00000000000000011100101110110101;
assign LUT_3[10188] = 32'b00000000000000010001001001101010;
assign LUT_3[10189] = 32'b00000000000000010111110101000111;
assign LUT_3[10190] = 32'b00000000000000010011010001001110;
assign LUT_3[10191] = 32'b00000000000000011001111100101011;
assign LUT_3[10192] = 32'b00000000000000010001110101110001;
assign LUT_3[10193] = 32'b00000000000000011000100001001110;
assign LUT_3[10194] = 32'b00000000000000010011111101010101;
assign LUT_3[10195] = 32'b00000000000000011010101000110010;
assign LUT_3[10196] = 32'b00000000000000001111000011100111;
assign LUT_3[10197] = 32'b00000000000000010101101111000100;
assign LUT_3[10198] = 32'b00000000000000010001001011001011;
assign LUT_3[10199] = 32'b00000000000000010111110110101000;
assign LUT_3[10200] = 32'b00000000000000010111001110110111;
assign LUT_3[10201] = 32'b00000000000000011101111010010100;
assign LUT_3[10202] = 32'b00000000000000011001010110011011;
assign LUT_3[10203] = 32'b00000000000000100000000001111000;
assign LUT_3[10204] = 32'b00000000000000010100011100101101;
assign LUT_3[10205] = 32'b00000000000000011011001000001010;
assign LUT_3[10206] = 32'b00000000000000010110100100010001;
assign LUT_3[10207] = 32'b00000000000000011101001111101110;
assign LUT_3[10208] = 32'b00000000000000001111110001001110;
assign LUT_3[10209] = 32'b00000000000000010110011100101011;
assign LUT_3[10210] = 32'b00000000000000010001111000110010;
assign LUT_3[10211] = 32'b00000000000000011000100100001111;
assign LUT_3[10212] = 32'b00000000000000001100111111000100;
assign LUT_3[10213] = 32'b00000000000000010011101010100001;
assign LUT_3[10214] = 32'b00000000000000001111000110101000;
assign LUT_3[10215] = 32'b00000000000000010101110010000101;
assign LUT_3[10216] = 32'b00000000000000010101001010010100;
assign LUT_3[10217] = 32'b00000000000000011011110101110001;
assign LUT_3[10218] = 32'b00000000000000010111010001111000;
assign LUT_3[10219] = 32'b00000000000000011101111101010101;
assign LUT_3[10220] = 32'b00000000000000010010011000001010;
assign LUT_3[10221] = 32'b00000000000000011001000011100111;
assign LUT_3[10222] = 32'b00000000000000010100011111101110;
assign LUT_3[10223] = 32'b00000000000000011011001011001011;
assign LUT_3[10224] = 32'b00000000000000010011000100010001;
assign LUT_3[10225] = 32'b00000000000000011001101111101110;
assign LUT_3[10226] = 32'b00000000000000010101001011110101;
assign LUT_3[10227] = 32'b00000000000000011011110111010010;
assign LUT_3[10228] = 32'b00000000000000010000010010000111;
assign LUT_3[10229] = 32'b00000000000000010110111101100100;
assign LUT_3[10230] = 32'b00000000000000010010011001101011;
assign LUT_3[10231] = 32'b00000000000000011001000101001000;
assign LUT_3[10232] = 32'b00000000000000011000011101010111;
assign LUT_3[10233] = 32'b00000000000000011111001000110100;
assign LUT_3[10234] = 32'b00000000000000011010100100111011;
assign LUT_3[10235] = 32'b00000000000000100001010000011000;
assign LUT_3[10236] = 32'b00000000000000010101101011001101;
assign LUT_3[10237] = 32'b00000000000000011100010110101010;
assign LUT_3[10238] = 32'b00000000000000010111110010110001;
assign LUT_3[10239] = 32'b00000000000000011110011110001110;
assign LUT_3[10240] = 32'b00000000000000001000001011101001;
assign LUT_3[10241] = 32'b00000000000000001110110111000110;
assign LUT_3[10242] = 32'b00000000000000001010010011001101;
assign LUT_3[10243] = 32'b00000000000000010000111110101010;
assign LUT_3[10244] = 32'b00000000000000000101011001011111;
assign LUT_3[10245] = 32'b00000000000000001100000100111100;
assign LUT_3[10246] = 32'b00000000000000000111100001000011;
assign LUT_3[10247] = 32'b00000000000000001110001100100000;
assign LUT_3[10248] = 32'b00000000000000001101100100101111;
assign LUT_3[10249] = 32'b00000000000000010100010000001100;
assign LUT_3[10250] = 32'b00000000000000001111101100010011;
assign LUT_3[10251] = 32'b00000000000000010110010111110000;
assign LUT_3[10252] = 32'b00000000000000001010110010100101;
assign LUT_3[10253] = 32'b00000000000000010001011110000010;
assign LUT_3[10254] = 32'b00000000000000001100111010001001;
assign LUT_3[10255] = 32'b00000000000000010011100101100110;
assign LUT_3[10256] = 32'b00000000000000001011011110101100;
assign LUT_3[10257] = 32'b00000000000000010010001010001001;
assign LUT_3[10258] = 32'b00000000000000001101100110010000;
assign LUT_3[10259] = 32'b00000000000000010100010001101101;
assign LUT_3[10260] = 32'b00000000000000001000101100100010;
assign LUT_3[10261] = 32'b00000000000000001111010111111111;
assign LUT_3[10262] = 32'b00000000000000001010110100000110;
assign LUT_3[10263] = 32'b00000000000000010001011111100011;
assign LUT_3[10264] = 32'b00000000000000010000110111110010;
assign LUT_3[10265] = 32'b00000000000000010111100011001111;
assign LUT_3[10266] = 32'b00000000000000010010111111010110;
assign LUT_3[10267] = 32'b00000000000000011001101010110011;
assign LUT_3[10268] = 32'b00000000000000001110000101101000;
assign LUT_3[10269] = 32'b00000000000000010100110001000101;
assign LUT_3[10270] = 32'b00000000000000010000001101001100;
assign LUT_3[10271] = 32'b00000000000000010110111000101001;
assign LUT_3[10272] = 32'b00000000000000001001011010001001;
assign LUT_3[10273] = 32'b00000000000000010000000101100110;
assign LUT_3[10274] = 32'b00000000000000001011100001101101;
assign LUT_3[10275] = 32'b00000000000000010010001101001010;
assign LUT_3[10276] = 32'b00000000000000000110100111111111;
assign LUT_3[10277] = 32'b00000000000000001101010011011100;
assign LUT_3[10278] = 32'b00000000000000001000101111100011;
assign LUT_3[10279] = 32'b00000000000000001111011011000000;
assign LUT_3[10280] = 32'b00000000000000001110110011001111;
assign LUT_3[10281] = 32'b00000000000000010101011110101100;
assign LUT_3[10282] = 32'b00000000000000010000111010110011;
assign LUT_3[10283] = 32'b00000000000000010111100110010000;
assign LUT_3[10284] = 32'b00000000000000001100000001000101;
assign LUT_3[10285] = 32'b00000000000000010010101100100010;
assign LUT_3[10286] = 32'b00000000000000001110001000101001;
assign LUT_3[10287] = 32'b00000000000000010100110100000110;
assign LUT_3[10288] = 32'b00000000000000001100101101001100;
assign LUT_3[10289] = 32'b00000000000000010011011000101001;
assign LUT_3[10290] = 32'b00000000000000001110110100110000;
assign LUT_3[10291] = 32'b00000000000000010101100000001101;
assign LUT_3[10292] = 32'b00000000000000001001111011000010;
assign LUT_3[10293] = 32'b00000000000000010000100110011111;
assign LUT_3[10294] = 32'b00000000000000001100000010100110;
assign LUT_3[10295] = 32'b00000000000000010010101110000011;
assign LUT_3[10296] = 32'b00000000000000010010000110010010;
assign LUT_3[10297] = 32'b00000000000000011000110001101111;
assign LUT_3[10298] = 32'b00000000000000010100001101110110;
assign LUT_3[10299] = 32'b00000000000000011010111001010011;
assign LUT_3[10300] = 32'b00000000000000001111010100001000;
assign LUT_3[10301] = 32'b00000000000000010101111111100101;
assign LUT_3[10302] = 32'b00000000000000010001011011101100;
assign LUT_3[10303] = 32'b00000000000000011000000111001001;
assign LUT_3[10304] = 32'b00000000000000001000000100010100;
assign LUT_3[10305] = 32'b00000000000000001110101111110001;
assign LUT_3[10306] = 32'b00000000000000001010001011111000;
assign LUT_3[10307] = 32'b00000000000000010000110111010101;
assign LUT_3[10308] = 32'b00000000000000000101010010001010;
assign LUT_3[10309] = 32'b00000000000000001011111101100111;
assign LUT_3[10310] = 32'b00000000000000000111011001101110;
assign LUT_3[10311] = 32'b00000000000000001110000101001011;
assign LUT_3[10312] = 32'b00000000000000001101011101011010;
assign LUT_3[10313] = 32'b00000000000000010100001000110111;
assign LUT_3[10314] = 32'b00000000000000001111100100111110;
assign LUT_3[10315] = 32'b00000000000000010110010000011011;
assign LUT_3[10316] = 32'b00000000000000001010101011010000;
assign LUT_3[10317] = 32'b00000000000000010001010110101101;
assign LUT_3[10318] = 32'b00000000000000001100110010110100;
assign LUT_3[10319] = 32'b00000000000000010011011110010001;
assign LUT_3[10320] = 32'b00000000000000001011010111010111;
assign LUT_3[10321] = 32'b00000000000000010010000010110100;
assign LUT_3[10322] = 32'b00000000000000001101011110111011;
assign LUT_3[10323] = 32'b00000000000000010100001010011000;
assign LUT_3[10324] = 32'b00000000000000001000100101001101;
assign LUT_3[10325] = 32'b00000000000000001111010000101010;
assign LUT_3[10326] = 32'b00000000000000001010101100110001;
assign LUT_3[10327] = 32'b00000000000000010001011000001110;
assign LUT_3[10328] = 32'b00000000000000010000110000011101;
assign LUT_3[10329] = 32'b00000000000000010111011011111010;
assign LUT_3[10330] = 32'b00000000000000010010111000000001;
assign LUT_3[10331] = 32'b00000000000000011001100011011110;
assign LUT_3[10332] = 32'b00000000000000001101111110010011;
assign LUT_3[10333] = 32'b00000000000000010100101001110000;
assign LUT_3[10334] = 32'b00000000000000010000000101110111;
assign LUT_3[10335] = 32'b00000000000000010110110001010100;
assign LUT_3[10336] = 32'b00000000000000001001010010110100;
assign LUT_3[10337] = 32'b00000000000000001111111110010001;
assign LUT_3[10338] = 32'b00000000000000001011011010011000;
assign LUT_3[10339] = 32'b00000000000000010010000101110101;
assign LUT_3[10340] = 32'b00000000000000000110100000101010;
assign LUT_3[10341] = 32'b00000000000000001101001100000111;
assign LUT_3[10342] = 32'b00000000000000001000101000001110;
assign LUT_3[10343] = 32'b00000000000000001111010011101011;
assign LUT_3[10344] = 32'b00000000000000001110101011111010;
assign LUT_3[10345] = 32'b00000000000000010101010111010111;
assign LUT_3[10346] = 32'b00000000000000010000110011011110;
assign LUT_3[10347] = 32'b00000000000000010111011110111011;
assign LUT_3[10348] = 32'b00000000000000001011111001110000;
assign LUT_3[10349] = 32'b00000000000000010010100101001101;
assign LUT_3[10350] = 32'b00000000000000001110000001010100;
assign LUT_3[10351] = 32'b00000000000000010100101100110001;
assign LUT_3[10352] = 32'b00000000000000001100100101110111;
assign LUT_3[10353] = 32'b00000000000000010011010001010100;
assign LUT_3[10354] = 32'b00000000000000001110101101011011;
assign LUT_3[10355] = 32'b00000000000000010101011000111000;
assign LUT_3[10356] = 32'b00000000000000001001110011101101;
assign LUT_3[10357] = 32'b00000000000000010000011111001010;
assign LUT_3[10358] = 32'b00000000000000001011111011010001;
assign LUT_3[10359] = 32'b00000000000000010010100110101110;
assign LUT_3[10360] = 32'b00000000000000010001111110111101;
assign LUT_3[10361] = 32'b00000000000000011000101010011010;
assign LUT_3[10362] = 32'b00000000000000010100000110100001;
assign LUT_3[10363] = 32'b00000000000000011010110001111110;
assign LUT_3[10364] = 32'b00000000000000001111001100110011;
assign LUT_3[10365] = 32'b00000000000000010101111000010000;
assign LUT_3[10366] = 32'b00000000000000010001010100010111;
assign LUT_3[10367] = 32'b00000000000000010111111111110100;
assign LUT_3[10368] = 32'b00000000000000001010010110100111;
assign LUT_3[10369] = 32'b00000000000000010001000010000100;
assign LUT_3[10370] = 32'b00000000000000001100011110001011;
assign LUT_3[10371] = 32'b00000000000000010011001001101000;
assign LUT_3[10372] = 32'b00000000000000000111100100011101;
assign LUT_3[10373] = 32'b00000000000000001110001111111010;
assign LUT_3[10374] = 32'b00000000000000001001101100000001;
assign LUT_3[10375] = 32'b00000000000000010000010111011110;
assign LUT_3[10376] = 32'b00000000000000001111101111101101;
assign LUT_3[10377] = 32'b00000000000000010110011011001010;
assign LUT_3[10378] = 32'b00000000000000010001110111010001;
assign LUT_3[10379] = 32'b00000000000000011000100010101110;
assign LUT_3[10380] = 32'b00000000000000001100111101100011;
assign LUT_3[10381] = 32'b00000000000000010011101001000000;
assign LUT_3[10382] = 32'b00000000000000001111000101000111;
assign LUT_3[10383] = 32'b00000000000000010101110000100100;
assign LUT_3[10384] = 32'b00000000000000001101101001101010;
assign LUT_3[10385] = 32'b00000000000000010100010101000111;
assign LUT_3[10386] = 32'b00000000000000001111110001001110;
assign LUT_3[10387] = 32'b00000000000000010110011100101011;
assign LUT_3[10388] = 32'b00000000000000001010110111100000;
assign LUT_3[10389] = 32'b00000000000000010001100010111101;
assign LUT_3[10390] = 32'b00000000000000001100111111000100;
assign LUT_3[10391] = 32'b00000000000000010011101010100001;
assign LUT_3[10392] = 32'b00000000000000010011000010110000;
assign LUT_3[10393] = 32'b00000000000000011001101110001101;
assign LUT_3[10394] = 32'b00000000000000010101001010010100;
assign LUT_3[10395] = 32'b00000000000000011011110101110001;
assign LUT_3[10396] = 32'b00000000000000010000010000100110;
assign LUT_3[10397] = 32'b00000000000000010110111100000011;
assign LUT_3[10398] = 32'b00000000000000010010011000001010;
assign LUT_3[10399] = 32'b00000000000000011001000011100111;
assign LUT_3[10400] = 32'b00000000000000001011100101000111;
assign LUT_3[10401] = 32'b00000000000000010010010000100100;
assign LUT_3[10402] = 32'b00000000000000001101101100101011;
assign LUT_3[10403] = 32'b00000000000000010100011000001000;
assign LUT_3[10404] = 32'b00000000000000001000110010111101;
assign LUT_3[10405] = 32'b00000000000000001111011110011010;
assign LUT_3[10406] = 32'b00000000000000001010111010100001;
assign LUT_3[10407] = 32'b00000000000000010001100101111110;
assign LUT_3[10408] = 32'b00000000000000010000111110001101;
assign LUT_3[10409] = 32'b00000000000000010111101001101010;
assign LUT_3[10410] = 32'b00000000000000010011000101110001;
assign LUT_3[10411] = 32'b00000000000000011001110001001110;
assign LUT_3[10412] = 32'b00000000000000001110001100000011;
assign LUT_3[10413] = 32'b00000000000000010100110111100000;
assign LUT_3[10414] = 32'b00000000000000010000010011100111;
assign LUT_3[10415] = 32'b00000000000000010110111111000100;
assign LUT_3[10416] = 32'b00000000000000001110111000001010;
assign LUT_3[10417] = 32'b00000000000000010101100011100111;
assign LUT_3[10418] = 32'b00000000000000010000111111101110;
assign LUT_3[10419] = 32'b00000000000000010111101011001011;
assign LUT_3[10420] = 32'b00000000000000001100000110000000;
assign LUT_3[10421] = 32'b00000000000000010010110001011101;
assign LUT_3[10422] = 32'b00000000000000001110001101100100;
assign LUT_3[10423] = 32'b00000000000000010100111001000001;
assign LUT_3[10424] = 32'b00000000000000010100010001010000;
assign LUT_3[10425] = 32'b00000000000000011010111100101101;
assign LUT_3[10426] = 32'b00000000000000010110011000110100;
assign LUT_3[10427] = 32'b00000000000000011101000100010001;
assign LUT_3[10428] = 32'b00000000000000010001011111000110;
assign LUT_3[10429] = 32'b00000000000000011000001010100011;
assign LUT_3[10430] = 32'b00000000000000010011100110101010;
assign LUT_3[10431] = 32'b00000000000000011010010010000111;
assign LUT_3[10432] = 32'b00000000000000001010001111010010;
assign LUT_3[10433] = 32'b00000000000000010000111010101111;
assign LUT_3[10434] = 32'b00000000000000001100010110110110;
assign LUT_3[10435] = 32'b00000000000000010011000010010011;
assign LUT_3[10436] = 32'b00000000000000000111011101001000;
assign LUT_3[10437] = 32'b00000000000000001110001000100101;
assign LUT_3[10438] = 32'b00000000000000001001100100101100;
assign LUT_3[10439] = 32'b00000000000000010000010000001001;
assign LUT_3[10440] = 32'b00000000000000001111101000011000;
assign LUT_3[10441] = 32'b00000000000000010110010011110101;
assign LUT_3[10442] = 32'b00000000000000010001101111111100;
assign LUT_3[10443] = 32'b00000000000000011000011011011001;
assign LUT_3[10444] = 32'b00000000000000001100110110001110;
assign LUT_3[10445] = 32'b00000000000000010011100001101011;
assign LUT_3[10446] = 32'b00000000000000001110111101110010;
assign LUT_3[10447] = 32'b00000000000000010101101001001111;
assign LUT_3[10448] = 32'b00000000000000001101100010010101;
assign LUT_3[10449] = 32'b00000000000000010100001101110010;
assign LUT_3[10450] = 32'b00000000000000001111101001111001;
assign LUT_3[10451] = 32'b00000000000000010110010101010110;
assign LUT_3[10452] = 32'b00000000000000001010110000001011;
assign LUT_3[10453] = 32'b00000000000000010001011011101000;
assign LUT_3[10454] = 32'b00000000000000001100110111101111;
assign LUT_3[10455] = 32'b00000000000000010011100011001100;
assign LUT_3[10456] = 32'b00000000000000010010111011011011;
assign LUT_3[10457] = 32'b00000000000000011001100110111000;
assign LUT_3[10458] = 32'b00000000000000010101000010111111;
assign LUT_3[10459] = 32'b00000000000000011011101110011100;
assign LUT_3[10460] = 32'b00000000000000010000001001010001;
assign LUT_3[10461] = 32'b00000000000000010110110100101110;
assign LUT_3[10462] = 32'b00000000000000010010010000110101;
assign LUT_3[10463] = 32'b00000000000000011000111100010010;
assign LUT_3[10464] = 32'b00000000000000001011011101110010;
assign LUT_3[10465] = 32'b00000000000000010010001001001111;
assign LUT_3[10466] = 32'b00000000000000001101100101010110;
assign LUT_3[10467] = 32'b00000000000000010100010000110011;
assign LUT_3[10468] = 32'b00000000000000001000101011101000;
assign LUT_3[10469] = 32'b00000000000000001111010111000101;
assign LUT_3[10470] = 32'b00000000000000001010110011001100;
assign LUT_3[10471] = 32'b00000000000000010001011110101001;
assign LUT_3[10472] = 32'b00000000000000010000110110111000;
assign LUT_3[10473] = 32'b00000000000000010111100010010101;
assign LUT_3[10474] = 32'b00000000000000010010111110011100;
assign LUT_3[10475] = 32'b00000000000000011001101001111001;
assign LUT_3[10476] = 32'b00000000000000001110000100101110;
assign LUT_3[10477] = 32'b00000000000000010100110000001011;
assign LUT_3[10478] = 32'b00000000000000010000001100010010;
assign LUT_3[10479] = 32'b00000000000000010110110111101111;
assign LUT_3[10480] = 32'b00000000000000001110110000110101;
assign LUT_3[10481] = 32'b00000000000000010101011100010010;
assign LUT_3[10482] = 32'b00000000000000010000111000011001;
assign LUT_3[10483] = 32'b00000000000000010111100011110110;
assign LUT_3[10484] = 32'b00000000000000001011111110101011;
assign LUT_3[10485] = 32'b00000000000000010010101010001000;
assign LUT_3[10486] = 32'b00000000000000001110000110001111;
assign LUT_3[10487] = 32'b00000000000000010100110001101100;
assign LUT_3[10488] = 32'b00000000000000010100001001111011;
assign LUT_3[10489] = 32'b00000000000000011010110101011000;
assign LUT_3[10490] = 32'b00000000000000010110010001011111;
assign LUT_3[10491] = 32'b00000000000000011100111100111100;
assign LUT_3[10492] = 32'b00000000000000010001010111110001;
assign LUT_3[10493] = 32'b00000000000000011000000011001110;
assign LUT_3[10494] = 32'b00000000000000010011011111010101;
assign LUT_3[10495] = 32'b00000000000000011010001010110010;
assign LUT_3[10496] = 32'b00000000000000000100011011001010;
assign LUT_3[10497] = 32'b00000000000000001011000110100111;
assign LUT_3[10498] = 32'b00000000000000000110100010101110;
assign LUT_3[10499] = 32'b00000000000000001101001110001011;
assign LUT_3[10500] = 32'b00000000000000000001101001000000;
assign LUT_3[10501] = 32'b00000000000000001000010100011101;
assign LUT_3[10502] = 32'b00000000000000000011110000100100;
assign LUT_3[10503] = 32'b00000000000000001010011100000001;
assign LUT_3[10504] = 32'b00000000000000001001110100010000;
assign LUT_3[10505] = 32'b00000000000000010000011111101101;
assign LUT_3[10506] = 32'b00000000000000001011111011110100;
assign LUT_3[10507] = 32'b00000000000000010010100111010001;
assign LUT_3[10508] = 32'b00000000000000000111000010000110;
assign LUT_3[10509] = 32'b00000000000000001101101101100011;
assign LUT_3[10510] = 32'b00000000000000001001001001101010;
assign LUT_3[10511] = 32'b00000000000000001111110101000111;
assign LUT_3[10512] = 32'b00000000000000000111101110001101;
assign LUT_3[10513] = 32'b00000000000000001110011001101010;
assign LUT_3[10514] = 32'b00000000000000001001110101110001;
assign LUT_3[10515] = 32'b00000000000000010000100001001110;
assign LUT_3[10516] = 32'b00000000000000000100111100000011;
assign LUT_3[10517] = 32'b00000000000000001011100111100000;
assign LUT_3[10518] = 32'b00000000000000000111000011100111;
assign LUT_3[10519] = 32'b00000000000000001101101111000100;
assign LUT_3[10520] = 32'b00000000000000001101000111010011;
assign LUT_3[10521] = 32'b00000000000000010011110010110000;
assign LUT_3[10522] = 32'b00000000000000001111001110110111;
assign LUT_3[10523] = 32'b00000000000000010101111010010100;
assign LUT_3[10524] = 32'b00000000000000001010010101001001;
assign LUT_3[10525] = 32'b00000000000000010001000000100110;
assign LUT_3[10526] = 32'b00000000000000001100011100101101;
assign LUT_3[10527] = 32'b00000000000000010011001000001010;
assign LUT_3[10528] = 32'b00000000000000000101101001101010;
assign LUT_3[10529] = 32'b00000000000000001100010101000111;
assign LUT_3[10530] = 32'b00000000000000000111110001001110;
assign LUT_3[10531] = 32'b00000000000000001110011100101011;
assign LUT_3[10532] = 32'b00000000000000000010110111100000;
assign LUT_3[10533] = 32'b00000000000000001001100010111101;
assign LUT_3[10534] = 32'b00000000000000000100111111000100;
assign LUT_3[10535] = 32'b00000000000000001011101010100001;
assign LUT_3[10536] = 32'b00000000000000001011000010110000;
assign LUT_3[10537] = 32'b00000000000000010001101110001101;
assign LUT_3[10538] = 32'b00000000000000001101001010010100;
assign LUT_3[10539] = 32'b00000000000000010011110101110001;
assign LUT_3[10540] = 32'b00000000000000001000010000100110;
assign LUT_3[10541] = 32'b00000000000000001110111100000011;
assign LUT_3[10542] = 32'b00000000000000001010011000001010;
assign LUT_3[10543] = 32'b00000000000000010001000011100111;
assign LUT_3[10544] = 32'b00000000000000001000111100101101;
assign LUT_3[10545] = 32'b00000000000000001111101000001010;
assign LUT_3[10546] = 32'b00000000000000001011000100010001;
assign LUT_3[10547] = 32'b00000000000000010001101111101110;
assign LUT_3[10548] = 32'b00000000000000000110001010100011;
assign LUT_3[10549] = 32'b00000000000000001100110110000000;
assign LUT_3[10550] = 32'b00000000000000001000010010000111;
assign LUT_3[10551] = 32'b00000000000000001110111101100100;
assign LUT_3[10552] = 32'b00000000000000001110010101110011;
assign LUT_3[10553] = 32'b00000000000000010101000001010000;
assign LUT_3[10554] = 32'b00000000000000010000011101010111;
assign LUT_3[10555] = 32'b00000000000000010111001000110100;
assign LUT_3[10556] = 32'b00000000000000001011100011101001;
assign LUT_3[10557] = 32'b00000000000000010010001111000110;
assign LUT_3[10558] = 32'b00000000000000001101101011001101;
assign LUT_3[10559] = 32'b00000000000000010100010110101010;
assign LUT_3[10560] = 32'b00000000000000000100010011110101;
assign LUT_3[10561] = 32'b00000000000000001010111111010010;
assign LUT_3[10562] = 32'b00000000000000000110011011011001;
assign LUT_3[10563] = 32'b00000000000000001101000110110110;
assign LUT_3[10564] = 32'b00000000000000000001100001101011;
assign LUT_3[10565] = 32'b00000000000000001000001101001000;
assign LUT_3[10566] = 32'b00000000000000000011101001001111;
assign LUT_3[10567] = 32'b00000000000000001010010100101100;
assign LUT_3[10568] = 32'b00000000000000001001101100111011;
assign LUT_3[10569] = 32'b00000000000000010000011000011000;
assign LUT_3[10570] = 32'b00000000000000001011110100011111;
assign LUT_3[10571] = 32'b00000000000000010010011111111100;
assign LUT_3[10572] = 32'b00000000000000000110111010110001;
assign LUT_3[10573] = 32'b00000000000000001101100110001110;
assign LUT_3[10574] = 32'b00000000000000001001000010010101;
assign LUT_3[10575] = 32'b00000000000000001111101101110010;
assign LUT_3[10576] = 32'b00000000000000000111100110111000;
assign LUT_3[10577] = 32'b00000000000000001110010010010101;
assign LUT_3[10578] = 32'b00000000000000001001101110011100;
assign LUT_3[10579] = 32'b00000000000000010000011001111001;
assign LUT_3[10580] = 32'b00000000000000000100110100101110;
assign LUT_3[10581] = 32'b00000000000000001011100000001011;
assign LUT_3[10582] = 32'b00000000000000000110111100010010;
assign LUT_3[10583] = 32'b00000000000000001101100111101111;
assign LUT_3[10584] = 32'b00000000000000001100111111111110;
assign LUT_3[10585] = 32'b00000000000000010011101011011011;
assign LUT_3[10586] = 32'b00000000000000001111000111100010;
assign LUT_3[10587] = 32'b00000000000000010101110010111111;
assign LUT_3[10588] = 32'b00000000000000001010001101110100;
assign LUT_3[10589] = 32'b00000000000000010000111001010001;
assign LUT_3[10590] = 32'b00000000000000001100010101011000;
assign LUT_3[10591] = 32'b00000000000000010011000000110101;
assign LUT_3[10592] = 32'b00000000000000000101100010010101;
assign LUT_3[10593] = 32'b00000000000000001100001101110010;
assign LUT_3[10594] = 32'b00000000000000000111101001111001;
assign LUT_3[10595] = 32'b00000000000000001110010101010110;
assign LUT_3[10596] = 32'b00000000000000000010110000001011;
assign LUT_3[10597] = 32'b00000000000000001001011011101000;
assign LUT_3[10598] = 32'b00000000000000000100110111101111;
assign LUT_3[10599] = 32'b00000000000000001011100011001100;
assign LUT_3[10600] = 32'b00000000000000001010111011011011;
assign LUT_3[10601] = 32'b00000000000000010001100110111000;
assign LUT_3[10602] = 32'b00000000000000001101000010111111;
assign LUT_3[10603] = 32'b00000000000000010011101110011100;
assign LUT_3[10604] = 32'b00000000000000001000001001010001;
assign LUT_3[10605] = 32'b00000000000000001110110100101110;
assign LUT_3[10606] = 32'b00000000000000001010010000110101;
assign LUT_3[10607] = 32'b00000000000000010000111100010010;
assign LUT_3[10608] = 32'b00000000000000001000110101011000;
assign LUT_3[10609] = 32'b00000000000000001111100000110101;
assign LUT_3[10610] = 32'b00000000000000001010111100111100;
assign LUT_3[10611] = 32'b00000000000000010001101000011001;
assign LUT_3[10612] = 32'b00000000000000000110000011001110;
assign LUT_3[10613] = 32'b00000000000000001100101110101011;
assign LUT_3[10614] = 32'b00000000000000001000001010110010;
assign LUT_3[10615] = 32'b00000000000000001110110110001111;
assign LUT_3[10616] = 32'b00000000000000001110001110011110;
assign LUT_3[10617] = 32'b00000000000000010100111001111011;
assign LUT_3[10618] = 32'b00000000000000010000010110000010;
assign LUT_3[10619] = 32'b00000000000000010111000001011111;
assign LUT_3[10620] = 32'b00000000000000001011011100010100;
assign LUT_3[10621] = 32'b00000000000000010010000111110001;
assign LUT_3[10622] = 32'b00000000000000001101100011111000;
assign LUT_3[10623] = 32'b00000000000000010100001111010101;
assign LUT_3[10624] = 32'b00000000000000000110100110001000;
assign LUT_3[10625] = 32'b00000000000000001101010001100101;
assign LUT_3[10626] = 32'b00000000000000001000101101101100;
assign LUT_3[10627] = 32'b00000000000000001111011001001001;
assign LUT_3[10628] = 32'b00000000000000000011110011111110;
assign LUT_3[10629] = 32'b00000000000000001010011111011011;
assign LUT_3[10630] = 32'b00000000000000000101111011100010;
assign LUT_3[10631] = 32'b00000000000000001100100110111111;
assign LUT_3[10632] = 32'b00000000000000001011111111001110;
assign LUT_3[10633] = 32'b00000000000000010010101010101011;
assign LUT_3[10634] = 32'b00000000000000001110000110110010;
assign LUT_3[10635] = 32'b00000000000000010100110010001111;
assign LUT_3[10636] = 32'b00000000000000001001001101000100;
assign LUT_3[10637] = 32'b00000000000000001111111000100001;
assign LUT_3[10638] = 32'b00000000000000001011010100101000;
assign LUT_3[10639] = 32'b00000000000000010010000000000101;
assign LUT_3[10640] = 32'b00000000000000001001111001001011;
assign LUT_3[10641] = 32'b00000000000000010000100100101000;
assign LUT_3[10642] = 32'b00000000000000001100000000101111;
assign LUT_3[10643] = 32'b00000000000000010010101100001100;
assign LUT_3[10644] = 32'b00000000000000000111000111000001;
assign LUT_3[10645] = 32'b00000000000000001101110010011110;
assign LUT_3[10646] = 32'b00000000000000001001001110100101;
assign LUT_3[10647] = 32'b00000000000000001111111010000010;
assign LUT_3[10648] = 32'b00000000000000001111010010010001;
assign LUT_3[10649] = 32'b00000000000000010101111101101110;
assign LUT_3[10650] = 32'b00000000000000010001011001110101;
assign LUT_3[10651] = 32'b00000000000000011000000101010010;
assign LUT_3[10652] = 32'b00000000000000001100100000000111;
assign LUT_3[10653] = 32'b00000000000000010011001011100100;
assign LUT_3[10654] = 32'b00000000000000001110100111101011;
assign LUT_3[10655] = 32'b00000000000000010101010011001000;
assign LUT_3[10656] = 32'b00000000000000000111110100101000;
assign LUT_3[10657] = 32'b00000000000000001110100000000101;
assign LUT_3[10658] = 32'b00000000000000001001111100001100;
assign LUT_3[10659] = 32'b00000000000000010000100111101001;
assign LUT_3[10660] = 32'b00000000000000000101000010011110;
assign LUT_3[10661] = 32'b00000000000000001011101101111011;
assign LUT_3[10662] = 32'b00000000000000000111001010000010;
assign LUT_3[10663] = 32'b00000000000000001101110101011111;
assign LUT_3[10664] = 32'b00000000000000001101001101101110;
assign LUT_3[10665] = 32'b00000000000000010011111001001011;
assign LUT_3[10666] = 32'b00000000000000001111010101010010;
assign LUT_3[10667] = 32'b00000000000000010110000000101111;
assign LUT_3[10668] = 32'b00000000000000001010011011100100;
assign LUT_3[10669] = 32'b00000000000000010001000111000001;
assign LUT_3[10670] = 32'b00000000000000001100100011001000;
assign LUT_3[10671] = 32'b00000000000000010011001110100101;
assign LUT_3[10672] = 32'b00000000000000001011000111101011;
assign LUT_3[10673] = 32'b00000000000000010001110011001000;
assign LUT_3[10674] = 32'b00000000000000001101001111001111;
assign LUT_3[10675] = 32'b00000000000000010011111010101100;
assign LUT_3[10676] = 32'b00000000000000001000010101100001;
assign LUT_3[10677] = 32'b00000000000000001111000000111110;
assign LUT_3[10678] = 32'b00000000000000001010011101000101;
assign LUT_3[10679] = 32'b00000000000000010001001000100010;
assign LUT_3[10680] = 32'b00000000000000010000100000110001;
assign LUT_3[10681] = 32'b00000000000000010111001100001110;
assign LUT_3[10682] = 32'b00000000000000010010101000010101;
assign LUT_3[10683] = 32'b00000000000000011001010011110010;
assign LUT_3[10684] = 32'b00000000000000001101101110100111;
assign LUT_3[10685] = 32'b00000000000000010100011010000100;
assign LUT_3[10686] = 32'b00000000000000001111110110001011;
assign LUT_3[10687] = 32'b00000000000000010110100001101000;
assign LUT_3[10688] = 32'b00000000000000000110011110110011;
assign LUT_3[10689] = 32'b00000000000000001101001010010000;
assign LUT_3[10690] = 32'b00000000000000001000100110010111;
assign LUT_3[10691] = 32'b00000000000000001111010001110100;
assign LUT_3[10692] = 32'b00000000000000000011101100101001;
assign LUT_3[10693] = 32'b00000000000000001010011000000110;
assign LUT_3[10694] = 32'b00000000000000000101110100001101;
assign LUT_3[10695] = 32'b00000000000000001100011111101010;
assign LUT_3[10696] = 32'b00000000000000001011110111111001;
assign LUT_3[10697] = 32'b00000000000000010010100011010110;
assign LUT_3[10698] = 32'b00000000000000001101111111011101;
assign LUT_3[10699] = 32'b00000000000000010100101010111010;
assign LUT_3[10700] = 32'b00000000000000001001000101101111;
assign LUT_3[10701] = 32'b00000000000000001111110001001100;
assign LUT_3[10702] = 32'b00000000000000001011001101010011;
assign LUT_3[10703] = 32'b00000000000000010001111000110000;
assign LUT_3[10704] = 32'b00000000000000001001110001110110;
assign LUT_3[10705] = 32'b00000000000000010000011101010011;
assign LUT_3[10706] = 32'b00000000000000001011111001011010;
assign LUT_3[10707] = 32'b00000000000000010010100100110111;
assign LUT_3[10708] = 32'b00000000000000000110111111101100;
assign LUT_3[10709] = 32'b00000000000000001101101011001001;
assign LUT_3[10710] = 32'b00000000000000001001000111010000;
assign LUT_3[10711] = 32'b00000000000000001111110010101101;
assign LUT_3[10712] = 32'b00000000000000001111001010111100;
assign LUT_3[10713] = 32'b00000000000000010101110110011001;
assign LUT_3[10714] = 32'b00000000000000010001010010100000;
assign LUT_3[10715] = 32'b00000000000000010111111101111101;
assign LUT_3[10716] = 32'b00000000000000001100011000110010;
assign LUT_3[10717] = 32'b00000000000000010011000100001111;
assign LUT_3[10718] = 32'b00000000000000001110100000010110;
assign LUT_3[10719] = 32'b00000000000000010101001011110011;
assign LUT_3[10720] = 32'b00000000000000000111101101010011;
assign LUT_3[10721] = 32'b00000000000000001110011000110000;
assign LUT_3[10722] = 32'b00000000000000001001110100110111;
assign LUT_3[10723] = 32'b00000000000000010000100000010100;
assign LUT_3[10724] = 32'b00000000000000000100111011001001;
assign LUT_3[10725] = 32'b00000000000000001011100110100110;
assign LUT_3[10726] = 32'b00000000000000000111000010101101;
assign LUT_3[10727] = 32'b00000000000000001101101110001010;
assign LUT_3[10728] = 32'b00000000000000001101000110011001;
assign LUT_3[10729] = 32'b00000000000000010011110001110110;
assign LUT_3[10730] = 32'b00000000000000001111001101111101;
assign LUT_3[10731] = 32'b00000000000000010101111001011010;
assign LUT_3[10732] = 32'b00000000000000001010010100001111;
assign LUT_3[10733] = 32'b00000000000000010000111111101100;
assign LUT_3[10734] = 32'b00000000000000001100011011110011;
assign LUT_3[10735] = 32'b00000000000000010011000111010000;
assign LUT_3[10736] = 32'b00000000000000001011000000010110;
assign LUT_3[10737] = 32'b00000000000000010001101011110011;
assign LUT_3[10738] = 32'b00000000000000001101000111111010;
assign LUT_3[10739] = 32'b00000000000000010011110011010111;
assign LUT_3[10740] = 32'b00000000000000001000001110001100;
assign LUT_3[10741] = 32'b00000000000000001110111001101001;
assign LUT_3[10742] = 32'b00000000000000001010010101110000;
assign LUT_3[10743] = 32'b00000000000000010001000001001101;
assign LUT_3[10744] = 32'b00000000000000010000011001011100;
assign LUT_3[10745] = 32'b00000000000000010111000100111001;
assign LUT_3[10746] = 32'b00000000000000010010100001000000;
assign LUT_3[10747] = 32'b00000000000000011001001100011101;
assign LUT_3[10748] = 32'b00000000000000001101100111010010;
assign LUT_3[10749] = 32'b00000000000000010100010010101111;
assign LUT_3[10750] = 32'b00000000000000001111101110110110;
assign LUT_3[10751] = 32'b00000000000000010110011010010011;
assign LUT_3[10752] = 32'b00000000000000001011100000110101;
assign LUT_3[10753] = 32'b00000000000000010010001100010010;
assign LUT_3[10754] = 32'b00000000000000001101101000011001;
assign LUT_3[10755] = 32'b00000000000000010100010011110110;
assign LUT_3[10756] = 32'b00000000000000001000101110101011;
assign LUT_3[10757] = 32'b00000000000000001111011010001000;
assign LUT_3[10758] = 32'b00000000000000001010110110001111;
assign LUT_3[10759] = 32'b00000000000000010001100001101100;
assign LUT_3[10760] = 32'b00000000000000010000111001111011;
assign LUT_3[10761] = 32'b00000000000000010111100101011000;
assign LUT_3[10762] = 32'b00000000000000010011000001011111;
assign LUT_3[10763] = 32'b00000000000000011001101100111100;
assign LUT_3[10764] = 32'b00000000000000001110000111110001;
assign LUT_3[10765] = 32'b00000000000000010100110011001110;
assign LUT_3[10766] = 32'b00000000000000010000001111010101;
assign LUT_3[10767] = 32'b00000000000000010110111010110010;
assign LUT_3[10768] = 32'b00000000000000001110110011111000;
assign LUT_3[10769] = 32'b00000000000000010101011111010101;
assign LUT_3[10770] = 32'b00000000000000010000111011011100;
assign LUT_3[10771] = 32'b00000000000000010111100110111001;
assign LUT_3[10772] = 32'b00000000000000001100000001101110;
assign LUT_3[10773] = 32'b00000000000000010010101101001011;
assign LUT_3[10774] = 32'b00000000000000001110001001010010;
assign LUT_3[10775] = 32'b00000000000000010100110100101111;
assign LUT_3[10776] = 32'b00000000000000010100001100111110;
assign LUT_3[10777] = 32'b00000000000000011010111000011011;
assign LUT_3[10778] = 32'b00000000000000010110010100100010;
assign LUT_3[10779] = 32'b00000000000000011100111111111111;
assign LUT_3[10780] = 32'b00000000000000010001011010110100;
assign LUT_3[10781] = 32'b00000000000000011000000110010001;
assign LUT_3[10782] = 32'b00000000000000010011100010011000;
assign LUT_3[10783] = 32'b00000000000000011010001101110101;
assign LUT_3[10784] = 32'b00000000000000001100101111010101;
assign LUT_3[10785] = 32'b00000000000000010011011010110010;
assign LUT_3[10786] = 32'b00000000000000001110110110111001;
assign LUT_3[10787] = 32'b00000000000000010101100010010110;
assign LUT_3[10788] = 32'b00000000000000001001111101001011;
assign LUT_3[10789] = 32'b00000000000000010000101000101000;
assign LUT_3[10790] = 32'b00000000000000001100000100101111;
assign LUT_3[10791] = 32'b00000000000000010010110000001100;
assign LUT_3[10792] = 32'b00000000000000010010001000011011;
assign LUT_3[10793] = 32'b00000000000000011000110011111000;
assign LUT_3[10794] = 32'b00000000000000010100001111111111;
assign LUT_3[10795] = 32'b00000000000000011010111011011100;
assign LUT_3[10796] = 32'b00000000000000001111010110010001;
assign LUT_3[10797] = 32'b00000000000000010110000001101110;
assign LUT_3[10798] = 32'b00000000000000010001011101110101;
assign LUT_3[10799] = 32'b00000000000000011000001001010010;
assign LUT_3[10800] = 32'b00000000000000010000000010011000;
assign LUT_3[10801] = 32'b00000000000000010110101101110101;
assign LUT_3[10802] = 32'b00000000000000010010001001111100;
assign LUT_3[10803] = 32'b00000000000000011000110101011001;
assign LUT_3[10804] = 32'b00000000000000001101010000001110;
assign LUT_3[10805] = 32'b00000000000000010011111011101011;
assign LUT_3[10806] = 32'b00000000000000001111010111110010;
assign LUT_3[10807] = 32'b00000000000000010110000011001111;
assign LUT_3[10808] = 32'b00000000000000010101011011011110;
assign LUT_3[10809] = 32'b00000000000000011100000110111011;
assign LUT_3[10810] = 32'b00000000000000010111100011000010;
assign LUT_3[10811] = 32'b00000000000000011110001110011111;
assign LUT_3[10812] = 32'b00000000000000010010101001010100;
assign LUT_3[10813] = 32'b00000000000000011001010100110001;
assign LUT_3[10814] = 32'b00000000000000010100110000111000;
assign LUT_3[10815] = 32'b00000000000000011011011100010101;
assign LUT_3[10816] = 32'b00000000000000001011011001100000;
assign LUT_3[10817] = 32'b00000000000000010010000100111101;
assign LUT_3[10818] = 32'b00000000000000001101100001000100;
assign LUT_3[10819] = 32'b00000000000000010100001100100001;
assign LUT_3[10820] = 32'b00000000000000001000100111010110;
assign LUT_3[10821] = 32'b00000000000000001111010010110011;
assign LUT_3[10822] = 32'b00000000000000001010101110111010;
assign LUT_3[10823] = 32'b00000000000000010001011010010111;
assign LUT_3[10824] = 32'b00000000000000010000110010100110;
assign LUT_3[10825] = 32'b00000000000000010111011110000011;
assign LUT_3[10826] = 32'b00000000000000010010111010001010;
assign LUT_3[10827] = 32'b00000000000000011001100101100111;
assign LUT_3[10828] = 32'b00000000000000001110000000011100;
assign LUT_3[10829] = 32'b00000000000000010100101011111001;
assign LUT_3[10830] = 32'b00000000000000010000001000000000;
assign LUT_3[10831] = 32'b00000000000000010110110011011101;
assign LUT_3[10832] = 32'b00000000000000001110101100100011;
assign LUT_3[10833] = 32'b00000000000000010101011000000000;
assign LUT_3[10834] = 32'b00000000000000010000110100000111;
assign LUT_3[10835] = 32'b00000000000000010111011111100100;
assign LUT_3[10836] = 32'b00000000000000001011111010011001;
assign LUT_3[10837] = 32'b00000000000000010010100101110110;
assign LUT_3[10838] = 32'b00000000000000001110000001111101;
assign LUT_3[10839] = 32'b00000000000000010100101101011010;
assign LUT_3[10840] = 32'b00000000000000010100000101101001;
assign LUT_3[10841] = 32'b00000000000000011010110001000110;
assign LUT_3[10842] = 32'b00000000000000010110001101001101;
assign LUT_3[10843] = 32'b00000000000000011100111000101010;
assign LUT_3[10844] = 32'b00000000000000010001010011011111;
assign LUT_3[10845] = 32'b00000000000000010111111110111100;
assign LUT_3[10846] = 32'b00000000000000010011011011000011;
assign LUT_3[10847] = 32'b00000000000000011010000110100000;
assign LUT_3[10848] = 32'b00000000000000001100101000000000;
assign LUT_3[10849] = 32'b00000000000000010011010011011101;
assign LUT_3[10850] = 32'b00000000000000001110101111100100;
assign LUT_3[10851] = 32'b00000000000000010101011011000001;
assign LUT_3[10852] = 32'b00000000000000001001110101110110;
assign LUT_3[10853] = 32'b00000000000000010000100001010011;
assign LUT_3[10854] = 32'b00000000000000001011111101011010;
assign LUT_3[10855] = 32'b00000000000000010010101000110111;
assign LUT_3[10856] = 32'b00000000000000010010000001000110;
assign LUT_3[10857] = 32'b00000000000000011000101100100011;
assign LUT_3[10858] = 32'b00000000000000010100001000101010;
assign LUT_3[10859] = 32'b00000000000000011010110100000111;
assign LUT_3[10860] = 32'b00000000000000001111001110111100;
assign LUT_3[10861] = 32'b00000000000000010101111010011001;
assign LUT_3[10862] = 32'b00000000000000010001010110100000;
assign LUT_3[10863] = 32'b00000000000000011000000001111101;
assign LUT_3[10864] = 32'b00000000000000001111111011000011;
assign LUT_3[10865] = 32'b00000000000000010110100110100000;
assign LUT_3[10866] = 32'b00000000000000010010000010100111;
assign LUT_3[10867] = 32'b00000000000000011000101110000100;
assign LUT_3[10868] = 32'b00000000000000001101001000111001;
assign LUT_3[10869] = 32'b00000000000000010011110100010110;
assign LUT_3[10870] = 32'b00000000000000001111010000011101;
assign LUT_3[10871] = 32'b00000000000000010101111011111010;
assign LUT_3[10872] = 32'b00000000000000010101010100001001;
assign LUT_3[10873] = 32'b00000000000000011011111111100110;
assign LUT_3[10874] = 32'b00000000000000010111011011101101;
assign LUT_3[10875] = 32'b00000000000000011110000111001010;
assign LUT_3[10876] = 32'b00000000000000010010100001111111;
assign LUT_3[10877] = 32'b00000000000000011001001101011100;
assign LUT_3[10878] = 32'b00000000000000010100101001100011;
assign LUT_3[10879] = 32'b00000000000000011011010101000000;
assign LUT_3[10880] = 32'b00000000000000001101101011110011;
assign LUT_3[10881] = 32'b00000000000000010100010111010000;
assign LUT_3[10882] = 32'b00000000000000001111110011010111;
assign LUT_3[10883] = 32'b00000000000000010110011110110100;
assign LUT_3[10884] = 32'b00000000000000001010111001101001;
assign LUT_3[10885] = 32'b00000000000000010001100101000110;
assign LUT_3[10886] = 32'b00000000000000001101000001001101;
assign LUT_3[10887] = 32'b00000000000000010011101100101010;
assign LUT_3[10888] = 32'b00000000000000010011000100111001;
assign LUT_3[10889] = 32'b00000000000000011001110000010110;
assign LUT_3[10890] = 32'b00000000000000010101001100011101;
assign LUT_3[10891] = 32'b00000000000000011011110111111010;
assign LUT_3[10892] = 32'b00000000000000010000010010101111;
assign LUT_3[10893] = 32'b00000000000000010110111110001100;
assign LUT_3[10894] = 32'b00000000000000010010011010010011;
assign LUT_3[10895] = 32'b00000000000000011001000101110000;
assign LUT_3[10896] = 32'b00000000000000010000111110110110;
assign LUT_3[10897] = 32'b00000000000000010111101010010011;
assign LUT_3[10898] = 32'b00000000000000010011000110011010;
assign LUT_3[10899] = 32'b00000000000000011001110001110111;
assign LUT_3[10900] = 32'b00000000000000001110001100101100;
assign LUT_3[10901] = 32'b00000000000000010100111000001001;
assign LUT_3[10902] = 32'b00000000000000010000010100010000;
assign LUT_3[10903] = 32'b00000000000000010110111111101101;
assign LUT_3[10904] = 32'b00000000000000010110010111111100;
assign LUT_3[10905] = 32'b00000000000000011101000011011001;
assign LUT_3[10906] = 32'b00000000000000011000011111100000;
assign LUT_3[10907] = 32'b00000000000000011111001010111101;
assign LUT_3[10908] = 32'b00000000000000010011100101110010;
assign LUT_3[10909] = 32'b00000000000000011010010001001111;
assign LUT_3[10910] = 32'b00000000000000010101101101010110;
assign LUT_3[10911] = 32'b00000000000000011100011000110011;
assign LUT_3[10912] = 32'b00000000000000001110111010010011;
assign LUT_3[10913] = 32'b00000000000000010101100101110000;
assign LUT_3[10914] = 32'b00000000000000010001000001110111;
assign LUT_3[10915] = 32'b00000000000000010111101101010100;
assign LUT_3[10916] = 32'b00000000000000001100001000001001;
assign LUT_3[10917] = 32'b00000000000000010010110011100110;
assign LUT_3[10918] = 32'b00000000000000001110001111101101;
assign LUT_3[10919] = 32'b00000000000000010100111011001010;
assign LUT_3[10920] = 32'b00000000000000010100010011011001;
assign LUT_3[10921] = 32'b00000000000000011010111110110110;
assign LUT_3[10922] = 32'b00000000000000010110011010111101;
assign LUT_3[10923] = 32'b00000000000000011101000110011010;
assign LUT_3[10924] = 32'b00000000000000010001100001001111;
assign LUT_3[10925] = 32'b00000000000000011000001100101100;
assign LUT_3[10926] = 32'b00000000000000010011101000110011;
assign LUT_3[10927] = 32'b00000000000000011010010100010000;
assign LUT_3[10928] = 32'b00000000000000010010001101010110;
assign LUT_3[10929] = 32'b00000000000000011000111000110011;
assign LUT_3[10930] = 32'b00000000000000010100010100111010;
assign LUT_3[10931] = 32'b00000000000000011011000000010111;
assign LUT_3[10932] = 32'b00000000000000001111011011001100;
assign LUT_3[10933] = 32'b00000000000000010110000110101001;
assign LUT_3[10934] = 32'b00000000000000010001100010110000;
assign LUT_3[10935] = 32'b00000000000000011000001110001101;
assign LUT_3[10936] = 32'b00000000000000010111100110011100;
assign LUT_3[10937] = 32'b00000000000000011110010001111001;
assign LUT_3[10938] = 32'b00000000000000011001101110000000;
assign LUT_3[10939] = 32'b00000000000000100000011001011101;
assign LUT_3[10940] = 32'b00000000000000010100110100010010;
assign LUT_3[10941] = 32'b00000000000000011011011111101111;
assign LUT_3[10942] = 32'b00000000000000010110111011110110;
assign LUT_3[10943] = 32'b00000000000000011101100111010011;
assign LUT_3[10944] = 32'b00000000000000001101100100011110;
assign LUT_3[10945] = 32'b00000000000000010100001111111011;
assign LUT_3[10946] = 32'b00000000000000001111101100000010;
assign LUT_3[10947] = 32'b00000000000000010110010111011111;
assign LUT_3[10948] = 32'b00000000000000001010110010010100;
assign LUT_3[10949] = 32'b00000000000000010001011101110001;
assign LUT_3[10950] = 32'b00000000000000001100111001111000;
assign LUT_3[10951] = 32'b00000000000000010011100101010101;
assign LUT_3[10952] = 32'b00000000000000010010111101100100;
assign LUT_3[10953] = 32'b00000000000000011001101001000001;
assign LUT_3[10954] = 32'b00000000000000010101000101001000;
assign LUT_3[10955] = 32'b00000000000000011011110000100101;
assign LUT_3[10956] = 32'b00000000000000010000001011011010;
assign LUT_3[10957] = 32'b00000000000000010110110110110111;
assign LUT_3[10958] = 32'b00000000000000010010010010111110;
assign LUT_3[10959] = 32'b00000000000000011000111110011011;
assign LUT_3[10960] = 32'b00000000000000010000110111100001;
assign LUT_3[10961] = 32'b00000000000000010111100010111110;
assign LUT_3[10962] = 32'b00000000000000010010111111000101;
assign LUT_3[10963] = 32'b00000000000000011001101010100010;
assign LUT_3[10964] = 32'b00000000000000001110000101010111;
assign LUT_3[10965] = 32'b00000000000000010100110000110100;
assign LUT_3[10966] = 32'b00000000000000010000001100111011;
assign LUT_3[10967] = 32'b00000000000000010110111000011000;
assign LUT_3[10968] = 32'b00000000000000010110010000100111;
assign LUT_3[10969] = 32'b00000000000000011100111100000100;
assign LUT_3[10970] = 32'b00000000000000011000011000001011;
assign LUT_3[10971] = 32'b00000000000000011111000011101000;
assign LUT_3[10972] = 32'b00000000000000010011011110011101;
assign LUT_3[10973] = 32'b00000000000000011010001001111010;
assign LUT_3[10974] = 32'b00000000000000010101100110000001;
assign LUT_3[10975] = 32'b00000000000000011100010001011110;
assign LUT_3[10976] = 32'b00000000000000001110110010111110;
assign LUT_3[10977] = 32'b00000000000000010101011110011011;
assign LUT_3[10978] = 32'b00000000000000010000111010100010;
assign LUT_3[10979] = 32'b00000000000000010111100101111111;
assign LUT_3[10980] = 32'b00000000000000001100000000110100;
assign LUT_3[10981] = 32'b00000000000000010010101100010001;
assign LUT_3[10982] = 32'b00000000000000001110001000011000;
assign LUT_3[10983] = 32'b00000000000000010100110011110101;
assign LUT_3[10984] = 32'b00000000000000010100001100000100;
assign LUT_3[10985] = 32'b00000000000000011010110111100001;
assign LUT_3[10986] = 32'b00000000000000010110010011101000;
assign LUT_3[10987] = 32'b00000000000000011100111111000101;
assign LUT_3[10988] = 32'b00000000000000010001011001111010;
assign LUT_3[10989] = 32'b00000000000000011000000101010111;
assign LUT_3[10990] = 32'b00000000000000010011100001011110;
assign LUT_3[10991] = 32'b00000000000000011010001100111011;
assign LUT_3[10992] = 32'b00000000000000010010000110000001;
assign LUT_3[10993] = 32'b00000000000000011000110001011110;
assign LUT_3[10994] = 32'b00000000000000010100001101100101;
assign LUT_3[10995] = 32'b00000000000000011010111001000010;
assign LUT_3[10996] = 32'b00000000000000001111010011110111;
assign LUT_3[10997] = 32'b00000000000000010101111111010100;
assign LUT_3[10998] = 32'b00000000000000010001011011011011;
assign LUT_3[10999] = 32'b00000000000000011000000110111000;
assign LUT_3[11000] = 32'b00000000000000010111011111000111;
assign LUT_3[11001] = 32'b00000000000000011110001010100100;
assign LUT_3[11002] = 32'b00000000000000011001100110101011;
assign LUT_3[11003] = 32'b00000000000000100000010010001000;
assign LUT_3[11004] = 32'b00000000000000010100101100111101;
assign LUT_3[11005] = 32'b00000000000000011011011000011010;
assign LUT_3[11006] = 32'b00000000000000010110110100100001;
assign LUT_3[11007] = 32'b00000000000000011101011111111110;
assign LUT_3[11008] = 32'b00000000000000000111110000010110;
assign LUT_3[11009] = 32'b00000000000000001110011011110011;
assign LUT_3[11010] = 32'b00000000000000001001110111111010;
assign LUT_3[11011] = 32'b00000000000000010000100011010111;
assign LUT_3[11012] = 32'b00000000000000000100111110001100;
assign LUT_3[11013] = 32'b00000000000000001011101001101001;
assign LUT_3[11014] = 32'b00000000000000000111000101110000;
assign LUT_3[11015] = 32'b00000000000000001101110001001101;
assign LUT_3[11016] = 32'b00000000000000001101001001011100;
assign LUT_3[11017] = 32'b00000000000000010011110100111001;
assign LUT_3[11018] = 32'b00000000000000001111010001000000;
assign LUT_3[11019] = 32'b00000000000000010101111100011101;
assign LUT_3[11020] = 32'b00000000000000001010010111010010;
assign LUT_3[11021] = 32'b00000000000000010001000010101111;
assign LUT_3[11022] = 32'b00000000000000001100011110110110;
assign LUT_3[11023] = 32'b00000000000000010011001010010011;
assign LUT_3[11024] = 32'b00000000000000001011000011011001;
assign LUT_3[11025] = 32'b00000000000000010001101110110110;
assign LUT_3[11026] = 32'b00000000000000001101001010111101;
assign LUT_3[11027] = 32'b00000000000000010011110110011010;
assign LUT_3[11028] = 32'b00000000000000001000010001001111;
assign LUT_3[11029] = 32'b00000000000000001110111100101100;
assign LUT_3[11030] = 32'b00000000000000001010011000110011;
assign LUT_3[11031] = 32'b00000000000000010001000100010000;
assign LUT_3[11032] = 32'b00000000000000010000011100011111;
assign LUT_3[11033] = 32'b00000000000000010111000111111100;
assign LUT_3[11034] = 32'b00000000000000010010100100000011;
assign LUT_3[11035] = 32'b00000000000000011001001111100000;
assign LUT_3[11036] = 32'b00000000000000001101101010010101;
assign LUT_3[11037] = 32'b00000000000000010100010101110010;
assign LUT_3[11038] = 32'b00000000000000001111110001111001;
assign LUT_3[11039] = 32'b00000000000000010110011101010110;
assign LUT_3[11040] = 32'b00000000000000001000111110110110;
assign LUT_3[11041] = 32'b00000000000000001111101010010011;
assign LUT_3[11042] = 32'b00000000000000001011000110011010;
assign LUT_3[11043] = 32'b00000000000000010001110001110111;
assign LUT_3[11044] = 32'b00000000000000000110001100101100;
assign LUT_3[11045] = 32'b00000000000000001100111000001001;
assign LUT_3[11046] = 32'b00000000000000001000010100010000;
assign LUT_3[11047] = 32'b00000000000000001110111111101101;
assign LUT_3[11048] = 32'b00000000000000001110010111111100;
assign LUT_3[11049] = 32'b00000000000000010101000011011001;
assign LUT_3[11050] = 32'b00000000000000010000011111100000;
assign LUT_3[11051] = 32'b00000000000000010111001010111101;
assign LUT_3[11052] = 32'b00000000000000001011100101110010;
assign LUT_3[11053] = 32'b00000000000000010010010001001111;
assign LUT_3[11054] = 32'b00000000000000001101101101010110;
assign LUT_3[11055] = 32'b00000000000000010100011000110011;
assign LUT_3[11056] = 32'b00000000000000001100010001111001;
assign LUT_3[11057] = 32'b00000000000000010010111101010110;
assign LUT_3[11058] = 32'b00000000000000001110011001011101;
assign LUT_3[11059] = 32'b00000000000000010101000100111010;
assign LUT_3[11060] = 32'b00000000000000001001011111101111;
assign LUT_3[11061] = 32'b00000000000000010000001011001100;
assign LUT_3[11062] = 32'b00000000000000001011100111010011;
assign LUT_3[11063] = 32'b00000000000000010010010010110000;
assign LUT_3[11064] = 32'b00000000000000010001101010111111;
assign LUT_3[11065] = 32'b00000000000000011000010110011100;
assign LUT_3[11066] = 32'b00000000000000010011110010100011;
assign LUT_3[11067] = 32'b00000000000000011010011110000000;
assign LUT_3[11068] = 32'b00000000000000001110111000110101;
assign LUT_3[11069] = 32'b00000000000000010101100100010010;
assign LUT_3[11070] = 32'b00000000000000010001000000011001;
assign LUT_3[11071] = 32'b00000000000000010111101011110110;
assign LUT_3[11072] = 32'b00000000000000000111101001000001;
assign LUT_3[11073] = 32'b00000000000000001110010100011110;
assign LUT_3[11074] = 32'b00000000000000001001110000100101;
assign LUT_3[11075] = 32'b00000000000000010000011100000010;
assign LUT_3[11076] = 32'b00000000000000000100110110110111;
assign LUT_3[11077] = 32'b00000000000000001011100010010100;
assign LUT_3[11078] = 32'b00000000000000000110111110011011;
assign LUT_3[11079] = 32'b00000000000000001101101001111000;
assign LUT_3[11080] = 32'b00000000000000001101000010000111;
assign LUT_3[11081] = 32'b00000000000000010011101101100100;
assign LUT_3[11082] = 32'b00000000000000001111001001101011;
assign LUT_3[11083] = 32'b00000000000000010101110101001000;
assign LUT_3[11084] = 32'b00000000000000001010001111111101;
assign LUT_3[11085] = 32'b00000000000000010000111011011010;
assign LUT_3[11086] = 32'b00000000000000001100010111100001;
assign LUT_3[11087] = 32'b00000000000000010011000010111110;
assign LUT_3[11088] = 32'b00000000000000001010111100000100;
assign LUT_3[11089] = 32'b00000000000000010001100111100001;
assign LUT_3[11090] = 32'b00000000000000001101000011101000;
assign LUT_3[11091] = 32'b00000000000000010011101111000101;
assign LUT_3[11092] = 32'b00000000000000001000001001111010;
assign LUT_3[11093] = 32'b00000000000000001110110101010111;
assign LUT_3[11094] = 32'b00000000000000001010010001011110;
assign LUT_3[11095] = 32'b00000000000000010000111100111011;
assign LUT_3[11096] = 32'b00000000000000010000010101001010;
assign LUT_3[11097] = 32'b00000000000000010111000000100111;
assign LUT_3[11098] = 32'b00000000000000010010011100101110;
assign LUT_3[11099] = 32'b00000000000000011001001000001011;
assign LUT_3[11100] = 32'b00000000000000001101100011000000;
assign LUT_3[11101] = 32'b00000000000000010100001110011101;
assign LUT_3[11102] = 32'b00000000000000001111101010100100;
assign LUT_3[11103] = 32'b00000000000000010110010110000001;
assign LUT_3[11104] = 32'b00000000000000001000110111100001;
assign LUT_3[11105] = 32'b00000000000000001111100010111110;
assign LUT_3[11106] = 32'b00000000000000001010111111000101;
assign LUT_3[11107] = 32'b00000000000000010001101010100010;
assign LUT_3[11108] = 32'b00000000000000000110000101010111;
assign LUT_3[11109] = 32'b00000000000000001100110000110100;
assign LUT_3[11110] = 32'b00000000000000001000001100111011;
assign LUT_3[11111] = 32'b00000000000000001110111000011000;
assign LUT_3[11112] = 32'b00000000000000001110010000100111;
assign LUT_3[11113] = 32'b00000000000000010100111100000100;
assign LUT_3[11114] = 32'b00000000000000010000011000001011;
assign LUT_3[11115] = 32'b00000000000000010111000011101000;
assign LUT_3[11116] = 32'b00000000000000001011011110011101;
assign LUT_3[11117] = 32'b00000000000000010010001001111010;
assign LUT_3[11118] = 32'b00000000000000001101100110000001;
assign LUT_3[11119] = 32'b00000000000000010100010001011110;
assign LUT_3[11120] = 32'b00000000000000001100001010100100;
assign LUT_3[11121] = 32'b00000000000000010010110110000001;
assign LUT_3[11122] = 32'b00000000000000001110010010001000;
assign LUT_3[11123] = 32'b00000000000000010100111101100101;
assign LUT_3[11124] = 32'b00000000000000001001011000011010;
assign LUT_3[11125] = 32'b00000000000000010000000011110111;
assign LUT_3[11126] = 32'b00000000000000001011011111111110;
assign LUT_3[11127] = 32'b00000000000000010010001011011011;
assign LUT_3[11128] = 32'b00000000000000010001100011101010;
assign LUT_3[11129] = 32'b00000000000000011000001111000111;
assign LUT_3[11130] = 32'b00000000000000010011101011001110;
assign LUT_3[11131] = 32'b00000000000000011010010110101011;
assign LUT_3[11132] = 32'b00000000000000001110110001100000;
assign LUT_3[11133] = 32'b00000000000000010101011100111101;
assign LUT_3[11134] = 32'b00000000000000010000111001000100;
assign LUT_3[11135] = 32'b00000000000000010111100100100001;
assign LUT_3[11136] = 32'b00000000000000001001111011010100;
assign LUT_3[11137] = 32'b00000000000000010000100110110001;
assign LUT_3[11138] = 32'b00000000000000001100000010111000;
assign LUT_3[11139] = 32'b00000000000000010010101110010101;
assign LUT_3[11140] = 32'b00000000000000000111001001001010;
assign LUT_3[11141] = 32'b00000000000000001101110100100111;
assign LUT_3[11142] = 32'b00000000000000001001010000101110;
assign LUT_3[11143] = 32'b00000000000000001111111100001011;
assign LUT_3[11144] = 32'b00000000000000001111010100011010;
assign LUT_3[11145] = 32'b00000000000000010101111111110111;
assign LUT_3[11146] = 32'b00000000000000010001011011111110;
assign LUT_3[11147] = 32'b00000000000000011000000111011011;
assign LUT_3[11148] = 32'b00000000000000001100100010010000;
assign LUT_3[11149] = 32'b00000000000000010011001101101101;
assign LUT_3[11150] = 32'b00000000000000001110101001110100;
assign LUT_3[11151] = 32'b00000000000000010101010101010001;
assign LUT_3[11152] = 32'b00000000000000001101001110010111;
assign LUT_3[11153] = 32'b00000000000000010011111001110100;
assign LUT_3[11154] = 32'b00000000000000001111010101111011;
assign LUT_3[11155] = 32'b00000000000000010110000001011000;
assign LUT_3[11156] = 32'b00000000000000001010011100001101;
assign LUT_3[11157] = 32'b00000000000000010001000111101010;
assign LUT_3[11158] = 32'b00000000000000001100100011110001;
assign LUT_3[11159] = 32'b00000000000000010011001111001110;
assign LUT_3[11160] = 32'b00000000000000010010100111011101;
assign LUT_3[11161] = 32'b00000000000000011001010010111010;
assign LUT_3[11162] = 32'b00000000000000010100101111000001;
assign LUT_3[11163] = 32'b00000000000000011011011010011110;
assign LUT_3[11164] = 32'b00000000000000001111110101010011;
assign LUT_3[11165] = 32'b00000000000000010110100000110000;
assign LUT_3[11166] = 32'b00000000000000010001111100110111;
assign LUT_3[11167] = 32'b00000000000000011000101000010100;
assign LUT_3[11168] = 32'b00000000000000001011001001110100;
assign LUT_3[11169] = 32'b00000000000000010001110101010001;
assign LUT_3[11170] = 32'b00000000000000001101010001011000;
assign LUT_3[11171] = 32'b00000000000000010011111100110101;
assign LUT_3[11172] = 32'b00000000000000001000010111101010;
assign LUT_3[11173] = 32'b00000000000000001111000011000111;
assign LUT_3[11174] = 32'b00000000000000001010011111001110;
assign LUT_3[11175] = 32'b00000000000000010001001010101011;
assign LUT_3[11176] = 32'b00000000000000010000100010111010;
assign LUT_3[11177] = 32'b00000000000000010111001110010111;
assign LUT_3[11178] = 32'b00000000000000010010101010011110;
assign LUT_3[11179] = 32'b00000000000000011001010101111011;
assign LUT_3[11180] = 32'b00000000000000001101110000110000;
assign LUT_3[11181] = 32'b00000000000000010100011100001101;
assign LUT_3[11182] = 32'b00000000000000001111111000010100;
assign LUT_3[11183] = 32'b00000000000000010110100011110001;
assign LUT_3[11184] = 32'b00000000000000001110011100110111;
assign LUT_3[11185] = 32'b00000000000000010101001000010100;
assign LUT_3[11186] = 32'b00000000000000010000100100011011;
assign LUT_3[11187] = 32'b00000000000000010111001111111000;
assign LUT_3[11188] = 32'b00000000000000001011101010101101;
assign LUT_3[11189] = 32'b00000000000000010010010110001010;
assign LUT_3[11190] = 32'b00000000000000001101110010010001;
assign LUT_3[11191] = 32'b00000000000000010100011101101110;
assign LUT_3[11192] = 32'b00000000000000010011110101111101;
assign LUT_3[11193] = 32'b00000000000000011010100001011010;
assign LUT_3[11194] = 32'b00000000000000010101111101100001;
assign LUT_3[11195] = 32'b00000000000000011100101000111110;
assign LUT_3[11196] = 32'b00000000000000010001000011110011;
assign LUT_3[11197] = 32'b00000000000000010111101111010000;
assign LUT_3[11198] = 32'b00000000000000010011001011010111;
assign LUT_3[11199] = 32'b00000000000000011001110110110100;
assign LUT_3[11200] = 32'b00000000000000001001110011111111;
assign LUT_3[11201] = 32'b00000000000000010000011111011100;
assign LUT_3[11202] = 32'b00000000000000001011111011100011;
assign LUT_3[11203] = 32'b00000000000000010010100111000000;
assign LUT_3[11204] = 32'b00000000000000000111000001110101;
assign LUT_3[11205] = 32'b00000000000000001101101101010010;
assign LUT_3[11206] = 32'b00000000000000001001001001011001;
assign LUT_3[11207] = 32'b00000000000000001111110100110110;
assign LUT_3[11208] = 32'b00000000000000001111001101000101;
assign LUT_3[11209] = 32'b00000000000000010101111000100010;
assign LUT_3[11210] = 32'b00000000000000010001010100101001;
assign LUT_3[11211] = 32'b00000000000000011000000000000110;
assign LUT_3[11212] = 32'b00000000000000001100011010111011;
assign LUT_3[11213] = 32'b00000000000000010011000110011000;
assign LUT_3[11214] = 32'b00000000000000001110100010011111;
assign LUT_3[11215] = 32'b00000000000000010101001101111100;
assign LUT_3[11216] = 32'b00000000000000001101000111000010;
assign LUT_3[11217] = 32'b00000000000000010011110010011111;
assign LUT_3[11218] = 32'b00000000000000001111001110100110;
assign LUT_3[11219] = 32'b00000000000000010101111010000011;
assign LUT_3[11220] = 32'b00000000000000001010010100111000;
assign LUT_3[11221] = 32'b00000000000000010001000000010101;
assign LUT_3[11222] = 32'b00000000000000001100011100011100;
assign LUT_3[11223] = 32'b00000000000000010011000111111001;
assign LUT_3[11224] = 32'b00000000000000010010100000001000;
assign LUT_3[11225] = 32'b00000000000000011001001011100101;
assign LUT_3[11226] = 32'b00000000000000010100100111101100;
assign LUT_3[11227] = 32'b00000000000000011011010011001001;
assign LUT_3[11228] = 32'b00000000000000001111101101111110;
assign LUT_3[11229] = 32'b00000000000000010110011001011011;
assign LUT_3[11230] = 32'b00000000000000010001110101100010;
assign LUT_3[11231] = 32'b00000000000000011000100000111111;
assign LUT_3[11232] = 32'b00000000000000001011000010011111;
assign LUT_3[11233] = 32'b00000000000000010001101101111100;
assign LUT_3[11234] = 32'b00000000000000001101001010000011;
assign LUT_3[11235] = 32'b00000000000000010011110101100000;
assign LUT_3[11236] = 32'b00000000000000001000010000010101;
assign LUT_3[11237] = 32'b00000000000000001110111011110010;
assign LUT_3[11238] = 32'b00000000000000001010010111111001;
assign LUT_3[11239] = 32'b00000000000000010001000011010110;
assign LUT_3[11240] = 32'b00000000000000010000011011100101;
assign LUT_3[11241] = 32'b00000000000000010111000111000010;
assign LUT_3[11242] = 32'b00000000000000010010100011001001;
assign LUT_3[11243] = 32'b00000000000000011001001110100110;
assign LUT_3[11244] = 32'b00000000000000001101101001011011;
assign LUT_3[11245] = 32'b00000000000000010100010100111000;
assign LUT_3[11246] = 32'b00000000000000001111110000111111;
assign LUT_3[11247] = 32'b00000000000000010110011100011100;
assign LUT_3[11248] = 32'b00000000000000001110010101100010;
assign LUT_3[11249] = 32'b00000000000000010101000000111111;
assign LUT_3[11250] = 32'b00000000000000010000011101000110;
assign LUT_3[11251] = 32'b00000000000000010111001000100011;
assign LUT_3[11252] = 32'b00000000000000001011100011011000;
assign LUT_3[11253] = 32'b00000000000000010010001110110101;
assign LUT_3[11254] = 32'b00000000000000001101101010111100;
assign LUT_3[11255] = 32'b00000000000000010100010110011001;
assign LUT_3[11256] = 32'b00000000000000010011101110101000;
assign LUT_3[11257] = 32'b00000000000000011010011010000101;
assign LUT_3[11258] = 32'b00000000000000010101110110001100;
assign LUT_3[11259] = 32'b00000000000000011100100001101001;
assign LUT_3[11260] = 32'b00000000000000010000111100011110;
assign LUT_3[11261] = 32'b00000000000000010111100111111011;
assign LUT_3[11262] = 32'b00000000000000010011000100000010;
assign LUT_3[11263] = 32'b00000000000000011001101111011111;
assign LUT_3[11264] = 32'b00000000000000001110110000100110;
assign LUT_3[11265] = 32'b00000000000000010101011100000011;
assign LUT_3[11266] = 32'b00000000000000010000111000001010;
assign LUT_3[11267] = 32'b00000000000000010111100011100111;
assign LUT_3[11268] = 32'b00000000000000001011111110011100;
assign LUT_3[11269] = 32'b00000000000000010010101001111001;
assign LUT_3[11270] = 32'b00000000000000001110000110000000;
assign LUT_3[11271] = 32'b00000000000000010100110001011101;
assign LUT_3[11272] = 32'b00000000000000010100001001101100;
assign LUT_3[11273] = 32'b00000000000000011010110101001001;
assign LUT_3[11274] = 32'b00000000000000010110010001010000;
assign LUT_3[11275] = 32'b00000000000000011100111100101101;
assign LUT_3[11276] = 32'b00000000000000010001010111100010;
assign LUT_3[11277] = 32'b00000000000000011000000010111111;
assign LUT_3[11278] = 32'b00000000000000010011011111000110;
assign LUT_3[11279] = 32'b00000000000000011010001010100011;
assign LUT_3[11280] = 32'b00000000000000010010000011101001;
assign LUT_3[11281] = 32'b00000000000000011000101111000110;
assign LUT_3[11282] = 32'b00000000000000010100001011001101;
assign LUT_3[11283] = 32'b00000000000000011010110110101010;
assign LUT_3[11284] = 32'b00000000000000001111010001011111;
assign LUT_3[11285] = 32'b00000000000000010101111100111100;
assign LUT_3[11286] = 32'b00000000000000010001011001000011;
assign LUT_3[11287] = 32'b00000000000000011000000100100000;
assign LUT_3[11288] = 32'b00000000000000010111011100101111;
assign LUT_3[11289] = 32'b00000000000000011110001000001100;
assign LUT_3[11290] = 32'b00000000000000011001100100010011;
assign LUT_3[11291] = 32'b00000000000000100000001111110000;
assign LUT_3[11292] = 32'b00000000000000010100101010100101;
assign LUT_3[11293] = 32'b00000000000000011011010110000010;
assign LUT_3[11294] = 32'b00000000000000010110110010001001;
assign LUT_3[11295] = 32'b00000000000000011101011101100110;
assign LUT_3[11296] = 32'b00000000000000001111111111000110;
assign LUT_3[11297] = 32'b00000000000000010110101010100011;
assign LUT_3[11298] = 32'b00000000000000010010000110101010;
assign LUT_3[11299] = 32'b00000000000000011000110010000111;
assign LUT_3[11300] = 32'b00000000000000001101001100111100;
assign LUT_3[11301] = 32'b00000000000000010011111000011001;
assign LUT_3[11302] = 32'b00000000000000001111010100100000;
assign LUT_3[11303] = 32'b00000000000000010101111111111101;
assign LUT_3[11304] = 32'b00000000000000010101011000001100;
assign LUT_3[11305] = 32'b00000000000000011100000011101001;
assign LUT_3[11306] = 32'b00000000000000010111011111110000;
assign LUT_3[11307] = 32'b00000000000000011110001011001101;
assign LUT_3[11308] = 32'b00000000000000010010100110000010;
assign LUT_3[11309] = 32'b00000000000000011001010001011111;
assign LUT_3[11310] = 32'b00000000000000010100101101100110;
assign LUT_3[11311] = 32'b00000000000000011011011001000011;
assign LUT_3[11312] = 32'b00000000000000010011010010001001;
assign LUT_3[11313] = 32'b00000000000000011001111101100110;
assign LUT_3[11314] = 32'b00000000000000010101011001101101;
assign LUT_3[11315] = 32'b00000000000000011100000101001010;
assign LUT_3[11316] = 32'b00000000000000010000011111111111;
assign LUT_3[11317] = 32'b00000000000000010111001011011100;
assign LUT_3[11318] = 32'b00000000000000010010100111100011;
assign LUT_3[11319] = 32'b00000000000000011001010011000000;
assign LUT_3[11320] = 32'b00000000000000011000101011001111;
assign LUT_3[11321] = 32'b00000000000000011111010110101100;
assign LUT_3[11322] = 32'b00000000000000011010110010110011;
assign LUT_3[11323] = 32'b00000000000000100001011110010000;
assign LUT_3[11324] = 32'b00000000000000010101111001000101;
assign LUT_3[11325] = 32'b00000000000000011100100100100010;
assign LUT_3[11326] = 32'b00000000000000011000000000101001;
assign LUT_3[11327] = 32'b00000000000000011110101100000110;
assign LUT_3[11328] = 32'b00000000000000001110101001010001;
assign LUT_3[11329] = 32'b00000000000000010101010100101110;
assign LUT_3[11330] = 32'b00000000000000010000110000110101;
assign LUT_3[11331] = 32'b00000000000000010111011100010010;
assign LUT_3[11332] = 32'b00000000000000001011110111000111;
assign LUT_3[11333] = 32'b00000000000000010010100010100100;
assign LUT_3[11334] = 32'b00000000000000001101111110101011;
assign LUT_3[11335] = 32'b00000000000000010100101010001000;
assign LUT_3[11336] = 32'b00000000000000010100000010010111;
assign LUT_3[11337] = 32'b00000000000000011010101101110100;
assign LUT_3[11338] = 32'b00000000000000010110001001111011;
assign LUT_3[11339] = 32'b00000000000000011100110101011000;
assign LUT_3[11340] = 32'b00000000000000010001010000001101;
assign LUT_3[11341] = 32'b00000000000000010111111011101010;
assign LUT_3[11342] = 32'b00000000000000010011010111110001;
assign LUT_3[11343] = 32'b00000000000000011010000011001110;
assign LUT_3[11344] = 32'b00000000000000010001111100010100;
assign LUT_3[11345] = 32'b00000000000000011000100111110001;
assign LUT_3[11346] = 32'b00000000000000010100000011111000;
assign LUT_3[11347] = 32'b00000000000000011010101111010101;
assign LUT_3[11348] = 32'b00000000000000001111001010001010;
assign LUT_3[11349] = 32'b00000000000000010101110101100111;
assign LUT_3[11350] = 32'b00000000000000010001010001101110;
assign LUT_3[11351] = 32'b00000000000000010111111101001011;
assign LUT_3[11352] = 32'b00000000000000010111010101011010;
assign LUT_3[11353] = 32'b00000000000000011110000000110111;
assign LUT_3[11354] = 32'b00000000000000011001011100111110;
assign LUT_3[11355] = 32'b00000000000000100000001000011011;
assign LUT_3[11356] = 32'b00000000000000010100100011010000;
assign LUT_3[11357] = 32'b00000000000000011011001110101101;
assign LUT_3[11358] = 32'b00000000000000010110101010110100;
assign LUT_3[11359] = 32'b00000000000000011101010110010001;
assign LUT_3[11360] = 32'b00000000000000001111110111110001;
assign LUT_3[11361] = 32'b00000000000000010110100011001110;
assign LUT_3[11362] = 32'b00000000000000010001111111010101;
assign LUT_3[11363] = 32'b00000000000000011000101010110010;
assign LUT_3[11364] = 32'b00000000000000001101000101100111;
assign LUT_3[11365] = 32'b00000000000000010011110001000100;
assign LUT_3[11366] = 32'b00000000000000001111001101001011;
assign LUT_3[11367] = 32'b00000000000000010101111000101000;
assign LUT_3[11368] = 32'b00000000000000010101010000110111;
assign LUT_3[11369] = 32'b00000000000000011011111100010100;
assign LUT_3[11370] = 32'b00000000000000010111011000011011;
assign LUT_3[11371] = 32'b00000000000000011110000011111000;
assign LUT_3[11372] = 32'b00000000000000010010011110101101;
assign LUT_3[11373] = 32'b00000000000000011001001010001010;
assign LUT_3[11374] = 32'b00000000000000010100100110010001;
assign LUT_3[11375] = 32'b00000000000000011011010001101110;
assign LUT_3[11376] = 32'b00000000000000010011001010110100;
assign LUT_3[11377] = 32'b00000000000000011001110110010001;
assign LUT_3[11378] = 32'b00000000000000010101010010011000;
assign LUT_3[11379] = 32'b00000000000000011011111101110101;
assign LUT_3[11380] = 32'b00000000000000010000011000101010;
assign LUT_3[11381] = 32'b00000000000000010111000100000111;
assign LUT_3[11382] = 32'b00000000000000010010100000001110;
assign LUT_3[11383] = 32'b00000000000000011001001011101011;
assign LUT_3[11384] = 32'b00000000000000011000100011111010;
assign LUT_3[11385] = 32'b00000000000000011111001111010111;
assign LUT_3[11386] = 32'b00000000000000011010101011011110;
assign LUT_3[11387] = 32'b00000000000000100001010110111011;
assign LUT_3[11388] = 32'b00000000000000010101110001110000;
assign LUT_3[11389] = 32'b00000000000000011100011101001101;
assign LUT_3[11390] = 32'b00000000000000010111111001010100;
assign LUT_3[11391] = 32'b00000000000000011110100100110001;
assign LUT_3[11392] = 32'b00000000000000010000111011100100;
assign LUT_3[11393] = 32'b00000000000000010111100111000001;
assign LUT_3[11394] = 32'b00000000000000010011000011001000;
assign LUT_3[11395] = 32'b00000000000000011001101110100101;
assign LUT_3[11396] = 32'b00000000000000001110001001011010;
assign LUT_3[11397] = 32'b00000000000000010100110100110111;
assign LUT_3[11398] = 32'b00000000000000010000010000111110;
assign LUT_3[11399] = 32'b00000000000000010110111100011011;
assign LUT_3[11400] = 32'b00000000000000010110010100101010;
assign LUT_3[11401] = 32'b00000000000000011101000000000111;
assign LUT_3[11402] = 32'b00000000000000011000011100001110;
assign LUT_3[11403] = 32'b00000000000000011111000111101011;
assign LUT_3[11404] = 32'b00000000000000010011100010100000;
assign LUT_3[11405] = 32'b00000000000000011010001101111101;
assign LUT_3[11406] = 32'b00000000000000010101101010000100;
assign LUT_3[11407] = 32'b00000000000000011100010101100001;
assign LUT_3[11408] = 32'b00000000000000010100001110100111;
assign LUT_3[11409] = 32'b00000000000000011010111010000100;
assign LUT_3[11410] = 32'b00000000000000010110010110001011;
assign LUT_3[11411] = 32'b00000000000000011101000001101000;
assign LUT_3[11412] = 32'b00000000000000010001011100011101;
assign LUT_3[11413] = 32'b00000000000000011000000111111010;
assign LUT_3[11414] = 32'b00000000000000010011100100000001;
assign LUT_3[11415] = 32'b00000000000000011010001111011110;
assign LUT_3[11416] = 32'b00000000000000011001100111101101;
assign LUT_3[11417] = 32'b00000000000000100000010011001010;
assign LUT_3[11418] = 32'b00000000000000011011101111010001;
assign LUT_3[11419] = 32'b00000000000000100010011010101110;
assign LUT_3[11420] = 32'b00000000000000010110110101100011;
assign LUT_3[11421] = 32'b00000000000000011101100001000000;
assign LUT_3[11422] = 32'b00000000000000011000111101000111;
assign LUT_3[11423] = 32'b00000000000000011111101000100100;
assign LUT_3[11424] = 32'b00000000000000010010001010000100;
assign LUT_3[11425] = 32'b00000000000000011000110101100001;
assign LUT_3[11426] = 32'b00000000000000010100010001101000;
assign LUT_3[11427] = 32'b00000000000000011010111101000101;
assign LUT_3[11428] = 32'b00000000000000001111010111111010;
assign LUT_3[11429] = 32'b00000000000000010110000011010111;
assign LUT_3[11430] = 32'b00000000000000010001011111011110;
assign LUT_3[11431] = 32'b00000000000000011000001010111011;
assign LUT_3[11432] = 32'b00000000000000010111100011001010;
assign LUT_3[11433] = 32'b00000000000000011110001110100111;
assign LUT_3[11434] = 32'b00000000000000011001101010101110;
assign LUT_3[11435] = 32'b00000000000000100000010110001011;
assign LUT_3[11436] = 32'b00000000000000010100110001000000;
assign LUT_3[11437] = 32'b00000000000000011011011100011101;
assign LUT_3[11438] = 32'b00000000000000010110111000100100;
assign LUT_3[11439] = 32'b00000000000000011101100100000001;
assign LUT_3[11440] = 32'b00000000000000010101011101000111;
assign LUT_3[11441] = 32'b00000000000000011100001000100100;
assign LUT_3[11442] = 32'b00000000000000010111100100101011;
assign LUT_3[11443] = 32'b00000000000000011110010000001000;
assign LUT_3[11444] = 32'b00000000000000010010101010111101;
assign LUT_3[11445] = 32'b00000000000000011001010110011010;
assign LUT_3[11446] = 32'b00000000000000010100110010100001;
assign LUT_3[11447] = 32'b00000000000000011011011101111110;
assign LUT_3[11448] = 32'b00000000000000011010110110001101;
assign LUT_3[11449] = 32'b00000000000000100001100001101010;
assign LUT_3[11450] = 32'b00000000000000011100111101110001;
assign LUT_3[11451] = 32'b00000000000000100011101001001110;
assign LUT_3[11452] = 32'b00000000000000011000000100000011;
assign LUT_3[11453] = 32'b00000000000000011110101111100000;
assign LUT_3[11454] = 32'b00000000000000011010001011100111;
assign LUT_3[11455] = 32'b00000000000000100000110111000100;
assign LUT_3[11456] = 32'b00000000000000010000110100001111;
assign LUT_3[11457] = 32'b00000000000000010111011111101100;
assign LUT_3[11458] = 32'b00000000000000010010111011110011;
assign LUT_3[11459] = 32'b00000000000000011001100111010000;
assign LUT_3[11460] = 32'b00000000000000001110000010000101;
assign LUT_3[11461] = 32'b00000000000000010100101101100010;
assign LUT_3[11462] = 32'b00000000000000010000001001101001;
assign LUT_3[11463] = 32'b00000000000000010110110101000110;
assign LUT_3[11464] = 32'b00000000000000010110001101010101;
assign LUT_3[11465] = 32'b00000000000000011100111000110010;
assign LUT_3[11466] = 32'b00000000000000011000010100111001;
assign LUT_3[11467] = 32'b00000000000000011111000000010110;
assign LUT_3[11468] = 32'b00000000000000010011011011001011;
assign LUT_3[11469] = 32'b00000000000000011010000110101000;
assign LUT_3[11470] = 32'b00000000000000010101100010101111;
assign LUT_3[11471] = 32'b00000000000000011100001110001100;
assign LUT_3[11472] = 32'b00000000000000010100000111010010;
assign LUT_3[11473] = 32'b00000000000000011010110010101111;
assign LUT_3[11474] = 32'b00000000000000010110001110110110;
assign LUT_3[11475] = 32'b00000000000000011100111010010011;
assign LUT_3[11476] = 32'b00000000000000010001010101001000;
assign LUT_3[11477] = 32'b00000000000000011000000000100101;
assign LUT_3[11478] = 32'b00000000000000010011011100101100;
assign LUT_3[11479] = 32'b00000000000000011010001000001001;
assign LUT_3[11480] = 32'b00000000000000011001100000011000;
assign LUT_3[11481] = 32'b00000000000000100000001011110101;
assign LUT_3[11482] = 32'b00000000000000011011100111111100;
assign LUT_3[11483] = 32'b00000000000000100010010011011001;
assign LUT_3[11484] = 32'b00000000000000010110101110001110;
assign LUT_3[11485] = 32'b00000000000000011101011001101011;
assign LUT_3[11486] = 32'b00000000000000011000110101110010;
assign LUT_3[11487] = 32'b00000000000000011111100001001111;
assign LUT_3[11488] = 32'b00000000000000010010000010101111;
assign LUT_3[11489] = 32'b00000000000000011000101110001100;
assign LUT_3[11490] = 32'b00000000000000010100001010010011;
assign LUT_3[11491] = 32'b00000000000000011010110101110000;
assign LUT_3[11492] = 32'b00000000000000001111010000100101;
assign LUT_3[11493] = 32'b00000000000000010101111100000010;
assign LUT_3[11494] = 32'b00000000000000010001011000001001;
assign LUT_3[11495] = 32'b00000000000000011000000011100110;
assign LUT_3[11496] = 32'b00000000000000010111011011110101;
assign LUT_3[11497] = 32'b00000000000000011110000111010010;
assign LUT_3[11498] = 32'b00000000000000011001100011011001;
assign LUT_3[11499] = 32'b00000000000000100000001110110110;
assign LUT_3[11500] = 32'b00000000000000010100101001101011;
assign LUT_3[11501] = 32'b00000000000000011011010101001000;
assign LUT_3[11502] = 32'b00000000000000010110110001001111;
assign LUT_3[11503] = 32'b00000000000000011101011100101100;
assign LUT_3[11504] = 32'b00000000000000010101010101110010;
assign LUT_3[11505] = 32'b00000000000000011100000001001111;
assign LUT_3[11506] = 32'b00000000000000010111011101010110;
assign LUT_3[11507] = 32'b00000000000000011110001000110011;
assign LUT_3[11508] = 32'b00000000000000010010100011101000;
assign LUT_3[11509] = 32'b00000000000000011001001111000101;
assign LUT_3[11510] = 32'b00000000000000010100101011001100;
assign LUT_3[11511] = 32'b00000000000000011011010110101001;
assign LUT_3[11512] = 32'b00000000000000011010101110111000;
assign LUT_3[11513] = 32'b00000000000000100001011010010101;
assign LUT_3[11514] = 32'b00000000000000011100110110011100;
assign LUT_3[11515] = 32'b00000000000000100011100001111001;
assign LUT_3[11516] = 32'b00000000000000010111111100101110;
assign LUT_3[11517] = 32'b00000000000000011110101000001011;
assign LUT_3[11518] = 32'b00000000000000011010000100010010;
assign LUT_3[11519] = 32'b00000000000000100000101111101111;
assign LUT_3[11520] = 32'b00000000000000001011000000000111;
assign LUT_3[11521] = 32'b00000000000000010001101011100100;
assign LUT_3[11522] = 32'b00000000000000001101000111101011;
assign LUT_3[11523] = 32'b00000000000000010011110011001000;
assign LUT_3[11524] = 32'b00000000000000001000001101111101;
assign LUT_3[11525] = 32'b00000000000000001110111001011010;
assign LUT_3[11526] = 32'b00000000000000001010010101100001;
assign LUT_3[11527] = 32'b00000000000000010001000000111110;
assign LUT_3[11528] = 32'b00000000000000010000011001001101;
assign LUT_3[11529] = 32'b00000000000000010111000100101010;
assign LUT_3[11530] = 32'b00000000000000010010100000110001;
assign LUT_3[11531] = 32'b00000000000000011001001100001110;
assign LUT_3[11532] = 32'b00000000000000001101100111000011;
assign LUT_3[11533] = 32'b00000000000000010100010010100000;
assign LUT_3[11534] = 32'b00000000000000001111101110100111;
assign LUT_3[11535] = 32'b00000000000000010110011010000100;
assign LUT_3[11536] = 32'b00000000000000001110010011001010;
assign LUT_3[11537] = 32'b00000000000000010100111110100111;
assign LUT_3[11538] = 32'b00000000000000010000011010101110;
assign LUT_3[11539] = 32'b00000000000000010111000110001011;
assign LUT_3[11540] = 32'b00000000000000001011100001000000;
assign LUT_3[11541] = 32'b00000000000000010010001100011101;
assign LUT_3[11542] = 32'b00000000000000001101101000100100;
assign LUT_3[11543] = 32'b00000000000000010100010100000001;
assign LUT_3[11544] = 32'b00000000000000010011101100010000;
assign LUT_3[11545] = 32'b00000000000000011010010111101101;
assign LUT_3[11546] = 32'b00000000000000010101110011110100;
assign LUT_3[11547] = 32'b00000000000000011100011111010001;
assign LUT_3[11548] = 32'b00000000000000010000111010000110;
assign LUT_3[11549] = 32'b00000000000000010111100101100011;
assign LUT_3[11550] = 32'b00000000000000010011000001101010;
assign LUT_3[11551] = 32'b00000000000000011001101101000111;
assign LUT_3[11552] = 32'b00000000000000001100001110100111;
assign LUT_3[11553] = 32'b00000000000000010010111010000100;
assign LUT_3[11554] = 32'b00000000000000001110010110001011;
assign LUT_3[11555] = 32'b00000000000000010101000001101000;
assign LUT_3[11556] = 32'b00000000000000001001011100011101;
assign LUT_3[11557] = 32'b00000000000000010000000111111010;
assign LUT_3[11558] = 32'b00000000000000001011100100000001;
assign LUT_3[11559] = 32'b00000000000000010010001111011110;
assign LUT_3[11560] = 32'b00000000000000010001100111101101;
assign LUT_3[11561] = 32'b00000000000000011000010011001010;
assign LUT_3[11562] = 32'b00000000000000010011101111010001;
assign LUT_3[11563] = 32'b00000000000000011010011010101110;
assign LUT_3[11564] = 32'b00000000000000001110110101100011;
assign LUT_3[11565] = 32'b00000000000000010101100001000000;
assign LUT_3[11566] = 32'b00000000000000010000111101000111;
assign LUT_3[11567] = 32'b00000000000000010111101000100100;
assign LUT_3[11568] = 32'b00000000000000001111100001101010;
assign LUT_3[11569] = 32'b00000000000000010110001101000111;
assign LUT_3[11570] = 32'b00000000000000010001101001001110;
assign LUT_3[11571] = 32'b00000000000000011000010100101011;
assign LUT_3[11572] = 32'b00000000000000001100101111100000;
assign LUT_3[11573] = 32'b00000000000000010011011010111101;
assign LUT_3[11574] = 32'b00000000000000001110110111000100;
assign LUT_3[11575] = 32'b00000000000000010101100010100001;
assign LUT_3[11576] = 32'b00000000000000010100111010110000;
assign LUT_3[11577] = 32'b00000000000000011011100110001101;
assign LUT_3[11578] = 32'b00000000000000010111000010010100;
assign LUT_3[11579] = 32'b00000000000000011101101101110001;
assign LUT_3[11580] = 32'b00000000000000010010001000100110;
assign LUT_3[11581] = 32'b00000000000000011000110100000011;
assign LUT_3[11582] = 32'b00000000000000010100010000001010;
assign LUT_3[11583] = 32'b00000000000000011010111011100111;
assign LUT_3[11584] = 32'b00000000000000001010111000110010;
assign LUT_3[11585] = 32'b00000000000000010001100100001111;
assign LUT_3[11586] = 32'b00000000000000001101000000010110;
assign LUT_3[11587] = 32'b00000000000000010011101011110011;
assign LUT_3[11588] = 32'b00000000000000001000000110101000;
assign LUT_3[11589] = 32'b00000000000000001110110010000101;
assign LUT_3[11590] = 32'b00000000000000001010001110001100;
assign LUT_3[11591] = 32'b00000000000000010000111001101001;
assign LUT_3[11592] = 32'b00000000000000010000010001111000;
assign LUT_3[11593] = 32'b00000000000000010110111101010101;
assign LUT_3[11594] = 32'b00000000000000010010011001011100;
assign LUT_3[11595] = 32'b00000000000000011001000100111001;
assign LUT_3[11596] = 32'b00000000000000001101011111101110;
assign LUT_3[11597] = 32'b00000000000000010100001011001011;
assign LUT_3[11598] = 32'b00000000000000001111100111010010;
assign LUT_3[11599] = 32'b00000000000000010110010010101111;
assign LUT_3[11600] = 32'b00000000000000001110001011110101;
assign LUT_3[11601] = 32'b00000000000000010100110111010010;
assign LUT_3[11602] = 32'b00000000000000010000010011011001;
assign LUT_3[11603] = 32'b00000000000000010110111110110110;
assign LUT_3[11604] = 32'b00000000000000001011011001101011;
assign LUT_3[11605] = 32'b00000000000000010010000101001000;
assign LUT_3[11606] = 32'b00000000000000001101100001001111;
assign LUT_3[11607] = 32'b00000000000000010100001100101100;
assign LUT_3[11608] = 32'b00000000000000010011100100111011;
assign LUT_3[11609] = 32'b00000000000000011010010000011000;
assign LUT_3[11610] = 32'b00000000000000010101101100011111;
assign LUT_3[11611] = 32'b00000000000000011100010111111100;
assign LUT_3[11612] = 32'b00000000000000010000110010110001;
assign LUT_3[11613] = 32'b00000000000000010111011110001110;
assign LUT_3[11614] = 32'b00000000000000010010111010010101;
assign LUT_3[11615] = 32'b00000000000000011001100101110010;
assign LUT_3[11616] = 32'b00000000000000001100000111010010;
assign LUT_3[11617] = 32'b00000000000000010010110010101111;
assign LUT_3[11618] = 32'b00000000000000001110001110110110;
assign LUT_3[11619] = 32'b00000000000000010100111010010011;
assign LUT_3[11620] = 32'b00000000000000001001010101001000;
assign LUT_3[11621] = 32'b00000000000000010000000000100101;
assign LUT_3[11622] = 32'b00000000000000001011011100101100;
assign LUT_3[11623] = 32'b00000000000000010010001000001001;
assign LUT_3[11624] = 32'b00000000000000010001100000011000;
assign LUT_3[11625] = 32'b00000000000000011000001011110101;
assign LUT_3[11626] = 32'b00000000000000010011100111111100;
assign LUT_3[11627] = 32'b00000000000000011010010011011001;
assign LUT_3[11628] = 32'b00000000000000001110101110001110;
assign LUT_3[11629] = 32'b00000000000000010101011001101011;
assign LUT_3[11630] = 32'b00000000000000010000110101110010;
assign LUT_3[11631] = 32'b00000000000000010111100001001111;
assign LUT_3[11632] = 32'b00000000000000001111011010010101;
assign LUT_3[11633] = 32'b00000000000000010110000101110010;
assign LUT_3[11634] = 32'b00000000000000010001100001111001;
assign LUT_3[11635] = 32'b00000000000000011000001101010110;
assign LUT_3[11636] = 32'b00000000000000001100101000001011;
assign LUT_3[11637] = 32'b00000000000000010011010011101000;
assign LUT_3[11638] = 32'b00000000000000001110101111101111;
assign LUT_3[11639] = 32'b00000000000000010101011011001100;
assign LUT_3[11640] = 32'b00000000000000010100110011011011;
assign LUT_3[11641] = 32'b00000000000000011011011110111000;
assign LUT_3[11642] = 32'b00000000000000010110111010111111;
assign LUT_3[11643] = 32'b00000000000000011101100110011100;
assign LUT_3[11644] = 32'b00000000000000010010000001010001;
assign LUT_3[11645] = 32'b00000000000000011000101100101110;
assign LUT_3[11646] = 32'b00000000000000010100001000110101;
assign LUT_3[11647] = 32'b00000000000000011010110100010010;
assign LUT_3[11648] = 32'b00000000000000001101001011000101;
assign LUT_3[11649] = 32'b00000000000000010011110110100010;
assign LUT_3[11650] = 32'b00000000000000001111010010101001;
assign LUT_3[11651] = 32'b00000000000000010101111110000110;
assign LUT_3[11652] = 32'b00000000000000001010011000111011;
assign LUT_3[11653] = 32'b00000000000000010001000100011000;
assign LUT_3[11654] = 32'b00000000000000001100100000011111;
assign LUT_3[11655] = 32'b00000000000000010011001011111100;
assign LUT_3[11656] = 32'b00000000000000010010100100001011;
assign LUT_3[11657] = 32'b00000000000000011001001111101000;
assign LUT_3[11658] = 32'b00000000000000010100101011101111;
assign LUT_3[11659] = 32'b00000000000000011011010111001100;
assign LUT_3[11660] = 32'b00000000000000001111110010000001;
assign LUT_3[11661] = 32'b00000000000000010110011101011110;
assign LUT_3[11662] = 32'b00000000000000010001111001100101;
assign LUT_3[11663] = 32'b00000000000000011000100101000010;
assign LUT_3[11664] = 32'b00000000000000010000011110001000;
assign LUT_3[11665] = 32'b00000000000000010111001001100101;
assign LUT_3[11666] = 32'b00000000000000010010100101101100;
assign LUT_3[11667] = 32'b00000000000000011001010001001001;
assign LUT_3[11668] = 32'b00000000000000001101101011111110;
assign LUT_3[11669] = 32'b00000000000000010100010111011011;
assign LUT_3[11670] = 32'b00000000000000001111110011100010;
assign LUT_3[11671] = 32'b00000000000000010110011110111111;
assign LUT_3[11672] = 32'b00000000000000010101110111001110;
assign LUT_3[11673] = 32'b00000000000000011100100010101011;
assign LUT_3[11674] = 32'b00000000000000010111111110110010;
assign LUT_3[11675] = 32'b00000000000000011110101010001111;
assign LUT_3[11676] = 32'b00000000000000010011000101000100;
assign LUT_3[11677] = 32'b00000000000000011001110000100001;
assign LUT_3[11678] = 32'b00000000000000010101001100101000;
assign LUT_3[11679] = 32'b00000000000000011011111000000101;
assign LUT_3[11680] = 32'b00000000000000001110011001100101;
assign LUT_3[11681] = 32'b00000000000000010101000101000010;
assign LUT_3[11682] = 32'b00000000000000010000100001001001;
assign LUT_3[11683] = 32'b00000000000000010111001100100110;
assign LUT_3[11684] = 32'b00000000000000001011100111011011;
assign LUT_3[11685] = 32'b00000000000000010010010010111000;
assign LUT_3[11686] = 32'b00000000000000001101101110111111;
assign LUT_3[11687] = 32'b00000000000000010100011010011100;
assign LUT_3[11688] = 32'b00000000000000010011110010101011;
assign LUT_3[11689] = 32'b00000000000000011010011110001000;
assign LUT_3[11690] = 32'b00000000000000010101111010001111;
assign LUT_3[11691] = 32'b00000000000000011100100101101100;
assign LUT_3[11692] = 32'b00000000000000010001000000100001;
assign LUT_3[11693] = 32'b00000000000000010111101011111110;
assign LUT_3[11694] = 32'b00000000000000010011001000000101;
assign LUT_3[11695] = 32'b00000000000000011001110011100010;
assign LUT_3[11696] = 32'b00000000000000010001101100101000;
assign LUT_3[11697] = 32'b00000000000000011000011000000101;
assign LUT_3[11698] = 32'b00000000000000010011110100001100;
assign LUT_3[11699] = 32'b00000000000000011010011111101001;
assign LUT_3[11700] = 32'b00000000000000001110111010011110;
assign LUT_3[11701] = 32'b00000000000000010101100101111011;
assign LUT_3[11702] = 32'b00000000000000010001000010000010;
assign LUT_3[11703] = 32'b00000000000000010111101101011111;
assign LUT_3[11704] = 32'b00000000000000010111000101101110;
assign LUT_3[11705] = 32'b00000000000000011101110001001011;
assign LUT_3[11706] = 32'b00000000000000011001001101010010;
assign LUT_3[11707] = 32'b00000000000000011111111000101111;
assign LUT_3[11708] = 32'b00000000000000010100010011100100;
assign LUT_3[11709] = 32'b00000000000000011010111111000001;
assign LUT_3[11710] = 32'b00000000000000010110011011001000;
assign LUT_3[11711] = 32'b00000000000000011101000110100101;
assign LUT_3[11712] = 32'b00000000000000001101000011110000;
assign LUT_3[11713] = 32'b00000000000000010011101111001101;
assign LUT_3[11714] = 32'b00000000000000001111001011010100;
assign LUT_3[11715] = 32'b00000000000000010101110110110001;
assign LUT_3[11716] = 32'b00000000000000001010010001100110;
assign LUT_3[11717] = 32'b00000000000000010000111101000011;
assign LUT_3[11718] = 32'b00000000000000001100011001001010;
assign LUT_3[11719] = 32'b00000000000000010011000100100111;
assign LUT_3[11720] = 32'b00000000000000010010011100110110;
assign LUT_3[11721] = 32'b00000000000000011001001000010011;
assign LUT_3[11722] = 32'b00000000000000010100100100011010;
assign LUT_3[11723] = 32'b00000000000000011011001111110111;
assign LUT_3[11724] = 32'b00000000000000001111101010101100;
assign LUT_3[11725] = 32'b00000000000000010110010110001001;
assign LUT_3[11726] = 32'b00000000000000010001110010010000;
assign LUT_3[11727] = 32'b00000000000000011000011101101101;
assign LUT_3[11728] = 32'b00000000000000010000010110110011;
assign LUT_3[11729] = 32'b00000000000000010111000010010000;
assign LUT_3[11730] = 32'b00000000000000010010011110010111;
assign LUT_3[11731] = 32'b00000000000000011001001001110100;
assign LUT_3[11732] = 32'b00000000000000001101100100101001;
assign LUT_3[11733] = 32'b00000000000000010100010000000110;
assign LUT_3[11734] = 32'b00000000000000001111101100001101;
assign LUT_3[11735] = 32'b00000000000000010110010111101010;
assign LUT_3[11736] = 32'b00000000000000010101101111111001;
assign LUT_3[11737] = 32'b00000000000000011100011011010110;
assign LUT_3[11738] = 32'b00000000000000010111110111011101;
assign LUT_3[11739] = 32'b00000000000000011110100010111010;
assign LUT_3[11740] = 32'b00000000000000010010111101101111;
assign LUT_3[11741] = 32'b00000000000000011001101001001100;
assign LUT_3[11742] = 32'b00000000000000010101000101010011;
assign LUT_3[11743] = 32'b00000000000000011011110000110000;
assign LUT_3[11744] = 32'b00000000000000001110010010010000;
assign LUT_3[11745] = 32'b00000000000000010100111101101101;
assign LUT_3[11746] = 32'b00000000000000010000011001110100;
assign LUT_3[11747] = 32'b00000000000000010111000101010001;
assign LUT_3[11748] = 32'b00000000000000001011100000000110;
assign LUT_3[11749] = 32'b00000000000000010010001011100011;
assign LUT_3[11750] = 32'b00000000000000001101100111101010;
assign LUT_3[11751] = 32'b00000000000000010100010011000111;
assign LUT_3[11752] = 32'b00000000000000010011101011010110;
assign LUT_3[11753] = 32'b00000000000000011010010110110011;
assign LUT_3[11754] = 32'b00000000000000010101110010111010;
assign LUT_3[11755] = 32'b00000000000000011100011110010111;
assign LUT_3[11756] = 32'b00000000000000010000111001001100;
assign LUT_3[11757] = 32'b00000000000000010111100100101001;
assign LUT_3[11758] = 32'b00000000000000010011000000110000;
assign LUT_3[11759] = 32'b00000000000000011001101100001101;
assign LUT_3[11760] = 32'b00000000000000010001100101010011;
assign LUT_3[11761] = 32'b00000000000000011000010000110000;
assign LUT_3[11762] = 32'b00000000000000010011101100110111;
assign LUT_3[11763] = 32'b00000000000000011010011000010100;
assign LUT_3[11764] = 32'b00000000000000001110110011001001;
assign LUT_3[11765] = 32'b00000000000000010101011110100110;
assign LUT_3[11766] = 32'b00000000000000010000111010101101;
assign LUT_3[11767] = 32'b00000000000000010111100110001010;
assign LUT_3[11768] = 32'b00000000000000010110111110011001;
assign LUT_3[11769] = 32'b00000000000000011101101001110110;
assign LUT_3[11770] = 32'b00000000000000011001000101111101;
assign LUT_3[11771] = 32'b00000000000000011111110001011010;
assign LUT_3[11772] = 32'b00000000000000010100001100001111;
assign LUT_3[11773] = 32'b00000000000000011010110111101100;
assign LUT_3[11774] = 32'b00000000000000010110010011110011;
assign LUT_3[11775] = 32'b00000000000000011100111111010000;
assign LUT_3[11776] = 32'b00000000000000010010000101110010;
assign LUT_3[11777] = 32'b00000000000000011000110001001111;
assign LUT_3[11778] = 32'b00000000000000010100001101010110;
assign LUT_3[11779] = 32'b00000000000000011010111000110011;
assign LUT_3[11780] = 32'b00000000000000001111010011101000;
assign LUT_3[11781] = 32'b00000000000000010101111111000101;
assign LUT_3[11782] = 32'b00000000000000010001011011001100;
assign LUT_3[11783] = 32'b00000000000000011000000110101001;
assign LUT_3[11784] = 32'b00000000000000010111011110111000;
assign LUT_3[11785] = 32'b00000000000000011110001010010101;
assign LUT_3[11786] = 32'b00000000000000011001100110011100;
assign LUT_3[11787] = 32'b00000000000000100000010001111001;
assign LUT_3[11788] = 32'b00000000000000010100101100101110;
assign LUT_3[11789] = 32'b00000000000000011011011000001011;
assign LUT_3[11790] = 32'b00000000000000010110110100010010;
assign LUT_3[11791] = 32'b00000000000000011101011111101111;
assign LUT_3[11792] = 32'b00000000000000010101011000110101;
assign LUT_3[11793] = 32'b00000000000000011100000100010010;
assign LUT_3[11794] = 32'b00000000000000010111100000011001;
assign LUT_3[11795] = 32'b00000000000000011110001011110110;
assign LUT_3[11796] = 32'b00000000000000010010100110101011;
assign LUT_3[11797] = 32'b00000000000000011001010010001000;
assign LUT_3[11798] = 32'b00000000000000010100101110001111;
assign LUT_3[11799] = 32'b00000000000000011011011001101100;
assign LUT_3[11800] = 32'b00000000000000011010110001111011;
assign LUT_3[11801] = 32'b00000000000000100001011101011000;
assign LUT_3[11802] = 32'b00000000000000011100111001011111;
assign LUT_3[11803] = 32'b00000000000000100011100100111100;
assign LUT_3[11804] = 32'b00000000000000010111111111110001;
assign LUT_3[11805] = 32'b00000000000000011110101011001110;
assign LUT_3[11806] = 32'b00000000000000011010000111010101;
assign LUT_3[11807] = 32'b00000000000000100000110010110010;
assign LUT_3[11808] = 32'b00000000000000010011010100010010;
assign LUT_3[11809] = 32'b00000000000000011001111111101111;
assign LUT_3[11810] = 32'b00000000000000010101011011110110;
assign LUT_3[11811] = 32'b00000000000000011100000111010011;
assign LUT_3[11812] = 32'b00000000000000010000100010001000;
assign LUT_3[11813] = 32'b00000000000000010111001101100101;
assign LUT_3[11814] = 32'b00000000000000010010101001101100;
assign LUT_3[11815] = 32'b00000000000000011001010101001001;
assign LUT_3[11816] = 32'b00000000000000011000101101011000;
assign LUT_3[11817] = 32'b00000000000000011111011000110101;
assign LUT_3[11818] = 32'b00000000000000011010110100111100;
assign LUT_3[11819] = 32'b00000000000000100001100000011001;
assign LUT_3[11820] = 32'b00000000000000010101111011001110;
assign LUT_3[11821] = 32'b00000000000000011100100110101011;
assign LUT_3[11822] = 32'b00000000000000011000000010110010;
assign LUT_3[11823] = 32'b00000000000000011110101110001111;
assign LUT_3[11824] = 32'b00000000000000010110100111010101;
assign LUT_3[11825] = 32'b00000000000000011101010010110010;
assign LUT_3[11826] = 32'b00000000000000011000101110111001;
assign LUT_3[11827] = 32'b00000000000000011111011010010110;
assign LUT_3[11828] = 32'b00000000000000010011110101001011;
assign LUT_3[11829] = 32'b00000000000000011010100000101000;
assign LUT_3[11830] = 32'b00000000000000010101111100101111;
assign LUT_3[11831] = 32'b00000000000000011100101000001100;
assign LUT_3[11832] = 32'b00000000000000011100000000011011;
assign LUT_3[11833] = 32'b00000000000000100010101011111000;
assign LUT_3[11834] = 32'b00000000000000011110000111111111;
assign LUT_3[11835] = 32'b00000000000000100100110011011100;
assign LUT_3[11836] = 32'b00000000000000011001001110010001;
assign LUT_3[11837] = 32'b00000000000000011111111001101110;
assign LUT_3[11838] = 32'b00000000000000011011010101110101;
assign LUT_3[11839] = 32'b00000000000000100010000001010010;
assign LUT_3[11840] = 32'b00000000000000010001111110011101;
assign LUT_3[11841] = 32'b00000000000000011000101001111010;
assign LUT_3[11842] = 32'b00000000000000010100000110000001;
assign LUT_3[11843] = 32'b00000000000000011010110001011110;
assign LUT_3[11844] = 32'b00000000000000001111001100010011;
assign LUT_3[11845] = 32'b00000000000000010101110111110000;
assign LUT_3[11846] = 32'b00000000000000010001010011110111;
assign LUT_3[11847] = 32'b00000000000000010111111111010100;
assign LUT_3[11848] = 32'b00000000000000010111010111100011;
assign LUT_3[11849] = 32'b00000000000000011110000011000000;
assign LUT_3[11850] = 32'b00000000000000011001011111000111;
assign LUT_3[11851] = 32'b00000000000000100000001010100100;
assign LUT_3[11852] = 32'b00000000000000010100100101011001;
assign LUT_3[11853] = 32'b00000000000000011011010000110110;
assign LUT_3[11854] = 32'b00000000000000010110101100111101;
assign LUT_3[11855] = 32'b00000000000000011101011000011010;
assign LUT_3[11856] = 32'b00000000000000010101010001100000;
assign LUT_3[11857] = 32'b00000000000000011011111100111101;
assign LUT_3[11858] = 32'b00000000000000010111011001000100;
assign LUT_3[11859] = 32'b00000000000000011110000100100001;
assign LUT_3[11860] = 32'b00000000000000010010011111010110;
assign LUT_3[11861] = 32'b00000000000000011001001010110011;
assign LUT_3[11862] = 32'b00000000000000010100100110111010;
assign LUT_3[11863] = 32'b00000000000000011011010010010111;
assign LUT_3[11864] = 32'b00000000000000011010101010100110;
assign LUT_3[11865] = 32'b00000000000000100001010110000011;
assign LUT_3[11866] = 32'b00000000000000011100110010001010;
assign LUT_3[11867] = 32'b00000000000000100011011101100111;
assign LUT_3[11868] = 32'b00000000000000010111111000011100;
assign LUT_3[11869] = 32'b00000000000000011110100011111001;
assign LUT_3[11870] = 32'b00000000000000011010000000000000;
assign LUT_3[11871] = 32'b00000000000000100000101011011101;
assign LUT_3[11872] = 32'b00000000000000010011001100111101;
assign LUT_3[11873] = 32'b00000000000000011001111000011010;
assign LUT_3[11874] = 32'b00000000000000010101010100100001;
assign LUT_3[11875] = 32'b00000000000000011011111111111110;
assign LUT_3[11876] = 32'b00000000000000010000011010110011;
assign LUT_3[11877] = 32'b00000000000000010111000110010000;
assign LUT_3[11878] = 32'b00000000000000010010100010010111;
assign LUT_3[11879] = 32'b00000000000000011001001101110100;
assign LUT_3[11880] = 32'b00000000000000011000100110000011;
assign LUT_3[11881] = 32'b00000000000000011111010001100000;
assign LUT_3[11882] = 32'b00000000000000011010101101100111;
assign LUT_3[11883] = 32'b00000000000000100001011001000100;
assign LUT_3[11884] = 32'b00000000000000010101110011111001;
assign LUT_3[11885] = 32'b00000000000000011100011111010110;
assign LUT_3[11886] = 32'b00000000000000010111111011011101;
assign LUT_3[11887] = 32'b00000000000000011110100110111010;
assign LUT_3[11888] = 32'b00000000000000010110100000000000;
assign LUT_3[11889] = 32'b00000000000000011101001011011101;
assign LUT_3[11890] = 32'b00000000000000011000100111100100;
assign LUT_3[11891] = 32'b00000000000000011111010011000001;
assign LUT_3[11892] = 32'b00000000000000010011101101110110;
assign LUT_3[11893] = 32'b00000000000000011010011001010011;
assign LUT_3[11894] = 32'b00000000000000010101110101011010;
assign LUT_3[11895] = 32'b00000000000000011100100000110111;
assign LUT_3[11896] = 32'b00000000000000011011111001000110;
assign LUT_3[11897] = 32'b00000000000000100010100100100011;
assign LUT_3[11898] = 32'b00000000000000011110000000101010;
assign LUT_3[11899] = 32'b00000000000000100100101100000111;
assign LUT_3[11900] = 32'b00000000000000011001000110111100;
assign LUT_3[11901] = 32'b00000000000000011111110010011001;
assign LUT_3[11902] = 32'b00000000000000011011001110100000;
assign LUT_3[11903] = 32'b00000000000000100001111001111101;
assign LUT_3[11904] = 32'b00000000000000010100010000110000;
assign LUT_3[11905] = 32'b00000000000000011010111100001101;
assign LUT_3[11906] = 32'b00000000000000010110011000010100;
assign LUT_3[11907] = 32'b00000000000000011101000011110001;
assign LUT_3[11908] = 32'b00000000000000010001011110100110;
assign LUT_3[11909] = 32'b00000000000000011000001010000011;
assign LUT_3[11910] = 32'b00000000000000010011100110001010;
assign LUT_3[11911] = 32'b00000000000000011010010001100111;
assign LUT_3[11912] = 32'b00000000000000011001101001110110;
assign LUT_3[11913] = 32'b00000000000000100000010101010011;
assign LUT_3[11914] = 32'b00000000000000011011110001011010;
assign LUT_3[11915] = 32'b00000000000000100010011100110111;
assign LUT_3[11916] = 32'b00000000000000010110110111101100;
assign LUT_3[11917] = 32'b00000000000000011101100011001001;
assign LUT_3[11918] = 32'b00000000000000011000111111010000;
assign LUT_3[11919] = 32'b00000000000000011111101010101101;
assign LUT_3[11920] = 32'b00000000000000010111100011110011;
assign LUT_3[11921] = 32'b00000000000000011110001111010000;
assign LUT_3[11922] = 32'b00000000000000011001101011010111;
assign LUT_3[11923] = 32'b00000000000000100000010110110100;
assign LUT_3[11924] = 32'b00000000000000010100110001101001;
assign LUT_3[11925] = 32'b00000000000000011011011101000110;
assign LUT_3[11926] = 32'b00000000000000010110111001001101;
assign LUT_3[11927] = 32'b00000000000000011101100100101010;
assign LUT_3[11928] = 32'b00000000000000011100111100111001;
assign LUT_3[11929] = 32'b00000000000000100011101000010110;
assign LUT_3[11930] = 32'b00000000000000011111000100011101;
assign LUT_3[11931] = 32'b00000000000000100101101111111010;
assign LUT_3[11932] = 32'b00000000000000011010001010101111;
assign LUT_3[11933] = 32'b00000000000000100000110110001100;
assign LUT_3[11934] = 32'b00000000000000011100010010010011;
assign LUT_3[11935] = 32'b00000000000000100010111101110000;
assign LUT_3[11936] = 32'b00000000000000010101011111010000;
assign LUT_3[11937] = 32'b00000000000000011100001010101101;
assign LUT_3[11938] = 32'b00000000000000010111100110110100;
assign LUT_3[11939] = 32'b00000000000000011110010010010001;
assign LUT_3[11940] = 32'b00000000000000010010101101000110;
assign LUT_3[11941] = 32'b00000000000000011001011000100011;
assign LUT_3[11942] = 32'b00000000000000010100110100101010;
assign LUT_3[11943] = 32'b00000000000000011011100000000111;
assign LUT_3[11944] = 32'b00000000000000011010111000010110;
assign LUT_3[11945] = 32'b00000000000000100001100011110011;
assign LUT_3[11946] = 32'b00000000000000011100111111111010;
assign LUT_3[11947] = 32'b00000000000000100011101011010111;
assign LUT_3[11948] = 32'b00000000000000011000000110001100;
assign LUT_3[11949] = 32'b00000000000000011110110001101001;
assign LUT_3[11950] = 32'b00000000000000011010001101110000;
assign LUT_3[11951] = 32'b00000000000000100000111001001101;
assign LUT_3[11952] = 32'b00000000000000011000110010010011;
assign LUT_3[11953] = 32'b00000000000000011111011101110000;
assign LUT_3[11954] = 32'b00000000000000011010111001110111;
assign LUT_3[11955] = 32'b00000000000000100001100101010100;
assign LUT_3[11956] = 32'b00000000000000010110000000001001;
assign LUT_3[11957] = 32'b00000000000000011100101011100110;
assign LUT_3[11958] = 32'b00000000000000011000000111101101;
assign LUT_3[11959] = 32'b00000000000000011110110011001010;
assign LUT_3[11960] = 32'b00000000000000011110001011011001;
assign LUT_3[11961] = 32'b00000000000000100100110110110110;
assign LUT_3[11962] = 32'b00000000000000100000010010111101;
assign LUT_3[11963] = 32'b00000000000000100110111110011010;
assign LUT_3[11964] = 32'b00000000000000011011011001001111;
assign LUT_3[11965] = 32'b00000000000000100010000100101100;
assign LUT_3[11966] = 32'b00000000000000011101100000110011;
assign LUT_3[11967] = 32'b00000000000000100100001100010000;
assign LUT_3[11968] = 32'b00000000000000010100001001011011;
assign LUT_3[11969] = 32'b00000000000000011010110100111000;
assign LUT_3[11970] = 32'b00000000000000010110010000111111;
assign LUT_3[11971] = 32'b00000000000000011100111100011100;
assign LUT_3[11972] = 32'b00000000000000010001010111010001;
assign LUT_3[11973] = 32'b00000000000000011000000010101110;
assign LUT_3[11974] = 32'b00000000000000010011011110110101;
assign LUT_3[11975] = 32'b00000000000000011010001010010010;
assign LUT_3[11976] = 32'b00000000000000011001100010100001;
assign LUT_3[11977] = 32'b00000000000000100000001101111110;
assign LUT_3[11978] = 32'b00000000000000011011101010000101;
assign LUT_3[11979] = 32'b00000000000000100010010101100010;
assign LUT_3[11980] = 32'b00000000000000010110110000010111;
assign LUT_3[11981] = 32'b00000000000000011101011011110100;
assign LUT_3[11982] = 32'b00000000000000011000110111111011;
assign LUT_3[11983] = 32'b00000000000000011111100011011000;
assign LUT_3[11984] = 32'b00000000000000010111011100011110;
assign LUT_3[11985] = 32'b00000000000000011110000111111011;
assign LUT_3[11986] = 32'b00000000000000011001100100000010;
assign LUT_3[11987] = 32'b00000000000000100000001111011111;
assign LUT_3[11988] = 32'b00000000000000010100101010010100;
assign LUT_3[11989] = 32'b00000000000000011011010101110001;
assign LUT_3[11990] = 32'b00000000000000010110110001111000;
assign LUT_3[11991] = 32'b00000000000000011101011101010101;
assign LUT_3[11992] = 32'b00000000000000011100110101100100;
assign LUT_3[11993] = 32'b00000000000000100011100001000001;
assign LUT_3[11994] = 32'b00000000000000011110111101001000;
assign LUT_3[11995] = 32'b00000000000000100101101000100101;
assign LUT_3[11996] = 32'b00000000000000011010000011011010;
assign LUT_3[11997] = 32'b00000000000000100000101110110111;
assign LUT_3[11998] = 32'b00000000000000011100001010111110;
assign LUT_3[11999] = 32'b00000000000000100010110110011011;
assign LUT_3[12000] = 32'b00000000000000010101010111111011;
assign LUT_3[12001] = 32'b00000000000000011100000011011000;
assign LUT_3[12002] = 32'b00000000000000010111011111011111;
assign LUT_3[12003] = 32'b00000000000000011110001010111100;
assign LUT_3[12004] = 32'b00000000000000010010100101110001;
assign LUT_3[12005] = 32'b00000000000000011001010001001110;
assign LUT_3[12006] = 32'b00000000000000010100101101010101;
assign LUT_3[12007] = 32'b00000000000000011011011000110010;
assign LUT_3[12008] = 32'b00000000000000011010110001000001;
assign LUT_3[12009] = 32'b00000000000000100001011100011110;
assign LUT_3[12010] = 32'b00000000000000011100111000100101;
assign LUT_3[12011] = 32'b00000000000000100011100100000010;
assign LUT_3[12012] = 32'b00000000000000010111111110110111;
assign LUT_3[12013] = 32'b00000000000000011110101010010100;
assign LUT_3[12014] = 32'b00000000000000011010000110011011;
assign LUT_3[12015] = 32'b00000000000000100000110001111000;
assign LUT_3[12016] = 32'b00000000000000011000101010111110;
assign LUT_3[12017] = 32'b00000000000000011111010110011011;
assign LUT_3[12018] = 32'b00000000000000011010110010100010;
assign LUT_3[12019] = 32'b00000000000000100001011101111111;
assign LUT_3[12020] = 32'b00000000000000010101111000110100;
assign LUT_3[12021] = 32'b00000000000000011100100100010001;
assign LUT_3[12022] = 32'b00000000000000011000000000011000;
assign LUT_3[12023] = 32'b00000000000000011110101011110101;
assign LUT_3[12024] = 32'b00000000000000011110000100000100;
assign LUT_3[12025] = 32'b00000000000000100100101111100001;
assign LUT_3[12026] = 32'b00000000000000100000001011101000;
assign LUT_3[12027] = 32'b00000000000000100110110111000101;
assign LUT_3[12028] = 32'b00000000000000011011010001111010;
assign LUT_3[12029] = 32'b00000000000000100001111101010111;
assign LUT_3[12030] = 32'b00000000000000011101011001011110;
assign LUT_3[12031] = 32'b00000000000000100100000100111011;
assign LUT_3[12032] = 32'b00000000000000001110010101010011;
assign LUT_3[12033] = 32'b00000000000000010101000000110000;
assign LUT_3[12034] = 32'b00000000000000010000011100110111;
assign LUT_3[12035] = 32'b00000000000000010111001000010100;
assign LUT_3[12036] = 32'b00000000000000001011100011001001;
assign LUT_3[12037] = 32'b00000000000000010010001110100110;
assign LUT_3[12038] = 32'b00000000000000001101101010101101;
assign LUT_3[12039] = 32'b00000000000000010100010110001010;
assign LUT_3[12040] = 32'b00000000000000010011101110011001;
assign LUT_3[12041] = 32'b00000000000000011010011001110110;
assign LUT_3[12042] = 32'b00000000000000010101110101111101;
assign LUT_3[12043] = 32'b00000000000000011100100001011010;
assign LUT_3[12044] = 32'b00000000000000010000111100001111;
assign LUT_3[12045] = 32'b00000000000000010111100111101100;
assign LUT_3[12046] = 32'b00000000000000010011000011110011;
assign LUT_3[12047] = 32'b00000000000000011001101111010000;
assign LUT_3[12048] = 32'b00000000000000010001101000010110;
assign LUT_3[12049] = 32'b00000000000000011000010011110011;
assign LUT_3[12050] = 32'b00000000000000010011101111111010;
assign LUT_3[12051] = 32'b00000000000000011010011011010111;
assign LUT_3[12052] = 32'b00000000000000001110110110001100;
assign LUT_3[12053] = 32'b00000000000000010101100001101001;
assign LUT_3[12054] = 32'b00000000000000010000111101110000;
assign LUT_3[12055] = 32'b00000000000000010111101001001101;
assign LUT_3[12056] = 32'b00000000000000010111000001011100;
assign LUT_3[12057] = 32'b00000000000000011101101100111001;
assign LUT_3[12058] = 32'b00000000000000011001001001000000;
assign LUT_3[12059] = 32'b00000000000000011111110100011101;
assign LUT_3[12060] = 32'b00000000000000010100001111010010;
assign LUT_3[12061] = 32'b00000000000000011010111010101111;
assign LUT_3[12062] = 32'b00000000000000010110010110110110;
assign LUT_3[12063] = 32'b00000000000000011101000010010011;
assign LUT_3[12064] = 32'b00000000000000001111100011110011;
assign LUT_3[12065] = 32'b00000000000000010110001111010000;
assign LUT_3[12066] = 32'b00000000000000010001101011010111;
assign LUT_3[12067] = 32'b00000000000000011000010110110100;
assign LUT_3[12068] = 32'b00000000000000001100110001101001;
assign LUT_3[12069] = 32'b00000000000000010011011101000110;
assign LUT_3[12070] = 32'b00000000000000001110111001001101;
assign LUT_3[12071] = 32'b00000000000000010101100100101010;
assign LUT_3[12072] = 32'b00000000000000010100111100111001;
assign LUT_3[12073] = 32'b00000000000000011011101000010110;
assign LUT_3[12074] = 32'b00000000000000010111000100011101;
assign LUT_3[12075] = 32'b00000000000000011101101111111010;
assign LUT_3[12076] = 32'b00000000000000010010001010101111;
assign LUT_3[12077] = 32'b00000000000000011000110110001100;
assign LUT_3[12078] = 32'b00000000000000010100010010010011;
assign LUT_3[12079] = 32'b00000000000000011010111101110000;
assign LUT_3[12080] = 32'b00000000000000010010110110110110;
assign LUT_3[12081] = 32'b00000000000000011001100010010011;
assign LUT_3[12082] = 32'b00000000000000010100111110011010;
assign LUT_3[12083] = 32'b00000000000000011011101001110111;
assign LUT_3[12084] = 32'b00000000000000010000000100101100;
assign LUT_3[12085] = 32'b00000000000000010110110000001001;
assign LUT_3[12086] = 32'b00000000000000010010001100010000;
assign LUT_3[12087] = 32'b00000000000000011000110111101101;
assign LUT_3[12088] = 32'b00000000000000011000001111111100;
assign LUT_3[12089] = 32'b00000000000000011110111011011001;
assign LUT_3[12090] = 32'b00000000000000011010010111100000;
assign LUT_3[12091] = 32'b00000000000000100001000010111101;
assign LUT_3[12092] = 32'b00000000000000010101011101110010;
assign LUT_3[12093] = 32'b00000000000000011100001001001111;
assign LUT_3[12094] = 32'b00000000000000010111100101010110;
assign LUT_3[12095] = 32'b00000000000000011110010000110011;
assign LUT_3[12096] = 32'b00000000000000001110001101111110;
assign LUT_3[12097] = 32'b00000000000000010100111001011011;
assign LUT_3[12098] = 32'b00000000000000010000010101100010;
assign LUT_3[12099] = 32'b00000000000000010111000000111111;
assign LUT_3[12100] = 32'b00000000000000001011011011110100;
assign LUT_3[12101] = 32'b00000000000000010010000111010001;
assign LUT_3[12102] = 32'b00000000000000001101100011011000;
assign LUT_3[12103] = 32'b00000000000000010100001110110101;
assign LUT_3[12104] = 32'b00000000000000010011100111000100;
assign LUT_3[12105] = 32'b00000000000000011010010010100001;
assign LUT_3[12106] = 32'b00000000000000010101101110101000;
assign LUT_3[12107] = 32'b00000000000000011100011010000101;
assign LUT_3[12108] = 32'b00000000000000010000110100111010;
assign LUT_3[12109] = 32'b00000000000000010111100000010111;
assign LUT_3[12110] = 32'b00000000000000010010111100011110;
assign LUT_3[12111] = 32'b00000000000000011001100111111011;
assign LUT_3[12112] = 32'b00000000000000010001100001000001;
assign LUT_3[12113] = 32'b00000000000000011000001100011110;
assign LUT_3[12114] = 32'b00000000000000010011101000100101;
assign LUT_3[12115] = 32'b00000000000000011010010100000010;
assign LUT_3[12116] = 32'b00000000000000001110101110110111;
assign LUT_3[12117] = 32'b00000000000000010101011010010100;
assign LUT_3[12118] = 32'b00000000000000010000110110011011;
assign LUT_3[12119] = 32'b00000000000000010111100001111000;
assign LUT_3[12120] = 32'b00000000000000010110111010000111;
assign LUT_3[12121] = 32'b00000000000000011101100101100100;
assign LUT_3[12122] = 32'b00000000000000011001000001101011;
assign LUT_3[12123] = 32'b00000000000000011111101101001000;
assign LUT_3[12124] = 32'b00000000000000010100000111111101;
assign LUT_3[12125] = 32'b00000000000000011010110011011010;
assign LUT_3[12126] = 32'b00000000000000010110001111100001;
assign LUT_3[12127] = 32'b00000000000000011100111010111110;
assign LUT_3[12128] = 32'b00000000000000001111011100011110;
assign LUT_3[12129] = 32'b00000000000000010110000111111011;
assign LUT_3[12130] = 32'b00000000000000010001100100000010;
assign LUT_3[12131] = 32'b00000000000000011000001111011111;
assign LUT_3[12132] = 32'b00000000000000001100101010010100;
assign LUT_3[12133] = 32'b00000000000000010011010101110001;
assign LUT_3[12134] = 32'b00000000000000001110110001111000;
assign LUT_3[12135] = 32'b00000000000000010101011101010101;
assign LUT_3[12136] = 32'b00000000000000010100110101100100;
assign LUT_3[12137] = 32'b00000000000000011011100001000001;
assign LUT_3[12138] = 32'b00000000000000010110111101001000;
assign LUT_3[12139] = 32'b00000000000000011101101000100101;
assign LUT_3[12140] = 32'b00000000000000010010000011011010;
assign LUT_3[12141] = 32'b00000000000000011000101110110111;
assign LUT_3[12142] = 32'b00000000000000010100001010111110;
assign LUT_3[12143] = 32'b00000000000000011010110110011011;
assign LUT_3[12144] = 32'b00000000000000010010101111100001;
assign LUT_3[12145] = 32'b00000000000000011001011010111110;
assign LUT_3[12146] = 32'b00000000000000010100110111000101;
assign LUT_3[12147] = 32'b00000000000000011011100010100010;
assign LUT_3[12148] = 32'b00000000000000001111111101010111;
assign LUT_3[12149] = 32'b00000000000000010110101000110100;
assign LUT_3[12150] = 32'b00000000000000010010000100111011;
assign LUT_3[12151] = 32'b00000000000000011000110000011000;
assign LUT_3[12152] = 32'b00000000000000011000001000100111;
assign LUT_3[12153] = 32'b00000000000000011110110100000100;
assign LUT_3[12154] = 32'b00000000000000011010010000001011;
assign LUT_3[12155] = 32'b00000000000000100000111011101000;
assign LUT_3[12156] = 32'b00000000000000010101010110011101;
assign LUT_3[12157] = 32'b00000000000000011100000001111010;
assign LUT_3[12158] = 32'b00000000000000010111011110000001;
assign LUT_3[12159] = 32'b00000000000000011110001001011110;
assign LUT_3[12160] = 32'b00000000000000010000100000010001;
assign LUT_3[12161] = 32'b00000000000000010111001011101110;
assign LUT_3[12162] = 32'b00000000000000010010100111110101;
assign LUT_3[12163] = 32'b00000000000000011001010011010010;
assign LUT_3[12164] = 32'b00000000000000001101101110000111;
assign LUT_3[12165] = 32'b00000000000000010100011001100100;
assign LUT_3[12166] = 32'b00000000000000001111110101101011;
assign LUT_3[12167] = 32'b00000000000000010110100001001000;
assign LUT_3[12168] = 32'b00000000000000010101111001010111;
assign LUT_3[12169] = 32'b00000000000000011100100100110100;
assign LUT_3[12170] = 32'b00000000000000011000000000111011;
assign LUT_3[12171] = 32'b00000000000000011110101100011000;
assign LUT_3[12172] = 32'b00000000000000010011000111001101;
assign LUT_3[12173] = 32'b00000000000000011001110010101010;
assign LUT_3[12174] = 32'b00000000000000010101001110110001;
assign LUT_3[12175] = 32'b00000000000000011011111010001110;
assign LUT_3[12176] = 32'b00000000000000010011110011010100;
assign LUT_3[12177] = 32'b00000000000000011010011110110001;
assign LUT_3[12178] = 32'b00000000000000010101111010111000;
assign LUT_3[12179] = 32'b00000000000000011100100110010101;
assign LUT_3[12180] = 32'b00000000000000010001000001001010;
assign LUT_3[12181] = 32'b00000000000000010111101100100111;
assign LUT_3[12182] = 32'b00000000000000010011001000101110;
assign LUT_3[12183] = 32'b00000000000000011001110100001011;
assign LUT_3[12184] = 32'b00000000000000011001001100011010;
assign LUT_3[12185] = 32'b00000000000000011111110111110111;
assign LUT_3[12186] = 32'b00000000000000011011010011111110;
assign LUT_3[12187] = 32'b00000000000000100001111111011011;
assign LUT_3[12188] = 32'b00000000000000010110011010010000;
assign LUT_3[12189] = 32'b00000000000000011101000101101101;
assign LUT_3[12190] = 32'b00000000000000011000100001110100;
assign LUT_3[12191] = 32'b00000000000000011111001101010001;
assign LUT_3[12192] = 32'b00000000000000010001101110110001;
assign LUT_3[12193] = 32'b00000000000000011000011010001110;
assign LUT_3[12194] = 32'b00000000000000010011110110010101;
assign LUT_3[12195] = 32'b00000000000000011010100001110010;
assign LUT_3[12196] = 32'b00000000000000001110111100100111;
assign LUT_3[12197] = 32'b00000000000000010101101000000100;
assign LUT_3[12198] = 32'b00000000000000010001000100001011;
assign LUT_3[12199] = 32'b00000000000000010111101111101000;
assign LUT_3[12200] = 32'b00000000000000010111000111110111;
assign LUT_3[12201] = 32'b00000000000000011101110011010100;
assign LUT_3[12202] = 32'b00000000000000011001001111011011;
assign LUT_3[12203] = 32'b00000000000000011111111010111000;
assign LUT_3[12204] = 32'b00000000000000010100010101101101;
assign LUT_3[12205] = 32'b00000000000000011011000001001010;
assign LUT_3[12206] = 32'b00000000000000010110011101010001;
assign LUT_3[12207] = 32'b00000000000000011101001000101110;
assign LUT_3[12208] = 32'b00000000000000010101000001110100;
assign LUT_3[12209] = 32'b00000000000000011011101101010001;
assign LUT_3[12210] = 32'b00000000000000010111001001011000;
assign LUT_3[12211] = 32'b00000000000000011101110100110101;
assign LUT_3[12212] = 32'b00000000000000010010001111101010;
assign LUT_3[12213] = 32'b00000000000000011000111011000111;
assign LUT_3[12214] = 32'b00000000000000010100010111001110;
assign LUT_3[12215] = 32'b00000000000000011011000010101011;
assign LUT_3[12216] = 32'b00000000000000011010011010111010;
assign LUT_3[12217] = 32'b00000000000000100001000110010111;
assign LUT_3[12218] = 32'b00000000000000011100100010011110;
assign LUT_3[12219] = 32'b00000000000000100011001101111011;
assign LUT_3[12220] = 32'b00000000000000010111101000110000;
assign LUT_3[12221] = 32'b00000000000000011110010100001101;
assign LUT_3[12222] = 32'b00000000000000011001110000010100;
assign LUT_3[12223] = 32'b00000000000000100000011011110001;
assign LUT_3[12224] = 32'b00000000000000010000011000111100;
assign LUT_3[12225] = 32'b00000000000000010111000100011001;
assign LUT_3[12226] = 32'b00000000000000010010100000100000;
assign LUT_3[12227] = 32'b00000000000000011001001011111101;
assign LUT_3[12228] = 32'b00000000000000001101100110110010;
assign LUT_3[12229] = 32'b00000000000000010100010010001111;
assign LUT_3[12230] = 32'b00000000000000001111101110010110;
assign LUT_3[12231] = 32'b00000000000000010110011001110011;
assign LUT_3[12232] = 32'b00000000000000010101110010000010;
assign LUT_3[12233] = 32'b00000000000000011100011101011111;
assign LUT_3[12234] = 32'b00000000000000010111111001100110;
assign LUT_3[12235] = 32'b00000000000000011110100101000011;
assign LUT_3[12236] = 32'b00000000000000010010111111111000;
assign LUT_3[12237] = 32'b00000000000000011001101011010101;
assign LUT_3[12238] = 32'b00000000000000010101000111011100;
assign LUT_3[12239] = 32'b00000000000000011011110010111001;
assign LUT_3[12240] = 32'b00000000000000010011101011111111;
assign LUT_3[12241] = 32'b00000000000000011010010111011100;
assign LUT_3[12242] = 32'b00000000000000010101110011100011;
assign LUT_3[12243] = 32'b00000000000000011100011111000000;
assign LUT_3[12244] = 32'b00000000000000010000111001110101;
assign LUT_3[12245] = 32'b00000000000000010111100101010010;
assign LUT_3[12246] = 32'b00000000000000010011000001011001;
assign LUT_3[12247] = 32'b00000000000000011001101100110110;
assign LUT_3[12248] = 32'b00000000000000011001000101000101;
assign LUT_3[12249] = 32'b00000000000000011111110000100010;
assign LUT_3[12250] = 32'b00000000000000011011001100101001;
assign LUT_3[12251] = 32'b00000000000000100001111000000110;
assign LUT_3[12252] = 32'b00000000000000010110010010111011;
assign LUT_3[12253] = 32'b00000000000000011100111110011000;
assign LUT_3[12254] = 32'b00000000000000011000011010011111;
assign LUT_3[12255] = 32'b00000000000000011111000101111100;
assign LUT_3[12256] = 32'b00000000000000010001100111011100;
assign LUT_3[12257] = 32'b00000000000000011000010010111001;
assign LUT_3[12258] = 32'b00000000000000010011101111000000;
assign LUT_3[12259] = 32'b00000000000000011010011010011101;
assign LUT_3[12260] = 32'b00000000000000001110110101010010;
assign LUT_3[12261] = 32'b00000000000000010101100000101111;
assign LUT_3[12262] = 32'b00000000000000010000111100110110;
assign LUT_3[12263] = 32'b00000000000000010111101000010011;
assign LUT_3[12264] = 32'b00000000000000010111000000100010;
assign LUT_3[12265] = 32'b00000000000000011101101011111111;
assign LUT_3[12266] = 32'b00000000000000011001001000000110;
assign LUT_3[12267] = 32'b00000000000000011111110011100011;
assign LUT_3[12268] = 32'b00000000000000010100001110011000;
assign LUT_3[12269] = 32'b00000000000000011010111001110101;
assign LUT_3[12270] = 32'b00000000000000010110010101111100;
assign LUT_3[12271] = 32'b00000000000000011101000001011001;
assign LUT_3[12272] = 32'b00000000000000010100111010011111;
assign LUT_3[12273] = 32'b00000000000000011011100101111100;
assign LUT_3[12274] = 32'b00000000000000010111000010000011;
assign LUT_3[12275] = 32'b00000000000000011101101101100000;
assign LUT_3[12276] = 32'b00000000000000010010001000010101;
assign LUT_3[12277] = 32'b00000000000000011000110011110010;
assign LUT_3[12278] = 32'b00000000000000010100001111111001;
assign LUT_3[12279] = 32'b00000000000000011010111011010110;
assign LUT_3[12280] = 32'b00000000000000011010010011100101;
assign LUT_3[12281] = 32'b00000000000000100000111111000010;
assign LUT_3[12282] = 32'b00000000000000011100011011001001;
assign LUT_3[12283] = 32'b00000000000000100011000110100110;
assign LUT_3[12284] = 32'b00000000000000010111100001011011;
assign LUT_3[12285] = 32'b00000000000000011110001100111000;
assign LUT_3[12286] = 32'b00000000000000011001101000111111;
assign LUT_3[12287] = 32'b00000000000000100000010100011100;
assign LUT_3[12288] = 32'b00000000000000001010100110110110;
assign LUT_3[12289] = 32'b00000000000000010001010010010011;
assign LUT_3[12290] = 32'b00000000000000001100101110011010;
assign LUT_3[12291] = 32'b00000000000000010011011001110111;
assign LUT_3[12292] = 32'b00000000000000000111110100101100;
assign LUT_3[12293] = 32'b00000000000000001110100000001001;
assign LUT_3[12294] = 32'b00000000000000001001111100010000;
assign LUT_3[12295] = 32'b00000000000000010000100111101101;
assign LUT_3[12296] = 32'b00000000000000001111111111111100;
assign LUT_3[12297] = 32'b00000000000000010110101011011001;
assign LUT_3[12298] = 32'b00000000000000010010000111100000;
assign LUT_3[12299] = 32'b00000000000000011000110010111101;
assign LUT_3[12300] = 32'b00000000000000001101001101110010;
assign LUT_3[12301] = 32'b00000000000000010011111001001111;
assign LUT_3[12302] = 32'b00000000000000001111010101010110;
assign LUT_3[12303] = 32'b00000000000000010110000000110011;
assign LUT_3[12304] = 32'b00000000000000001101111001111001;
assign LUT_3[12305] = 32'b00000000000000010100100101010110;
assign LUT_3[12306] = 32'b00000000000000010000000001011101;
assign LUT_3[12307] = 32'b00000000000000010110101100111010;
assign LUT_3[12308] = 32'b00000000000000001011000111101111;
assign LUT_3[12309] = 32'b00000000000000010001110011001100;
assign LUT_3[12310] = 32'b00000000000000001101001111010011;
assign LUT_3[12311] = 32'b00000000000000010011111010110000;
assign LUT_3[12312] = 32'b00000000000000010011010010111111;
assign LUT_3[12313] = 32'b00000000000000011001111110011100;
assign LUT_3[12314] = 32'b00000000000000010101011010100011;
assign LUT_3[12315] = 32'b00000000000000011100000110000000;
assign LUT_3[12316] = 32'b00000000000000010000100000110101;
assign LUT_3[12317] = 32'b00000000000000010111001100010010;
assign LUT_3[12318] = 32'b00000000000000010010101000011001;
assign LUT_3[12319] = 32'b00000000000000011001010011110110;
assign LUT_3[12320] = 32'b00000000000000001011110101010110;
assign LUT_3[12321] = 32'b00000000000000010010100000110011;
assign LUT_3[12322] = 32'b00000000000000001101111100111010;
assign LUT_3[12323] = 32'b00000000000000010100101000010111;
assign LUT_3[12324] = 32'b00000000000000001001000011001100;
assign LUT_3[12325] = 32'b00000000000000001111101110101001;
assign LUT_3[12326] = 32'b00000000000000001011001010110000;
assign LUT_3[12327] = 32'b00000000000000010001110110001101;
assign LUT_3[12328] = 32'b00000000000000010001001110011100;
assign LUT_3[12329] = 32'b00000000000000010111111001111001;
assign LUT_3[12330] = 32'b00000000000000010011010110000000;
assign LUT_3[12331] = 32'b00000000000000011010000001011101;
assign LUT_3[12332] = 32'b00000000000000001110011100010010;
assign LUT_3[12333] = 32'b00000000000000010101000111101111;
assign LUT_3[12334] = 32'b00000000000000010000100011110110;
assign LUT_3[12335] = 32'b00000000000000010111001111010011;
assign LUT_3[12336] = 32'b00000000000000001111001000011001;
assign LUT_3[12337] = 32'b00000000000000010101110011110110;
assign LUT_3[12338] = 32'b00000000000000010001001111111101;
assign LUT_3[12339] = 32'b00000000000000010111111011011010;
assign LUT_3[12340] = 32'b00000000000000001100010110001111;
assign LUT_3[12341] = 32'b00000000000000010011000001101100;
assign LUT_3[12342] = 32'b00000000000000001110011101110011;
assign LUT_3[12343] = 32'b00000000000000010101001001010000;
assign LUT_3[12344] = 32'b00000000000000010100100001011111;
assign LUT_3[12345] = 32'b00000000000000011011001100111100;
assign LUT_3[12346] = 32'b00000000000000010110101001000011;
assign LUT_3[12347] = 32'b00000000000000011101010100100000;
assign LUT_3[12348] = 32'b00000000000000010001101111010101;
assign LUT_3[12349] = 32'b00000000000000011000011010110010;
assign LUT_3[12350] = 32'b00000000000000010011110110111001;
assign LUT_3[12351] = 32'b00000000000000011010100010010110;
assign LUT_3[12352] = 32'b00000000000000001010011111100001;
assign LUT_3[12353] = 32'b00000000000000010001001010111110;
assign LUT_3[12354] = 32'b00000000000000001100100111000101;
assign LUT_3[12355] = 32'b00000000000000010011010010100010;
assign LUT_3[12356] = 32'b00000000000000000111101101010111;
assign LUT_3[12357] = 32'b00000000000000001110011000110100;
assign LUT_3[12358] = 32'b00000000000000001001110100111011;
assign LUT_3[12359] = 32'b00000000000000010000100000011000;
assign LUT_3[12360] = 32'b00000000000000001111111000100111;
assign LUT_3[12361] = 32'b00000000000000010110100100000100;
assign LUT_3[12362] = 32'b00000000000000010010000000001011;
assign LUT_3[12363] = 32'b00000000000000011000101011101000;
assign LUT_3[12364] = 32'b00000000000000001101000110011101;
assign LUT_3[12365] = 32'b00000000000000010011110001111010;
assign LUT_3[12366] = 32'b00000000000000001111001110000001;
assign LUT_3[12367] = 32'b00000000000000010101111001011110;
assign LUT_3[12368] = 32'b00000000000000001101110010100100;
assign LUT_3[12369] = 32'b00000000000000010100011110000001;
assign LUT_3[12370] = 32'b00000000000000001111111010001000;
assign LUT_3[12371] = 32'b00000000000000010110100101100101;
assign LUT_3[12372] = 32'b00000000000000001011000000011010;
assign LUT_3[12373] = 32'b00000000000000010001101011110111;
assign LUT_3[12374] = 32'b00000000000000001101000111111110;
assign LUT_3[12375] = 32'b00000000000000010011110011011011;
assign LUT_3[12376] = 32'b00000000000000010011001011101010;
assign LUT_3[12377] = 32'b00000000000000011001110111000111;
assign LUT_3[12378] = 32'b00000000000000010101010011001110;
assign LUT_3[12379] = 32'b00000000000000011011111110101011;
assign LUT_3[12380] = 32'b00000000000000010000011001100000;
assign LUT_3[12381] = 32'b00000000000000010111000100111101;
assign LUT_3[12382] = 32'b00000000000000010010100001000100;
assign LUT_3[12383] = 32'b00000000000000011001001100100001;
assign LUT_3[12384] = 32'b00000000000000001011101110000001;
assign LUT_3[12385] = 32'b00000000000000010010011001011110;
assign LUT_3[12386] = 32'b00000000000000001101110101100101;
assign LUT_3[12387] = 32'b00000000000000010100100001000010;
assign LUT_3[12388] = 32'b00000000000000001000111011110111;
assign LUT_3[12389] = 32'b00000000000000001111100111010100;
assign LUT_3[12390] = 32'b00000000000000001011000011011011;
assign LUT_3[12391] = 32'b00000000000000010001101110111000;
assign LUT_3[12392] = 32'b00000000000000010001000111000111;
assign LUT_3[12393] = 32'b00000000000000010111110010100100;
assign LUT_3[12394] = 32'b00000000000000010011001110101011;
assign LUT_3[12395] = 32'b00000000000000011001111010001000;
assign LUT_3[12396] = 32'b00000000000000001110010100111101;
assign LUT_3[12397] = 32'b00000000000000010101000000011010;
assign LUT_3[12398] = 32'b00000000000000010000011100100001;
assign LUT_3[12399] = 32'b00000000000000010111000111111110;
assign LUT_3[12400] = 32'b00000000000000001111000001000100;
assign LUT_3[12401] = 32'b00000000000000010101101100100001;
assign LUT_3[12402] = 32'b00000000000000010001001000101000;
assign LUT_3[12403] = 32'b00000000000000010111110100000101;
assign LUT_3[12404] = 32'b00000000000000001100001110111010;
assign LUT_3[12405] = 32'b00000000000000010010111010010111;
assign LUT_3[12406] = 32'b00000000000000001110010110011110;
assign LUT_3[12407] = 32'b00000000000000010101000001111011;
assign LUT_3[12408] = 32'b00000000000000010100011010001010;
assign LUT_3[12409] = 32'b00000000000000011011000101100111;
assign LUT_3[12410] = 32'b00000000000000010110100001101110;
assign LUT_3[12411] = 32'b00000000000000011101001101001011;
assign LUT_3[12412] = 32'b00000000000000010001101000000000;
assign LUT_3[12413] = 32'b00000000000000011000010011011101;
assign LUT_3[12414] = 32'b00000000000000010011101111100100;
assign LUT_3[12415] = 32'b00000000000000011010011011000001;
assign LUT_3[12416] = 32'b00000000000000001100110001110100;
assign LUT_3[12417] = 32'b00000000000000010011011101010001;
assign LUT_3[12418] = 32'b00000000000000001110111001011000;
assign LUT_3[12419] = 32'b00000000000000010101100100110101;
assign LUT_3[12420] = 32'b00000000000000001001111111101010;
assign LUT_3[12421] = 32'b00000000000000010000101011000111;
assign LUT_3[12422] = 32'b00000000000000001100000111001110;
assign LUT_3[12423] = 32'b00000000000000010010110010101011;
assign LUT_3[12424] = 32'b00000000000000010010001010111010;
assign LUT_3[12425] = 32'b00000000000000011000110110010111;
assign LUT_3[12426] = 32'b00000000000000010100010010011110;
assign LUT_3[12427] = 32'b00000000000000011010111101111011;
assign LUT_3[12428] = 32'b00000000000000001111011000110000;
assign LUT_3[12429] = 32'b00000000000000010110000100001101;
assign LUT_3[12430] = 32'b00000000000000010001100000010100;
assign LUT_3[12431] = 32'b00000000000000011000001011110001;
assign LUT_3[12432] = 32'b00000000000000010000000100110111;
assign LUT_3[12433] = 32'b00000000000000010110110000010100;
assign LUT_3[12434] = 32'b00000000000000010010001100011011;
assign LUT_3[12435] = 32'b00000000000000011000110111111000;
assign LUT_3[12436] = 32'b00000000000000001101010010101101;
assign LUT_3[12437] = 32'b00000000000000010011111110001010;
assign LUT_3[12438] = 32'b00000000000000001111011010010001;
assign LUT_3[12439] = 32'b00000000000000010110000101101110;
assign LUT_3[12440] = 32'b00000000000000010101011101111101;
assign LUT_3[12441] = 32'b00000000000000011100001001011010;
assign LUT_3[12442] = 32'b00000000000000010111100101100001;
assign LUT_3[12443] = 32'b00000000000000011110010000111110;
assign LUT_3[12444] = 32'b00000000000000010010101011110011;
assign LUT_3[12445] = 32'b00000000000000011001010111010000;
assign LUT_3[12446] = 32'b00000000000000010100110011010111;
assign LUT_3[12447] = 32'b00000000000000011011011110110100;
assign LUT_3[12448] = 32'b00000000000000001110000000010100;
assign LUT_3[12449] = 32'b00000000000000010100101011110001;
assign LUT_3[12450] = 32'b00000000000000010000000111111000;
assign LUT_3[12451] = 32'b00000000000000010110110011010101;
assign LUT_3[12452] = 32'b00000000000000001011001110001010;
assign LUT_3[12453] = 32'b00000000000000010001111001100111;
assign LUT_3[12454] = 32'b00000000000000001101010101101110;
assign LUT_3[12455] = 32'b00000000000000010100000001001011;
assign LUT_3[12456] = 32'b00000000000000010011011001011010;
assign LUT_3[12457] = 32'b00000000000000011010000100110111;
assign LUT_3[12458] = 32'b00000000000000010101100000111110;
assign LUT_3[12459] = 32'b00000000000000011100001100011011;
assign LUT_3[12460] = 32'b00000000000000010000100111010000;
assign LUT_3[12461] = 32'b00000000000000010111010010101101;
assign LUT_3[12462] = 32'b00000000000000010010101110110100;
assign LUT_3[12463] = 32'b00000000000000011001011010010001;
assign LUT_3[12464] = 32'b00000000000000010001010011010111;
assign LUT_3[12465] = 32'b00000000000000010111111110110100;
assign LUT_3[12466] = 32'b00000000000000010011011010111011;
assign LUT_3[12467] = 32'b00000000000000011010000110011000;
assign LUT_3[12468] = 32'b00000000000000001110100001001101;
assign LUT_3[12469] = 32'b00000000000000010101001100101010;
assign LUT_3[12470] = 32'b00000000000000010000101000110001;
assign LUT_3[12471] = 32'b00000000000000010111010100001110;
assign LUT_3[12472] = 32'b00000000000000010110101100011101;
assign LUT_3[12473] = 32'b00000000000000011101010111111010;
assign LUT_3[12474] = 32'b00000000000000011000110100000001;
assign LUT_3[12475] = 32'b00000000000000011111011111011110;
assign LUT_3[12476] = 32'b00000000000000010011111010010011;
assign LUT_3[12477] = 32'b00000000000000011010100101110000;
assign LUT_3[12478] = 32'b00000000000000010110000001110111;
assign LUT_3[12479] = 32'b00000000000000011100101101010100;
assign LUT_3[12480] = 32'b00000000000000001100101010011111;
assign LUT_3[12481] = 32'b00000000000000010011010101111100;
assign LUT_3[12482] = 32'b00000000000000001110110010000011;
assign LUT_3[12483] = 32'b00000000000000010101011101100000;
assign LUT_3[12484] = 32'b00000000000000001001111000010101;
assign LUT_3[12485] = 32'b00000000000000010000100011110010;
assign LUT_3[12486] = 32'b00000000000000001011111111111001;
assign LUT_3[12487] = 32'b00000000000000010010101011010110;
assign LUT_3[12488] = 32'b00000000000000010010000011100101;
assign LUT_3[12489] = 32'b00000000000000011000101111000010;
assign LUT_3[12490] = 32'b00000000000000010100001011001001;
assign LUT_3[12491] = 32'b00000000000000011010110110100110;
assign LUT_3[12492] = 32'b00000000000000001111010001011011;
assign LUT_3[12493] = 32'b00000000000000010101111100111000;
assign LUT_3[12494] = 32'b00000000000000010001011000111111;
assign LUT_3[12495] = 32'b00000000000000011000000100011100;
assign LUT_3[12496] = 32'b00000000000000001111111101100010;
assign LUT_3[12497] = 32'b00000000000000010110101000111111;
assign LUT_3[12498] = 32'b00000000000000010010000101000110;
assign LUT_3[12499] = 32'b00000000000000011000110000100011;
assign LUT_3[12500] = 32'b00000000000000001101001011011000;
assign LUT_3[12501] = 32'b00000000000000010011110110110101;
assign LUT_3[12502] = 32'b00000000000000001111010010111100;
assign LUT_3[12503] = 32'b00000000000000010101111110011001;
assign LUT_3[12504] = 32'b00000000000000010101010110101000;
assign LUT_3[12505] = 32'b00000000000000011100000010000101;
assign LUT_3[12506] = 32'b00000000000000010111011110001100;
assign LUT_3[12507] = 32'b00000000000000011110001001101001;
assign LUT_3[12508] = 32'b00000000000000010010100100011110;
assign LUT_3[12509] = 32'b00000000000000011001001111111011;
assign LUT_3[12510] = 32'b00000000000000010100101100000010;
assign LUT_3[12511] = 32'b00000000000000011011010111011111;
assign LUT_3[12512] = 32'b00000000000000001101111000111111;
assign LUT_3[12513] = 32'b00000000000000010100100100011100;
assign LUT_3[12514] = 32'b00000000000000010000000000100011;
assign LUT_3[12515] = 32'b00000000000000010110101100000000;
assign LUT_3[12516] = 32'b00000000000000001011000110110101;
assign LUT_3[12517] = 32'b00000000000000010001110010010010;
assign LUT_3[12518] = 32'b00000000000000001101001110011001;
assign LUT_3[12519] = 32'b00000000000000010011111001110110;
assign LUT_3[12520] = 32'b00000000000000010011010010000101;
assign LUT_3[12521] = 32'b00000000000000011001111101100010;
assign LUT_3[12522] = 32'b00000000000000010101011001101001;
assign LUT_3[12523] = 32'b00000000000000011100000101000110;
assign LUT_3[12524] = 32'b00000000000000010000011111111011;
assign LUT_3[12525] = 32'b00000000000000010111001011011000;
assign LUT_3[12526] = 32'b00000000000000010010100111011111;
assign LUT_3[12527] = 32'b00000000000000011001010010111100;
assign LUT_3[12528] = 32'b00000000000000010001001100000010;
assign LUT_3[12529] = 32'b00000000000000010111110111011111;
assign LUT_3[12530] = 32'b00000000000000010011010011100110;
assign LUT_3[12531] = 32'b00000000000000011001111111000011;
assign LUT_3[12532] = 32'b00000000000000001110011001111000;
assign LUT_3[12533] = 32'b00000000000000010101000101010101;
assign LUT_3[12534] = 32'b00000000000000010000100001011100;
assign LUT_3[12535] = 32'b00000000000000010111001100111001;
assign LUT_3[12536] = 32'b00000000000000010110100101001000;
assign LUT_3[12537] = 32'b00000000000000011101010000100101;
assign LUT_3[12538] = 32'b00000000000000011000101100101100;
assign LUT_3[12539] = 32'b00000000000000011111011000001001;
assign LUT_3[12540] = 32'b00000000000000010011110010111110;
assign LUT_3[12541] = 32'b00000000000000011010011110011011;
assign LUT_3[12542] = 32'b00000000000000010101111010100010;
assign LUT_3[12543] = 32'b00000000000000011100100101111111;
assign LUT_3[12544] = 32'b00000000000000000110110110010111;
assign LUT_3[12545] = 32'b00000000000000001101100001110100;
assign LUT_3[12546] = 32'b00000000000000001000111101111011;
assign LUT_3[12547] = 32'b00000000000000001111101001011000;
assign LUT_3[12548] = 32'b00000000000000000100000100001101;
assign LUT_3[12549] = 32'b00000000000000001010101111101010;
assign LUT_3[12550] = 32'b00000000000000000110001011110001;
assign LUT_3[12551] = 32'b00000000000000001100110111001110;
assign LUT_3[12552] = 32'b00000000000000001100001111011101;
assign LUT_3[12553] = 32'b00000000000000010010111010111010;
assign LUT_3[12554] = 32'b00000000000000001110010111000001;
assign LUT_3[12555] = 32'b00000000000000010101000010011110;
assign LUT_3[12556] = 32'b00000000000000001001011101010011;
assign LUT_3[12557] = 32'b00000000000000010000001000110000;
assign LUT_3[12558] = 32'b00000000000000001011100100110111;
assign LUT_3[12559] = 32'b00000000000000010010010000010100;
assign LUT_3[12560] = 32'b00000000000000001010001001011010;
assign LUT_3[12561] = 32'b00000000000000010000110100110111;
assign LUT_3[12562] = 32'b00000000000000001100010000111110;
assign LUT_3[12563] = 32'b00000000000000010010111100011011;
assign LUT_3[12564] = 32'b00000000000000000111010111010000;
assign LUT_3[12565] = 32'b00000000000000001110000010101101;
assign LUT_3[12566] = 32'b00000000000000001001011110110100;
assign LUT_3[12567] = 32'b00000000000000010000001010010001;
assign LUT_3[12568] = 32'b00000000000000001111100010100000;
assign LUT_3[12569] = 32'b00000000000000010110001101111101;
assign LUT_3[12570] = 32'b00000000000000010001101010000100;
assign LUT_3[12571] = 32'b00000000000000011000010101100001;
assign LUT_3[12572] = 32'b00000000000000001100110000010110;
assign LUT_3[12573] = 32'b00000000000000010011011011110011;
assign LUT_3[12574] = 32'b00000000000000001110110111111010;
assign LUT_3[12575] = 32'b00000000000000010101100011010111;
assign LUT_3[12576] = 32'b00000000000000001000000100110111;
assign LUT_3[12577] = 32'b00000000000000001110110000010100;
assign LUT_3[12578] = 32'b00000000000000001010001100011011;
assign LUT_3[12579] = 32'b00000000000000010000110111111000;
assign LUT_3[12580] = 32'b00000000000000000101010010101101;
assign LUT_3[12581] = 32'b00000000000000001011111110001010;
assign LUT_3[12582] = 32'b00000000000000000111011010010001;
assign LUT_3[12583] = 32'b00000000000000001110000101101110;
assign LUT_3[12584] = 32'b00000000000000001101011101111101;
assign LUT_3[12585] = 32'b00000000000000010100001001011010;
assign LUT_3[12586] = 32'b00000000000000001111100101100001;
assign LUT_3[12587] = 32'b00000000000000010110010000111110;
assign LUT_3[12588] = 32'b00000000000000001010101011110011;
assign LUT_3[12589] = 32'b00000000000000010001010111010000;
assign LUT_3[12590] = 32'b00000000000000001100110011010111;
assign LUT_3[12591] = 32'b00000000000000010011011110110100;
assign LUT_3[12592] = 32'b00000000000000001011010111111010;
assign LUT_3[12593] = 32'b00000000000000010010000011010111;
assign LUT_3[12594] = 32'b00000000000000001101011111011110;
assign LUT_3[12595] = 32'b00000000000000010100001010111011;
assign LUT_3[12596] = 32'b00000000000000001000100101110000;
assign LUT_3[12597] = 32'b00000000000000001111010001001101;
assign LUT_3[12598] = 32'b00000000000000001010101101010100;
assign LUT_3[12599] = 32'b00000000000000010001011000110001;
assign LUT_3[12600] = 32'b00000000000000010000110001000000;
assign LUT_3[12601] = 32'b00000000000000010111011100011101;
assign LUT_3[12602] = 32'b00000000000000010010111000100100;
assign LUT_3[12603] = 32'b00000000000000011001100100000001;
assign LUT_3[12604] = 32'b00000000000000001101111110110110;
assign LUT_3[12605] = 32'b00000000000000010100101010010011;
assign LUT_3[12606] = 32'b00000000000000010000000110011010;
assign LUT_3[12607] = 32'b00000000000000010110110001110111;
assign LUT_3[12608] = 32'b00000000000000000110101111000010;
assign LUT_3[12609] = 32'b00000000000000001101011010011111;
assign LUT_3[12610] = 32'b00000000000000001000110110100110;
assign LUT_3[12611] = 32'b00000000000000001111100010000011;
assign LUT_3[12612] = 32'b00000000000000000011111100111000;
assign LUT_3[12613] = 32'b00000000000000001010101000010101;
assign LUT_3[12614] = 32'b00000000000000000110000100011100;
assign LUT_3[12615] = 32'b00000000000000001100101111111001;
assign LUT_3[12616] = 32'b00000000000000001100001000001000;
assign LUT_3[12617] = 32'b00000000000000010010110011100101;
assign LUT_3[12618] = 32'b00000000000000001110001111101100;
assign LUT_3[12619] = 32'b00000000000000010100111011001001;
assign LUT_3[12620] = 32'b00000000000000001001010101111110;
assign LUT_3[12621] = 32'b00000000000000010000000001011011;
assign LUT_3[12622] = 32'b00000000000000001011011101100010;
assign LUT_3[12623] = 32'b00000000000000010010001000111111;
assign LUT_3[12624] = 32'b00000000000000001010000010000101;
assign LUT_3[12625] = 32'b00000000000000010000101101100010;
assign LUT_3[12626] = 32'b00000000000000001100001001101001;
assign LUT_3[12627] = 32'b00000000000000010010110101000110;
assign LUT_3[12628] = 32'b00000000000000000111001111111011;
assign LUT_3[12629] = 32'b00000000000000001101111011011000;
assign LUT_3[12630] = 32'b00000000000000001001010111011111;
assign LUT_3[12631] = 32'b00000000000000010000000010111100;
assign LUT_3[12632] = 32'b00000000000000001111011011001011;
assign LUT_3[12633] = 32'b00000000000000010110000110101000;
assign LUT_3[12634] = 32'b00000000000000010001100010101111;
assign LUT_3[12635] = 32'b00000000000000011000001110001100;
assign LUT_3[12636] = 32'b00000000000000001100101001000001;
assign LUT_3[12637] = 32'b00000000000000010011010100011110;
assign LUT_3[12638] = 32'b00000000000000001110110000100101;
assign LUT_3[12639] = 32'b00000000000000010101011100000010;
assign LUT_3[12640] = 32'b00000000000000000111111101100010;
assign LUT_3[12641] = 32'b00000000000000001110101000111111;
assign LUT_3[12642] = 32'b00000000000000001010000101000110;
assign LUT_3[12643] = 32'b00000000000000010000110000100011;
assign LUT_3[12644] = 32'b00000000000000000101001011011000;
assign LUT_3[12645] = 32'b00000000000000001011110110110101;
assign LUT_3[12646] = 32'b00000000000000000111010010111100;
assign LUT_3[12647] = 32'b00000000000000001101111110011001;
assign LUT_3[12648] = 32'b00000000000000001101010110101000;
assign LUT_3[12649] = 32'b00000000000000010100000010000101;
assign LUT_3[12650] = 32'b00000000000000001111011110001100;
assign LUT_3[12651] = 32'b00000000000000010110001001101001;
assign LUT_3[12652] = 32'b00000000000000001010100100011110;
assign LUT_3[12653] = 32'b00000000000000010001001111111011;
assign LUT_3[12654] = 32'b00000000000000001100101100000010;
assign LUT_3[12655] = 32'b00000000000000010011010111011111;
assign LUT_3[12656] = 32'b00000000000000001011010000100101;
assign LUT_3[12657] = 32'b00000000000000010001111100000010;
assign LUT_3[12658] = 32'b00000000000000001101011000001001;
assign LUT_3[12659] = 32'b00000000000000010100000011100110;
assign LUT_3[12660] = 32'b00000000000000001000011110011011;
assign LUT_3[12661] = 32'b00000000000000001111001001111000;
assign LUT_3[12662] = 32'b00000000000000001010100101111111;
assign LUT_3[12663] = 32'b00000000000000010001010001011100;
assign LUT_3[12664] = 32'b00000000000000010000101001101011;
assign LUT_3[12665] = 32'b00000000000000010111010101001000;
assign LUT_3[12666] = 32'b00000000000000010010110001001111;
assign LUT_3[12667] = 32'b00000000000000011001011100101100;
assign LUT_3[12668] = 32'b00000000000000001101110111100001;
assign LUT_3[12669] = 32'b00000000000000010100100010111110;
assign LUT_3[12670] = 32'b00000000000000001111111111000101;
assign LUT_3[12671] = 32'b00000000000000010110101010100010;
assign LUT_3[12672] = 32'b00000000000000001001000001010101;
assign LUT_3[12673] = 32'b00000000000000001111101100110010;
assign LUT_3[12674] = 32'b00000000000000001011001000111001;
assign LUT_3[12675] = 32'b00000000000000010001110100010110;
assign LUT_3[12676] = 32'b00000000000000000110001111001011;
assign LUT_3[12677] = 32'b00000000000000001100111010101000;
assign LUT_3[12678] = 32'b00000000000000001000010110101111;
assign LUT_3[12679] = 32'b00000000000000001111000010001100;
assign LUT_3[12680] = 32'b00000000000000001110011010011011;
assign LUT_3[12681] = 32'b00000000000000010101000101111000;
assign LUT_3[12682] = 32'b00000000000000010000100001111111;
assign LUT_3[12683] = 32'b00000000000000010111001101011100;
assign LUT_3[12684] = 32'b00000000000000001011101000010001;
assign LUT_3[12685] = 32'b00000000000000010010010011101110;
assign LUT_3[12686] = 32'b00000000000000001101101111110101;
assign LUT_3[12687] = 32'b00000000000000010100011011010010;
assign LUT_3[12688] = 32'b00000000000000001100010100011000;
assign LUT_3[12689] = 32'b00000000000000010010111111110101;
assign LUT_3[12690] = 32'b00000000000000001110011011111100;
assign LUT_3[12691] = 32'b00000000000000010101000111011001;
assign LUT_3[12692] = 32'b00000000000000001001100010001110;
assign LUT_3[12693] = 32'b00000000000000010000001101101011;
assign LUT_3[12694] = 32'b00000000000000001011101001110010;
assign LUT_3[12695] = 32'b00000000000000010010010101001111;
assign LUT_3[12696] = 32'b00000000000000010001101101011110;
assign LUT_3[12697] = 32'b00000000000000011000011000111011;
assign LUT_3[12698] = 32'b00000000000000010011110101000010;
assign LUT_3[12699] = 32'b00000000000000011010100000011111;
assign LUT_3[12700] = 32'b00000000000000001110111011010100;
assign LUT_3[12701] = 32'b00000000000000010101100110110001;
assign LUT_3[12702] = 32'b00000000000000010001000010111000;
assign LUT_3[12703] = 32'b00000000000000010111101110010101;
assign LUT_3[12704] = 32'b00000000000000001010001111110101;
assign LUT_3[12705] = 32'b00000000000000010000111011010010;
assign LUT_3[12706] = 32'b00000000000000001100010111011001;
assign LUT_3[12707] = 32'b00000000000000010011000010110110;
assign LUT_3[12708] = 32'b00000000000000000111011101101011;
assign LUT_3[12709] = 32'b00000000000000001110001001001000;
assign LUT_3[12710] = 32'b00000000000000001001100101001111;
assign LUT_3[12711] = 32'b00000000000000010000010000101100;
assign LUT_3[12712] = 32'b00000000000000001111101000111011;
assign LUT_3[12713] = 32'b00000000000000010110010100011000;
assign LUT_3[12714] = 32'b00000000000000010001110000011111;
assign LUT_3[12715] = 32'b00000000000000011000011011111100;
assign LUT_3[12716] = 32'b00000000000000001100110110110001;
assign LUT_3[12717] = 32'b00000000000000010011100010001110;
assign LUT_3[12718] = 32'b00000000000000001110111110010101;
assign LUT_3[12719] = 32'b00000000000000010101101001110010;
assign LUT_3[12720] = 32'b00000000000000001101100010111000;
assign LUT_3[12721] = 32'b00000000000000010100001110010101;
assign LUT_3[12722] = 32'b00000000000000001111101010011100;
assign LUT_3[12723] = 32'b00000000000000010110010101111001;
assign LUT_3[12724] = 32'b00000000000000001010110000101110;
assign LUT_3[12725] = 32'b00000000000000010001011100001011;
assign LUT_3[12726] = 32'b00000000000000001100111000010010;
assign LUT_3[12727] = 32'b00000000000000010011100011101111;
assign LUT_3[12728] = 32'b00000000000000010010111011111110;
assign LUT_3[12729] = 32'b00000000000000011001100111011011;
assign LUT_3[12730] = 32'b00000000000000010101000011100010;
assign LUT_3[12731] = 32'b00000000000000011011101110111111;
assign LUT_3[12732] = 32'b00000000000000010000001001110100;
assign LUT_3[12733] = 32'b00000000000000010110110101010001;
assign LUT_3[12734] = 32'b00000000000000010010010001011000;
assign LUT_3[12735] = 32'b00000000000000011000111100110101;
assign LUT_3[12736] = 32'b00000000000000001000111010000000;
assign LUT_3[12737] = 32'b00000000000000001111100101011101;
assign LUT_3[12738] = 32'b00000000000000001011000001100100;
assign LUT_3[12739] = 32'b00000000000000010001101101000001;
assign LUT_3[12740] = 32'b00000000000000000110000111110110;
assign LUT_3[12741] = 32'b00000000000000001100110011010011;
assign LUT_3[12742] = 32'b00000000000000001000001111011010;
assign LUT_3[12743] = 32'b00000000000000001110111010110111;
assign LUT_3[12744] = 32'b00000000000000001110010011000110;
assign LUT_3[12745] = 32'b00000000000000010100111110100011;
assign LUT_3[12746] = 32'b00000000000000010000011010101010;
assign LUT_3[12747] = 32'b00000000000000010111000110000111;
assign LUT_3[12748] = 32'b00000000000000001011100000111100;
assign LUT_3[12749] = 32'b00000000000000010010001100011001;
assign LUT_3[12750] = 32'b00000000000000001101101000100000;
assign LUT_3[12751] = 32'b00000000000000010100010011111101;
assign LUT_3[12752] = 32'b00000000000000001100001101000011;
assign LUT_3[12753] = 32'b00000000000000010010111000100000;
assign LUT_3[12754] = 32'b00000000000000001110010100100111;
assign LUT_3[12755] = 32'b00000000000000010101000000000100;
assign LUT_3[12756] = 32'b00000000000000001001011010111001;
assign LUT_3[12757] = 32'b00000000000000010000000110010110;
assign LUT_3[12758] = 32'b00000000000000001011100010011101;
assign LUT_3[12759] = 32'b00000000000000010010001101111010;
assign LUT_3[12760] = 32'b00000000000000010001100110001001;
assign LUT_3[12761] = 32'b00000000000000011000010001100110;
assign LUT_3[12762] = 32'b00000000000000010011101101101101;
assign LUT_3[12763] = 32'b00000000000000011010011001001010;
assign LUT_3[12764] = 32'b00000000000000001110110011111111;
assign LUT_3[12765] = 32'b00000000000000010101011111011100;
assign LUT_3[12766] = 32'b00000000000000010000111011100011;
assign LUT_3[12767] = 32'b00000000000000010111100111000000;
assign LUT_3[12768] = 32'b00000000000000001010001000100000;
assign LUT_3[12769] = 32'b00000000000000010000110011111101;
assign LUT_3[12770] = 32'b00000000000000001100010000000100;
assign LUT_3[12771] = 32'b00000000000000010010111011100001;
assign LUT_3[12772] = 32'b00000000000000000111010110010110;
assign LUT_3[12773] = 32'b00000000000000001110000001110011;
assign LUT_3[12774] = 32'b00000000000000001001011101111010;
assign LUT_3[12775] = 32'b00000000000000010000001001010111;
assign LUT_3[12776] = 32'b00000000000000001111100001100110;
assign LUT_3[12777] = 32'b00000000000000010110001101000011;
assign LUT_3[12778] = 32'b00000000000000010001101001001010;
assign LUT_3[12779] = 32'b00000000000000011000010100100111;
assign LUT_3[12780] = 32'b00000000000000001100101111011100;
assign LUT_3[12781] = 32'b00000000000000010011011010111001;
assign LUT_3[12782] = 32'b00000000000000001110110111000000;
assign LUT_3[12783] = 32'b00000000000000010101100010011101;
assign LUT_3[12784] = 32'b00000000000000001101011011100011;
assign LUT_3[12785] = 32'b00000000000000010100000111000000;
assign LUT_3[12786] = 32'b00000000000000001111100011000111;
assign LUT_3[12787] = 32'b00000000000000010110001110100100;
assign LUT_3[12788] = 32'b00000000000000001010101001011001;
assign LUT_3[12789] = 32'b00000000000000010001010100110110;
assign LUT_3[12790] = 32'b00000000000000001100110000111101;
assign LUT_3[12791] = 32'b00000000000000010011011100011010;
assign LUT_3[12792] = 32'b00000000000000010010110100101001;
assign LUT_3[12793] = 32'b00000000000000011001100000000110;
assign LUT_3[12794] = 32'b00000000000000010100111100001101;
assign LUT_3[12795] = 32'b00000000000000011011100111101010;
assign LUT_3[12796] = 32'b00000000000000010000000010011111;
assign LUT_3[12797] = 32'b00000000000000010110101101111100;
assign LUT_3[12798] = 32'b00000000000000010010001010000011;
assign LUT_3[12799] = 32'b00000000000000011000110101100000;
assign LUT_3[12800] = 32'b00000000000000001101111100000010;
assign LUT_3[12801] = 32'b00000000000000010100100111011111;
assign LUT_3[12802] = 32'b00000000000000010000000011100110;
assign LUT_3[12803] = 32'b00000000000000010110101111000011;
assign LUT_3[12804] = 32'b00000000000000001011001001111000;
assign LUT_3[12805] = 32'b00000000000000010001110101010101;
assign LUT_3[12806] = 32'b00000000000000001101010001011100;
assign LUT_3[12807] = 32'b00000000000000010011111100111001;
assign LUT_3[12808] = 32'b00000000000000010011010101001000;
assign LUT_3[12809] = 32'b00000000000000011010000000100101;
assign LUT_3[12810] = 32'b00000000000000010101011100101100;
assign LUT_3[12811] = 32'b00000000000000011100001000001001;
assign LUT_3[12812] = 32'b00000000000000010000100010111110;
assign LUT_3[12813] = 32'b00000000000000010111001110011011;
assign LUT_3[12814] = 32'b00000000000000010010101010100010;
assign LUT_3[12815] = 32'b00000000000000011001010101111111;
assign LUT_3[12816] = 32'b00000000000000010001001111000101;
assign LUT_3[12817] = 32'b00000000000000010111111010100010;
assign LUT_3[12818] = 32'b00000000000000010011010110101001;
assign LUT_3[12819] = 32'b00000000000000011010000010000110;
assign LUT_3[12820] = 32'b00000000000000001110011100111011;
assign LUT_3[12821] = 32'b00000000000000010101001000011000;
assign LUT_3[12822] = 32'b00000000000000010000100100011111;
assign LUT_3[12823] = 32'b00000000000000010111001111111100;
assign LUT_3[12824] = 32'b00000000000000010110101000001011;
assign LUT_3[12825] = 32'b00000000000000011101010011101000;
assign LUT_3[12826] = 32'b00000000000000011000101111101111;
assign LUT_3[12827] = 32'b00000000000000011111011011001100;
assign LUT_3[12828] = 32'b00000000000000010011110110000001;
assign LUT_3[12829] = 32'b00000000000000011010100001011110;
assign LUT_3[12830] = 32'b00000000000000010101111101100101;
assign LUT_3[12831] = 32'b00000000000000011100101001000010;
assign LUT_3[12832] = 32'b00000000000000001111001010100010;
assign LUT_3[12833] = 32'b00000000000000010101110101111111;
assign LUT_3[12834] = 32'b00000000000000010001010010000110;
assign LUT_3[12835] = 32'b00000000000000010111111101100011;
assign LUT_3[12836] = 32'b00000000000000001100011000011000;
assign LUT_3[12837] = 32'b00000000000000010011000011110101;
assign LUT_3[12838] = 32'b00000000000000001110011111111100;
assign LUT_3[12839] = 32'b00000000000000010101001011011001;
assign LUT_3[12840] = 32'b00000000000000010100100011101000;
assign LUT_3[12841] = 32'b00000000000000011011001111000101;
assign LUT_3[12842] = 32'b00000000000000010110101011001100;
assign LUT_3[12843] = 32'b00000000000000011101010110101001;
assign LUT_3[12844] = 32'b00000000000000010001110001011110;
assign LUT_3[12845] = 32'b00000000000000011000011100111011;
assign LUT_3[12846] = 32'b00000000000000010011111001000010;
assign LUT_3[12847] = 32'b00000000000000011010100100011111;
assign LUT_3[12848] = 32'b00000000000000010010011101100101;
assign LUT_3[12849] = 32'b00000000000000011001001001000010;
assign LUT_3[12850] = 32'b00000000000000010100100101001001;
assign LUT_3[12851] = 32'b00000000000000011011010000100110;
assign LUT_3[12852] = 32'b00000000000000001111101011011011;
assign LUT_3[12853] = 32'b00000000000000010110010110111000;
assign LUT_3[12854] = 32'b00000000000000010001110010111111;
assign LUT_3[12855] = 32'b00000000000000011000011110011100;
assign LUT_3[12856] = 32'b00000000000000010111110110101011;
assign LUT_3[12857] = 32'b00000000000000011110100010001000;
assign LUT_3[12858] = 32'b00000000000000011001111110001111;
assign LUT_3[12859] = 32'b00000000000000100000101001101100;
assign LUT_3[12860] = 32'b00000000000000010101000100100001;
assign LUT_3[12861] = 32'b00000000000000011011101111111110;
assign LUT_3[12862] = 32'b00000000000000010111001100000101;
assign LUT_3[12863] = 32'b00000000000000011101110111100010;
assign LUT_3[12864] = 32'b00000000000000001101110100101101;
assign LUT_3[12865] = 32'b00000000000000010100100000001010;
assign LUT_3[12866] = 32'b00000000000000001111111100010001;
assign LUT_3[12867] = 32'b00000000000000010110100111101110;
assign LUT_3[12868] = 32'b00000000000000001011000010100011;
assign LUT_3[12869] = 32'b00000000000000010001101110000000;
assign LUT_3[12870] = 32'b00000000000000001101001010000111;
assign LUT_3[12871] = 32'b00000000000000010011110101100100;
assign LUT_3[12872] = 32'b00000000000000010011001101110011;
assign LUT_3[12873] = 32'b00000000000000011001111001010000;
assign LUT_3[12874] = 32'b00000000000000010101010101010111;
assign LUT_3[12875] = 32'b00000000000000011100000000110100;
assign LUT_3[12876] = 32'b00000000000000010000011011101001;
assign LUT_3[12877] = 32'b00000000000000010111000111000110;
assign LUT_3[12878] = 32'b00000000000000010010100011001101;
assign LUT_3[12879] = 32'b00000000000000011001001110101010;
assign LUT_3[12880] = 32'b00000000000000010001000111110000;
assign LUT_3[12881] = 32'b00000000000000010111110011001101;
assign LUT_3[12882] = 32'b00000000000000010011001111010100;
assign LUT_3[12883] = 32'b00000000000000011001111010110001;
assign LUT_3[12884] = 32'b00000000000000001110010101100110;
assign LUT_3[12885] = 32'b00000000000000010101000001000011;
assign LUT_3[12886] = 32'b00000000000000010000011101001010;
assign LUT_3[12887] = 32'b00000000000000010111001000100111;
assign LUT_3[12888] = 32'b00000000000000010110100000110110;
assign LUT_3[12889] = 32'b00000000000000011101001100010011;
assign LUT_3[12890] = 32'b00000000000000011000101000011010;
assign LUT_3[12891] = 32'b00000000000000011111010011110111;
assign LUT_3[12892] = 32'b00000000000000010011101110101100;
assign LUT_3[12893] = 32'b00000000000000011010011010001001;
assign LUT_3[12894] = 32'b00000000000000010101110110010000;
assign LUT_3[12895] = 32'b00000000000000011100100001101101;
assign LUT_3[12896] = 32'b00000000000000001111000011001101;
assign LUT_3[12897] = 32'b00000000000000010101101110101010;
assign LUT_3[12898] = 32'b00000000000000010001001010110001;
assign LUT_3[12899] = 32'b00000000000000010111110110001110;
assign LUT_3[12900] = 32'b00000000000000001100010001000011;
assign LUT_3[12901] = 32'b00000000000000010010111100100000;
assign LUT_3[12902] = 32'b00000000000000001110011000100111;
assign LUT_3[12903] = 32'b00000000000000010101000100000100;
assign LUT_3[12904] = 32'b00000000000000010100011100010011;
assign LUT_3[12905] = 32'b00000000000000011011000111110000;
assign LUT_3[12906] = 32'b00000000000000010110100011110111;
assign LUT_3[12907] = 32'b00000000000000011101001111010100;
assign LUT_3[12908] = 32'b00000000000000010001101010001001;
assign LUT_3[12909] = 32'b00000000000000011000010101100110;
assign LUT_3[12910] = 32'b00000000000000010011110001101101;
assign LUT_3[12911] = 32'b00000000000000011010011101001010;
assign LUT_3[12912] = 32'b00000000000000010010010110010000;
assign LUT_3[12913] = 32'b00000000000000011001000001101101;
assign LUT_3[12914] = 32'b00000000000000010100011101110100;
assign LUT_3[12915] = 32'b00000000000000011011001001010001;
assign LUT_3[12916] = 32'b00000000000000001111100100000110;
assign LUT_3[12917] = 32'b00000000000000010110001111100011;
assign LUT_3[12918] = 32'b00000000000000010001101011101010;
assign LUT_3[12919] = 32'b00000000000000011000010111000111;
assign LUT_3[12920] = 32'b00000000000000010111101111010110;
assign LUT_3[12921] = 32'b00000000000000011110011010110011;
assign LUT_3[12922] = 32'b00000000000000011001110110111010;
assign LUT_3[12923] = 32'b00000000000000100000100010010111;
assign LUT_3[12924] = 32'b00000000000000010100111101001100;
assign LUT_3[12925] = 32'b00000000000000011011101000101001;
assign LUT_3[12926] = 32'b00000000000000010111000100110000;
assign LUT_3[12927] = 32'b00000000000000011101110000001101;
assign LUT_3[12928] = 32'b00000000000000010000000111000000;
assign LUT_3[12929] = 32'b00000000000000010110110010011101;
assign LUT_3[12930] = 32'b00000000000000010010001110100100;
assign LUT_3[12931] = 32'b00000000000000011000111010000001;
assign LUT_3[12932] = 32'b00000000000000001101010100110110;
assign LUT_3[12933] = 32'b00000000000000010100000000010011;
assign LUT_3[12934] = 32'b00000000000000001111011100011010;
assign LUT_3[12935] = 32'b00000000000000010110000111110111;
assign LUT_3[12936] = 32'b00000000000000010101100000000110;
assign LUT_3[12937] = 32'b00000000000000011100001011100011;
assign LUT_3[12938] = 32'b00000000000000010111100111101010;
assign LUT_3[12939] = 32'b00000000000000011110010011000111;
assign LUT_3[12940] = 32'b00000000000000010010101101111100;
assign LUT_3[12941] = 32'b00000000000000011001011001011001;
assign LUT_3[12942] = 32'b00000000000000010100110101100000;
assign LUT_3[12943] = 32'b00000000000000011011100000111101;
assign LUT_3[12944] = 32'b00000000000000010011011010000011;
assign LUT_3[12945] = 32'b00000000000000011010000101100000;
assign LUT_3[12946] = 32'b00000000000000010101100001100111;
assign LUT_3[12947] = 32'b00000000000000011100001101000100;
assign LUT_3[12948] = 32'b00000000000000010000100111111001;
assign LUT_3[12949] = 32'b00000000000000010111010011010110;
assign LUT_3[12950] = 32'b00000000000000010010101111011101;
assign LUT_3[12951] = 32'b00000000000000011001011010111010;
assign LUT_3[12952] = 32'b00000000000000011000110011001001;
assign LUT_3[12953] = 32'b00000000000000011111011110100110;
assign LUT_3[12954] = 32'b00000000000000011010111010101101;
assign LUT_3[12955] = 32'b00000000000000100001100110001010;
assign LUT_3[12956] = 32'b00000000000000010110000000111111;
assign LUT_3[12957] = 32'b00000000000000011100101100011100;
assign LUT_3[12958] = 32'b00000000000000011000001000100011;
assign LUT_3[12959] = 32'b00000000000000011110110100000000;
assign LUT_3[12960] = 32'b00000000000000010001010101100000;
assign LUT_3[12961] = 32'b00000000000000011000000000111101;
assign LUT_3[12962] = 32'b00000000000000010011011101000100;
assign LUT_3[12963] = 32'b00000000000000011010001000100001;
assign LUT_3[12964] = 32'b00000000000000001110100011010110;
assign LUT_3[12965] = 32'b00000000000000010101001110110011;
assign LUT_3[12966] = 32'b00000000000000010000101010111010;
assign LUT_3[12967] = 32'b00000000000000010111010110010111;
assign LUT_3[12968] = 32'b00000000000000010110101110100110;
assign LUT_3[12969] = 32'b00000000000000011101011010000011;
assign LUT_3[12970] = 32'b00000000000000011000110110001010;
assign LUT_3[12971] = 32'b00000000000000011111100001100111;
assign LUT_3[12972] = 32'b00000000000000010011111100011100;
assign LUT_3[12973] = 32'b00000000000000011010100111111001;
assign LUT_3[12974] = 32'b00000000000000010110000100000000;
assign LUT_3[12975] = 32'b00000000000000011100101111011101;
assign LUT_3[12976] = 32'b00000000000000010100101000100011;
assign LUT_3[12977] = 32'b00000000000000011011010100000000;
assign LUT_3[12978] = 32'b00000000000000010110110000000111;
assign LUT_3[12979] = 32'b00000000000000011101011011100100;
assign LUT_3[12980] = 32'b00000000000000010001110110011001;
assign LUT_3[12981] = 32'b00000000000000011000100001110110;
assign LUT_3[12982] = 32'b00000000000000010011111101111101;
assign LUT_3[12983] = 32'b00000000000000011010101001011010;
assign LUT_3[12984] = 32'b00000000000000011010000001101001;
assign LUT_3[12985] = 32'b00000000000000100000101101000110;
assign LUT_3[12986] = 32'b00000000000000011100001001001101;
assign LUT_3[12987] = 32'b00000000000000100010110100101010;
assign LUT_3[12988] = 32'b00000000000000010111001111011111;
assign LUT_3[12989] = 32'b00000000000000011101111010111100;
assign LUT_3[12990] = 32'b00000000000000011001010111000011;
assign LUT_3[12991] = 32'b00000000000000100000000010100000;
assign LUT_3[12992] = 32'b00000000000000001111111111101011;
assign LUT_3[12993] = 32'b00000000000000010110101011001000;
assign LUT_3[12994] = 32'b00000000000000010010000111001111;
assign LUT_3[12995] = 32'b00000000000000011000110010101100;
assign LUT_3[12996] = 32'b00000000000000001101001101100001;
assign LUT_3[12997] = 32'b00000000000000010011111000111110;
assign LUT_3[12998] = 32'b00000000000000001111010101000101;
assign LUT_3[12999] = 32'b00000000000000010110000000100010;
assign LUT_3[13000] = 32'b00000000000000010101011000110001;
assign LUT_3[13001] = 32'b00000000000000011100000100001110;
assign LUT_3[13002] = 32'b00000000000000010111100000010101;
assign LUT_3[13003] = 32'b00000000000000011110001011110010;
assign LUT_3[13004] = 32'b00000000000000010010100110100111;
assign LUT_3[13005] = 32'b00000000000000011001010010000100;
assign LUT_3[13006] = 32'b00000000000000010100101110001011;
assign LUT_3[13007] = 32'b00000000000000011011011001101000;
assign LUT_3[13008] = 32'b00000000000000010011010010101110;
assign LUT_3[13009] = 32'b00000000000000011001111110001011;
assign LUT_3[13010] = 32'b00000000000000010101011010010010;
assign LUT_3[13011] = 32'b00000000000000011100000101101111;
assign LUT_3[13012] = 32'b00000000000000010000100000100100;
assign LUT_3[13013] = 32'b00000000000000010111001100000001;
assign LUT_3[13014] = 32'b00000000000000010010101000001000;
assign LUT_3[13015] = 32'b00000000000000011001010011100101;
assign LUT_3[13016] = 32'b00000000000000011000101011110100;
assign LUT_3[13017] = 32'b00000000000000011111010111010001;
assign LUT_3[13018] = 32'b00000000000000011010110011011000;
assign LUT_3[13019] = 32'b00000000000000100001011110110101;
assign LUT_3[13020] = 32'b00000000000000010101111001101010;
assign LUT_3[13021] = 32'b00000000000000011100100101000111;
assign LUT_3[13022] = 32'b00000000000000011000000001001110;
assign LUT_3[13023] = 32'b00000000000000011110101100101011;
assign LUT_3[13024] = 32'b00000000000000010001001110001011;
assign LUT_3[13025] = 32'b00000000000000010111111001101000;
assign LUT_3[13026] = 32'b00000000000000010011010101101111;
assign LUT_3[13027] = 32'b00000000000000011010000001001100;
assign LUT_3[13028] = 32'b00000000000000001110011100000001;
assign LUT_3[13029] = 32'b00000000000000010101000111011110;
assign LUT_3[13030] = 32'b00000000000000010000100011100101;
assign LUT_3[13031] = 32'b00000000000000010111001111000010;
assign LUT_3[13032] = 32'b00000000000000010110100111010001;
assign LUT_3[13033] = 32'b00000000000000011101010010101110;
assign LUT_3[13034] = 32'b00000000000000011000101110110101;
assign LUT_3[13035] = 32'b00000000000000011111011010010010;
assign LUT_3[13036] = 32'b00000000000000010011110101000111;
assign LUT_3[13037] = 32'b00000000000000011010100000100100;
assign LUT_3[13038] = 32'b00000000000000010101111100101011;
assign LUT_3[13039] = 32'b00000000000000011100101000001000;
assign LUT_3[13040] = 32'b00000000000000010100100001001110;
assign LUT_3[13041] = 32'b00000000000000011011001100101011;
assign LUT_3[13042] = 32'b00000000000000010110101000110010;
assign LUT_3[13043] = 32'b00000000000000011101010100001111;
assign LUT_3[13044] = 32'b00000000000000010001101111000100;
assign LUT_3[13045] = 32'b00000000000000011000011010100001;
assign LUT_3[13046] = 32'b00000000000000010011110110101000;
assign LUT_3[13047] = 32'b00000000000000011010100010000101;
assign LUT_3[13048] = 32'b00000000000000011001111010010100;
assign LUT_3[13049] = 32'b00000000000000100000100101110001;
assign LUT_3[13050] = 32'b00000000000000011100000001111000;
assign LUT_3[13051] = 32'b00000000000000100010101101010101;
assign LUT_3[13052] = 32'b00000000000000010111001000001010;
assign LUT_3[13053] = 32'b00000000000000011101110011100111;
assign LUT_3[13054] = 32'b00000000000000011001001111101110;
assign LUT_3[13055] = 32'b00000000000000011111111011001011;
assign LUT_3[13056] = 32'b00000000000000001010001011100011;
assign LUT_3[13057] = 32'b00000000000000010000110111000000;
assign LUT_3[13058] = 32'b00000000000000001100010011000111;
assign LUT_3[13059] = 32'b00000000000000010010111110100100;
assign LUT_3[13060] = 32'b00000000000000000111011001011001;
assign LUT_3[13061] = 32'b00000000000000001110000100110110;
assign LUT_3[13062] = 32'b00000000000000001001100000111101;
assign LUT_3[13063] = 32'b00000000000000010000001100011010;
assign LUT_3[13064] = 32'b00000000000000001111100100101001;
assign LUT_3[13065] = 32'b00000000000000010110010000000110;
assign LUT_3[13066] = 32'b00000000000000010001101100001101;
assign LUT_3[13067] = 32'b00000000000000011000010111101010;
assign LUT_3[13068] = 32'b00000000000000001100110010011111;
assign LUT_3[13069] = 32'b00000000000000010011011101111100;
assign LUT_3[13070] = 32'b00000000000000001110111010000011;
assign LUT_3[13071] = 32'b00000000000000010101100101100000;
assign LUT_3[13072] = 32'b00000000000000001101011110100110;
assign LUT_3[13073] = 32'b00000000000000010100001010000011;
assign LUT_3[13074] = 32'b00000000000000001111100110001010;
assign LUT_3[13075] = 32'b00000000000000010110010001100111;
assign LUT_3[13076] = 32'b00000000000000001010101100011100;
assign LUT_3[13077] = 32'b00000000000000010001010111111001;
assign LUT_3[13078] = 32'b00000000000000001100110100000000;
assign LUT_3[13079] = 32'b00000000000000010011011111011101;
assign LUT_3[13080] = 32'b00000000000000010010110111101100;
assign LUT_3[13081] = 32'b00000000000000011001100011001001;
assign LUT_3[13082] = 32'b00000000000000010100111111010000;
assign LUT_3[13083] = 32'b00000000000000011011101010101101;
assign LUT_3[13084] = 32'b00000000000000010000000101100010;
assign LUT_3[13085] = 32'b00000000000000010110110000111111;
assign LUT_3[13086] = 32'b00000000000000010010001101000110;
assign LUT_3[13087] = 32'b00000000000000011000111000100011;
assign LUT_3[13088] = 32'b00000000000000001011011010000011;
assign LUT_3[13089] = 32'b00000000000000010010000101100000;
assign LUT_3[13090] = 32'b00000000000000001101100001100111;
assign LUT_3[13091] = 32'b00000000000000010100001101000100;
assign LUT_3[13092] = 32'b00000000000000001000100111111001;
assign LUT_3[13093] = 32'b00000000000000001111010011010110;
assign LUT_3[13094] = 32'b00000000000000001010101111011101;
assign LUT_3[13095] = 32'b00000000000000010001011010111010;
assign LUT_3[13096] = 32'b00000000000000010000110011001001;
assign LUT_3[13097] = 32'b00000000000000010111011110100110;
assign LUT_3[13098] = 32'b00000000000000010010111010101101;
assign LUT_3[13099] = 32'b00000000000000011001100110001010;
assign LUT_3[13100] = 32'b00000000000000001110000000111111;
assign LUT_3[13101] = 32'b00000000000000010100101100011100;
assign LUT_3[13102] = 32'b00000000000000010000001000100011;
assign LUT_3[13103] = 32'b00000000000000010110110100000000;
assign LUT_3[13104] = 32'b00000000000000001110101101000110;
assign LUT_3[13105] = 32'b00000000000000010101011000100011;
assign LUT_3[13106] = 32'b00000000000000010000110100101010;
assign LUT_3[13107] = 32'b00000000000000010111100000000111;
assign LUT_3[13108] = 32'b00000000000000001011111010111100;
assign LUT_3[13109] = 32'b00000000000000010010100110011001;
assign LUT_3[13110] = 32'b00000000000000001110000010100000;
assign LUT_3[13111] = 32'b00000000000000010100101101111101;
assign LUT_3[13112] = 32'b00000000000000010100000110001100;
assign LUT_3[13113] = 32'b00000000000000011010110001101001;
assign LUT_3[13114] = 32'b00000000000000010110001101110000;
assign LUT_3[13115] = 32'b00000000000000011100111001001101;
assign LUT_3[13116] = 32'b00000000000000010001010100000010;
assign LUT_3[13117] = 32'b00000000000000010111111111011111;
assign LUT_3[13118] = 32'b00000000000000010011011011100110;
assign LUT_3[13119] = 32'b00000000000000011010000111000011;
assign LUT_3[13120] = 32'b00000000000000001010000100001110;
assign LUT_3[13121] = 32'b00000000000000010000101111101011;
assign LUT_3[13122] = 32'b00000000000000001100001011110010;
assign LUT_3[13123] = 32'b00000000000000010010110111001111;
assign LUT_3[13124] = 32'b00000000000000000111010010000100;
assign LUT_3[13125] = 32'b00000000000000001101111101100001;
assign LUT_3[13126] = 32'b00000000000000001001011001101000;
assign LUT_3[13127] = 32'b00000000000000010000000101000101;
assign LUT_3[13128] = 32'b00000000000000001111011101010100;
assign LUT_3[13129] = 32'b00000000000000010110001000110001;
assign LUT_3[13130] = 32'b00000000000000010001100100111000;
assign LUT_3[13131] = 32'b00000000000000011000010000010101;
assign LUT_3[13132] = 32'b00000000000000001100101011001010;
assign LUT_3[13133] = 32'b00000000000000010011010110100111;
assign LUT_3[13134] = 32'b00000000000000001110110010101110;
assign LUT_3[13135] = 32'b00000000000000010101011110001011;
assign LUT_3[13136] = 32'b00000000000000001101010111010001;
assign LUT_3[13137] = 32'b00000000000000010100000010101110;
assign LUT_3[13138] = 32'b00000000000000001111011110110101;
assign LUT_3[13139] = 32'b00000000000000010110001010010010;
assign LUT_3[13140] = 32'b00000000000000001010100101000111;
assign LUT_3[13141] = 32'b00000000000000010001010000100100;
assign LUT_3[13142] = 32'b00000000000000001100101100101011;
assign LUT_3[13143] = 32'b00000000000000010011011000001000;
assign LUT_3[13144] = 32'b00000000000000010010110000010111;
assign LUT_3[13145] = 32'b00000000000000011001011011110100;
assign LUT_3[13146] = 32'b00000000000000010100110111111011;
assign LUT_3[13147] = 32'b00000000000000011011100011011000;
assign LUT_3[13148] = 32'b00000000000000001111111110001101;
assign LUT_3[13149] = 32'b00000000000000010110101001101010;
assign LUT_3[13150] = 32'b00000000000000010010000101110001;
assign LUT_3[13151] = 32'b00000000000000011000110001001110;
assign LUT_3[13152] = 32'b00000000000000001011010010101110;
assign LUT_3[13153] = 32'b00000000000000010001111110001011;
assign LUT_3[13154] = 32'b00000000000000001101011010010010;
assign LUT_3[13155] = 32'b00000000000000010100000101101111;
assign LUT_3[13156] = 32'b00000000000000001000100000100100;
assign LUT_3[13157] = 32'b00000000000000001111001100000001;
assign LUT_3[13158] = 32'b00000000000000001010101000001000;
assign LUT_3[13159] = 32'b00000000000000010001010011100101;
assign LUT_3[13160] = 32'b00000000000000010000101011110100;
assign LUT_3[13161] = 32'b00000000000000010111010111010001;
assign LUT_3[13162] = 32'b00000000000000010010110011011000;
assign LUT_3[13163] = 32'b00000000000000011001011110110101;
assign LUT_3[13164] = 32'b00000000000000001101111001101010;
assign LUT_3[13165] = 32'b00000000000000010100100101000111;
assign LUT_3[13166] = 32'b00000000000000010000000001001110;
assign LUT_3[13167] = 32'b00000000000000010110101100101011;
assign LUT_3[13168] = 32'b00000000000000001110100101110001;
assign LUT_3[13169] = 32'b00000000000000010101010001001110;
assign LUT_3[13170] = 32'b00000000000000010000101101010101;
assign LUT_3[13171] = 32'b00000000000000010111011000110010;
assign LUT_3[13172] = 32'b00000000000000001011110011100111;
assign LUT_3[13173] = 32'b00000000000000010010011111000100;
assign LUT_3[13174] = 32'b00000000000000001101111011001011;
assign LUT_3[13175] = 32'b00000000000000010100100110101000;
assign LUT_3[13176] = 32'b00000000000000010011111110110111;
assign LUT_3[13177] = 32'b00000000000000011010101010010100;
assign LUT_3[13178] = 32'b00000000000000010110000110011011;
assign LUT_3[13179] = 32'b00000000000000011100110001111000;
assign LUT_3[13180] = 32'b00000000000000010001001100101101;
assign LUT_3[13181] = 32'b00000000000000010111111000001010;
assign LUT_3[13182] = 32'b00000000000000010011010100010001;
assign LUT_3[13183] = 32'b00000000000000011001111111101110;
assign LUT_3[13184] = 32'b00000000000000001100010110100001;
assign LUT_3[13185] = 32'b00000000000000010011000001111110;
assign LUT_3[13186] = 32'b00000000000000001110011110000101;
assign LUT_3[13187] = 32'b00000000000000010101001001100010;
assign LUT_3[13188] = 32'b00000000000000001001100100010111;
assign LUT_3[13189] = 32'b00000000000000010000001111110100;
assign LUT_3[13190] = 32'b00000000000000001011101011111011;
assign LUT_3[13191] = 32'b00000000000000010010010111011000;
assign LUT_3[13192] = 32'b00000000000000010001101111100111;
assign LUT_3[13193] = 32'b00000000000000011000011011000100;
assign LUT_3[13194] = 32'b00000000000000010011110111001011;
assign LUT_3[13195] = 32'b00000000000000011010100010101000;
assign LUT_3[13196] = 32'b00000000000000001110111101011101;
assign LUT_3[13197] = 32'b00000000000000010101101000111010;
assign LUT_3[13198] = 32'b00000000000000010001000101000001;
assign LUT_3[13199] = 32'b00000000000000010111110000011110;
assign LUT_3[13200] = 32'b00000000000000001111101001100100;
assign LUT_3[13201] = 32'b00000000000000010110010101000001;
assign LUT_3[13202] = 32'b00000000000000010001110001001000;
assign LUT_3[13203] = 32'b00000000000000011000011100100101;
assign LUT_3[13204] = 32'b00000000000000001100110111011010;
assign LUT_3[13205] = 32'b00000000000000010011100010110111;
assign LUT_3[13206] = 32'b00000000000000001110111110111110;
assign LUT_3[13207] = 32'b00000000000000010101101010011011;
assign LUT_3[13208] = 32'b00000000000000010101000010101010;
assign LUT_3[13209] = 32'b00000000000000011011101110000111;
assign LUT_3[13210] = 32'b00000000000000010111001010001110;
assign LUT_3[13211] = 32'b00000000000000011101110101101011;
assign LUT_3[13212] = 32'b00000000000000010010010000100000;
assign LUT_3[13213] = 32'b00000000000000011000111011111101;
assign LUT_3[13214] = 32'b00000000000000010100011000000100;
assign LUT_3[13215] = 32'b00000000000000011011000011100001;
assign LUT_3[13216] = 32'b00000000000000001101100101000001;
assign LUT_3[13217] = 32'b00000000000000010100010000011110;
assign LUT_3[13218] = 32'b00000000000000001111101100100101;
assign LUT_3[13219] = 32'b00000000000000010110011000000010;
assign LUT_3[13220] = 32'b00000000000000001010110010110111;
assign LUT_3[13221] = 32'b00000000000000010001011110010100;
assign LUT_3[13222] = 32'b00000000000000001100111010011011;
assign LUT_3[13223] = 32'b00000000000000010011100101111000;
assign LUT_3[13224] = 32'b00000000000000010010111110000111;
assign LUT_3[13225] = 32'b00000000000000011001101001100100;
assign LUT_3[13226] = 32'b00000000000000010101000101101011;
assign LUT_3[13227] = 32'b00000000000000011011110001001000;
assign LUT_3[13228] = 32'b00000000000000010000001011111101;
assign LUT_3[13229] = 32'b00000000000000010110110111011010;
assign LUT_3[13230] = 32'b00000000000000010010010011100001;
assign LUT_3[13231] = 32'b00000000000000011000111110111110;
assign LUT_3[13232] = 32'b00000000000000010000111000000100;
assign LUT_3[13233] = 32'b00000000000000010111100011100001;
assign LUT_3[13234] = 32'b00000000000000010010111111101000;
assign LUT_3[13235] = 32'b00000000000000011001101011000101;
assign LUT_3[13236] = 32'b00000000000000001110000101111010;
assign LUT_3[13237] = 32'b00000000000000010100110001010111;
assign LUT_3[13238] = 32'b00000000000000010000001101011110;
assign LUT_3[13239] = 32'b00000000000000010110111000111011;
assign LUT_3[13240] = 32'b00000000000000010110010001001010;
assign LUT_3[13241] = 32'b00000000000000011100111100100111;
assign LUT_3[13242] = 32'b00000000000000011000011000101110;
assign LUT_3[13243] = 32'b00000000000000011111000100001011;
assign LUT_3[13244] = 32'b00000000000000010011011111000000;
assign LUT_3[13245] = 32'b00000000000000011010001010011101;
assign LUT_3[13246] = 32'b00000000000000010101100110100100;
assign LUT_3[13247] = 32'b00000000000000011100010010000001;
assign LUT_3[13248] = 32'b00000000000000001100001111001100;
assign LUT_3[13249] = 32'b00000000000000010010111010101001;
assign LUT_3[13250] = 32'b00000000000000001110010110110000;
assign LUT_3[13251] = 32'b00000000000000010101000010001101;
assign LUT_3[13252] = 32'b00000000000000001001011101000010;
assign LUT_3[13253] = 32'b00000000000000010000001000011111;
assign LUT_3[13254] = 32'b00000000000000001011100100100110;
assign LUT_3[13255] = 32'b00000000000000010010010000000011;
assign LUT_3[13256] = 32'b00000000000000010001101000010010;
assign LUT_3[13257] = 32'b00000000000000011000010011101111;
assign LUT_3[13258] = 32'b00000000000000010011101111110110;
assign LUT_3[13259] = 32'b00000000000000011010011011010011;
assign LUT_3[13260] = 32'b00000000000000001110110110001000;
assign LUT_3[13261] = 32'b00000000000000010101100001100101;
assign LUT_3[13262] = 32'b00000000000000010000111101101100;
assign LUT_3[13263] = 32'b00000000000000010111101001001001;
assign LUT_3[13264] = 32'b00000000000000001111100010001111;
assign LUT_3[13265] = 32'b00000000000000010110001101101100;
assign LUT_3[13266] = 32'b00000000000000010001101001110011;
assign LUT_3[13267] = 32'b00000000000000011000010101010000;
assign LUT_3[13268] = 32'b00000000000000001100110000000101;
assign LUT_3[13269] = 32'b00000000000000010011011011100010;
assign LUT_3[13270] = 32'b00000000000000001110110111101001;
assign LUT_3[13271] = 32'b00000000000000010101100011000110;
assign LUT_3[13272] = 32'b00000000000000010100111011010101;
assign LUT_3[13273] = 32'b00000000000000011011100110110010;
assign LUT_3[13274] = 32'b00000000000000010111000010111001;
assign LUT_3[13275] = 32'b00000000000000011101101110010110;
assign LUT_3[13276] = 32'b00000000000000010010001001001011;
assign LUT_3[13277] = 32'b00000000000000011000110100101000;
assign LUT_3[13278] = 32'b00000000000000010100010000101111;
assign LUT_3[13279] = 32'b00000000000000011010111100001100;
assign LUT_3[13280] = 32'b00000000000000001101011101101100;
assign LUT_3[13281] = 32'b00000000000000010100001001001001;
assign LUT_3[13282] = 32'b00000000000000001111100101010000;
assign LUT_3[13283] = 32'b00000000000000010110010000101101;
assign LUT_3[13284] = 32'b00000000000000001010101011100010;
assign LUT_3[13285] = 32'b00000000000000010001010110111111;
assign LUT_3[13286] = 32'b00000000000000001100110011000110;
assign LUT_3[13287] = 32'b00000000000000010011011110100011;
assign LUT_3[13288] = 32'b00000000000000010010110110110010;
assign LUT_3[13289] = 32'b00000000000000011001100010001111;
assign LUT_3[13290] = 32'b00000000000000010100111110010110;
assign LUT_3[13291] = 32'b00000000000000011011101001110011;
assign LUT_3[13292] = 32'b00000000000000010000000100101000;
assign LUT_3[13293] = 32'b00000000000000010110110000000101;
assign LUT_3[13294] = 32'b00000000000000010010001100001100;
assign LUT_3[13295] = 32'b00000000000000011000110111101001;
assign LUT_3[13296] = 32'b00000000000000010000110000101111;
assign LUT_3[13297] = 32'b00000000000000010111011100001100;
assign LUT_3[13298] = 32'b00000000000000010010111000010011;
assign LUT_3[13299] = 32'b00000000000000011001100011110000;
assign LUT_3[13300] = 32'b00000000000000001101111110100101;
assign LUT_3[13301] = 32'b00000000000000010100101010000010;
assign LUT_3[13302] = 32'b00000000000000010000000110001001;
assign LUT_3[13303] = 32'b00000000000000010110110001100110;
assign LUT_3[13304] = 32'b00000000000000010110001001110101;
assign LUT_3[13305] = 32'b00000000000000011100110101010010;
assign LUT_3[13306] = 32'b00000000000000011000010001011001;
assign LUT_3[13307] = 32'b00000000000000011110111100110110;
assign LUT_3[13308] = 32'b00000000000000010011010111101011;
assign LUT_3[13309] = 32'b00000000000000011010000011001000;
assign LUT_3[13310] = 32'b00000000000000010101011111001111;
assign LUT_3[13311] = 32'b00000000000000011100001010101100;
assign LUT_3[13312] = 32'b00000000000000010001001011110011;
assign LUT_3[13313] = 32'b00000000000000010111110111010000;
assign LUT_3[13314] = 32'b00000000000000010011010011010111;
assign LUT_3[13315] = 32'b00000000000000011001111110110100;
assign LUT_3[13316] = 32'b00000000000000001110011001101001;
assign LUT_3[13317] = 32'b00000000000000010101000101000110;
assign LUT_3[13318] = 32'b00000000000000010000100001001101;
assign LUT_3[13319] = 32'b00000000000000010111001100101010;
assign LUT_3[13320] = 32'b00000000000000010110100100111001;
assign LUT_3[13321] = 32'b00000000000000011101010000010110;
assign LUT_3[13322] = 32'b00000000000000011000101100011101;
assign LUT_3[13323] = 32'b00000000000000011111010111111010;
assign LUT_3[13324] = 32'b00000000000000010011110010101111;
assign LUT_3[13325] = 32'b00000000000000011010011110001100;
assign LUT_3[13326] = 32'b00000000000000010101111010010011;
assign LUT_3[13327] = 32'b00000000000000011100100101110000;
assign LUT_3[13328] = 32'b00000000000000010100011110110110;
assign LUT_3[13329] = 32'b00000000000000011011001010010011;
assign LUT_3[13330] = 32'b00000000000000010110100110011010;
assign LUT_3[13331] = 32'b00000000000000011101010001110111;
assign LUT_3[13332] = 32'b00000000000000010001101100101100;
assign LUT_3[13333] = 32'b00000000000000011000011000001001;
assign LUT_3[13334] = 32'b00000000000000010011110100010000;
assign LUT_3[13335] = 32'b00000000000000011010011111101101;
assign LUT_3[13336] = 32'b00000000000000011001110111111100;
assign LUT_3[13337] = 32'b00000000000000100000100011011001;
assign LUT_3[13338] = 32'b00000000000000011011111111100000;
assign LUT_3[13339] = 32'b00000000000000100010101010111101;
assign LUT_3[13340] = 32'b00000000000000010111000101110010;
assign LUT_3[13341] = 32'b00000000000000011101110001001111;
assign LUT_3[13342] = 32'b00000000000000011001001101010110;
assign LUT_3[13343] = 32'b00000000000000011111111000110011;
assign LUT_3[13344] = 32'b00000000000000010010011010010011;
assign LUT_3[13345] = 32'b00000000000000011001000101110000;
assign LUT_3[13346] = 32'b00000000000000010100100001110111;
assign LUT_3[13347] = 32'b00000000000000011011001101010100;
assign LUT_3[13348] = 32'b00000000000000001111101000001001;
assign LUT_3[13349] = 32'b00000000000000010110010011100110;
assign LUT_3[13350] = 32'b00000000000000010001101111101101;
assign LUT_3[13351] = 32'b00000000000000011000011011001010;
assign LUT_3[13352] = 32'b00000000000000010111110011011001;
assign LUT_3[13353] = 32'b00000000000000011110011110110110;
assign LUT_3[13354] = 32'b00000000000000011001111010111101;
assign LUT_3[13355] = 32'b00000000000000100000100110011010;
assign LUT_3[13356] = 32'b00000000000000010101000001001111;
assign LUT_3[13357] = 32'b00000000000000011011101100101100;
assign LUT_3[13358] = 32'b00000000000000010111001000110011;
assign LUT_3[13359] = 32'b00000000000000011101110100010000;
assign LUT_3[13360] = 32'b00000000000000010101101101010110;
assign LUT_3[13361] = 32'b00000000000000011100011000110011;
assign LUT_3[13362] = 32'b00000000000000010111110100111010;
assign LUT_3[13363] = 32'b00000000000000011110100000010111;
assign LUT_3[13364] = 32'b00000000000000010010111011001100;
assign LUT_3[13365] = 32'b00000000000000011001100110101001;
assign LUT_3[13366] = 32'b00000000000000010101000010110000;
assign LUT_3[13367] = 32'b00000000000000011011101110001101;
assign LUT_3[13368] = 32'b00000000000000011011000110011100;
assign LUT_3[13369] = 32'b00000000000000100001110001111001;
assign LUT_3[13370] = 32'b00000000000000011101001110000000;
assign LUT_3[13371] = 32'b00000000000000100011111001011101;
assign LUT_3[13372] = 32'b00000000000000011000010100010010;
assign LUT_3[13373] = 32'b00000000000000011110111111101111;
assign LUT_3[13374] = 32'b00000000000000011010011011110110;
assign LUT_3[13375] = 32'b00000000000000100001000111010011;
assign LUT_3[13376] = 32'b00000000000000010001000100011110;
assign LUT_3[13377] = 32'b00000000000000010111101111111011;
assign LUT_3[13378] = 32'b00000000000000010011001100000010;
assign LUT_3[13379] = 32'b00000000000000011001110111011111;
assign LUT_3[13380] = 32'b00000000000000001110010010010100;
assign LUT_3[13381] = 32'b00000000000000010100111101110001;
assign LUT_3[13382] = 32'b00000000000000010000011001111000;
assign LUT_3[13383] = 32'b00000000000000010111000101010101;
assign LUT_3[13384] = 32'b00000000000000010110011101100100;
assign LUT_3[13385] = 32'b00000000000000011101001001000001;
assign LUT_3[13386] = 32'b00000000000000011000100101001000;
assign LUT_3[13387] = 32'b00000000000000011111010000100101;
assign LUT_3[13388] = 32'b00000000000000010011101011011010;
assign LUT_3[13389] = 32'b00000000000000011010010110110111;
assign LUT_3[13390] = 32'b00000000000000010101110010111110;
assign LUT_3[13391] = 32'b00000000000000011100011110011011;
assign LUT_3[13392] = 32'b00000000000000010100010111100001;
assign LUT_3[13393] = 32'b00000000000000011011000010111110;
assign LUT_3[13394] = 32'b00000000000000010110011111000101;
assign LUT_3[13395] = 32'b00000000000000011101001010100010;
assign LUT_3[13396] = 32'b00000000000000010001100101010111;
assign LUT_3[13397] = 32'b00000000000000011000010000110100;
assign LUT_3[13398] = 32'b00000000000000010011101100111011;
assign LUT_3[13399] = 32'b00000000000000011010011000011000;
assign LUT_3[13400] = 32'b00000000000000011001110000100111;
assign LUT_3[13401] = 32'b00000000000000100000011100000100;
assign LUT_3[13402] = 32'b00000000000000011011111000001011;
assign LUT_3[13403] = 32'b00000000000000100010100011101000;
assign LUT_3[13404] = 32'b00000000000000010110111110011101;
assign LUT_3[13405] = 32'b00000000000000011101101001111010;
assign LUT_3[13406] = 32'b00000000000000011001000110000001;
assign LUT_3[13407] = 32'b00000000000000011111110001011110;
assign LUT_3[13408] = 32'b00000000000000010010010010111110;
assign LUT_3[13409] = 32'b00000000000000011000111110011011;
assign LUT_3[13410] = 32'b00000000000000010100011010100010;
assign LUT_3[13411] = 32'b00000000000000011011000101111111;
assign LUT_3[13412] = 32'b00000000000000001111100000110100;
assign LUT_3[13413] = 32'b00000000000000010110001100010001;
assign LUT_3[13414] = 32'b00000000000000010001101000011000;
assign LUT_3[13415] = 32'b00000000000000011000010011110101;
assign LUT_3[13416] = 32'b00000000000000010111101100000100;
assign LUT_3[13417] = 32'b00000000000000011110010111100001;
assign LUT_3[13418] = 32'b00000000000000011001110011101000;
assign LUT_3[13419] = 32'b00000000000000100000011111000101;
assign LUT_3[13420] = 32'b00000000000000010100111001111010;
assign LUT_3[13421] = 32'b00000000000000011011100101010111;
assign LUT_3[13422] = 32'b00000000000000010111000001011110;
assign LUT_3[13423] = 32'b00000000000000011101101100111011;
assign LUT_3[13424] = 32'b00000000000000010101100110000001;
assign LUT_3[13425] = 32'b00000000000000011100010001011110;
assign LUT_3[13426] = 32'b00000000000000010111101101100101;
assign LUT_3[13427] = 32'b00000000000000011110011001000010;
assign LUT_3[13428] = 32'b00000000000000010010110011110111;
assign LUT_3[13429] = 32'b00000000000000011001011111010100;
assign LUT_3[13430] = 32'b00000000000000010100111011011011;
assign LUT_3[13431] = 32'b00000000000000011011100110111000;
assign LUT_3[13432] = 32'b00000000000000011010111111000111;
assign LUT_3[13433] = 32'b00000000000000100001101010100100;
assign LUT_3[13434] = 32'b00000000000000011101000110101011;
assign LUT_3[13435] = 32'b00000000000000100011110010001000;
assign LUT_3[13436] = 32'b00000000000000011000001100111101;
assign LUT_3[13437] = 32'b00000000000000011110111000011010;
assign LUT_3[13438] = 32'b00000000000000011010010100100001;
assign LUT_3[13439] = 32'b00000000000000100000111111111110;
assign LUT_3[13440] = 32'b00000000000000010011010110110001;
assign LUT_3[13441] = 32'b00000000000000011010000010001110;
assign LUT_3[13442] = 32'b00000000000000010101011110010101;
assign LUT_3[13443] = 32'b00000000000000011100001001110010;
assign LUT_3[13444] = 32'b00000000000000010000100100100111;
assign LUT_3[13445] = 32'b00000000000000010111010000000100;
assign LUT_3[13446] = 32'b00000000000000010010101100001011;
assign LUT_3[13447] = 32'b00000000000000011001010111101000;
assign LUT_3[13448] = 32'b00000000000000011000101111110111;
assign LUT_3[13449] = 32'b00000000000000011111011011010100;
assign LUT_3[13450] = 32'b00000000000000011010110111011011;
assign LUT_3[13451] = 32'b00000000000000100001100010111000;
assign LUT_3[13452] = 32'b00000000000000010101111101101101;
assign LUT_3[13453] = 32'b00000000000000011100101001001010;
assign LUT_3[13454] = 32'b00000000000000011000000101010001;
assign LUT_3[13455] = 32'b00000000000000011110110000101110;
assign LUT_3[13456] = 32'b00000000000000010110101001110100;
assign LUT_3[13457] = 32'b00000000000000011101010101010001;
assign LUT_3[13458] = 32'b00000000000000011000110001011000;
assign LUT_3[13459] = 32'b00000000000000011111011100110101;
assign LUT_3[13460] = 32'b00000000000000010011110111101010;
assign LUT_3[13461] = 32'b00000000000000011010100011000111;
assign LUT_3[13462] = 32'b00000000000000010101111111001110;
assign LUT_3[13463] = 32'b00000000000000011100101010101011;
assign LUT_3[13464] = 32'b00000000000000011100000010111010;
assign LUT_3[13465] = 32'b00000000000000100010101110010111;
assign LUT_3[13466] = 32'b00000000000000011110001010011110;
assign LUT_3[13467] = 32'b00000000000000100100110101111011;
assign LUT_3[13468] = 32'b00000000000000011001010000110000;
assign LUT_3[13469] = 32'b00000000000000011111111100001101;
assign LUT_3[13470] = 32'b00000000000000011011011000010100;
assign LUT_3[13471] = 32'b00000000000000100010000011110001;
assign LUT_3[13472] = 32'b00000000000000010100100101010001;
assign LUT_3[13473] = 32'b00000000000000011011010000101110;
assign LUT_3[13474] = 32'b00000000000000010110101100110101;
assign LUT_3[13475] = 32'b00000000000000011101011000010010;
assign LUT_3[13476] = 32'b00000000000000010001110011000111;
assign LUT_3[13477] = 32'b00000000000000011000011110100100;
assign LUT_3[13478] = 32'b00000000000000010011111010101011;
assign LUT_3[13479] = 32'b00000000000000011010100110001000;
assign LUT_3[13480] = 32'b00000000000000011001111110010111;
assign LUT_3[13481] = 32'b00000000000000100000101001110100;
assign LUT_3[13482] = 32'b00000000000000011100000101111011;
assign LUT_3[13483] = 32'b00000000000000100010110001011000;
assign LUT_3[13484] = 32'b00000000000000010111001100001101;
assign LUT_3[13485] = 32'b00000000000000011101110111101010;
assign LUT_3[13486] = 32'b00000000000000011001010011110001;
assign LUT_3[13487] = 32'b00000000000000011111111111001110;
assign LUT_3[13488] = 32'b00000000000000010111111000010100;
assign LUT_3[13489] = 32'b00000000000000011110100011110001;
assign LUT_3[13490] = 32'b00000000000000011001111111111000;
assign LUT_3[13491] = 32'b00000000000000100000101011010101;
assign LUT_3[13492] = 32'b00000000000000010101000110001010;
assign LUT_3[13493] = 32'b00000000000000011011110001100111;
assign LUT_3[13494] = 32'b00000000000000010111001101101110;
assign LUT_3[13495] = 32'b00000000000000011101111001001011;
assign LUT_3[13496] = 32'b00000000000000011101010001011010;
assign LUT_3[13497] = 32'b00000000000000100011111100110111;
assign LUT_3[13498] = 32'b00000000000000011111011000111110;
assign LUT_3[13499] = 32'b00000000000000100110000100011011;
assign LUT_3[13500] = 32'b00000000000000011010011111010000;
assign LUT_3[13501] = 32'b00000000000000100001001010101101;
assign LUT_3[13502] = 32'b00000000000000011100100110110100;
assign LUT_3[13503] = 32'b00000000000000100011010010010001;
assign LUT_3[13504] = 32'b00000000000000010011001111011100;
assign LUT_3[13505] = 32'b00000000000000011001111010111001;
assign LUT_3[13506] = 32'b00000000000000010101010111000000;
assign LUT_3[13507] = 32'b00000000000000011100000010011101;
assign LUT_3[13508] = 32'b00000000000000010000011101010010;
assign LUT_3[13509] = 32'b00000000000000010111001000101111;
assign LUT_3[13510] = 32'b00000000000000010010100100110110;
assign LUT_3[13511] = 32'b00000000000000011001010000010011;
assign LUT_3[13512] = 32'b00000000000000011000101000100010;
assign LUT_3[13513] = 32'b00000000000000011111010011111111;
assign LUT_3[13514] = 32'b00000000000000011010110000000110;
assign LUT_3[13515] = 32'b00000000000000100001011011100011;
assign LUT_3[13516] = 32'b00000000000000010101110110011000;
assign LUT_3[13517] = 32'b00000000000000011100100001110101;
assign LUT_3[13518] = 32'b00000000000000010111111101111100;
assign LUT_3[13519] = 32'b00000000000000011110101001011001;
assign LUT_3[13520] = 32'b00000000000000010110100010011111;
assign LUT_3[13521] = 32'b00000000000000011101001101111100;
assign LUT_3[13522] = 32'b00000000000000011000101010000011;
assign LUT_3[13523] = 32'b00000000000000011111010101100000;
assign LUT_3[13524] = 32'b00000000000000010011110000010101;
assign LUT_3[13525] = 32'b00000000000000011010011011110010;
assign LUT_3[13526] = 32'b00000000000000010101110111111001;
assign LUT_3[13527] = 32'b00000000000000011100100011010110;
assign LUT_3[13528] = 32'b00000000000000011011111011100101;
assign LUT_3[13529] = 32'b00000000000000100010100111000010;
assign LUT_3[13530] = 32'b00000000000000011110000011001001;
assign LUT_3[13531] = 32'b00000000000000100100101110100110;
assign LUT_3[13532] = 32'b00000000000000011001001001011011;
assign LUT_3[13533] = 32'b00000000000000011111110100111000;
assign LUT_3[13534] = 32'b00000000000000011011010000111111;
assign LUT_3[13535] = 32'b00000000000000100001111100011100;
assign LUT_3[13536] = 32'b00000000000000010100011101111100;
assign LUT_3[13537] = 32'b00000000000000011011001001011001;
assign LUT_3[13538] = 32'b00000000000000010110100101100000;
assign LUT_3[13539] = 32'b00000000000000011101010000111101;
assign LUT_3[13540] = 32'b00000000000000010001101011110010;
assign LUT_3[13541] = 32'b00000000000000011000010111001111;
assign LUT_3[13542] = 32'b00000000000000010011110011010110;
assign LUT_3[13543] = 32'b00000000000000011010011110110011;
assign LUT_3[13544] = 32'b00000000000000011001110111000010;
assign LUT_3[13545] = 32'b00000000000000100000100010011111;
assign LUT_3[13546] = 32'b00000000000000011011111110100110;
assign LUT_3[13547] = 32'b00000000000000100010101010000011;
assign LUT_3[13548] = 32'b00000000000000010111000100111000;
assign LUT_3[13549] = 32'b00000000000000011101110000010101;
assign LUT_3[13550] = 32'b00000000000000011001001100011100;
assign LUT_3[13551] = 32'b00000000000000011111110111111001;
assign LUT_3[13552] = 32'b00000000000000010111110000111111;
assign LUT_3[13553] = 32'b00000000000000011110011100011100;
assign LUT_3[13554] = 32'b00000000000000011001111000100011;
assign LUT_3[13555] = 32'b00000000000000100000100100000000;
assign LUT_3[13556] = 32'b00000000000000010100111110110101;
assign LUT_3[13557] = 32'b00000000000000011011101010010010;
assign LUT_3[13558] = 32'b00000000000000010111000110011001;
assign LUT_3[13559] = 32'b00000000000000011101110001110110;
assign LUT_3[13560] = 32'b00000000000000011101001010000101;
assign LUT_3[13561] = 32'b00000000000000100011110101100010;
assign LUT_3[13562] = 32'b00000000000000011111010001101001;
assign LUT_3[13563] = 32'b00000000000000100101111101000110;
assign LUT_3[13564] = 32'b00000000000000011010010111111011;
assign LUT_3[13565] = 32'b00000000000000100001000011011000;
assign LUT_3[13566] = 32'b00000000000000011100011111011111;
assign LUT_3[13567] = 32'b00000000000000100011001010111100;
assign LUT_3[13568] = 32'b00000000000000001101011011010100;
assign LUT_3[13569] = 32'b00000000000000010100000110110001;
assign LUT_3[13570] = 32'b00000000000000001111100010111000;
assign LUT_3[13571] = 32'b00000000000000010110001110010101;
assign LUT_3[13572] = 32'b00000000000000001010101001001010;
assign LUT_3[13573] = 32'b00000000000000010001010100100111;
assign LUT_3[13574] = 32'b00000000000000001100110000101110;
assign LUT_3[13575] = 32'b00000000000000010011011100001011;
assign LUT_3[13576] = 32'b00000000000000010010110100011010;
assign LUT_3[13577] = 32'b00000000000000011001011111110111;
assign LUT_3[13578] = 32'b00000000000000010100111011111110;
assign LUT_3[13579] = 32'b00000000000000011011100111011011;
assign LUT_3[13580] = 32'b00000000000000010000000010010000;
assign LUT_3[13581] = 32'b00000000000000010110101101101101;
assign LUT_3[13582] = 32'b00000000000000010010001001110100;
assign LUT_3[13583] = 32'b00000000000000011000110101010001;
assign LUT_3[13584] = 32'b00000000000000010000101110010111;
assign LUT_3[13585] = 32'b00000000000000010111011001110100;
assign LUT_3[13586] = 32'b00000000000000010010110101111011;
assign LUT_3[13587] = 32'b00000000000000011001100001011000;
assign LUT_3[13588] = 32'b00000000000000001101111100001101;
assign LUT_3[13589] = 32'b00000000000000010100100111101010;
assign LUT_3[13590] = 32'b00000000000000010000000011110001;
assign LUT_3[13591] = 32'b00000000000000010110101111001110;
assign LUT_3[13592] = 32'b00000000000000010110000111011101;
assign LUT_3[13593] = 32'b00000000000000011100110010111010;
assign LUT_3[13594] = 32'b00000000000000011000001111000001;
assign LUT_3[13595] = 32'b00000000000000011110111010011110;
assign LUT_3[13596] = 32'b00000000000000010011010101010011;
assign LUT_3[13597] = 32'b00000000000000011010000000110000;
assign LUT_3[13598] = 32'b00000000000000010101011100110111;
assign LUT_3[13599] = 32'b00000000000000011100001000010100;
assign LUT_3[13600] = 32'b00000000000000001110101001110100;
assign LUT_3[13601] = 32'b00000000000000010101010101010001;
assign LUT_3[13602] = 32'b00000000000000010000110001011000;
assign LUT_3[13603] = 32'b00000000000000010111011100110101;
assign LUT_3[13604] = 32'b00000000000000001011110111101010;
assign LUT_3[13605] = 32'b00000000000000010010100011000111;
assign LUT_3[13606] = 32'b00000000000000001101111111001110;
assign LUT_3[13607] = 32'b00000000000000010100101010101011;
assign LUT_3[13608] = 32'b00000000000000010100000010111010;
assign LUT_3[13609] = 32'b00000000000000011010101110010111;
assign LUT_3[13610] = 32'b00000000000000010110001010011110;
assign LUT_3[13611] = 32'b00000000000000011100110101111011;
assign LUT_3[13612] = 32'b00000000000000010001010000110000;
assign LUT_3[13613] = 32'b00000000000000010111111100001101;
assign LUT_3[13614] = 32'b00000000000000010011011000010100;
assign LUT_3[13615] = 32'b00000000000000011010000011110001;
assign LUT_3[13616] = 32'b00000000000000010001111100110111;
assign LUT_3[13617] = 32'b00000000000000011000101000010100;
assign LUT_3[13618] = 32'b00000000000000010100000100011011;
assign LUT_3[13619] = 32'b00000000000000011010101111111000;
assign LUT_3[13620] = 32'b00000000000000001111001010101101;
assign LUT_3[13621] = 32'b00000000000000010101110110001010;
assign LUT_3[13622] = 32'b00000000000000010001010010010001;
assign LUT_3[13623] = 32'b00000000000000010111111101101110;
assign LUT_3[13624] = 32'b00000000000000010111010101111101;
assign LUT_3[13625] = 32'b00000000000000011110000001011010;
assign LUT_3[13626] = 32'b00000000000000011001011101100001;
assign LUT_3[13627] = 32'b00000000000000100000001000111110;
assign LUT_3[13628] = 32'b00000000000000010100100011110011;
assign LUT_3[13629] = 32'b00000000000000011011001111010000;
assign LUT_3[13630] = 32'b00000000000000010110101011010111;
assign LUT_3[13631] = 32'b00000000000000011101010110110100;
assign LUT_3[13632] = 32'b00000000000000001101010011111111;
assign LUT_3[13633] = 32'b00000000000000010011111111011100;
assign LUT_3[13634] = 32'b00000000000000001111011011100011;
assign LUT_3[13635] = 32'b00000000000000010110000111000000;
assign LUT_3[13636] = 32'b00000000000000001010100001110101;
assign LUT_3[13637] = 32'b00000000000000010001001101010010;
assign LUT_3[13638] = 32'b00000000000000001100101001011001;
assign LUT_3[13639] = 32'b00000000000000010011010100110110;
assign LUT_3[13640] = 32'b00000000000000010010101101000101;
assign LUT_3[13641] = 32'b00000000000000011001011000100010;
assign LUT_3[13642] = 32'b00000000000000010100110100101001;
assign LUT_3[13643] = 32'b00000000000000011011100000000110;
assign LUT_3[13644] = 32'b00000000000000001111111010111011;
assign LUT_3[13645] = 32'b00000000000000010110100110011000;
assign LUT_3[13646] = 32'b00000000000000010010000010011111;
assign LUT_3[13647] = 32'b00000000000000011000101101111100;
assign LUT_3[13648] = 32'b00000000000000010000100111000010;
assign LUT_3[13649] = 32'b00000000000000010111010010011111;
assign LUT_3[13650] = 32'b00000000000000010010101110100110;
assign LUT_3[13651] = 32'b00000000000000011001011010000011;
assign LUT_3[13652] = 32'b00000000000000001101110100111000;
assign LUT_3[13653] = 32'b00000000000000010100100000010101;
assign LUT_3[13654] = 32'b00000000000000001111111100011100;
assign LUT_3[13655] = 32'b00000000000000010110100111111001;
assign LUT_3[13656] = 32'b00000000000000010110000000001000;
assign LUT_3[13657] = 32'b00000000000000011100101011100101;
assign LUT_3[13658] = 32'b00000000000000011000000111101100;
assign LUT_3[13659] = 32'b00000000000000011110110011001001;
assign LUT_3[13660] = 32'b00000000000000010011001101111110;
assign LUT_3[13661] = 32'b00000000000000011001111001011011;
assign LUT_3[13662] = 32'b00000000000000010101010101100010;
assign LUT_3[13663] = 32'b00000000000000011100000000111111;
assign LUT_3[13664] = 32'b00000000000000001110100010011111;
assign LUT_3[13665] = 32'b00000000000000010101001101111100;
assign LUT_3[13666] = 32'b00000000000000010000101010000011;
assign LUT_3[13667] = 32'b00000000000000010111010101100000;
assign LUT_3[13668] = 32'b00000000000000001011110000010101;
assign LUT_3[13669] = 32'b00000000000000010010011011110010;
assign LUT_3[13670] = 32'b00000000000000001101110111111001;
assign LUT_3[13671] = 32'b00000000000000010100100011010110;
assign LUT_3[13672] = 32'b00000000000000010011111011100101;
assign LUT_3[13673] = 32'b00000000000000011010100111000010;
assign LUT_3[13674] = 32'b00000000000000010110000011001001;
assign LUT_3[13675] = 32'b00000000000000011100101110100110;
assign LUT_3[13676] = 32'b00000000000000010001001001011011;
assign LUT_3[13677] = 32'b00000000000000010111110100111000;
assign LUT_3[13678] = 32'b00000000000000010011010000111111;
assign LUT_3[13679] = 32'b00000000000000011001111100011100;
assign LUT_3[13680] = 32'b00000000000000010001110101100010;
assign LUT_3[13681] = 32'b00000000000000011000100000111111;
assign LUT_3[13682] = 32'b00000000000000010011111101000110;
assign LUT_3[13683] = 32'b00000000000000011010101000100011;
assign LUT_3[13684] = 32'b00000000000000001111000011011000;
assign LUT_3[13685] = 32'b00000000000000010101101110110101;
assign LUT_3[13686] = 32'b00000000000000010001001010111100;
assign LUT_3[13687] = 32'b00000000000000010111110110011001;
assign LUT_3[13688] = 32'b00000000000000010111001110101000;
assign LUT_3[13689] = 32'b00000000000000011101111010000101;
assign LUT_3[13690] = 32'b00000000000000011001010110001100;
assign LUT_3[13691] = 32'b00000000000000100000000001101001;
assign LUT_3[13692] = 32'b00000000000000010100011100011110;
assign LUT_3[13693] = 32'b00000000000000011011000111111011;
assign LUT_3[13694] = 32'b00000000000000010110100100000010;
assign LUT_3[13695] = 32'b00000000000000011101001111011111;
assign LUT_3[13696] = 32'b00000000000000001111100110010010;
assign LUT_3[13697] = 32'b00000000000000010110010001101111;
assign LUT_3[13698] = 32'b00000000000000010001101101110110;
assign LUT_3[13699] = 32'b00000000000000011000011001010011;
assign LUT_3[13700] = 32'b00000000000000001100110100001000;
assign LUT_3[13701] = 32'b00000000000000010011011111100101;
assign LUT_3[13702] = 32'b00000000000000001110111011101100;
assign LUT_3[13703] = 32'b00000000000000010101100111001001;
assign LUT_3[13704] = 32'b00000000000000010100111111011000;
assign LUT_3[13705] = 32'b00000000000000011011101010110101;
assign LUT_3[13706] = 32'b00000000000000010111000110111100;
assign LUT_3[13707] = 32'b00000000000000011101110010011001;
assign LUT_3[13708] = 32'b00000000000000010010001101001110;
assign LUT_3[13709] = 32'b00000000000000011000111000101011;
assign LUT_3[13710] = 32'b00000000000000010100010100110010;
assign LUT_3[13711] = 32'b00000000000000011011000000001111;
assign LUT_3[13712] = 32'b00000000000000010010111001010101;
assign LUT_3[13713] = 32'b00000000000000011001100100110010;
assign LUT_3[13714] = 32'b00000000000000010101000000111001;
assign LUT_3[13715] = 32'b00000000000000011011101100010110;
assign LUT_3[13716] = 32'b00000000000000010000000111001011;
assign LUT_3[13717] = 32'b00000000000000010110110010101000;
assign LUT_3[13718] = 32'b00000000000000010010001110101111;
assign LUT_3[13719] = 32'b00000000000000011000111010001100;
assign LUT_3[13720] = 32'b00000000000000011000010010011011;
assign LUT_3[13721] = 32'b00000000000000011110111101111000;
assign LUT_3[13722] = 32'b00000000000000011010011001111111;
assign LUT_3[13723] = 32'b00000000000000100001000101011100;
assign LUT_3[13724] = 32'b00000000000000010101100000010001;
assign LUT_3[13725] = 32'b00000000000000011100001011101110;
assign LUT_3[13726] = 32'b00000000000000010111100111110101;
assign LUT_3[13727] = 32'b00000000000000011110010011010010;
assign LUT_3[13728] = 32'b00000000000000010000110100110010;
assign LUT_3[13729] = 32'b00000000000000010111100000001111;
assign LUT_3[13730] = 32'b00000000000000010010111100010110;
assign LUT_3[13731] = 32'b00000000000000011001100111110011;
assign LUT_3[13732] = 32'b00000000000000001110000010101000;
assign LUT_3[13733] = 32'b00000000000000010100101110000101;
assign LUT_3[13734] = 32'b00000000000000010000001010001100;
assign LUT_3[13735] = 32'b00000000000000010110110101101001;
assign LUT_3[13736] = 32'b00000000000000010110001101111000;
assign LUT_3[13737] = 32'b00000000000000011100111001010101;
assign LUT_3[13738] = 32'b00000000000000011000010101011100;
assign LUT_3[13739] = 32'b00000000000000011111000000111001;
assign LUT_3[13740] = 32'b00000000000000010011011011101110;
assign LUT_3[13741] = 32'b00000000000000011010000111001011;
assign LUT_3[13742] = 32'b00000000000000010101100011010010;
assign LUT_3[13743] = 32'b00000000000000011100001110101111;
assign LUT_3[13744] = 32'b00000000000000010100000111110101;
assign LUT_3[13745] = 32'b00000000000000011010110011010010;
assign LUT_3[13746] = 32'b00000000000000010110001111011001;
assign LUT_3[13747] = 32'b00000000000000011100111010110110;
assign LUT_3[13748] = 32'b00000000000000010001010101101011;
assign LUT_3[13749] = 32'b00000000000000011000000001001000;
assign LUT_3[13750] = 32'b00000000000000010011011101001111;
assign LUT_3[13751] = 32'b00000000000000011010001000101100;
assign LUT_3[13752] = 32'b00000000000000011001100000111011;
assign LUT_3[13753] = 32'b00000000000000100000001100011000;
assign LUT_3[13754] = 32'b00000000000000011011101000011111;
assign LUT_3[13755] = 32'b00000000000000100010010011111100;
assign LUT_3[13756] = 32'b00000000000000010110101110110001;
assign LUT_3[13757] = 32'b00000000000000011101011010001110;
assign LUT_3[13758] = 32'b00000000000000011000110110010101;
assign LUT_3[13759] = 32'b00000000000000011111100001110010;
assign LUT_3[13760] = 32'b00000000000000001111011110111101;
assign LUT_3[13761] = 32'b00000000000000010110001010011010;
assign LUT_3[13762] = 32'b00000000000000010001100110100001;
assign LUT_3[13763] = 32'b00000000000000011000010001111110;
assign LUT_3[13764] = 32'b00000000000000001100101100110011;
assign LUT_3[13765] = 32'b00000000000000010011011000010000;
assign LUT_3[13766] = 32'b00000000000000001110110100010111;
assign LUT_3[13767] = 32'b00000000000000010101011111110100;
assign LUT_3[13768] = 32'b00000000000000010100111000000011;
assign LUT_3[13769] = 32'b00000000000000011011100011100000;
assign LUT_3[13770] = 32'b00000000000000010110111111100111;
assign LUT_3[13771] = 32'b00000000000000011101101011000100;
assign LUT_3[13772] = 32'b00000000000000010010000101111001;
assign LUT_3[13773] = 32'b00000000000000011000110001010110;
assign LUT_3[13774] = 32'b00000000000000010100001101011101;
assign LUT_3[13775] = 32'b00000000000000011010111000111010;
assign LUT_3[13776] = 32'b00000000000000010010110010000000;
assign LUT_3[13777] = 32'b00000000000000011001011101011101;
assign LUT_3[13778] = 32'b00000000000000010100111001100100;
assign LUT_3[13779] = 32'b00000000000000011011100101000001;
assign LUT_3[13780] = 32'b00000000000000001111111111110110;
assign LUT_3[13781] = 32'b00000000000000010110101011010011;
assign LUT_3[13782] = 32'b00000000000000010010000111011010;
assign LUT_3[13783] = 32'b00000000000000011000110010110111;
assign LUT_3[13784] = 32'b00000000000000011000001011000110;
assign LUT_3[13785] = 32'b00000000000000011110110110100011;
assign LUT_3[13786] = 32'b00000000000000011010010010101010;
assign LUT_3[13787] = 32'b00000000000000100000111110000111;
assign LUT_3[13788] = 32'b00000000000000010101011000111100;
assign LUT_3[13789] = 32'b00000000000000011100000100011001;
assign LUT_3[13790] = 32'b00000000000000010111100000100000;
assign LUT_3[13791] = 32'b00000000000000011110001011111101;
assign LUT_3[13792] = 32'b00000000000000010000101101011101;
assign LUT_3[13793] = 32'b00000000000000010111011000111010;
assign LUT_3[13794] = 32'b00000000000000010010110101000001;
assign LUT_3[13795] = 32'b00000000000000011001100000011110;
assign LUT_3[13796] = 32'b00000000000000001101111011010011;
assign LUT_3[13797] = 32'b00000000000000010100100110110000;
assign LUT_3[13798] = 32'b00000000000000010000000010110111;
assign LUT_3[13799] = 32'b00000000000000010110101110010100;
assign LUT_3[13800] = 32'b00000000000000010110000110100011;
assign LUT_3[13801] = 32'b00000000000000011100110010000000;
assign LUT_3[13802] = 32'b00000000000000011000001110000111;
assign LUT_3[13803] = 32'b00000000000000011110111001100100;
assign LUT_3[13804] = 32'b00000000000000010011010100011001;
assign LUT_3[13805] = 32'b00000000000000011001111111110110;
assign LUT_3[13806] = 32'b00000000000000010101011011111101;
assign LUT_3[13807] = 32'b00000000000000011100000111011010;
assign LUT_3[13808] = 32'b00000000000000010100000000100000;
assign LUT_3[13809] = 32'b00000000000000011010101011111101;
assign LUT_3[13810] = 32'b00000000000000010110001000000100;
assign LUT_3[13811] = 32'b00000000000000011100110011100001;
assign LUT_3[13812] = 32'b00000000000000010001001110010110;
assign LUT_3[13813] = 32'b00000000000000010111111001110011;
assign LUT_3[13814] = 32'b00000000000000010011010101111010;
assign LUT_3[13815] = 32'b00000000000000011010000001010111;
assign LUT_3[13816] = 32'b00000000000000011001011001100110;
assign LUT_3[13817] = 32'b00000000000000100000000101000011;
assign LUT_3[13818] = 32'b00000000000000011011100001001010;
assign LUT_3[13819] = 32'b00000000000000100010001100100111;
assign LUT_3[13820] = 32'b00000000000000010110100111011100;
assign LUT_3[13821] = 32'b00000000000000011101010010111001;
assign LUT_3[13822] = 32'b00000000000000011000101111000000;
assign LUT_3[13823] = 32'b00000000000000011111011010011101;
assign LUT_3[13824] = 32'b00000000000000010100100000111111;
assign LUT_3[13825] = 32'b00000000000000011011001100011100;
assign LUT_3[13826] = 32'b00000000000000010110101000100011;
assign LUT_3[13827] = 32'b00000000000000011101010100000000;
assign LUT_3[13828] = 32'b00000000000000010001101110110101;
assign LUT_3[13829] = 32'b00000000000000011000011010010010;
assign LUT_3[13830] = 32'b00000000000000010011110110011001;
assign LUT_3[13831] = 32'b00000000000000011010100001110110;
assign LUT_3[13832] = 32'b00000000000000011001111010000101;
assign LUT_3[13833] = 32'b00000000000000100000100101100010;
assign LUT_3[13834] = 32'b00000000000000011100000001101001;
assign LUT_3[13835] = 32'b00000000000000100010101101000110;
assign LUT_3[13836] = 32'b00000000000000010111000111111011;
assign LUT_3[13837] = 32'b00000000000000011101110011011000;
assign LUT_3[13838] = 32'b00000000000000011001001111011111;
assign LUT_3[13839] = 32'b00000000000000011111111010111100;
assign LUT_3[13840] = 32'b00000000000000010111110100000010;
assign LUT_3[13841] = 32'b00000000000000011110011111011111;
assign LUT_3[13842] = 32'b00000000000000011001111011100110;
assign LUT_3[13843] = 32'b00000000000000100000100111000011;
assign LUT_3[13844] = 32'b00000000000000010101000001111000;
assign LUT_3[13845] = 32'b00000000000000011011101101010101;
assign LUT_3[13846] = 32'b00000000000000010111001001011100;
assign LUT_3[13847] = 32'b00000000000000011101110100111001;
assign LUT_3[13848] = 32'b00000000000000011101001101001000;
assign LUT_3[13849] = 32'b00000000000000100011111000100101;
assign LUT_3[13850] = 32'b00000000000000011111010100101100;
assign LUT_3[13851] = 32'b00000000000000100110000000001001;
assign LUT_3[13852] = 32'b00000000000000011010011010111110;
assign LUT_3[13853] = 32'b00000000000000100001000110011011;
assign LUT_3[13854] = 32'b00000000000000011100100010100010;
assign LUT_3[13855] = 32'b00000000000000100011001101111111;
assign LUT_3[13856] = 32'b00000000000000010101101111011111;
assign LUT_3[13857] = 32'b00000000000000011100011010111100;
assign LUT_3[13858] = 32'b00000000000000010111110111000011;
assign LUT_3[13859] = 32'b00000000000000011110100010100000;
assign LUT_3[13860] = 32'b00000000000000010010111101010101;
assign LUT_3[13861] = 32'b00000000000000011001101000110010;
assign LUT_3[13862] = 32'b00000000000000010101000100111001;
assign LUT_3[13863] = 32'b00000000000000011011110000010110;
assign LUT_3[13864] = 32'b00000000000000011011001000100101;
assign LUT_3[13865] = 32'b00000000000000100001110100000010;
assign LUT_3[13866] = 32'b00000000000000011101010000001001;
assign LUT_3[13867] = 32'b00000000000000100011111011100110;
assign LUT_3[13868] = 32'b00000000000000011000010110011011;
assign LUT_3[13869] = 32'b00000000000000011111000001111000;
assign LUT_3[13870] = 32'b00000000000000011010011101111111;
assign LUT_3[13871] = 32'b00000000000000100001001001011100;
assign LUT_3[13872] = 32'b00000000000000011001000010100010;
assign LUT_3[13873] = 32'b00000000000000011111101101111111;
assign LUT_3[13874] = 32'b00000000000000011011001010000110;
assign LUT_3[13875] = 32'b00000000000000100001110101100011;
assign LUT_3[13876] = 32'b00000000000000010110010000011000;
assign LUT_3[13877] = 32'b00000000000000011100111011110101;
assign LUT_3[13878] = 32'b00000000000000011000010111111100;
assign LUT_3[13879] = 32'b00000000000000011111000011011001;
assign LUT_3[13880] = 32'b00000000000000011110011011101000;
assign LUT_3[13881] = 32'b00000000000000100101000111000101;
assign LUT_3[13882] = 32'b00000000000000100000100011001100;
assign LUT_3[13883] = 32'b00000000000000100111001110101001;
assign LUT_3[13884] = 32'b00000000000000011011101001011110;
assign LUT_3[13885] = 32'b00000000000000100010010100111011;
assign LUT_3[13886] = 32'b00000000000000011101110001000010;
assign LUT_3[13887] = 32'b00000000000000100100011100011111;
assign LUT_3[13888] = 32'b00000000000000010100011001101010;
assign LUT_3[13889] = 32'b00000000000000011011000101000111;
assign LUT_3[13890] = 32'b00000000000000010110100001001110;
assign LUT_3[13891] = 32'b00000000000000011101001100101011;
assign LUT_3[13892] = 32'b00000000000000010001100111100000;
assign LUT_3[13893] = 32'b00000000000000011000010010111101;
assign LUT_3[13894] = 32'b00000000000000010011101111000100;
assign LUT_3[13895] = 32'b00000000000000011010011010100001;
assign LUT_3[13896] = 32'b00000000000000011001110010110000;
assign LUT_3[13897] = 32'b00000000000000100000011110001101;
assign LUT_3[13898] = 32'b00000000000000011011111010010100;
assign LUT_3[13899] = 32'b00000000000000100010100101110001;
assign LUT_3[13900] = 32'b00000000000000010111000000100110;
assign LUT_3[13901] = 32'b00000000000000011101101100000011;
assign LUT_3[13902] = 32'b00000000000000011001001000001010;
assign LUT_3[13903] = 32'b00000000000000011111110011100111;
assign LUT_3[13904] = 32'b00000000000000010111101100101101;
assign LUT_3[13905] = 32'b00000000000000011110011000001010;
assign LUT_3[13906] = 32'b00000000000000011001110100010001;
assign LUT_3[13907] = 32'b00000000000000100000011111101110;
assign LUT_3[13908] = 32'b00000000000000010100111010100011;
assign LUT_3[13909] = 32'b00000000000000011011100110000000;
assign LUT_3[13910] = 32'b00000000000000010111000010000111;
assign LUT_3[13911] = 32'b00000000000000011101101101100100;
assign LUT_3[13912] = 32'b00000000000000011101000101110011;
assign LUT_3[13913] = 32'b00000000000000100011110001010000;
assign LUT_3[13914] = 32'b00000000000000011111001101010111;
assign LUT_3[13915] = 32'b00000000000000100101111000110100;
assign LUT_3[13916] = 32'b00000000000000011010010011101001;
assign LUT_3[13917] = 32'b00000000000000100000111111000110;
assign LUT_3[13918] = 32'b00000000000000011100011011001101;
assign LUT_3[13919] = 32'b00000000000000100011000110101010;
assign LUT_3[13920] = 32'b00000000000000010101101000001010;
assign LUT_3[13921] = 32'b00000000000000011100010011100111;
assign LUT_3[13922] = 32'b00000000000000010111101111101110;
assign LUT_3[13923] = 32'b00000000000000011110011011001011;
assign LUT_3[13924] = 32'b00000000000000010010110110000000;
assign LUT_3[13925] = 32'b00000000000000011001100001011101;
assign LUT_3[13926] = 32'b00000000000000010100111101100100;
assign LUT_3[13927] = 32'b00000000000000011011101001000001;
assign LUT_3[13928] = 32'b00000000000000011011000001010000;
assign LUT_3[13929] = 32'b00000000000000100001101100101101;
assign LUT_3[13930] = 32'b00000000000000011101001000110100;
assign LUT_3[13931] = 32'b00000000000000100011110100010001;
assign LUT_3[13932] = 32'b00000000000000011000001111000110;
assign LUT_3[13933] = 32'b00000000000000011110111010100011;
assign LUT_3[13934] = 32'b00000000000000011010010110101010;
assign LUT_3[13935] = 32'b00000000000000100001000010000111;
assign LUT_3[13936] = 32'b00000000000000011000111011001101;
assign LUT_3[13937] = 32'b00000000000000011111100110101010;
assign LUT_3[13938] = 32'b00000000000000011011000010110001;
assign LUT_3[13939] = 32'b00000000000000100001101110001110;
assign LUT_3[13940] = 32'b00000000000000010110001001000011;
assign LUT_3[13941] = 32'b00000000000000011100110100100000;
assign LUT_3[13942] = 32'b00000000000000011000010000100111;
assign LUT_3[13943] = 32'b00000000000000011110111100000100;
assign LUT_3[13944] = 32'b00000000000000011110010100010011;
assign LUT_3[13945] = 32'b00000000000000100100111111110000;
assign LUT_3[13946] = 32'b00000000000000100000011011110111;
assign LUT_3[13947] = 32'b00000000000000100111000111010100;
assign LUT_3[13948] = 32'b00000000000000011011100010001001;
assign LUT_3[13949] = 32'b00000000000000100010001101100110;
assign LUT_3[13950] = 32'b00000000000000011101101001101101;
assign LUT_3[13951] = 32'b00000000000000100100010101001010;
assign LUT_3[13952] = 32'b00000000000000010110101011111101;
assign LUT_3[13953] = 32'b00000000000000011101010111011010;
assign LUT_3[13954] = 32'b00000000000000011000110011100001;
assign LUT_3[13955] = 32'b00000000000000011111011110111110;
assign LUT_3[13956] = 32'b00000000000000010011111001110011;
assign LUT_3[13957] = 32'b00000000000000011010100101010000;
assign LUT_3[13958] = 32'b00000000000000010110000001010111;
assign LUT_3[13959] = 32'b00000000000000011100101100110100;
assign LUT_3[13960] = 32'b00000000000000011100000101000011;
assign LUT_3[13961] = 32'b00000000000000100010110000100000;
assign LUT_3[13962] = 32'b00000000000000011110001100100111;
assign LUT_3[13963] = 32'b00000000000000100100111000000100;
assign LUT_3[13964] = 32'b00000000000000011001010010111001;
assign LUT_3[13965] = 32'b00000000000000011111111110010110;
assign LUT_3[13966] = 32'b00000000000000011011011010011101;
assign LUT_3[13967] = 32'b00000000000000100010000101111010;
assign LUT_3[13968] = 32'b00000000000000011001111111000000;
assign LUT_3[13969] = 32'b00000000000000100000101010011101;
assign LUT_3[13970] = 32'b00000000000000011100000110100100;
assign LUT_3[13971] = 32'b00000000000000100010110010000001;
assign LUT_3[13972] = 32'b00000000000000010111001100110110;
assign LUT_3[13973] = 32'b00000000000000011101111000010011;
assign LUT_3[13974] = 32'b00000000000000011001010100011010;
assign LUT_3[13975] = 32'b00000000000000011111111111110111;
assign LUT_3[13976] = 32'b00000000000000011111011000000110;
assign LUT_3[13977] = 32'b00000000000000100110000011100011;
assign LUT_3[13978] = 32'b00000000000000100001011111101010;
assign LUT_3[13979] = 32'b00000000000000101000001011000111;
assign LUT_3[13980] = 32'b00000000000000011100100101111100;
assign LUT_3[13981] = 32'b00000000000000100011010001011001;
assign LUT_3[13982] = 32'b00000000000000011110101101100000;
assign LUT_3[13983] = 32'b00000000000000100101011000111101;
assign LUT_3[13984] = 32'b00000000000000010111111010011101;
assign LUT_3[13985] = 32'b00000000000000011110100101111010;
assign LUT_3[13986] = 32'b00000000000000011010000010000001;
assign LUT_3[13987] = 32'b00000000000000100000101101011110;
assign LUT_3[13988] = 32'b00000000000000010101001000010011;
assign LUT_3[13989] = 32'b00000000000000011011110011110000;
assign LUT_3[13990] = 32'b00000000000000010111001111110111;
assign LUT_3[13991] = 32'b00000000000000011101111011010100;
assign LUT_3[13992] = 32'b00000000000000011101010011100011;
assign LUT_3[13993] = 32'b00000000000000100011111111000000;
assign LUT_3[13994] = 32'b00000000000000011111011011000111;
assign LUT_3[13995] = 32'b00000000000000100110000110100100;
assign LUT_3[13996] = 32'b00000000000000011010100001011001;
assign LUT_3[13997] = 32'b00000000000000100001001100110110;
assign LUT_3[13998] = 32'b00000000000000011100101000111101;
assign LUT_3[13999] = 32'b00000000000000100011010100011010;
assign LUT_3[14000] = 32'b00000000000000011011001101100000;
assign LUT_3[14001] = 32'b00000000000000100001111000111101;
assign LUT_3[14002] = 32'b00000000000000011101010101000100;
assign LUT_3[14003] = 32'b00000000000000100100000000100001;
assign LUT_3[14004] = 32'b00000000000000011000011011010110;
assign LUT_3[14005] = 32'b00000000000000011111000110110011;
assign LUT_3[14006] = 32'b00000000000000011010100010111010;
assign LUT_3[14007] = 32'b00000000000000100001001110010111;
assign LUT_3[14008] = 32'b00000000000000100000100110100110;
assign LUT_3[14009] = 32'b00000000000000100111010010000011;
assign LUT_3[14010] = 32'b00000000000000100010101110001010;
assign LUT_3[14011] = 32'b00000000000000101001011001100111;
assign LUT_3[14012] = 32'b00000000000000011101110100011100;
assign LUT_3[14013] = 32'b00000000000000100100011111111001;
assign LUT_3[14014] = 32'b00000000000000011111111100000000;
assign LUT_3[14015] = 32'b00000000000000100110100111011101;
assign LUT_3[14016] = 32'b00000000000000010110100100101000;
assign LUT_3[14017] = 32'b00000000000000011101010000000101;
assign LUT_3[14018] = 32'b00000000000000011000101100001100;
assign LUT_3[14019] = 32'b00000000000000011111010111101001;
assign LUT_3[14020] = 32'b00000000000000010011110010011110;
assign LUT_3[14021] = 32'b00000000000000011010011101111011;
assign LUT_3[14022] = 32'b00000000000000010101111010000010;
assign LUT_3[14023] = 32'b00000000000000011100100101011111;
assign LUT_3[14024] = 32'b00000000000000011011111101101110;
assign LUT_3[14025] = 32'b00000000000000100010101001001011;
assign LUT_3[14026] = 32'b00000000000000011110000101010010;
assign LUT_3[14027] = 32'b00000000000000100100110000101111;
assign LUT_3[14028] = 32'b00000000000000011001001011100100;
assign LUT_3[14029] = 32'b00000000000000011111110111000001;
assign LUT_3[14030] = 32'b00000000000000011011010011001000;
assign LUT_3[14031] = 32'b00000000000000100001111110100101;
assign LUT_3[14032] = 32'b00000000000000011001110111101011;
assign LUT_3[14033] = 32'b00000000000000100000100011001000;
assign LUT_3[14034] = 32'b00000000000000011011111111001111;
assign LUT_3[14035] = 32'b00000000000000100010101010101100;
assign LUT_3[14036] = 32'b00000000000000010111000101100001;
assign LUT_3[14037] = 32'b00000000000000011101110000111110;
assign LUT_3[14038] = 32'b00000000000000011001001101000101;
assign LUT_3[14039] = 32'b00000000000000011111111000100010;
assign LUT_3[14040] = 32'b00000000000000011111010000110001;
assign LUT_3[14041] = 32'b00000000000000100101111100001110;
assign LUT_3[14042] = 32'b00000000000000100001011000010101;
assign LUT_3[14043] = 32'b00000000000000101000000011110010;
assign LUT_3[14044] = 32'b00000000000000011100011110100111;
assign LUT_3[14045] = 32'b00000000000000100011001010000100;
assign LUT_3[14046] = 32'b00000000000000011110100110001011;
assign LUT_3[14047] = 32'b00000000000000100101010001101000;
assign LUT_3[14048] = 32'b00000000000000010111110011001000;
assign LUT_3[14049] = 32'b00000000000000011110011110100101;
assign LUT_3[14050] = 32'b00000000000000011001111010101100;
assign LUT_3[14051] = 32'b00000000000000100000100110001001;
assign LUT_3[14052] = 32'b00000000000000010101000000111110;
assign LUT_3[14053] = 32'b00000000000000011011101100011011;
assign LUT_3[14054] = 32'b00000000000000010111001000100010;
assign LUT_3[14055] = 32'b00000000000000011101110011111111;
assign LUT_3[14056] = 32'b00000000000000011101001100001110;
assign LUT_3[14057] = 32'b00000000000000100011110111101011;
assign LUT_3[14058] = 32'b00000000000000011111010011110010;
assign LUT_3[14059] = 32'b00000000000000100101111111001111;
assign LUT_3[14060] = 32'b00000000000000011010011010000100;
assign LUT_3[14061] = 32'b00000000000000100001000101100001;
assign LUT_3[14062] = 32'b00000000000000011100100001101000;
assign LUT_3[14063] = 32'b00000000000000100011001101000101;
assign LUT_3[14064] = 32'b00000000000000011011000110001011;
assign LUT_3[14065] = 32'b00000000000000100001110001101000;
assign LUT_3[14066] = 32'b00000000000000011101001101101111;
assign LUT_3[14067] = 32'b00000000000000100011111001001100;
assign LUT_3[14068] = 32'b00000000000000011000010100000001;
assign LUT_3[14069] = 32'b00000000000000011110111111011110;
assign LUT_3[14070] = 32'b00000000000000011010011011100101;
assign LUT_3[14071] = 32'b00000000000000100001000111000010;
assign LUT_3[14072] = 32'b00000000000000100000011111010001;
assign LUT_3[14073] = 32'b00000000000000100111001010101110;
assign LUT_3[14074] = 32'b00000000000000100010100110110101;
assign LUT_3[14075] = 32'b00000000000000101001010010010010;
assign LUT_3[14076] = 32'b00000000000000011101101101000111;
assign LUT_3[14077] = 32'b00000000000000100100011000100100;
assign LUT_3[14078] = 32'b00000000000000011111110100101011;
assign LUT_3[14079] = 32'b00000000000000100110100000001000;
assign LUT_3[14080] = 32'b00000000000000010000110000100000;
assign LUT_3[14081] = 32'b00000000000000010111011011111101;
assign LUT_3[14082] = 32'b00000000000000010010111000000100;
assign LUT_3[14083] = 32'b00000000000000011001100011100001;
assign LUT_3[14084] = 32'b00000000000000001101111110010110;
assign LUT_3[14085] = 32'b00000000000000010100101001110011;
assign LUT_3[14086] = 32'b00000000000000010000000101111010;
assign LUT_3[14087] = 32'b00000000000000010110110001010111;
assign LUT_3[14088] = 32'b00000000000000010110001001100110;
assign LUT_3[14089] = 32'b00000000000000011100110101000011;
assign LUT_3[14090] = 32'b00000000000000011000010001001010;
assign LUT_3[14091] = 32'b00000000000000011110111100100111;
assign LUT_3[14092] = 32'b00000000000000010011010111011100;
assign LUT_3[14093] = 32'b00000000000000011010000010111001;
assign LUT_3[14094] = 32'b00000000000000010101011111000000;
assign LUT_3[14095] = 32'b00000000000000011100001010011101;
assign LUT_3[14096] = 32'b00000000000000010100000011100011;
assign LUT_3[14097] = 32'b00000000000000011010101111000000;
assign LUT_3[14098] = 32'b00000000000000010110001011000111;
assign LUT_3[14099] = 32'b00000000000000011100110110100100;
assign LUT_3[14100] = 32'b00000000000000010001010001011001;
assign LUT_3[14101] = 32'b00000000000000010111111100110110;
assign LUT_3[14102] = 32'b00000000000000010011011000111101;
assign LUT_3[14103] = 32'b00000000000000011010000100011010;
assign LUT_3[14104] = 32'b00000000000000011001011100101001;
assign LUT_3[14105] = 32'b00000000000000100000001000000110;
assign LUT_3[14106] = 32'b00000000000000011011100100001101;
assign LUT_3[14107] = 32'b00000000000000100010001111101010;
assign LUT_3[14108] = 32'b00000000000000010110101010011111;
assign LUT_3[14109] = 32'b00000000000000011101010101111100;
assign LUT_3[14110] = 32'b00000000000000011000110010000011;
assign LUT_3[14111] = 32'b00000000000000011111011101100000;
assign LUT_3[14112] = 32'b00000000000000010001111111000000;
assign LUT_3[14113] = 32'b00000000000000011000101010011101;
assign LUT_3[14114] = 32'b00000000000000010100000110100100;
assign LUT_3[14115] = 32'b00000000000000011010110010000001;
assign LUT_3[14116] = 32'b00000000000000001111001100110110;
assign LUT_3[14117] = 32'b00000000000000010101111000010011;
assign LUT_3[14118] = 32'b00000000000000010001010100011010;
assign LUT_3[14119] = 32'b00000000000000010111111111110111;
assign LUT_3[14120] = 32'b00000000000000010111011000000110;
assign LUT_3[14121] = 32'b00000000000000011110000011100011;
assign LUT_3[14122] = 32'b00000000000000011001011111101010;
assign LUT_3[14123] = 32'b00000000000000100000001011000111;
assign LUT_3[14124] = 32'b00000000000000010100100101111100;
assign LUT_3[14125] = 32'b00000000000000011011010001011001;
assign LUT_3[14126] = 32'b00000000000000010110101101100000;
assign LUT_3[14127] = 32'b00000000000000011101011000111101;
assign LUT_3[14128] = 32'b00000000000000010101010010000011;
assign LUT_3[14129] = 32'b00000000000000011011111101100000;
assign LUT_3[14130] = 32'b00000000000000010111011001100111;
assign LUT_3[14131] = 32'b00000000000000011110000101000100;
assign LUT_3[14132] = 32'b00000000000000010010011111111001;
assign LUT_3[14133] = 32'b00000000000000011001001011010110;
assign LUT_3[14134] = 32'b00000000000000010100100111011101;
assign LUT_3[14135] = 32'b00000000000000011011010010111010;
assign LUT_3[14136] = 32'b00000000000000011010101011001001;
assign LUT_3[14137] = 32'b00000000000000100001010110100110;
assign LUT_3[14138] = 32'b00000000000000011100110010101101;
assign LUT_3[14139] = 32'b00000000000000100011011110001010;
assign LUT_3[14140] = 32'b00000000000000010111111000111111;
assign LUT_3[14141] = 32'b00000000000000011110100100011100;
assign LUT_3[14142] = 32'b00000000000000011010000000100011;
assign LUT_3[14143] = 32'b00000000000000100000101100000000;
assign LUT_3[14144] = 32'b00000000000000010000101001001011;
assign LUT_3[14145] = 32'b00000000000000010111010100101000;
assign LUT_3[14146] = 32'b00000000000000010010110000101111;
assign LUT_3[14147] = 32'b00000000000000011001011100001100;
assign LUT_3[14148] = 32'b00000000000000001101110111000001;
assign LUT_3[14149] = 32'b00000000000000010100100010011110;
assign LUT_3[14150] = 32'b00000000000000001111111110100101;
assign LUT_3[14151] = 32'b00000000000000010110101010000010;
assign LUT_3[14152] = 32'b00000000000000010110000010010001;
assign LUT_3[14153] = 32'b00000000000000011100101101101110;
assign LUT_3[14154] = 32'b00000000000000011000001001110101;
assign LUT_3[14155] = 32'b00000000000000011110110101010010;
assign LUT_3[14156] = 32'b00000000000000010011010000000111;
assign LUT_3[14157] = 32'b00000000000000011001111011100100;
assign LUT_3[14158] = 32'b00000000000000010101010111101011;
assign LUT_3[14159] = 32'b00000000000000011100000011001000;
assign LUT_3[14160] = 32'b00000000000000010011111100001110;
assign LUT_3[14161] = 32'b00000000000000011010100111101011;
assign LUT_3[14162] = 32'b00000000000000010110000011110010;
assign LUT_3[14163] = 32'b00000000000000011100101111001111;
assign LUT_3[14164] = 32'b00000000000000010001001010000100;
assign LUT_3[14165] = 32'b00000000000000010111110101100001;
assign LUT_3[14166] = 32'b00000000000000010011010001101000;
assign LUT_3[14167] = 32'b00000000000000011001111101000101;
assign LUT_3[14168] = 32'b00000000000000011001010101010100;
assign LUT_3[14169] = 32'b00000000000000100000000000110001;
assign LUT_3[14170] = 32'b00000000000000011011011100111000;
assign LUT_3[14171] = 32'b00000000000000100010001000010101;
assign LUT_3[14172] = 32'b00000000000000010110100011001010;
assign LUT_3[14173] = 32'b00000000000000011101001110100111;
assign LUT_3[14174] = 32'b00000000000000011000101010101110;
assign LUT_3[14175] = 32'b00000000000000011111010110001011;
assign LUT_3[14176] = 32'b00000000000000010001110111101011;
assign LUT_3[14177] = 32'b00000000000000011000100011001000;
assign LUT_3[14178] = 32'b00000000000000010011111111001111;
assign LUT_3[14179] = 32'b00000000000000011010101010101100;
assign LUT_3[14180] = 32'b00000000000000001111000101100001;
assign LUT_3[14181] = 32'b00000000000000010101110000111110;
assign LUT_3[14182] = 32'b00000000000000010001001101000101;
assign LUT_3[14183] = 32'b00000000000000010111111000100010;
assign LUT_3[14184] = 32'b00000000000000010111010000110001;
assign LUT_3[14185] = 32'b00000000000000011101111100001110;
assign LUT_3[14186] = 32'b00000000000000011001011000010101;
assign LUT_3[14187] = 32'b00000000000000100000000011110010;
assign LUT_3[14188] = 32'b00000000000000010100011110100111;
assign LUT_3[14189] = 32'b00000000000000011011001010000100;
assign LUT_3[14190] = 32'b00000000000000010110100110001011;
assign LUT_3[14191] = 32'b00000000000000011101010001101000;
assign LUT_3[14192] = 32'b00000000000000010101001010101110;
assign LUT_3[14193] = 32'b00000000000000011011110110001011;
assign LUT_3[14194] = 32'b00000000000000010111010010010010;
assign LUT_3[14195] = 32'b00000000000000011101111101101111;
assign LUT_3[14196] = 32'b00000000000000010010011000100100;
assign LUT_3[14197] = 32'b00000000000000011001000100000001;
assign LUT_3[14198] = 32'b00000000000000010100100000001000;
assign LUT_3[14199] = 32'b00000000000000011011001011100101;
assign LUT_3[14200] = 32'b00000000000000011010100011110100;
assign LUT_3[14201] = 32'b00000000000000100001001111010001;
assign LUT_3[14202] = 32'b00000000000000011100101011011000;
assign LUT_3[14203] = 32'b00000000000000100011010110110101;
assign LUT_3[14204] = 32'b00000000000000010111110001101010;
assign LUT_3[14205] = 32'b00000000000000011110011101000111;
assign LUT_3[14206] = 32'b00000000000000011001111001001110;
assign LUT_3[14207] = 32'b00000000000000100000100100101011;
assign LUT_3[14208] = 32'b00000000000000010010111011011110;
assign LUT_3[14209] = 32'b00000000000000011001100110111011;
assign LUT_3[14210] = 32'b00000000000000010101000011000010;
assign LUT_3[14211] = 32'b00000000000000011011101110011111;
assign LUT_3[14212] = 32'b00000000000000010000001001010100;
assign LUT_3[14213] = 32'b00000000000000010110110100110001;
assign LUT_3[14214] = 32'b00000000000000010010010000111000;
assign LUT_3[14215] = 32'b00000000000000011000111100010101;
assign LUT_3[14216] = 32'b00000000000000011000010100100100;
assign LUT_3[14217] = 32'b00000000000000011111000000000001;
assign LUT_3[14218] = 32'b00000000000000011010011100001000;
assign LUT_3[14219] = 32'b00000000000000100001000111100101;
assign LUT_3[14220] = 32'b00000000000000010101100010011010;
assign LUT_3[14221] = 32'b00000000000000011100001101110111;
assign LUT_3[14222] = 32'b00000000000000010111101001111110;
assign LUT_3[14223] = 32'b00000000000000011110010101011011;
assign LUT_3[14224] = 32'b00000000000000010110001110100001;
assign LUT_3[14225] = 32'b00000000000000011100111001111110;
assign LUT_3[14226] = 32'b00000000000000011000010110000101;
assign LUT_3[14227] = 32'b00000000000000011111000001100010;
assign LUT_3[14228] = 32'b00000000000000010011011100010111;
assign LUT_3[14229] = 32'b00000000000000011010000111110100;
assign LUT_3[14230] = 32'b00000000000000010101100011111011;
assign LUT_3[14231] = 32'b00000000000000011100001111011000;
assign LUT_3[14232] = 32'b00000000000000011011100111100111;
assign LUT_3[14233] = 32'b00000000000000100010010011000100;
assign LUT_3[14234] = 32'b00000000000000011101101111001011;
assign LUT_3[14235] = 32'b00000000000000100100011010101000;
assign LUT_3[14236] = 32'b00000000000000011000110101011101;
assign LUT_3[14237] = 32'b00000000000000011111100000111010;
assign LUT_3[14238] = 32'b00000000000000011010111101000001;
assign LUT_3[14239] = 32'b00000000000000100001101000011110;
assign LUT_3[14240] = 32'b00000000000000010100001001111110;
assign LUT_3[14241] = 32'b00000000000000011010110101011011;
assign LUT_3[14242] = 32'b00000000000000010110010001100010;
assign LUT_3[14243] = 32'b00000000000000011100111100111111;
assign LUT_3[14244] = 32'b00000000000000010001010111110100;
assign LUT_3[14245] = 32'b00000000000000011000000011010001;
assign LUT_3[14246] = 32'b00000000000000010011011111011000;
assign LUT_3[14247] = 32'b00000000000000011010001010110101;
assign LUT_3[14248] = 32'b00000000000000011001100011000100;
assign LUT_3[14249] = 32'b00000000000000100000001110100001;
assign LUT_3[14250] = 32'b00000000000000011011101010101000;
assign LUT_3[14251] = 32'b00000000000000100010010110000101;
assign LUT_3[14252] = 32'b00000000000000010110110000111010;
assign LUT_3[14253] = 32'b00000000000000011101011100010111;
assign LUT_3[14254] = 32'b00000000000000011000111000011110;
assign LUT_3[14255] = 32'b00000000000000011111100011111011;
assign LUT_3[14256] = 32'b00000000000000010111011101000001;
assign LUT_3[14257] = 32'b00000000000000011110001000011110;
assign LUT_3[14258] = 32'b00000000000000011001100100100101;
assign LUT_3[14259] = 32'b00000000000000100000010000000010;
assign LUT_3[14260] = 32'b00000000000000010100101010110111;
assign LUT_3[14261] = 32'b00000000000000011011010110010100;
assign LUT_3[14262] = 32'b00000000000000010110110010011011;
assign LUT_3[14263] = 32'b00000000000000011101011101111000;
assign LUT_3[14264] = 32'b00000000000000011100110110000111;
assign LUT_3[14265] = 32'b00000000000000100011100001100100;
assign LUT_3[14266] = 32'b00000000000000011110111101101011;
assign LUT_3[14267] = 32'b00000000000000100101101001001000;
assign LUT_3[14268] = 32'b00000000000000011010000011111101;
assign LUT_3[14269] = 32'b00000000000000100000101111011010;
assign LUT_3[14270] = 32'b00000000000000011100001011100001;
assign LUT_3[14271] = 32'b00000000000000100010110110111110;
assign LUT_3[14272] = 32'b00000000000000010010110100001001;
assign LUT_3[14273] = 32'b00000000000000011001011111100110;
assign LUT_3[14274] = 32'b00000000000000010100111011101101;
assign LUT_3[14275] = 32'b00000000000000011011100111001010;
assign LUT_3[14276] = 32'b00000000000000010000000001111111;
assign LUT_3[14277] = 32'b00000000000000010110101101011100;
assign LUT_3[14278] = 32'b00000000000000010010001001100011;
assign LUT_3[14279] = 32'b00000000000000011000110101000000;
assign LUT_3[14280] = 32'b00000000000000011000001101001111;
assign LUT_3[14281] = 32'b00000000000000011110111000101100;
assign LUT_3[14282] = 32'b00000000000000011010010100110011;
assign LUT_3[14283] = 32'b00000000000000100001000000010000;
assign LUT_3[14284] = 32'b00000000000000010101011011000101;
assign LUT_3[14285] = 32'b00000000000000011100000110100010;
assign LUT_3[14286] = 32'b00000000000000010111100010101001;
assign LUT_3[14287] = 32'b00000000000000011110001110000110;
assign LUT_3[14288] = 32'b00000000000000010110000111001100;
assign LUT_3[14289] = 32'b00000000000000011100110010101001;
assign LUT_3[14290] = 32'b00000000000000011000001110110000;
assign LUT_3[14291] = 32'b00000000000000011110111010001101;
assign LUT_3[14292] = 32'b00000000000000010011010101000010;
assign LUT_3[14293] = 32'b00000000000000011010000000011111;
assign LUT_3[14294] = 32'b00000000000000010101011100100110;
assign LUT_3[14295] = 32'b00000000000000011100001000000011;
assign LUT_3[14296] = 32'b00000000000000011011100000010010;
assign LUT_3[14297] = 32'b00000000000000100010001011101111;
assign LUT_3[14298] = 32'b00000000000000011101100111110110;
assign LUT_3[14299] = 32'b00000000000000100100010011010011;
assign LUT_3[14300] = 32'b00000000000000011000101110001000;
assign LUT_3[14301] = 32'b00000000000000011111011001100101;
assign LUT_3[14302] = 32'b00000000000000011010110101101100;
assign LUT_3[14303] = 32'b00000000000000100001100001001001;
assign LUT_3[14304] = 32'b00000000000000010100000010101001;
assign LUT_3[14305] = 32'b00000000000000011010101110000110;
assign LUT_3[14306] = 32'b00000000000000010110001010001101;
assign LUT_3[14307] = 32'b00000000000000011100110101101010;
assign LUT_3[14308] = 32'b00000000000000010001010000011111;
assign LUT_3[14309] = 32'b00000000000000010111111011111100;
assign LUT_3[14310] = 32'b00000000000000010011011000000011;
assign LUT_3[14311] = 32'b00000000000000011010000011100000;
assign LUT_3[14312] = 32'b00000000000000011001011011101111;
assign LUT_3[14313] = 32'b00000000000000100000000111001100;
assign LUT_3[14314] = 32'b00000000000000011011100011010011;
assign LUT_3[14315] = 32'b00000000000000100010001110110000;
assign LUT_3[14316] = 32'b00000000000000010110101001100101;
assign LUT_3[14317] = 32'b00000000000000011101010101000010;
assign LUT_3[14318] = 32'b00000000000000011000110001001001;
assign LUT_3[14319] = 32'b00000000000000011111011100100110;
assign LUT_3[14320] = 32'b00000000000000010111010101101100;
assign LUT_3[14321] = 32'b00000000000000011110000001001001;
assign LUT_3[14322] = 32'b00000000000000011001011101010000;
assign LUT_3[14323] = 32'b00000000000000100000001000101101;
assign LUT_3[14324] = 32'b00000000000000010100100011100010;
assign LUT_3[14325] = 32'b00000000000000011011001110111111;
assign LUT_3[14326] = 32'b00000000000000010110101011000110;
assign LUT_3[14327] = 32'b00000000000000011101010110100011;
assign LUT_3[14328] = 32'b00000000000000011100101110110010;
assign LUT_3[14329] = 32'b00000000000000100011011010001111;
assign LUT_3[14330] = 32'b00000000000000011110110110010110;
assign LUT_3[14331] = 32'b00000000000000100101100001110011;
assign LUT_3[14332] = 32'b00000000000000011001111100101000;
assign LUT_3[14333] = 32'b00000000000000100000101000000101;
assign LUT_3[14334] = 32'b00000000000000011100000100001100;
assign LUT_3[14335] = 32'b00000000000000100010101111101001;
assign LUT_3[14336] = 32'b00000000000000001100011101000100;
assign LUT_3[14337] = 32'b00000000000000010011001000100001;
assign LUT_3[14338] = 32'b00000000000000001110100100101000;
assign LUT_3[14339] = 32'b00000000000000010101010000000101;
assign LUT_3[14340] = 32'b00000000000000001001101010111010;
assign LUT_3[14341] = 32'b00000000000000010000010110010111;
assign LUT_3[14342] = 32'b00000000000000001011110010011110;
assign LUT_3[14343] = 32'b00000000000000010010011101111011;
assign LUT_3[14344] = 32'b00000000000000010001110110001010;
assign LUT_3[14345] = 32'b00000000000000011000100001100111;
assign LUT_3[14346] = 32'b00000000000000010011111101101110;
assign LUT_3[14347] = 32'b00000000000000011010101001001011;
assign LUT_3[14348] = 32'b00000000000000001111000100000000;
assign LUT_3[14349] = 32'b00000000000000010101101111011101;
assign LUT_3[14350] = 32'b00000000000000010001001011100100;
assign LUT_3[14351] = 32'b00000000000000010111110111000001;
assign LUT_3[14352] = 32'b00000000000000001111110000000111;
assign LUT_3[14353] = 32'b00000000000000010110011011100100;
assign LUT_3[14354] = 32'b00000000000000010001110111101011;
assign LUT_3[14355] = 32'b00000000000000011000100011001000;
assign LUT_3[14356] = 32'b00000000000000001100111101111101;
assign LUT_3[14357] = 32'b00000000000000010011101001011010;
assign LUT_3[14358] = 32'b00000000000000001111000101100001;
assign LUT_3[14359] = 32'b00000000000000010101110000111110;
assign LUT_3[14360] = 32'b00000000000000010101001001001101;
assign LUT_3[14361] = 32'b00000000000000011011110100101010;
assign LUT_3[14362] = 32'b00000000000000010111010000110001;
assign LUT_3[14363] = 32'b00000000000000011101111100001110;
assign LUT_3[14364] = 32'b00000000000000010010010111000011;
assign LUT_3[14365] = 32'b00000000000000011001000010100000;
assign LUT_3[14366] = 32'b00000000000000010100011110100111;
assign LUT_3[14367] = 32'b00000000000000011011001010000100;
assign LUT_3[14368] = 32'b00000000000000001101101011100100;
assign LUT_3[14369] = 32'b00000000000000010100010111000001;
assign LUT_3[14370] = 32'b00000000000000001111110011001000;
assign LUT_3[14371] = 32'b00000000000000010110011110100101;
assign LUT_3[14372] = 32'b00000000000000001010111001011010;
assign LUT_3[14373] = 32'b00000000000000010001100100110111;
assign LUT_3[14374] = 32'b00000000000000001101000000111110;
assign LUT_3[14375] = 32'b00000000000000010011101100011011;
assign LUT_3[14376] = 32'b00000000000000010011000100101010;
assign LUT_3[14377] = 32'b00000000000000011001110000000111;
assign LUT_3[14378] = 32'b00000000000000010101001100001110;
assign LUT_3[14379] = 32'b00000000000000011011110111101011;
assign LUT_3[14380] = 32'b00000000000000010000010010100000;
assign LUT_3[14381] = 32'b00000000000000010110111101111101;
assign LUT_3[14382] = 32'b00000000000000010010011010000100;
assign LUT_3[14383] = 32'b00000000000000011001000101100001;
assign LUT_3[14384] = 32'b00000000000000010000111110100111;
assign LUT_3[14385] = 32'b00000000000000010111101010000100;
assign LUT_3[14386] = 32'b00000000000000010011000110001011;
assign LUT_3[14387] = 32'b00000000000000011001110001101000;
assign LUT_3[14388] = 32'b00000000000000001110001100011101;
assign LUT_3[14389] = 32'b00000000000000010100110111111010;
assign LUT_3[14390] = 32'b00000000000000010000010100000001;
assign LUT_3[14391] = 32'b00000000000000010110111111011110;
assign LUT_3[14392] = 32'b00000000000000010110010111101101;
assign LUT_3[14393] = 32'b00000000000000011101000011001010;
assign LUT_3[14394] = 32'b00000000000000011000011111010001;
assign LUT_3[14395] = 32'b00000000000000011111001010101110;
assign LUT_3[14396] = 32'b00000000000000010011100101100011;
assign LUT_3[14397] = 32'b00000000000000011010010001000000;
assign LUT_3[14398] = 32'b00000000000000010101101101000111;
assign LUT_3[14399] = 32'b00000000000000011100011000100100;
assign LUT_3[14400] = 32'b00000000000000001100010101101111;
assign LUT_3[14401] = 32'b00000000000000010011000001001100;
assign LUT_3[14402] = 32'b00000000000000001110011101010011;
assign LUT_3[14403] = 32'b00000000000000010101001000110000;
assign LUT_3[14404] = 32'b00000000000000001001100011100101;
assign LUT_3[14405] = 32'b00000000000000010000001111000010;
assign LUT_3[14406] = 32'b00000000000000001011101011001001;
assign LUT_3[14407] = 32'b00000000000000010010010110100110;
assign LUT_3[14408] = 32'b00000000000000010001101110110101;
assign LUT_3[14409] = 32'b00000000000000011000011010010010;
assign LUT_3[14410] = 32'b00000000000000010011110110011001;
assign LUT_3[14411] = 32'b00000000000000011010100001110110;
assign LUT_3[14412] = 32'b00000000000000001110111100101011;
assign LUT_3[14413] = 32'b00000000000000010101101000001000;
assign LUT_3[14414] = 32'b00000000000000010001000100001111;
assign LUT_3[14415] = 32'b00000000000000010111101111101100;
assign LUT_3[14416] = 32'b00000000000000001111101000110010;
assign LUT_3[14417] = 32'b00000000000000010110010100001111;
assign LUT_3[14418] = 32'b00000000000000010001110000010110;
assign LUT_3[14419] = 32'b00000000000000011000011011110011;
assign LUT_3[14420] = 32'b00000000000000001100110110101000;
assign LUT_3[14421] = 32'b00000000000000010011100010000101;
assign LUT_3[14422] = 32'b00000000000000001110111110001100;
assign LUT_3[14423] = 32'b00000000000000010101101001101001;
assign LUT_3[14424] = 32'b00000000000000010101000001111000;
assign LUT_3[14425] = 32'b00000000000000011011101101010101;
assign LUT_3[14426] = 32'b00000000000000010111001001011100;
assign LUT_3[14427] = 32'b00000000000000011101110100111001;
assign LUT_3[14428] = 32'b00000000000000010010001111101110;
assign LUT_3[14429] = 32'b00000000000000011000111011001011;
assign LUT_3[14430] = 32'b00000000000000010100010111010010;
assign LUT_3[14431] = 32'b00000000000000011011000010101111;
assign LUT_3[14432] = 32'b00000000000000001101100100001111;
assign LUT_3[14433] = 32'b00000000000000010100001111101100;
assign LUT_3[14434] = 32'b00000000000000001111101011110011;
assign LUT_3[14435] = 32'b00000000000000010110010111010000;
assign LUT_3[14436] = 32'b00000000000000001010110010000101;
assign LUT_3[14437] = 32'b00000000000000010001011101100010;
assign LUT_3[14438] = 32'b00000000000000001100111001101001;
assign LUT_3[14439] = 32'b00000000000000010011100101000110;
assign LUT_3[14440] = 32'b00000000000000010010111101010101;
assign LUT_3[14441] = 32'b00000000000000011001101000110010;
assign LUT_3[14442] = 32'b00000000000000010101000100111001;
assign LUT_3[14443] = 32'b00000000000000011011110000010110;
assign LUT_3[14444] = 32'b00000000000000010000001011001011;
assign LUT_3[14445] = 32'b00000000000000010110110110101000;
assign LUT_3[14446] = 32'b00000000000000010010010010101111;
assign LUT_3[14447] = 32'b00000000000000011000111110001100;
assign LUT_3[14448] = 32'b00000000000000010000110111010010;
assign LUT_3[14449] = 32'b00000000000000010111100010101111;
assign LUT_3[14450] = 32'b00000000000000010010111110110110;
assign LUT_3[14451] = 32'b00000000000000011001101010010011;
assign LUT_3[14452] = 32'b00000000000000001110000101001000;
assign LUT_3[14453] = 32'b00000000000000010100110000100101;
assign LUT_3[14454] = 32'b00000000000000010000001100101100;
assign LUT_3[14455] = 32'b00000000000000010110111000001001;
assign LUT_3[14456] = 32'b00000000000000010110010000011000;
assign LUT_3[14457] = 32'b00000000000000011100111011110101;
assign LUT_3[14458] = 32'b00000000000000011000010111111100;
assign LUT_3[14459] = 32'b00000000000000011111000011011001;
assign LUT_3[14460] = 32'b00000000000000010011011110001110;
assign LUT_3[14461] = 32'b00000000000000011010001001101011;
assign LUT_3[14462] = 32'b00000000000000010101100101110010;
assign LUT_3[14463] = 32'b00000000000000011100010001001111;
assign LUT_3[14464] = 32'b00000000000000001110101000000010;
assign LUT_3[14465] = 32'b00000000000000010101010011011111;
assign LUT_3[14466] = 32'b00000000000000010000101111100110;
assign LUT_3[14467] = 32'b00000000000000010111011011000011;
assign LUT_3[14468] = 32'b00000000000000001011110101111000;
assign LUT_3[14469] = 32'b00000000000000010010100001010101;
assign LUT_3[14470] = 32'b00000000000000001101111101011100;
assign LUT_3[14471] = 32'b00000000000000010100101000111001;
assign LUT_3[14472] = 32'b00000000000000010100000001001000;
assign LUT_3[14473] = 32'b00000000000000011010101100100101;
assign LUT_3[14474] = 32'b00000000000000010110001000101100;
assign LUT_3[14475] = 32'b00000000000000011100110100001001;
assign LUT_3[14476] = 32'b00000000000000010001001110111110;
assign LUT_3[14477] = 32'b00000000000000010111111010011011;
assign LUT_3[14478] = 32'b00000000000000010011010110100010;
assign LUT_3[14479] = 32'b00000000000000011010000001111111;
assign LUT_3[14480] = 32'b00000000000000010001111011000101;
assign LUT_3[14481] = 32'b00000000000000011000100110100010;
assign LUT_3[14482] = 32'b00000000000000010100000010101001;
assign LUT_3[14483] = 32'b00000000000000011010101110000110;
assign LUT_3[14484] = 32'b00000000000000001111001000111011;
assign LUT_3[14485] = 32'b00000000000000010101110100011000;
assign LUT_3[14486] = 32'b00000000000000010001010000011111;
assign LUT_3[14487] = 32'b00000000000000010111111011111100;
assign LUT_3[14488] = 32'b00000000000000010111010100001011;
assign LUT_3[14489] = 32'b00000000000000011101111111101000;
assign LUT_3[14490] = 32'b00000000000000011001011011101111;
assign LUT_3[14491] = 32'b00000000000000100000000111001100;
assign LUT_3[14492] = 32'b00000000000000010100100010000001;
assign LUT_3[14493] = 32'b00000000000000011011001101011110;
assign LUT_3[14494] = 32'b00000000000000010110101001100101;
assign LUT_3[14495] = 32'b00000000000000011101010101000010;
assign LUT_3[14496] = 32'b00000000000000001111110110100010;
assign LUT_3[14497] = 32'b00000000000000010110100001111111;
assign LUT_3[14498] = 32'b00000000000000010001111110000110;
assign LUT_3[14499] = 32'b00000000000000011000101001100011;
assign LUT_3[14500] = 32'b00000000000000001101000100011000;
assign LUT_3[14501] = 32'b00000000000000010011101111110101;
assign LUT_3[14502] = 32'b00000000000000001111001011111100;
assign LUT_3[14503] = 32'b00000000000000010101110111011001;
assign LUT_3[14504] = 32'b00000000000000010101001111101000;
assign LUT_3[14505] = 32'b00000000000000011011111011000101;
assign LUT_3[14506] = 32'b00000000000000010111010111001100;
assign LUT_3[14507] = 32'b00000000000000011110000010101001;
assign LUT_3[14508] = 32'b00000000000000010010011101011110;
assign LUT_3[14509] = 32'b00000000000000011001001000111011;
assign LUT_3[14510] = 32'b00000000000000010100100101000010;
assign LUT_3[14511] = 32'b00000000000000011011010000011111;
assign LUT_3[14512] = 32'b00000000000000010011001001100101;
assign LUT_3[14513] = 32'b00000000000000011001110101000010;
assign LUT_3[14514] = 32'b00000000000000010101010001001001;
assign LUT_3[14515] = 32'b00000000000000011011111100100110;
assign LUT_3[14516] = 32'b00000000000000010000010111011011;
assign LUT_3[14517] = 32'b00000000000000010111000010111000;
assign LUT_3[14518] = 32'b00000000000000010010011110111111;
assign LUT_3[14519] = 32'b00000000000000011001001010011100;
assign LUT_3[14520] = 32'b00000000000000011000100010101011;
assign LUT_3[14521] = 32'b00000000000000011111001110001000;
assign LUT_3[14522] = 32'b00000000000000011010101010001111;
assign LUT_3[14523] = 32'b00000000000000100001010101101100;
assign LUT_3[14524] = 32'b00000000000000010101110000100001;
assign LUT_3[14525] = 32'b00000000000000011100011011111110;
assign LUT_3[14526] = 32'b00000000000000010111111000000101;
assign LUT_3[14527] = 32'b00000000000000011110100011100010;
assign LUT_3[14528] = 32'b00000000000000001110100000101101;
assign LUT_3[14529] = 32'b00000000000000010101001100001010;
assign LUT_3[14530] = 32'b00000000000000010000101000010001;
assign LUT_3[14531] = 32'b00000000000000010111010011101110;
assign LUT_3[14532] = 32'b00000000000000001011101110100011;
assign LUT_3[14533] = 32'b00000000000000010010011010000000;
assign LUT_3[14534] = 32'b00000000000000001101110110000111;
assign LUT_3[14535] = 32'b00000000000000010100100001100100;
assign LUT_3[14536] = 32'b00000000000000010011111001110011;
assign LUT_3[14537] = 32'b00000000000000011010100101010000;
assign LUT_3[14538] = 32'b00000000000000010110000001010111;
assign LUT_3[14539] = 32'b00000000000000011100101100110100;
assign LUT_3[14540] = 32'b00000000000000010001000111101001;
assign LUT_3[14541] = 32'b00000000000000010111110011000110;
assign LUT_3[14542] = 32'b00000000000000010011001111001101;
assign LUT_3[14543] = 32'b00000000000000011001111010101010;
assign LUT_3[14544] = 32'b00000000000000010001110011110000;
assign LUT_3[14545] = 32'b00000000000000011000011111001101;
assign LUT_3[14546] = 32'b00000000000000010011111011010100;
assign LUT_3[14547] = 32'b00000000000000011010100110110001;
assign LUT_3[14548] = 32'b00000000000000001111000001100110;
assign LUT_3[14549] = 32'b00000000000000010101101101000011;
assign LUT_3[14550] = 32'b00000000000000010001001001001010;
assign LUT_3[14551] = 32'b00000000000000010111110100100111;
assign LUT_3[14552] = 32'b00000000000000010111001100110110;
assign LUT_3[14553] = 32'b00000000000000011101111000010011;
assign LUT_3[14554] = 32'b00000000000000011001010100011010;
assign LUT_3[14555] = 32'b00000000000000011111111111110111;
assign LUT_3[14556] = 32'b00000000000000010100011010101100;
assign LUT_3[14557] = 32'b00000000000000011011000110001001;
assign LUT_3[14558] = 32'b00000000000000010110100010010000;
assign LUT_3[14559] = 32'b00000000000000011101001101101101;
assign LUT_3[14560] = 32'b00000000000000001111101111001101;
assign LUT_3[14561] = 32'b00000000000000010110011010101010;
assign LUT_3[14562] = 32'b00000000000000010001110110110001;
assign LUT_3[14563] = 32'b00000000000000011000100010001110;
assign LUT_3[14564] = 32'b00000000000000001100111101000011;
assign LUT_3[14565] = 32'b00000000000000010011101000100000;
assign LUT_3[14566] = 32'b00000000000000001111000100100111;
assign LUT_3[14567] = 32'b00000000000000010101110000000100;
assign LUT_3[14568] = 32'b00000000000000010101001000010011;
assign LUT_3[14569] = 32'b00000000000000011011110011110000;
assign LUT_3[14570] = 32'b00000000000000010111001111110111;
assign LUT_3[14571] = 32'b00000000000000011101111011010100;
assign LUT_3[14572] = 32'b00000000000000010010010110001001;
assign LUT_3[14573] = 32'b00000000000000011001000001100110;
assign LUT_3[14574] = 32'b00000000000000010100011101101101;
assign LUT_3[14575] = 32'b00000000000000011011001001001010;
assign LUT_3[14576] = 32'b00000000000000010011000010010000;
assign LUT_3[14577] = 32'b00000000000000011001101101101101;
assign LUT_3[14578] = 32'b00000000000000010101001001110100;
assign LUT_3[14579] = 32'b00000000000000011011110101010001;
assign LUT_3[14580] = 32'b00000000000000010000010000000110;
assign LUT_3[14581] = 32'b00000000000000010110111011100011;
assign LUT_3[14582] = 32'b00000000000000010010010111101010;
assign LUT_3[14583] = 32'b00000000000000011001000011000111;
assign LUT_3[14584] = 32'b00000000000000011000011011010110;
assign LUT_3[14585] = 32'b00000000000000011111000110110011;
assign LUT_3[14586] = 32'b00000000000000011010100010111010;
assign LUT_3[14587] = 32'b00000000000000100001001110010111;
assign LUT_3[14588] = 32'b00000000000000010101101001001100;
assign LUT_3[14589] = 32'b00000000000000011100010100101001;
assign LUT_3[14590] = 32'b00000000000000010111110000110000;
assign LUT_3[14591] = 32'b00000000000000011110011100001101;
assign LUT_3[14592] = 32'b00000000000000001000101100100101;
assign LUT_3[14593] = 32'b00000000000000001111011000000010;
assign LUT_3[14594] = 32'b00000000000000001010110100001001;
assign LUT_3[14595] = 32'b00000000000000010001011111100110;
assign LUT_3[14596] = 32'b00000000000000000101111010011011;
assign LUT_3[14597] = 32'b00000000000000001100100101111000;
assign LUT_3[14598] = 32'b00000000000000001000000001111111;
assign LUT_3[14599] = 32'b00000000000000001110101101011100;
assign LUT_3[14600] = 32'b00000000000000001110000101101011;
assign LUT_3[14601] = 32'b00000000000000010100110001001000;
assign LUT_3[14602] = 32'b00000000000000010000001101001111;
assign LUT_3[14603] = 32'b00000000000000010110111000101100;
assign LUT_3[14604] = 32'b00000000000000001011010011100001;
assign LUT_3[14605] = 32'b00000000000000010001111110111110;
assign LUT_3[14606] = 32'b00000000000000001101011011000101;
assign LUT_3[14607] = 32'b00000000000000010100000110100010;
assign LUT_3[14608] = 32'b00000000000000001011111111101000;
assign LUT_3[14609] = 32'b00000000000000010010101011000101;
assign LUT_3[14610] = 32'b00000000000000001110000111001100;
assign LUT_3[14611] = 32'b00000000000000010100110010101001;
assign LUT_3[14612] = 32'b00000000000000001001001101011110;
assign LUT_3[14613] = 32'b00000000000000001111111000111011;
assign LUT_3[14614] = 32'b00000000000000001011010101000010;
assign LUT_3[14615] = 32'b00000000000000010010000000011111;
assign LUT_3[14616] = 32'b00000000000000010001011000101110;
assign LUT_3[14617] = 32'b00000000000000011000000100001011;
assign LUT_3[14618] = 32'b00000000000000010011100000010010;
assign LUT_3[14619] = 32'b00000000000000011010001011101111;
assign LUT_3[14620] = 32'b00000000000000001110100110100100;
assign LUT_3[14621] = 32'b00000000000000010101010010000001;
assign LUT_3[14622] = 32'b00000000000000010000101110001000;
assign LUT_3[14623] = 32'b00000000000000010111011001100101;
assign LUT_3[14624] = 32'b00000000000000001001111011000101;
assign LUT_3[14625] = 32'b00000000000000010000100110100010;
assign LUT_3[14626] = 32'b00000000000000001100000010101001;
assign LUT_3[14627] = 32'b00000000000000010010101110000110;
assign LUT_3[14628] = 32'b00000000000000000111001000111011;
assign LUT_3[14629] = 32'b00000000000000001101110100011000;
assign LUT_3[14630] = 32'b00000000000000001001010000011111;
assign LUT_3[14631] = 32'b00000000000000001111111011111100;
assign LUT_3[14632] = 32'b00000000000000001111010100001011;
assign LUT_3[14633] = 32'b00000000000000010101111111101000;
assign LUT_3[14634] = 32'b00000000000000010001011011101111;
assign LUT_3[14635] = 32'b00000000000000011000000111001100;
assign LUT_3[14636] = 32'b00000000000000001100100010000001;
assign LUT_3[14637] = 32'b00000000000000010011001101011110;
assign LUT_3[14638] = 32'b00000000000000001110101001100101;
assign LUT_3[14639] = 32'b00000000000000010101010101000010;
assign LUT_3[14640] = 32'b00000000000000001101001110001000;
assign LUT_3[14641] = 32'b00000000000000010011111001100101;
assign LUT_3[14642] = 32'b00000000000000001111010101101100;
assign LUT_3[14643] = 32'b00000000000000010110000001001001;
assign LUT_3[14644] = 32'b00000000000000001010011011111110;
assign LUT_3[14645] = 32'b00000000000000010001000111011011;
assign LUT_3[14646] = 32'b00000000000000001100100011100010;
assign LUT_3[14647] = 32'b00000000000000010011001110111111;
assign LUT_3[14648] = 32'b00000000000000010010100111001110;
assign LUT_3[14649] = 32'b00000000000000011001010010101011;
assign LUT_3[14650] = 32'b00000000000000010100101110110010;
assign LUT_3[14651] = 32'b00000000000000011011011010001111;
assign LUT_3[14652] = 32'b00000000000000001111110101000100;
assign LUT_3[14653] = 32'b00000000000000010110100000100001;
assign LUT_3[14654] = 32'b00000000000000010001111100101000;
assign LUT_3[14655] = 32'b00000000000000011000101000000101;
assign LUT_3[14656] = 32'b00000000000000001000100101010000;
assign LUT_3[14657] = 32'b00000000000000001111010000101101;
assign LUT_3[14658] = 32'b00000000000000001010101100110100;
assign LUT_3[14659] = 32'b00000000000000010001011000010001;
assign LUT_3[14660] = 32'b00000000000000000101110011000110;
assign LUT_3[14661] = 32'b00000000000000001100011110100011;
assign LUT_3[14662] = 32'b00000000000000000111111010101010;
assign LUT_3[14663] = 32'b00000000000000001110100110000111;
assign LUT_3[14664] = 32'b00000000000000001101111110010110;
assign LUT_3[14665] = 32'b00000000000000010100101001110011;
assign LUT_3[14666] = 32'b00000000000000010000000101111010;
assign LUT_3[14667] = 32'b00000000000000010110110001010111;
assign LUT_3[14668] = 32'b00000000000000001011001100001100;
assign LUT_3[14669] = 32'b00000000000000010001110111101001;
assign LUT_3[14670] = 32'b00000000000000001101010011110000;
assign LUT_3[14671] = 32'b00000000000000010011111111001101;
assign LUT_3[14672] = 32'b00000000000000001011111000010011;
assign LUT_3[14673] = 32'b00000000000000010010100011110000;
assign LUT_3[14674] = 32'b00000000000000001101111111110111;
assign LUT_3[14675] = 32'b00000000000000010100101011010100;
assign LUT_3[14676] = 32'b00000000000000001001000110001001;
assign LUT_3[14677] = 32'b00000000000000001111110001100110;
assign LUT_3[14678] = 32'b00000000000000001011001101101101;
assign LUT_3[14679] = 32'b00000000000000010001111001001010;
assign LUT_3[14680] = 32'b00000000000000010001010001011001;
assign LUT_3[14681] = 32'b00000000000000010111111100110110;
assign LUT_3[14682] = 32'b00000000000000010011011000111101;
assign LUT_3[14683] = 32'b00000000000000011010000100011010;
assign LUT_3[14684] = 32'b00000000000000001110011111001111;
assign LUT_3[14685] = 32'b00000000000000010101001010101100;
assign LUT_3[14686] = 32'b00000000000000010000100110110011;
assign LUT_3[14687] = 32'b00000000000000010111010010010000;
assign LUT_3[14688] = 32'b00000000000000001001110011110000;
assign LUT_3[14689] = 32'b00000000000000010000011111001101;
assign LUT_3[14690] = 32'b00000000000000001011111011010100;
assign LUT_3[14691] = 32'b00000000000000010010100110110001;
assign LUT_3[14692] = 32'b00000000000000000111000001100110;
assign LUT_3[14693] = 32'b00000000000000001101101101000011;
assign LUT_3[14694] = 32'b00000000000000001001001001001010;
assign LUT_3[14695] = 32'b00000000000000001111110100100111;
assign LUT_3[14696] = 32'b00000000000000001111001100110110;
assign LUT_3[14697] = 32'b00000000000000010101111000010011;
assign LUT_3[14698] = 32'b00000000000000010001010100011010;
assign LUT_3[14699] = 32'b00000000000000010111111111110111;
assign LUT_3[14700] = 32'b00000000000000001100011010101100;
assign LUT_3[14701] = 32'b00000000000000010011000110001001;
assign LUT_3[14702] = 32'b00000000000000001110100010010000;
assign LUT_3[14703] = 32'b00000000000000010101001101101101;
assign LUT_3[14704] = 32'b00000000000000001101000110110011;
assign LUT_3[14705] = 32'b00000000000000010011110010010000;
assign LUT_3[14706] = 32'b00000000000000001111001110010111;
assign LUT_3[14707] = 32'b00000000000000010101111001110100;
assign LUT_3[14708] = 32'b00000000000000001010010100101001;
assign LUT_3[14709] = 32'b00000000000000010001000000000110;
assign LUT_3[14710] = 32'b00000000000000001100011100001101;
assign LUT_3[14711] = 32'b00000000000000010011000111101010;
assign LUT_3[14712] = 32'b00000000000000010010011111111001;
assign LUT_3[14713] = 32'b00000000000000011001001011010110;
assign LUT_3[14714] = 32'b00000000000000010100100111011101;
assign LUT_3[14715] = 32'b00000000000000011011010010111010;
assign LUT_3[14716] = 32'b00000000000000001111101101101111;
assign LUT_3[14717] = 32'b00000000000000010110011001001100;
assign LUT_3[14718] = 32'b00000000000000010001110101010011;
assign LUT_3[14719] = 32'b00000000000000011000100000110000;
assign LUT_3[14720] = 32'b00000000000000001010110111100011;
assign LUT_3[14721] = 32'b00000000000000010001100011000000;
assign LUT_3[14722] = 32'b00000000000000001100111111000111;
assign LUT_3[14723] = 32'b00000000000000010011101010100100;
assign LUT_3[14724] = 32'b00000000000000001000000101011001;
assign LUT_3[14725] = 32'b00000000000000001110110000110110;
assign LUT_3[14726] = 32'b00000000000000001010001100111101;
assign LUT_3[14727] = 32'b00000000000000010000111000011010;
assign LUT_3[14728] = 32'b00000000000000010000010000101001;
assign LUT_3[14729] = 32'b00000000000000010110111100000110;
assign LUT_3[14730] = 32'b00000000000000010010011000001101;
assign LUT_3[14731] = 32'b00000000000000011001000011101010;
assign LUT_3[14732] = 32'b00000000000000001101011110011111;
assign LUT_3[14733] = 32'b00000000000000010100001001111100;
assign LUT_3[14734] = 32'b00000000000000001111100110000011;
assign LUT_3[14735] = 32'b00000000000000010110010001100000;
assign LUT_3[14736] = 32'b00000000000000001110001010100110;
assign LUT_3[14737] = 32'b00000000000000010100110110000011;
assign LUT_3[14738] = 32'b00000000000000010000010010001010;
assign LUT_3[14739] = 32'b00000000000000010110111101100111;
assign LUT_3[14740] = 32'b00000000000000001011011000011100;
assign LUT_3[14741] = 32'b00000000000000010010000011111001;
assign LUT_3[14742] = 32'b00000000000000001101100000000000;
assign LUT_3[14743] = 32'b00000000000000010100001011011101;
assign LUT_3[14744] = 32'b00000000000000010011100011101100;
assign LUT_3[14745] = 32'b00000000000000011010001111001001;
assign LUT_3[14746] = 32'b00000000000000010101101011010000;
assign LUT_3[14747] = 32'b00000000000000011100010110101101;
assign LUT_3[14748] = 32'b00000000000000010000110001100010;
assign LUT_3[14749] = 32'b00000000000000010111011100111111;
assign LUT_3[14750] = 32'b00000000000000010010111001000110;
assign LUT_3[14751] = 32'b00000000000000011001100100100011;
assign LUT_3[14752] = 32'b00000000000000001100000110000011;
assign LUT_3[14753] = 32'b00000000000000010010110001100000;
assign LUT_3[14754] = 32'b00000000000000001110001101100111;
assign LUT_3[14755] = 32'b00000000000000010100111001000100;
assign LUT_3[14756] = 32'b00000000000000001001010011111001;
assign LUT_3[14757] = 32'b00000000000000001111111111010110;
assign LUT_3[14758] = 32'b00000000000000001011011011011101;
assign LUT_3[14759] = 32'b00000000000000010010000110111010;
assign LUT_3[14760] = 32'b00000000000000010001011111001001;
assign LUT_3[14761] = 32'b00000000000000011000001010100110;
assign LUT_3[14762] = 32'b00000000000000010011100110101101;
assign LUT_3[14763] = 32'b00000000000000011010010010001010;
assign LUT_3[14764] = 32'b00000000000000001110101100111111;
assign LUT_3[14765] = 32'b00000000000000010101011000011100;
assign LUT_3[14766] = 32'b00000000000000010000110100100011;
assign LUT_3[14767] = 32'b00000000000000010111100000000000;
assign LUT_3[14768] = 32'b00000000000000001111011001000110;
assign LUT_3[14769] = 32'b00000000000000010110000100100011;
assign LUT_3[14770] = 32'b00000000000000010001100000101010;
assign LUT_3[14771] = 32'b00000000000000011000001100000111;
assign LUT_3[14772] = 32'b00000000000000001100100110111100;
assign LUT_3[14773] = 32'b00000000000000010011010010011001;
assign LUT_3[14774] = 32'b00000000000000001110101110100000;
assign LUT_3[14775] = 32'b00000000000000010101011001111101;
assign LUT_3[14776] = 32'b00000000000000010100110010001100;
assign LUT_3[14777] = 32'b00000000000000011011011101101001;
assign LUT_3[14778] = 32'b00000000000000010110111001110000;
assign LUT_3[14779] = 32'b00000000000000011101100101001101;
assign LUT_3[14780] = 32'b00000000000000010010000000000010;
assign LUT_3[14781] = 32'b00000000000000011000101011011111;
assign LUT_3[14782] = 32'b00000000000000010100000111100110;
assign LUT_3[14783] = 32'b00000000000000011010110011000011;
assign LUT_3[14784] = 32'b00000000000000001010110000001110;
assign LUT_3[14785] = 32'b00000000000000010001011011101011;
assign LUT_3[14786] = 32'b00000000000000001100110111110010;
assign LUT_3[14787] = 32'b00000000000000010011100011001111;
assign LUT_3[14788] = 32'b00000000000000000111111110000100;
assign LUT_3[14789] = 32'b00000000000000001110101001100001;
assign LUT_3[14790] = 32'b00000000000000001010000101101000;
assign LUT_3[14791] = 32'b00000000000000010000110001000101;
assign LUT_3[14792] = 32'b00000000000000010000001001010100;
assign LUT_3[14793] = 32'b00000000000000010110110100110001;
assign LUT_3[14794] = 32'b00000000000000010010010000111000;
assign LUT_3[14795] = 32'b00000000000000011000111100010101;
assign LUT_3[14796] = 32'b00000000000000001101010111001010;
assign LUT_3[14797] = 32'b00000000000000010100000010100111;
assign LUT_3[14798] = 32'b00000000000000001111011110101110;
assign LUT_3[14799] = 32'b00000000000000010110001010001011;
assign LUT_3[14800] = 32'b00000000000000001110000011010001;
assign LUT_3[14801] = 32'b00000000000000010100101110101110;
assign LUT_3[14802] = 32'b00000000000000010000001010110101;
assign LUT_3[14803] = 32'b00000000000000010110110110010010;
assign LUT_3[14804] = 32'b00000000000000001011010001000111;
assign LUT_3[14805] = 32'b00000000000000010001111100100100;
assign LUT_3[14806] = 32'b00000000000000001101011000101011;
assign LUT_3[14807] = 32'b00000000000000010100000100001000;
assign LUT_3[14808] = 32'b00000000000000010011011100010111;
assign LUT_3[14809] = 32'b00000000000000011010000111110100;
assign LUT_3[14810] = 32'b00000000000000010101100011111011;
assign LUT_3[14811] = 32'b00000000000000011100001111011000;
assign LUT_3[14812] = 32'b00000000000000010000101010001101;
assign LUT_3[14813] = 32'b00000000000000010111010101101010;
assign LUT_3[14814] = 32'b00000000000000010010110001110001;
assign LUT_3[14815] = 32'b00000000000000011001011101001110;
assign LUT_3[14816] = 32'b00000000000000001011111110101110;
assign LUT_3[14817] = 32'b00000000000000010010101010001011;
assign LUT_3[14818] = 32'b00000000000000001110000110010010;
assign LUT_3[14819] = 32'b00000000000000010100110001101111;
assign LUT_3[14820] = 32'b00000000000000001001001100100100;
assign LUT_3[14821] = 32'b00000000000000001111111000000001;
assign LUT_3[14822] = 32'b00000000000000001011010100001000;
assign LUT_3[14823] = 32'b00000000000000010001111111100101;
assign LUT_3[14824] = 32'b00000000000000010001010111110100;
assign LUT_3[14825] = 32'b00000000000000011000000011010001;
assign LUT_3[14826] = 32'b00000000000000010011011111011000;
assign LUT_3[14827] = 32'b00000000000000011010001010110101;
assign LUT_3[14828] = 32'b00000000000000001110100101101010;
assign LUT_3[14829] = 32'b00000000000000010101010001000111;
assign LUT_3[14830] = 32'b00000000000000010000101101001110;
assign LUT_3[14831] = 32'b00000000000000010111011000101011;
assign LUT_3[14832] = 32'b00000000000000001111010001110001;
assign LUT_3[14833] = 32'b00000000000000010101111101001110;
assign LUT_3[14834] = 32'b00000000000000010001011001010101;
assign LUT_3[14835] = 32'b00000000000000011000000100110010;
assign LUT_3[14836] = 32'b00000000000000001100011111100111;
assign LUT_3[14837] = 32'b00000000000000010011001011000100;
assign LUT_3[14838] = 32'b00000000000000001110100111001011;
assign LUT_3[14839] = 32'b00000000000000010101010010101000;
assign LUT_3[14840] = 32'b00000000000000010100101010110111;
assign LUT_3[14841] = 32'b00000000000000011011010110010100;
assign LUT_3[14842] = 32'b00000000000000010110110010011011;
assign LUT_3[14843] = 32'b00000000000000011101011101111000;
assign LUT_3[14844] = 32'b00000000000000010001111000101101;
assign LUT_3[14845] = 32'b00000000000000011000100100001010;
assign LUT_3[14846] = 32'b00000000000000010100000000010001;
assign LUT_3[14847] = 32'b00000000000000011010101011101110;
assign LUT_3[14848] = 32'b00000000000000001111110010010000;
assign LUT_3[14849] = 32'b00000000000000010110011101101101;
assign LUT_3[14850] = 32'b00000000000000010001111001110100;
assign LUT_3[14851] = 32'b00000000000000011000100101010001;
assign LUT_3[14852] = 32'b00000000000000001101000000000110;
assign LUT_3[14853] = 32'b00000000000000010011101011100011;
assign LUT_3[14854] = 32'b00000000000000001111000111101010;
assign LUT_3[14855] = 32'b00000000000000010101110011000111;
assign LUT_3[14856] = 32'b00000000000000010101001011010110;
assign LUT_3[14857] = 32'b00000000000000011011110110110011;
assign LUT_3[14858] = 32'b00000000000000010111010010111010;
assign LUT_3[14859] = 32'b00000000000000011101111110010111;
assign LUT_3[14860] = 32'b00000000000000010010011001001100;
assign LUT_3[14861] = 32'b00000000000000011001000100101001;
assign LUT_3[14862] = 32'b00000000000000010100100000110000;
assign LUT_3[14863] = 32'b00000000000000011011001100001101;
assign LUT_3[14864] = 32'b00000000000000010011000101010011;
assign LUT_3[14865] = 32'b00000000000000011001110000110000;
assign LUT_3[14866] = 32'b00000000000000010101001100110111;
assign LUT_3[14867] = 32'b00000000000000011011111000010100;
assign LUT_3[14868] = 32'b00000000000000010000010011001001;
assign LUT_3[14869] = 32'b00000000000000010110111110100110;
assign LUT_3[14870] = 32'b00000000000000010010011010101101;
assign LUT_3[14871] = 32'b00000000000000011001000110001010;
assign LUT_3[14872] = 32'b00000000000000011000011110011001;
assign LUT_3[14873] = 32'b00000000000000011111001001110110;
assign LUT_3[14874] = 32'b00000000000000011010100101111101;
assign LUT_3[14875] = 32'b00000000000000100001010001011010;
assign LUT_3[14876] = 32'b00000000000000010101101100001111;
assign LUT_3[14877] = 32'b00000000000000011100010111101100;
assign LUT_3[14878] = 32'b00000000000000010111110011110011;
assign LUT_3[14879] = 32'b00000000000000011110011111010000;
assign LUT_3[14880] = 32'b00000000000000010001000000110000;
assign LUT_3[14881] = 32'b00000000000000010111101100001101;
assign LUT_3[14882] = 32'b00000000000000010011001000010100;
assign LUT_3[14883] = 32'b00000000000000011001110011110001;
assign LUT_3[14884] = 32'b00000000000000001110001110100110;
assign LUT_3[14885] = 32'b00000000000000010100111010000011;
assign LUT_3[14886] = 32'b00000000000000010000010110001010;
assign LUT_3[14887] = 32'b00000000000000010111000001100111;
assign LUT_3[14888] = 32'b00000000000000010110011001110110;
assign LUT_3[14889] = 32'b00000000000000011101000101010011;
assign LUT_3[14890] = 32'b00000000000000011000100001011010;
assign LUT_3[14891] = 32'b00000000000000011111001100110111;
assign LUT_3[14892] = 32'b00000000000000010011100111101100;
assign LUT_3[14893] = 32'b00000000000000011010010011001001;
assign LUT_3[14894] = 32'b00000000000000010101101111010000;
assign LUT_3[14895] = 32'b00000000000000011100011010101101;
assign LUT_3[14896] = 32'b00000000000000010100010011110011;
assign LUT_3[14897] = 32'b00000000000000011010111111010000;
assign LUT_3[14898] = 32'b00000000000000010110011011010111;
assign LUT_3[14899] = 32'b00000000000000011101000110110100;
assign LUT_3[14900] = 32'b00000000000000010001100001101001;
assign LUT_3[14901] = 32'b00000000000000011000001101000110;
assign LUT_3[14902] = 32'b00000000000000010011101001001101;
assign LUT_3[14903] = 32'b00000000000000011010010100101010;
assign LUT_3[14904] = 32'b00000000000000011001101100111001;
assign LUT_3[14905] = 32'b00000000000000100000011000010110;
assign LUT_3[14906] = 32'b00000000000000011011110100011101;
assign LUT_3[14907] = 32'b00000000000000100010011111111010;
assign LUT_3[14908] = 32'b00000000000000010110111010101111;
assign LUT_3[14909] = 32'b00000000000000011101100110001100;
assign LUT_3[14910] = 32'b00000000000000011001000010010011;
assign LUT_3[14911] = 32'b00000000000000011111101101110000;
assign LUT_3[14912] = 32'b00000000000000001111101010111011;
assign LUT_3[14913] = 32'b00000000000000010110010110011000;
assign LUT_3[14914] = 32'b00000000000000010001110010011111;
assign LUT_3[14915] = 32'b00000000000000011000011101111100;
assign LUT_3[14916] = 32'b00000000000000001100111000110001;
assign LUT_3[14917] = 32'b00000000000000010011100100001110;
assign LUT_3[14918] = 32'b00000000000000001111000000010101;
assign LUT_3[14919] = 32'b00000000000000010101101011110010;
assign LUT_3[14920] = 32'b00000000000000010101000100000001;
assign LUT_3[14921] = 32'b00000000000000011011101111011110;
assign LUT_3[14922] = 32'b00000000000000010111001011100101;
assign LUT_3[14923] = 32'b00000000000000011101110111000010;
assign LUT_3[14924] = 32'b00000000000000010010010001110111;
assign LUT_3[14925] = 32'b00000000000000011000111101010100;
assign LUT_3[14926] = 32'b00000000000000010100011001011011;
assign LUT_3[14927] = 32'b00000000000000011011000100111000;
assign LUT_3[14928] = 32'b00000000000000010010111101111110;
assign LUT_3[14929] = 32'b00000000000000011001101001011011;
assign LUT_3[14930] = 32'b00000000000000010101000101100010;
assign LUT_3[14931] = 32'b00000000000000011011110000111111;
assign LUT_3[14932] = 32'b00000000000000010000001011110100;
assign LUT_3[14933] = 32'b00000000000000010110110111010001;
assign LUT_3[14934] = 32'b00000000000000010010010011011000;
assign LUT_3[14935] = 32'b00000000000000011000111110110101;
assign LUT_3[14936] = 32'b00000000000000011000010111000100;
assign LUT_3[14937] = 32'b00000000000000011111000010100001;
assign LUT_3[14938] = 32'b00000000000000011010011110101000;
assign LUT_3[14939] = 32'b00000000000000100001001010000101;
assign LUT_3[14940] = 32'b00000000000000010101100100111010;
assign LUT_3[14941] = 32'b00000000000000011100010000010111;
assign LUT_3[14942] = 32'b00000000000000010111101100011110;
assign LUT_3[14943] = 32'b00000000000000011110010111111011;
assign LUT_3[14944] = 32'b00000000000000010000111001011011;
assign LUT_3[14945] = 32'b00000000000000010111100100111000;
assign LUT_3[14946] = 32'b00000000000000010011000000111111;
assign LUT_3[14947] = 32'b00000000000000011001101100011100;
assign LUT_3[14948] = 32'b00000000000000001110000111010001;
assign LUT_3[14949] = 32'b00000000000000010100110010101110;
assign LUT_3[14950] = 32'b00000000000000010000001110110101;
assign LUT_3[14951] = 32'b00000000000000010110111010010010;
assign LUT_3[14952] = 32'b00000000000000010110010010100001;
assign LUT_3[14953] = 32'b00000000000000011100111101111110;
assign LUT_3[14954] = 32'b00000000000000011000011010000101;
assign LUT_3[14955] = 32'b00000000000000011111000101100010;
assign LUT_3[14956] = 32'b00000000000000010011100000010111;
assign LUT_3[14957] = 32'b00000000000000011010001011110100;
assign LUT_3[14958] = 32'b00000000000000010101100111111011;
assign LUT_3[14959] = 32'b00000000000000011100010011011000;
assign LUT_3[14960] = 32'b00000000000000010100001100011110;
assign LUT_3[14961] = 32'b00000000000000011010110111111011;
assign LUT_3[14962] = 32'b00000000000000010110010100000010;
assign LUT_3[14963] = 32'b00000000000000011100111111011111;
assign LUT_3[14964] = 32'b00000000000000010001011010010100;
assign LUT_3[14965] = 32'b00000000000000011000000101110001;
assign LUT_3[14966] = 32'b00000000000000010011100001111000;
assign LUT_3[14967] = 32'b00000000000000011010001101010101;
assign LUT_3[14968] = 32'b00000000000000011001100101100100;
assign LUT_3[14969] = 32'b00000000000000100000010001000001;
assign LUT_3[14970] = 32'b00000000000000011011101101001000;
assign LUT_3[14971] = 32'b00000000000000100010011000100101;
assign LUT_3[14972] = 32'b00000000000000010110110011011010;
assign LUT_3[14973] = 32'b00000000000000011101011110110111;
assign LUT_3[14974] = 32'b00000000000000011000111010111110;
assign LUT_3[14975] = 32'b00000000000000011111100110011011;
assign LUT_3[14976] = 32'b00000000000000010001111101001110;
assign LUT_3[14977] = 32'b00000000000000011000101000101011;
assign LUT_3[14978] = 32'b00000000000000010100000100110010;
assign LUT_3[14979] = 32'b00000000000000011010110000001111;
assign LUT_3[14980] = 32'b00000000000000001111001011000100;
assign LUT_3[14981] = 32'b00000000000000010101110110100001;
assign LUT_3[14982] = 32'b00000000000000010001010010101000;
assign LUT_3[14983] = 32'b00000000000000010111111110000101;
assign LUT_3[14984] = 32'b00000000000000010111010110010100;
assign LUT_3[14985] = 32'b00000000000000011110000001110001;
assign LUT_3[14986] = 32'b00000000000000011001011101111000;
assign LUT_3[14987] = 32'b00000000000000100000001001010101;
assign LUT_3[14988] = 32'b00000000000000010100100100001010;
assign LUT_3[14989] = 32'b00000000000000011011001111100111;
assign LUT_3[14990] = 32'b00000000000000010110101011101110;
assign LUT_3[14991] = 32'b00000000000000011101010111001011;
assign LUT_3[14992] = 32'b00000000000000010101010000010001;
assign LUT_3[14993] = 32'b00000000000000011011111011101110;
assign LUT_3[14994] = 32'b00000000000000010111010111110101;
assign LUT_3[14995] = 32'b00000000000000011110000011010010;
assign LUT_3[14996] = 32'b00000000000000010010011110000111;
assign LUT_3[14997] = 32'b00000000000000011001001001100100;
assign LUT_3[14998] = 32'b00000000000000010100100101101011;
assign LUT_3[14999] = 32'b00000000000000011011010001001000;
assign LUT_3[15000] = 32'b00000000000000011010101001010111;
assign LUT_3[15001] = 32'b00000000000000100001010100110100;
assign LUT_3[15002] = 32'b00000000000000011100110000111011;
assign LUT_3[15003] = 32'b00000000000000100011011100011000;
assign LUT_3[15004] = 32'b00000000000000010111110111001101;
assign LUT_3[15005] = 32'b00000000000000011110100010101010;
assign LUT_3[15006] = 32'b00000000000000011001111110110001;
assign LUT_3[15007] = 32'b00000000000000100000101010001110;
assign LUT_3[15008] = 32'b00000000000000010011001011101110;
assign LUT_3[15009] = 32'b00000000000000011001110111001011;
assign LUT_3[15010] = 32'b00000000000000010101010011010010;
assign LUT_3[15011] = 32'b00000000000000011011111110101111;
assign LUT_3[15012] = 32'b00000000000000010000011001100100;
assign LUT_3[15013] = 32'b00000000000000010111000101000001;
assign LUT_3[15014] = 32'b00000000000000010010100001001000;
assign LUT_3[15015] = 32'b00000000000000011001001100100101;
assign LUT_3[15016] = 32'b00000000000000011000100100110100;
assign LUT_3[15017] = 32'b00000000000000011111010000010001;
assign LUT_3[15018] = 32'b00000000000000011010101100011000;
assign LUT_3[15019] = 32'b00000000000000100001010111110101;
assign LUT_3[15020] = 32'b00000000000000010101110010101010;
assign LUT_3[15021] = 32'b00000000000000011100011110000111;
assign LUT_3[15022] = 32'b00000000000000010111111010001110;
assign LUT_3[15023] = 32'b00000000000000011110100101101011;
assign LUT_3[15024] = 32'b00000000000000010110011110110001;
assign LUT_3[15025] = 32'b00000000000000011101001010001110;
assign LUT_3[15026] = 32'b00000000000000011000100110010101;
assign LUT_3[15027] = 32'b00000000000000011111010001110010;
assign LUT_3[15028] = 32'b00000000000000010011101100100111;
assign LUT_3[15029] = 32'b00000000000000011010011000000100;
assign LUT_3[15030] = 32'b00000000000000010101110100001011;
assign LUT_3[15031] = 32'b00000000000000011100011111101000;
assign LUT_3[15032] = 32'b00000000000000011011110111110111;
assign LUT_3[15033] = 32'b00000000000000100010100011010100;
assign LUT_3[15034] = 32'b00000000000000011101111111011011;
assign LUT_3[15035] = 32'b00000000000000100100101010111000;
assign LUT_3[15036] = 32'b00000000000000011001000101101101;
assign LUT_3[15037] = 32'b00000000000000011111110001001010;
assign LUT_3[15038] = 32'b00000000000000011011001101010001;
assign LUT_3[15039] = 32'b00000000000000100001111000101110;
assign LUT_3[15040] = 32'b00000000000000010001110101111001;
assign LUT_3[15041] = 32'b00000000000000011000100001010110;
assign LUT_3[15042] = 32'b00000000000000010011111101011101;
assign LUT_3[15043] = 32'b00000000000000011010101000111010;
assign LUT_3[15044] = 32'b00000000000000001111000011101111;
assign LUT_3[15045] = 32'b00000000000000010101101111001100;
assign LUT_3[15046] = 32'b00000000000000010001001011010011;
assign LUT_3[15047] = 32'b00000000000000010111110110110000;
assign LUT_3[15048] = 32'b00000000000000010111001110111111;
assign LUT_3[15049] = 32'b00000000000000011101111010011100;
assign LUT_3[15050] = 32'b00000000000000011001010110100011;
assign LUT_3[15051] = 32'b00000000000000100000000010000000;
assign LUT_3[15052] = 32'b00000000000000010100011100110101;
assign LUT_3[15053] = 32'b00000000000000011011001000010010;
assign LUT_3[15054] = 32'b00000000000000010110100100011001;
assign LUT_3[15055] = 32'b00000000000000011101001111110110;
assign LUT_3[15056] = 32'b00000000000000010101001000111100;
assign LUT_3[15057] = 32'b00000000000000011011110100011001;
assign LUT_3[15058] = 32'b00000000000000010111010000100000;
assign LUT_3[15059] = 32'b00000000000000011101111011111101;
assign LUT_3[15060] = 32'b00000000000000010010010110110010;
assign LUT_3[15061] = 32'b00000000000000011001000010001111;
assign LUT_3[15062] = 32'b00000000000000010100011110010110;
assign LUT_3[15063] = 32'b00000000000000011011001001110011;
assign LUT_3[15064] = 32'b00000000000000011010100010000010;
assign LUT_3[15065] = 32'b00000000000000100001001101011111;
assign LUT_3[15066] = 32'b00000000000000011100101001100110;
assign LUT_3[15067] = 32'b00000000000000100011010101000011;
assign LUT_3[15068] = 32'b00000000000000010111101111111000;
assign LUT_3[15069] = 32'b00000000000000011110011011010101;
assign LUT_3[15070] = 32'b00000000000000011001110111011100;
assign LUT_3[15071] = 32'b00000000000000100000100010111001;
assign LUT_3[15072] = 32'b00000000000000010011000100011001;
assign LUT_3[15073] = 32'b00000000000000011001101111110110;
assign LUT_3[15074] = 32'b00000000000000010101001011111101;
assign LUT_3[15075] = 32'b00000000000000011011110111011010;
assign LUT_3[15076] = 32'b00000000000000010000010010001111;
assign LUT_3[15077] = 32'b00000000000000010110111101101100;
assign LUT_3[15078] = 32'b00000000000000010010011001110011;
assign LUT_3[15079] = 32'b00000000000000011001000101010000;
assign LUT_3[15080] = 32'b00000000000000011000011101011111;
assign LUT_3[15081] = 32'b00000000000000011111001000111100;
assign LUT_3[15082] = 32'b00000000000000011010100101000011;
assign LUT_3[15083] = 32'b00000000000000100001010000100000;
assign LUT_3[15084] = 32'b00000000000000010101101011010101;
assign LUT_3[15085] = 32'b00000000000000011100010110110010;
assign LUT_3[15086] = 32'b00000000000000010111110010111001;
assign LUT_3[15087] = 32'b00000000000000011110011110010110;
assign LUT_3[15088] = 32'b00000000000000010110010111011100;
assign LUT_3[15089] = 32'b00000000000000011101000010111001;
assign LUT_3[15090] = 32'b00000000000000011000011111000000;
assign LUT_3[15091] = 32'b00000000000000011111001010011101;
assign LUT_3[15092] = 32'b00000000000000010011100101010010;
assign LUT_3[15093] = 32'b00000000000000011010010000101111;
assign LUT_3[15094] = 32'b00000000000000010101101100110110;
assign LUT_3[15095] = 32'b00000000000000011100011000010011;
assign LUT_3[15096] = 32'b00000000000000011011110000100010;
assign LUT_3[15097] = 32'b00000000000000100010011011111111;
assign LUT_3[15098] = 32'b00000000000000011101111000000110;
assign LUT_3[15099] = 32'b00000000000000100100100011100011;
assign LUT_3[15100] = 32'b00000000000000011000111110011000;
assign LUT_3[15101] = 32'b00000000000000011111101001110101;
assign LUT_3[15102] = 32'b00000000000000011011000101111100;
assign LUT_3[15103] = 32'b00000000000000100001110001011001;
assign LUT_3[15104] = 32'b00000000000000001100000001110001;
assign LUT_3[15105] = 32'b00000000000000010010101101001110;
assign LUT_3[15106] = 32'b00000000000000001110001001010101;
assign LUT_3[15107] = 32'b00000000000000010100110100110010;
assign LUT_3[15108] = 32'b00000000000000001001001111100111;
assign LUT_3[15109] = 32'b00000000000000001111111011000100;
assign LUT_3[15110] = 32'b00000000000000001011010111001011;
assign LUT_3[15111] = 32'b00000000000000010010000010101000;
assign LUT_3[15112] = 32'b00000000000000010001011010110111;
assign LUT_3[15113] = 32'b00000000000000011000000110010100;
assign LUT_3[15114] = 32'b00000000000000010011100010011011;
assign LUT_3[15115] = 32'b00000000000000011010001101111000;
assign LUT_3[15116] = 32'b00000000000000001110101000101101;
assign LUT_3[15117] = 32'b00000000000000010101010100001010;
assign LUT_3[15118] = 32'b00000000000000010000110000010001;
assign LUT_3[15119] = 32'b00000000000000010111011011101110;
assign LUT_3[15120] = 32'b00000000000000001111010100110100;
assign LUT_3[15121] = 32'b00000000000000010110000000010001;
assign LUT_3[15122] = 32'b00000000000000010001011100011000;
assign LUT_3[15123] = 32'b00000000000000011000000111110101;
assign LUT_3[15124] = 32'b00000000000000001100100010101010;
assign LUT_3[15125] = 32'b00000000000000010011001110000111;
assign LUT_3[15126] = 32'b00000000000000001110101010001110;
assign LUT_3[15127] = 32'b00000000000000010101010101101011;
assign LUT_3[15128] = 32'b00000000000000010100101101111010;
assign LUT_3[15129] = 32'b00000000000000011011011001010111;
assign LUT_3[15130] = 32'b00000000000000010110110101011110;
assign LUT_3[15131] = 32'b00000000000000011101100000111011;
assign LUT_3[15132] = 32'b00000000000000010001111011110000;
assign LUT_3[15133] = 32'b00000000000000011000100111001101;
assign LUT_3[15134] = 32'b00000000000000010100000011010100;
assign LUT_3[15135] = 32'b00000000000000011010101110110001;
assign LUT_3[15136] = 32'b00000000000000001101010000010001;
assign LUT_3[15137] = 32'b00000000000000010011111011101110;
assign LUT_3[15138] = 32'b00000000000000001111010111110101;
assign LUT_3[15139] = 32'b00000000000000010110000011010010;
assign LUT_3[15140] = 32'b00000000000000001010011110000111;
assign LUT_3[15141] = 32'b00000000000000010001001001100100;
assign LUT_3[15142] = 32'b00000000000000001100100101101011;
assign LUT_3[15143] = 32'b00000000000000010011010001001000;
assign LUT_3[15144] = 32'b00000000000000010010101001010111;
assign LUT_3[15145] = 32'b00000000000000011001010100110100;
assign LUT_3[15146] = 32'b00000000000000010100110000111011;
assign LUT_3[15147] = 32'b00000000000000011011011100011000;
assign LUT_3[15148] = 32'b00000000000000001111110111001101;
assign LUT_3[15149] = 32'b00000000000000010110100010101010;
assign LUT_3[15150] = 32'b00000000000000010001111110110001;
assign LUT_3[15151] = 32'b00000000000000011000101010001110;
assign LUT_3[15152] = 32'b00000000000000010000100011010100;
assign LUT_3[15153] = 32'b00000000000000010111001110110001;
assign LUT_3[15154] = 32'b00000000000000010010101010111000;
assign LUT_3[15155] = 32'b00000000000000011001010110010101;
assign LUT_3[15156] = 32'b00000000000000001101110001001010;
assign LUT_3[15157] = 32'b00000000000000010100011100100111;
assign LUT_3[15158] = 32'b00000000000000001111111000101110;
assign LUT_3[15159] = 32'b00000000000000010110100100001011;
assign LUT_3[15160] = 32'b00000000000000010101111100011010;
assign LUT_3[15161] = 32'b00000000000000011100100111110111;
assign LUT_3[15162] = 32'b00000000000000011000000011111110;
assign LUT_3[15163] = 32'b00000000000000011110101111011011;
assign LUT_3[15164] = 32'b00000000000000010011001010010000;
assign LUT_3[15165] = 32'b00000000000000011001110101101101;
assign LUT_3[15166] = 32'b00000000000000010101010001110100;
assign LUT_3[15167] = 32'b00000000000000011011111101010001;
assign LUT_3[15168] = 32'b00000000000000001011111010011100;
assign LUT_3[15169] = 32'b00000000000000010010100101111001;
assign LUT_3[15170] = 32'b00000000000000001110000010000000;
assign LUT_3[15171] = 32'b00000000000000010100101101011101;
assign LUT_3[15172] = 32'b00000000000000001001001000010010;
assign LUT_3[15173] = 32'b00000000000000001111110011101111;
assign LUT_3[15174] = 32'b00000000000000001011001111110110;
assign LUT_3[15175] = 32'b00000000000000010001111011010011;
assign LUT_3[15176] = 32'b00000000000000010001010011100010;
assign LUT_3[15177] = 32'b00000000000000010111111110111111;
assign LUT_3[15178] = 32'b00000000000000010011011011000110;
assign LUT_3[15179] = 32'b00000000000000011010000110100011;
assign LUT_3[15180] = 32'b00000000000000001110100001011000;
assign LUT_3[15181] = 32'b00000000000000010101001100110101;
assign LUT_3[15182] = 32'b00000000000000010000101000111100;
assign LUT_3[15183] = 32'b00000000000000010111010100011001;
assign LUT_3[15184] = 32'b00000000000000001111001101011111;
assign LUT_3[15185] = 32'b00000000000000010101111000111100;
assign LUT_3[15186] = 32'b00000000000000010001010101000011;
assign LUT_3[15187] = 32'b00000000000000011000000000100000;
assign LUT_3[15188] = 32'b00000000000000001100011011010101;
assign LUT_3[15189] = 32'b00000000000000010011000110110010;
assign LUT_3[15190] = 32'b00000000000000001110100010111001;
assign LUT_3[15191] = 32'b00000000000000010101001110010110;
assign LUT_3[15192] = 32'b00000000000000010100100110100101;
assign LUT_3[15193] = 32'b00000000000000011011010010000010;
assign LUT_3[15194] = 32'b00000000000000010110101110001001;
assign LUT_3[15195] = 32'b00000000000000011101011001100110;
assign LUT_3[15196] = 32'b00000000000000010001110100011011;
assign LUT_3[15197] = 32'b00000000000000011000011111111000;
assign LUT_3[15198] = 32'b00000000000000010011111011111111;
assign LUT_3[15199] = 32'b00000000000000011010100111011100;
assign LUT_3[15200] = 32'b00000000000000001101001000111100;
assign LUT_3[15201] = 32'b00000000000000010011110100011001;
assign LUT_3[15202] = 32'b00000000000000001111010000100000;
assign LUT_3[15203] = 32'b00000000000000010101111011111101;
assign LUT_3[15204] = 32'b00000000000000001010010110110010;
assign LUT_3[15205] = 32'b00000000000000010001000010001111;
assign LUT_3[15206] = 32'b00000000000000001100011110010110;
assign LUT_3[15207] = 32'b00000000000000010011001001110011;
assign LUT_3[15208] = 32'b00000000000000010010100010000010;
assign LUT_3[15209] = 32'b00000000000000011001001101011111;
assign LUT_3[15210] = 32'b00000000000000010100101001100110;
assign LUT_3[15211] = 32'b00000000000000011011010101000011;
assign LUT_3[15212] = 32'b00000000000000001111101111111000;
assign LUT_3[15213] = 32'b00000000000000010110011011010101;
assign LUT_3[15214] = 32'b00000000000000010001110111011100;
assign LUT_3[15215] = 32'b00000000000000011000100010111001;
assign LUT_3[15216] = 32'b00000000000000010000011011111111;
assign LUT_3[15217] = 32'b00000000000000010111000111011100;
assign LUT_3[15218] = 32'b00000000000000010010100011100011;
assign LUT_3[15219] = 32'b00000000000000011001001111000000;
assign LUT_3[15220] = 32'b00000000000000001101101001110101;
assign LUT_3[15221] = 32'b00000000000000010100010101010010;
assign LUT_3[15222] = 32'b00000000000000001111110001011001;
assign LUT_3[15223] = 32'b00000000000000010110011100110110;
assign LUT_3[15224] = 32'b00000000000000010101110101000101;
assign LUT_3[15225] = 32'b00000000000000011100100000100010;
assign LUT_3[15226] = 32'b00000000000000010111111100101001;
assign LUT_3[15227] = 32'b00000000000000011110101000000110;
assign LUT_3[15228] = 32'b00000000000000010011000010111011;
assign LUT_3[15229] = 32'b00000000000000011001101110011000;
assign LUT_3[15230] = 32'b00000000000000010101001010011111;
assign LUT_3[15231] = 32'b00000000000000011011110101111100;
assign LUT_3[15232] = 32'b00000000000000001110001100101111;
assign LUT_3[15233] = 32'b00000000000000010100111000001100;
assign LUT_3[15234] = 32'b00000000000000010000010100010011;
assign LUT_3[15235] = 32'b00000000000000010110111111110000;
assign LUT_3[15236] = 32'b00000000000000001011011010100101;
assign LUT_3[15237] = 32'b00000000000000010010000110000010;
assign LUT_3[15238] = 32'b00000000000000001101100010001001;
assign LUT_3[15239] = 32'b00000000000000010100001101100110;
assign LUT_3[15240] = 32'b00000000000000010011100101110101;
assign LUT_3[15241] = 32'b00000000000000011010010001010010;
assign LUT_3[15242] = 32'b00000000000000010101101101011001;
assign LUT_3[15243] = 32'b00000000000000011100011000110110;
assign LUT_3[15244] = 32'b00000000000000010000110011101011;
assign LUT_3[15245] = 32'b00000000000000010111011111001000;
assign LUT_3[15246] = 32'b00000000000000010010111011001111;
assign LUT_3[15247] = 32'b00000000000000011001100110101100;
assign LUT_3[15248] = 32'b00000000000000010001011111110010;
assign LUT_3[15249] = 32'b00000000000000011000001011001111;
assign LUT_3[15250] = 32'b00000000000000010011100111010110;
assign LUT_3[15251] = 32'b00000000000000011010010010110011;
assign LUT_3[15252] = 32'b00000000000000001110101101101000;
assign LUT_3[15253] = 32'b00000000000000010101011001000101;
assign LUT_3[15254] = 32'b00000000000000010000110101001100;
assign LUT_3[15255] = 32'b00000000000000010111100000101001;
assign LUT_3[15256] = 32'b00000000000000010110111000111000;
assign LUT_3[15257] = 32'b00000000000000011101100100010101;
assign LUT_3[15258] = 32'b00000000000000011001000000011100;
assign LUT_3[15259] = 32'b00000000000000011111101011111001;
assign LUT_3[15260] = 32'b00000000000000010100000110101110;
assign LUT_3[15261] = 32'b00000000000000011010110010001011;
assign LUT_3[15262] = 32'b00000000000000010110001110010010;
assign LUT_3[15263] = 32'b00000000000000011100111001101111;
assign LUT_3[15264] = 32'b00000000000000001111011011001111;
assign LUT_3[15265] = 32'b00000000000000010110000110101100;
assign LUT_3[15266] = 32'b00000000000000010001100010110011;
assign LUT_3[15267] = 32'b00000000000000011000001110010000;
assign LUT_3[15268] = 32'b00000000000000001100101001000101;
assign LUT_3[15269] = 32'b00000000000000010011010100100010;
assign LUT_3[15270] = 32'b00000000000000001110110000101001;
assign LUT_3[15271] = 32'b00000000000000010101011100000110;
assign LUT_3[15272] = 32'b00000000000000010100110100010101;
assign LUT_3[15273] = 32'b00000000000000011011011111110010;
assign LUT_3[15274] = 32'b00000000000000010110111011111001;
assign LUT_3[15275] = 32'b00000000000000011101100111010110;
assign LUT_3[15276] = 32'b00000000000000010010000010001011;
assign LUT_3[15277] = 32'b00000000000000011000101101101000;
assign LUT_3[15278] = 32'b00000000000000010100001001101111;
assign LUT_3[15279] = 32'b00000000000000011010110101001100;
assign LUT_3[15280] = 32'b00000000000000010010101110010010;
assign LUT_3[15281] = 32'b00000000000000011001011001101111;
assign LUT_3[15282] = 32'b00000000000000010100110101110110;
assign LUT_3[15283] = 32'b00000000000000011011100001010011;
assign LUT_3[15284] = 32'b00000000000000001111111100001000;
assign LUT_3[15285] = 32'b00000000000000010110100111100101;
assign LUT_3[15286] = 32'b00000000000000010010000011101100;
assign LUT_3[15287] = 32'b00000000000000011000101111001001;
assign LUT_3[15288] = 32'b00000000000000011000000111011000;
assign LUT_3[15289] = 32'b00000000000000011110110010110101;
assign LUT_3[15290] = 32'b00000000000000011010001110111100;
assign LUT_3[15291] = 32'b00000000000000100000111010011001;
assign LUT_3[15292] = 32'b00000000000000010101010101001110;
assign LUT_3[15293] = 32'b00000000000000011100000000101011;
assign LUT_3[15294] = 32'b00000000000000010111011100110010;
assign LUT_3[15295] = 32'b00000000000000011110001000001111;
assign LUT_3[15296] = 32'b00000000000000001110000101011010;
assign LUT_3[15297] = 32'b00000000000000010100110000110111;
assign LUT_3[15298] = 32'b00000000000000010000001100111110;
assign LUT_3[15299] = 32'b00000000000000010110111000011011;
assign LUT_3[15300] = 32'b00000000000000001011010011010000;
assign LUT_3[15301] = 32'b00000000000000010001111110101101;
assign LUT_3[15302] = 32'b00000000000000001101011010110100;
assign LUT_3[15303] = 32'b00000000000000010100000110010001;
assign LUT_3[15304] = 32'b00000000000000010011011110100000;
assign LUT_3[15305] = 32'b00000000000000011010001001111101;
assign LUT_3[15306] = 32'b00000000000000010101100110000100;
assign LUT_3[15307] = 32'b00000000000000011100010001100001;
assign LUT_3[15308] = 32'b00000000000000010000101100010110;
assign LUT_3[15309] = 32'b00000000000000010111010111110011;
assign LUT_3[15310] = 32'b00000000000000010010110011111010;
assign LUT_3[15311] = 32'b00000000000000011001011111010111;
assign LUT_3[15312] = 32'b00000000000000010001011000011101;
assign LUT_3[15313] = 32'b00000000000000011000000011111010;
assign LUT_3[15314] = 32'b00000000000000010011100000000001;
assign LUT_3[15315] = 32'b00000000000000011010001011011110;
assign LUT_3[15316] = 32'b00000000000000001110100110010011;
assign LUT_3[15317] = 32'b00000000000000010101010001110000;
assign LUT_3[15318] = 32'b00000000000000010000101101110111;
assign LUT_3[15319] = 32'b00000000000000010111011001010100;
assign LUT_3[15320] = 32'b00000000000000010110110001100011;
assign LUT_3[15321] = 32'b00000000000000011101011101000000;
assign LUT_3[15322] = 32'b00000000000000011000111001000111;
assign LUT_3[15323] = 32'b00000000000000011111100100100100;
assign LUT_3[15324] = 32'b00000000000000010011111111011001;
assign LUT_3[15325] = 32'b00000000000000011010101010110110;
assign LUT_3[15326] = 32'b00000000000000010110000110111101;
assign LUT_3[15327] = 32'b00000000000000011100110010011010;
assign LUT_3[15328] = 32'b00000000000000001111010011111010;
assign LUT_3[15329] = 32'b00000000000000010101111111010111;
assign LUT_3[15330] = 32'b00000000000000010001011011011110;
assign LUT_3[15331] = 32'b00000000000000011000000110111011;
assign LUT_3[15332] = 32'b00000000000000001100100001110000;
assign LUT_3[15333] = 32'b00000000000000010011001101001101;
assign LUT_3[15334] = 32'b00000000000000001110101001010100;
assign LUT_3[15335] = 32'b00000000000000010101010100110001;
assign LUT_3[15336] = 32'b00000000000000010100101101000000;
assign LUT_3[15337] = 32'b00000000000000011011011000011101;
assign LUT_3[15338] = 32'b00000000000000010110110100100100;
assign LUT_3[15339] = 32'b00000000000000011101100000000001;
assign LUT_3[15340] = 32'b00000000000000010001111010110110;
assign LUT_3[15341] = 32'b00000000000000011000100110010011;
assign LUT_3[15342] = 32'b00000000000000010100000010011010;
assign LUT_3[15343] = 32'b00000000000000011010101101110111;
assign LUT_3[15344] = 32'b00000000000000010010100110111101;
assign LUT_3[15345] = 32'b00000000000000011001010010011010;
assign LUT_3[15346] = 32'b00000000000000010100101110100001;
assign LUT_3[15347] = 32'b00000000000000011011011001111110;
assign LUT_3[15348] = 32'b00000000000000001111110100110011;
assign LUT_3[15349] = 32'b00000000000000010110100000010000;
assign LUT_3[15350] = 32'b00000000000000010001111100010111;
assign LUT_3[15351] = 32'b00000000000000011000100111110100;
assign LUT_3[15352] = 32'b00000000000000011000000000000011;
assign LUT_3[15353] = 32'b00000000000000011110101011100000;
assign LUT_3[15354] = 32'b00000000000000011010000111100111;
assign LUT_3[15355] = 32'b00000000000000100000110011000100;
assign LUT_3[15356] = 32'b00000000000000010101001101111001;
assign LUT_3[15357] = 32'b00000000000000011011111001010110;
assign LUT_3[15358] = 32'b00000000000000010111010101011101;
assign LUT_3[15359] = 32'b00000000000000011110000000111010;
assign LUT_3[15360] = 32'b00000000000000010011000010000001;
assign LUT_3[15361] = 32'b00000000000000011001101101011110;
assign LUT_3[15362] = 32'b00000000000000010101001001100101;
assign LUT_3[15363] = 32'b00000000000000011011110101000010;
assign LUT_3[15364] = 32'b00000000000000010000001111110111;
assign LUT_3[15365] = 32'b00000000000000010110111011010100;
assign LUT_3[15366] = 32'b00000000000000010010010111011011;
assign LUT_3[15367] = 32'b00000000000000011001000010111000;
assign LUT_3[15368] = 32'b00000000000000011000011011000111;
assign LUT_3[15369] = 32'b00000000000000011111000110100100;
assign LUT_3[15370] = 32'b00000000000000011010100010101011;
assign LUT_3[15371] = 32'b00000000000000100001001110001000;
assign LUT_3[15372] = 32'b00000000000000010101101000111101;
assign LUT_3[15373] = 32'b00000000000000011100010100011010;
assign LUT_3[15374] = 32'b00000000000000010111110000100001;
assign LUT_3[15375] = 32'b00000000000000011110011011111110;
assign LUT_3[15376] = 32'b00000000000000010110010101000100;
assign LUT_3[15377] = 32'b00000000000000011101000000100001;
assign LUT_3[15378] = 32'b00000000000000011000011100101000;
assign LUT_3[15379] = 32'b00000000000000011111001000000101;
assign LUT_3[15380] = 32'b00000000000000010011100010111010;
assign LUT_3[15381] = 32'b00000000000000011010001110010111;
assign LUT_3[15382] = 32'b00000000000000010101101010011110;
assign LUT_3[15383] = 32'b00000000000000011100010101111011;
assign LUT_3[15384] = 32'b00000000000000011011101110001010;
assign LUT_3[15385] = 32'b00000000000000100010011001100111;
assign LUT_3[15386] = 32'b00000000000000011101110101101110;
assign LUT_3[15387] = 32'b00000000000000100100100001001011;
assign LUT_3[15388] = 32'b00000000000000011000111100000000;
assign LUT_3[15389] = 32'b00000000000000011111100111011101;
assign LUT_3[15390] = 32'b00000000000000011011000011100100;
assign LUT_3[15391] = 32'b00000000000000100001101111000001;
assign LUT_3[15392] = 32'b00000000000000010100010000100001;
assign LUT_3[15393] = 32'b00000000000000011010111011111110;
assign LUT_3[15394] = 32'b00000000000000010110011000000101;
assign LUT_3[15395] = 32'b00000000000000011101000011100010;
assign LUT_3[15396] = 32'b00000000000000010001011110010111;
assign LUT_3[15397] = 32'b00000000000000011000001001110100;
assign LUT_3[15398] = 32'b00000000000000010011100101111011;
assign LUT_3[15399] = 32'b00000000000000011010010001011000;
assign LUT_3[15400] = 32'b00000000000000011001101001100111;
assign LUT_3[15401] = 32'b00000000000000100000010101000100;
assign LUT_3[15402] = 32'b00000000000000011011110001001011;
assign LUT_3[15403] = 32'b00000000000000100010011100101000;
assign LUT_3[15404] = 32'b00000000000000010110110111011101;
assign LUT_3[15405] = 32'b00000000000000011101100010111010;
assign LUT_3[15406] = 32'b00000000000000011000111111000001;
assign LUT_3[15407] = 32'b00000000000000011111101010011110;
assign LUT_3[15408] = 32'b00000000000000010111100011100100;
assign LUT_3[15409] = 32'b00000000000000011110001111000001;
assign LUT_3[15410] = 32'b00000000000000011001101011001000;
assign LUT_3[15411] = 32'b00000000000000100000010110100101;
assign LUT_3[15412] = 32'b00000000000000010100110001011010;
assign LUT_3[15413] = 32'b00000000000000011011011100110111;
assign LUT_3[15414] = 32'b00000000000000010110111000111110;
assign LUT_3[15415] = 32'b00000000000000011101100100011011;
assign LUT_3[15416] = 32'b00000000000000011100111100101010;
assign LUT_3[15417] = 32'b00000000000000100011101000000111;
assign LUT_3[15418] = 32'b00000000000000011111000100001110;
assign LUT_3[15419] = 32'b00000000000000100101101111101011;
assign LUT_3[15420] = 32'b00000000000000011010001010100000;
assign LUT_3[15421] = 32'b00000000000000100000110101111101;
assign LUT_3[15422] = 32'b00000000000000011100010010000100;
assign LUT_3[15423] = 32'b00000000000000100010111101100001;
assign LUT_3[15424] = 32'b00000000000000010010111010101100;
assign LUT_3[15425] = 32'b00000000000000011001100110001001;
assign LUT_3[15426] = 32'b00000000000000010101000010010000;
assign LUT_3[15427] = 32'b00000000000000011011101101101101;
assign LUT_3[15428] = 32'b00000000000000010000001000100010;
assign LUT_3[15429] = 32'b00000000000000010110110011111111;
assign LUT_3[15430] = 32'b00000000000000010010010000000110;
assign LUT_3[15431] = 32'b00000000000000011000111011100011;
assign LUT_3[15432] = 32'b00000000000000011000010011110010;
assign LUT_3[15433] = 32'b00000000000000011110111111001111;
assign LUT_3[15434] = 32'b00000000000000011010011011010110;
assign LUT_3[15435] = 32'b00000000000000100001000110110011;
assign LUT_3[15436] = 32'b00000000000000010101100001101000;
assign LUT_3[15437] = 32'b00000000000000011100001101000101;
assign LUT_3[15438] = 32'b00000000000000010111101001001100;
assign LUT_3[15439] = 32'b00000000000000011110010100101001;
assign LUT_3[15440] = 32'b00000000000000010110001101101111;
assign LUT_3[15441] = 32'b00000000000000011100111001001100;
assign LUT_3[15442] = 32'b00000000000000011000010101010011;
assign LUT_3[15443] = 32'b00000000000000011111000000110000;
assign LUT_3[15444] = 32'b00000000000000010011011011100101;
assign LUT_3[15445] = 32'b00000000000000011010000111000010;
assign LUT_3[15446] = 32'b00000000000000010101100011001001;
assign LUT_3[15447] = 32'b00000000000000011100001110100110;
assign LUT_3[15448] = 32'b00000000000000011011100110110101;
assign LUT_3[15449] = 32'b00000000000000100010010010010010;
assign LUT_3[15450] = 32'b00000000000000011101101110011001;
assign LUT_3[15451] = 32'b00000000000000100100011001110110;
assign LUT_3[15452] = 32'b00000000000000011000110100101011;
assign LUT_3[15453] = 32'b00000000000000011111100000001000;
assign LUT_3[15454] = 32'b00000000000000011010111100001111;
assign LUT_3[15455] = 32'b00000000000000100001100111101100;
assign LUT_3[15456] = 32'b00000000000000010100001001001100;
assign LUT_3[15457] = 32'b00000000000000011010110100101001;
assign LUT_3[15458] = 32'b00000000000000010110010000110000;
assign LUT_3[15459] = 32'b00000000000000011100111100001101;
assign LUT_3[15460] = 32'b00000000000000010001010111000010;
assign LUT_3[15461] = 32'b00000000000000011000000010011111;
assign LUT_3[15462] = 32'b00000000000000010011011110100110;
assign LUT_3[15463] = 32'b00000000000000011010001010000011;
assign LUT_3[15464] = 32'b00000000000000011001100010010010;
assign LUT_3[15465] = 32'b00000000000000100000001101101111;
assign LUT_3[15466] = 32'b00000000000000011011101001110110;
assign LUT_3[15467] = 32'b00000000000000100010010101010011;
assign LUT_3[15468] = 32'b00000000000000010110110000001000;
assign LUT_3[15469] = 32'b00000000000000011101011011100101;
assign LUT_3[15470] = 32'b00000000000000011000110111101100;
assign LUT_3[15471] = 32'b00000000000000011111100011001001;
assign LUT_3[15472] = 32'b00000000000000010111011100001111;
assign LUT_3[15473] = 32'b00000000000000011110000111101100;
assign LUT_3[15474] = 32'b00000000000000011001100011110011;
assign LUT_3[15475] = 32'b00000000000000100000001111010000;
assign LUT_3[15476] = 32'b00000000000000010100101010000101;
assign LUT_3[15477] = 32'b00000000000000011011010101100010;
assign LUT_3[15478] = 32'b00000000000000010110110001101001;
assign LUT_3[15479] = 32'b00000000000000011101011101000110;
assign LUT_3[15480] = 32'b00000000000000011100110101010101;
assign LUT_3[15481] = 32'b00000000000000100011100000110010;
assign LUT_3[15482] = 32'b00000000000000011110111100111001;
assign LUT_3[15483] = 32'b00000000000000100101101000010110;
assign LUT_3[15484] = 32'b00000000000000011010000011001011;
assign LUT_3[15485] = 32'b00000000000000100000101110101000;
assign LUT_3[15486] = 32'b00000000000000011100001010101111;
assign LUT_3[15487] = 32'b00000000000000100010110110001100;
assign LUT_3[15488] = 32'b00000000000000010101001100111111;
assign LUT_3[15489] = 32'b00000000000000011011111000011100;
assign LUT_3[15490] = 32'b00000000000000010111010100100011;
assign LUT_3[15491] = 32'b00000000000000011110000000000000;
assign LUT_3[15492] = 32'b00000000000000010010011010110101;
assign LUT_3[15493] = 32'b00000000000000011001000110010010;
assign LUT_3[15494] = 32'b00000000000000010100100010011001;
assign LUT_3[15495] = 32'b00000000000000011011001101110110;
assign LUT_3[15496] = 32'b00000000000000011010100110000101;
assign LUT_3[15497] = 32'b00000000000000100001010001100010;
assign LUT_3[15498] = 32'b00000000000000011100101101101001;
assign LUT_3[15499] = 32'b00000000000000100011011001000110;
assign LUT_3[15500] = 32'b00000000000000010111110011111011;
assign LUT_3[15501] = 32'b00000000000000011110011111011000;
assign LUT_3[15502] = 32'b00000000000000011001111011011111;
assign LUT_3[15503] = 32'b00000000000000100000100110111100;
assign LUT_3[15504] = 32'b00000000000000011000100000000010;
assign LUT_3[15505] = 32'b00000000000000011111001011011111;
assign LUT_3[15506] = 32'b00000000000000011010100111100110;
assign LUT_3[15507] = 32'b00000000000000100001010011000011;
assign LUT_3[15508] = 32'b00000000000000010101101101111000;
assign LUT_3[15509] = 32'b00000000000000011100011001010101;
assign LUT_3[15510] = 32'b00000000000000010111110101011100;
assign LUT_3[15511] = 32'b00000000000000011110100000111001;
assign LUT_3[15512] = 32'b00000000000000011101111001001000;
assign LUT_3[15513] = 32'b00000000000000100100100100100101;
assign LUT_3[15514] = 32'b00000000000000100000000000101100;
assign LUT_3[15515] = 32'b00000000000000100110101100001001;
assign LUT_3[15516] = 32'b00000000000000011011000110111110;
assign LUT_3[15517] = 32'b00000000000000100001110010011011;
assign LUT_3[15518] = 32'b00000000000000011101001110100010;
assign LUT_3[15519] = 32'b00000000000000100011111001111111;
assign LUT_3[15520] = 32'b00000000000000010110011011011111;
assign LUT_3[15521] = 32'b00000000000000011101000110111100;
assign LUT_3[15522] = 32'b00000000000000011000100011000011;
assign LUT_3[15523] = 32'b00000000000000011111001110100000;
assign LUT_3[15524] = 32'b00000000000000010011101001010101;
assign LUT_3[15525] = 32'b00000000000000011010010100110010;
assign LUT_3[15526] = 32'b00000000000000010101110000111001;
assign LUT_3[15527] = 32'b00000000000000011100011100010110;
assign LUT_3[15528] = 32'b00000000000000011011110100100101;
assign LUT_3[15529] = 32'b00000000000000100010100000000010;
assign LUT_3[15530] = 32'b00000000000000011101111100001001;
assign LUT_3[15531] = 32'b00000000000000100100100111100110;
assign LUT_3[15532] = 32'b00000000000000011001000010011011;
assign LUT_3[15533] = 32'b00000000000000011111101101111000;
assign LUT_3[15534] = 32'b00000000000000011011001001111111;
assign LUT_3[15535] = 32'b00000000000000100001110101011100;
assign LUT_3[15536] = 32'b00000000000000011001101110100010;
assign LUT_3[15537] = 32'b00000000000000100000011001111111;
assign LUT_3[15538] = 32'b00000000000000011011110110000110;
assign LUT_3[15539] = 32'b00000000000000100010100001100011;
assign LUT_3[15540] = 32'b00000000000000010110111100011000;
assign LUT_3[15541] = 32'b00000000000000011101100111110101;
assign LUT_3[15542] = 32'b00000000000000011001000011111100;
assign LUT_3[15543] = 32'b00000000000000011111101111011001;
assign LUT_3[15544] = 32'b00000000000000011111000111101000;
assign LUT_3[15545] = 32'b00000000000000100101110011000101;
assign LUT_3[15546] = 32'b00000000000000100001001111001100;
assign LUT_3[15547] = 32'b00000000000000100111111010101001;
assign LUT_3[15548] = 32'b00000000000000011100010101011110;
assign LUT_3[15549] = 32'b00000000000000100011000000111011;
assign LUT_3[15550] = 32'b00000000000000011110011101000010;
assign LUT_3[15551] = 32'b00000000000000100101001000011111;
assign LUT_3[15552] = 32'b00000000000000010101000101101010;
assign LUT_3[15553] = 32'b00000000000000011011110001000111;
assign LUT_3[15554] = 32'b00000000000000010111001101001110;
assign LUT_3[15555] = 32'b00000000000000011101111000101011;
assign LUT_3[15556] = 32'b00000000000000010010010011100000;
assign LUT_3[15557] = 32'b00000000000000011000111110111101;
assign LUT_3[15558] = 32'b00000000000000010100011011000100;
assign LUT_3[15559] = 32'b00000000000000011011000110100001;
assign LUT_3[15560] = 32'b00000000000000011010011110110000;
assign LUT_3[15561] = 32'b00000000000000100001001010001101;
assign LUT_3[15562] = 32'b00000000000000011100100110010100;
assign LUT_3[15563] = 32'b00000000000000100011010001110001;
assign LUT_3[15564] = 32'b00000000000000010111101100100110;
assign LUT_3[15565] = 32'b00000000000000011110011000000011;
assign LUT_3[15566] = 32'b00000000000000011001110100001010;
assign LUT_3[15567] = 32'b00000000000000100000011111100111;
assign LUT_3[15568] = 32'b00000000000000011000011000101101;
assign LUT_3[15569] = 32'b00000000000000011111000100001010;
assign LUT_3[15570] = 32'b00000000000000011010100000010001;
assign LUT_3[15571] = 32'b00000000000000100001001011101110;
assign LUT_3[15572] = 32'b00000000000000010101100110100011;
assign LUT_3[15573] = 32'b00000000000000011100010010000000;
assign LUT_3[15574] = 32'b00000000000000010111101110000111;
assign LUT_3[15575] = 32'b00000000000000011110011001100100;
assign LUT_3[15576] = 32'b00000000000000011101110001110011;
assign LUT_3[15577] = 32'b00000000000000100100011101010000;
assign LUT_3[15578] = 32'b00000000000000011111111001010111;
assign LUT_3[15579] = 32'b00000000000000100110100100110100;
assign LUT_3[15580] = 32'b00000000000000011010111111101001;
assign LUT_3[15581] = 32'b00000000000000100001101011000110;
assign LUT_3[15582] = 32'b00000000000000011101000111001101;
assign LUT_3[15583] = 32'b00000000000000100011110010101010;
assign LUT_3[15584] = 32'b00000000000000010110010100001010;
assign LUT_3[15585] = 32'b00000000000000011100111111100111;
assign LUT_3[15586] = 32'b00000000000000011000011011101110;
assign LUT_3[15587] = 32'b00000000000000011111000111001011;
assign LUT_3[15588] = 32'b00000000000000010011100010000000;
assign LUT_3[15589] = 32'b00000000000000011010001101011101;
assign LUT_3[15590] = 32'b00000000000000010101101001100100;
assign LUT_3[15591] = 32'b00000000000000011100010101000001;
assign LUT_3[15592] = 32'b00000000000000011011101101010000;
assign LUT_3[15593] = 32'b00000000000000100010011000101101;
assign LUT_3[15594] = 32'b00000000000000011101110100110100;
assign LUT_3[15595] = 32'b00000000000000100100100000010001;
assign LUT_3[15596] = 32'b00000000000000011000111011000110;
assign LUT_3[15597] = 32'b00000000000000011111100110100011;
assign LUT_3[15598] = 32'b00000000000000011011000010101010;
assign LUT_3[15599] = 32'b00000000000000100001101110000111;
assign LUT_3[15600] = 32'b00000000000000011001100111001101;
assign LUT_3[15601] = 32'b00000000000000100000010010101010;
assign LUT_3[15602] = 32'b00000000000000011011101110110001;
assign LUT_3[15603] = 32'b00000000000000100010011010001110;
assign LUT_3[15604] = 32'b00000000000000010110110101000011;
assign LUT_3[15605] = 32'b00000000000000011101100000100000;
assign LUT_3[15606] = 32'b00000000000000011000111100100111;
assign LUT_3[15607] = 32'b00000000000000011111101000000100;
assign LUT_3[15608] = 32'b00000000000000011111000000010011;
assign LUT_3[15609] = 32'b00000000000000100101101011110000;
assign LUT_3[15610] = 32'b00000000000000100001000111110111;
assign LUT_3[15611] = 32'b00000000000000100111110011010100;
assign LUT_3[15612] = 32'b00000000000000011100001110001001;
assign LUT_3[15613] = 32'b00000000000000100010111001100110;
assign LUT_3[15614] = 32'b00000000000000011110010101101101;
assign LUT_3[15615] = 32'b00000000000000100101000001001010;
assign LUT_3[15616] = 32'b00000000000000001111010001100010;
assign LUT_3[15617] = 32'b00000000000000010101111100111111;
assign LUT_3[15618] = 32'b00000000000000010001011001000110;
assign LUT_3[15619] = 32'b00000000000000011000000100100011;
assign LUT_3[15620] = 32'b00000000000000001100011111011000;
assign LUT_3[15621] = 32'b00000000000000010011001010110101;
assign LUT_3[15622] = 32'b00000000000000001110100110111100;
assign LUT_3[15623] = 32'b00000000000000010101010010011001;
assign LUT_3[15624] = 32'b00000000000000010100101010101000;
assign LUT_3[15625] = 32'b00000000000000011011010110000101;
assign LUT_3[15626] = 32'b00000000000000010110110010001100;
assign LUT_3[15627] = 32'b00000000000000011101011101101001;
assign LUT_3[15628] = 32'b00000000000000010001111000011110;
assign LUT_3[15629] = 32'b00000000000000011000100011111011;
assign LUT_3[15630] = 32'b00000000000000010100000000000010;
assign LUT_3[15631] = 32'b00000000000000011010101011011111;
assign LUT_3[15632] = 32'b00000000000000010010100100100101;
assign LUT_3[15633] = 32'b00000000000000011001010000000010;
assign LUT_3[15634] = 32'b00000000000000010100101100001001;
assign LUT_3[15635] = 32'b00000000000000011011010111100110;
assign LUT_3[15636] = 32'b00000000000000001111110010011011;
assign LUT_3[15637] = 32'b00000000000000010110011101111000;
assign LUT_3[15638] = 32'b00000000000000010001111001111111;
assign LUT_3[15639] = 32'b00000000000000011000100101011100;
assign LUT_3[15640] = 32'b00000000000000010111111101101011;
assign LUT_3[15641] = 32'b00000000000000011110101001001000;
assign LUT_3[15642] = 32'b00000000000000011010000101001111;
assign LUT_3[15643] = 32'b00000000000000100000110000101100;
assign LUT_3[15644] = 32'b00000000000000010101001011100001;
assign LUT_3[15645] = 32'b00000000000000011011110110111110;
assign LUT_3[15646] = 32'b00000000000000010111010011000101;
assign LUT_3[15647] = 32'b00000000000000011101111110100010;
assign LUT_3[15648] = 32'b00000000000000010000100000000010;
assign LUT_3[15649] = 32'b00000000000000010111001011011111;
assign LUT_3[15650] = 32'b00000000000000010010100111100110;
assign LUT_3[15651] = 32'b00000000000000011001010011000011;
assign LUT_3[15652] = 32'b00000000000000001101101101111000;
assign LUT_3[15653] = 32'b00000000000000010100011001010101;
assign LUT_3[15654] = 32'b00000000000000001111110101011100;
assign LUT_3[15655] = 32'b00000000000000010110100000111001;
assign LUT_3[15656] = 32'b00000000000000010101111001001000;
assign LUT_3[15657] = 32'b00000000000000011100100100100101;
assign LUT_3[15658] = 32'b00000000000000011000000000101100;
assign LUT_3[15659] = 32'b00000000000000011110101100001001;
assign LUT_3[15660] = 32'b00000000000000010011000110111110;
assign LUT_3[15661] = 32'b00000000000000011001110010011011;
assign LUT_3[15662] = 32'b00000000000000010101001110100010;
assign LUT_3[15663] = 32'b00000000000000011011111001111111;
assign LUT_3[15664] = 32'b00000000000000010011110011000101;
assign LUT_3[15665] = 32'b00000000000000011010011110100010;
assign LUT_3[15666] = 32'b00000000000000010101111010101001;
assign LUT_3[15667] = 32'b00000000000000011100100110000110;
assign LUT_3[15668] = 32'b00000000000000010001000000111011;
assign LUT_3[15669] = 32'b00000000000000010111101100011000;
assign LUT_3[15670] = 32'b00000000000000010011001000011111;
assign LUT_3[15671] = 32'b00000000000000011001110011111100;
assign LUT_3[15672] = 32'b00000000000000011001001100001011;
assign LUT_3[15673] = 32'b00000000000000011111110111101000;
assign LUT_3[15674] = 32'b00000000000000011011010011101111;
assign LUT_3[15675] = 32'b00000000000000100001111111001100;
assign LUT_3[15676] = 32'b00000000000000010110011010000001;
assign LUT_3[15677] = 32'b00000000000000011101000101011110;
assign LUT_3[15678] = 32'b00000000000000011000100001100101;
assign LUT_3[15679] = 32'b00000000000000011111001101000010;
assign LUT_3[15680] = 32'b00000000000000001111001010001101;
assign LUT_3[15681] = 32'b00000000000000010101110101101010;
assign LUT_3[15682] = 32'b00000000000000010001010001110001;
assign LUT_3[15683] = 32'b00000000000000010111111101001110;
assign LUT_3[15684] = 32'b00000000000000001100011000000011;
assign LUT_3[15685] = 32'b00000000000000010011000011100000;
assign LUT_3[15686] = 32'b00000000000000001110011111100111;
assign LUT_3[15687] = 32'b00000000000000010101001011000100;
assign LUT_3[15688] = 32'b00000000000000010100100011010011;
assign LUT_3[15689] = 32'b00000000000000011011001110110000;
assign LUT_3[15690] = 32'b00000000000000010110101010110111;
assign LUT_3[15691] = 32'b00000000000000011101010110010100;
assign LUT_3[15692] = 32'b00000000000000010001110001001001;
assign LUT_3[15693] = 32'b00000000000000011000011100100110;
assign LUT_3[15694] = 32'b00000000000000010011111000101101;
assign LUT_3[15695] = 32'b00000000000000011010100100001010;
assign LUT_3[15696] = 32'b00000000000000010010011101010000;
assign LUT_3[15697] = 32'b00000000000000011001001000101101;
assign LUT_3[15698] = 32'b00000000000000010100100100110100;
assign LUT_3[15699] = 32'b00000000000000011011010000010001;
assign LUT_3[15700] = 32'b00000000000000001111101011000110;
assign LUT_3[15701] = 32'b00000000000000010110010110100011;
assign LUT_3[15702] = 32'b00000000000000010001110010101010;
assign LUT_3[15703] = 32'b00000000000000011000011110000111;
assign LUT_3[15704] = 32'b00000000000000010111110110010110;
assign LUT_3[15705] = 32'b00000000000000011110100001110011;
assign LUT_3[15706] = 32'b00000000000000011001111101111010;
assign LUT_3[15707] = 32'b00000000000000100000101001010111;
assign LUT_3[15708] = 32'b00000000000000010101000100001100;
assign LUT_3[15709] = 32'b00000000000000011011101111101001;
assign LUT_3[15710] = 32'b00000000000000010111001011110000;
assign LUT_3[15711] = 32'b00000000000000011101110111001101;
assign LUT_3[15712] = 32'b00000000000000010000011000101101;
assign LUT_3[15713] = 32'b00000000000000010111000100001010;
assign LUT_3[15714] = 32'b00000000000000010010100000010001;
assign LUT_3[15715] = 32'b00000000000000011001001011101110;
assign LUT_3[15716] = 32'b00000000000000001101100110100011;
assign LUT_3[15717] = 32'b00000000000000010100010010000000;
assign LUT_3[15718] = 32'b00000000000000001111101110000111;
assign LUT_3[15719] = 32'b00000000000000010110011001100100;
assign LUT_3[15720] = 32'b00000000000000010101110001110011;
assign LUT_3[15721] = 32'b00000000000000011100011101010000;
assign LUT_3[15722] = 32'b00000000000000010111111001010111;
assign LUT_3[15723] = 32'b00000000000000011110100100110100;
assign LUT_3[15724] = 32'b00000000000000010010111111101001;
assign LUT_3[15725] = 32'b00000000000000011001101011000110;
assign LUT_3[15726] = 32'b00000000000000010101000111001101;
assign LUT_3[15727] = 32'b00000000000000011011110010101010;
assign LUT_3[15728] = 32'b00000000000000010011101011110000;
assign LUT_3[15729] = 32'b00000000000000011010010111001101;
assign LUT_3[15730] = 32'b00000000000000010101110011010100;
assign LUT_3[15731] = 32'b00000000000000011100011110110001;
assign LUT_3[15732] = 32'b00000000000000010000111001100110;
assign LUT_3[15733] = 32'b00000000000000010111100101000011;
assign LUT_3[15734] = 32'b00000000000000010011000001001010;
assign LUT_3[15735] = 32'b00000000000000011001101100100111;
assign LUT_3[15736] = 32'b00000000000000011001000100110110;
assign LUT_3[15737] = 32'b00000000000000011111110000010011;
assign LUT_3[15738] = 32'b00000000000000011011001100011010;
assign LUT_3[15739] = 32'b00000000000000100001110111110111;
assign LUT_3[15740] = 32'b00000000000000010110010010101100;
assign LUT_3[15741] = 32'b00000000000000011100111110001001;
assign LUT_3[15742] = 32'b00000000000000011000011010010000;
assign LUT_3[15743] = 32'b00000000000000011111000101101101;
assign LUT_3[15744] = 32'b00000000000000010001011100100000;
assign LUT_3[15745] = 32'b00000000000000011000000111111101;
assign LUT_3[15746] = 32'b00000000000000010011100100000100;
assign LUT_3[15747] = 32'b00000000000000011010001111100001;
assign LUT_3[15748] = 32'b00000000000000001110101010010110;
assign LUT_3[15749] = 32'b00000000000000010101010101110011;
assign LUT_3[15750] = 32'b00000000000000010000110001111010;
assign LUT_3[15751] = 32'b00000000000000010111011101010111;
assign LUT_3[15752] = 32'b00000000000000010110110101100110;
assign LUT_3[15753] = 32'b00000000000000011101100001000011;
assign LUT_3[15754] = 32'b00000000000000011000111101001010;
assign LUT_3[15755] = 32'b00000000000000011111101000100111;
assign LUT_3[15756] = 32'b00000000000000010100000011011100;
assign LUT_3[15757] = 32'b00000000000000011010101110111001;
assign LUT_3[15758] = 32'b00000000000000010110001011000000;
assign LUT_3[15759] = 32'b00000000000000011100110110011101;
assign LUT_3[15760] = 32'b00000000000000010100101111100011;
assign LUT_3[15761] = 32'b00000000000000011011011011000000;
assign LUT_3[15762] = 32'b00000000000000010110110111000111;
assign LUT_3[15763] = 32'b00000000000000011101100010100100;
assign LUT_3[15764] = 32'b00000000000000010001111101011001;
assign LUT_3[15765] = 32'b00000000000000011000101000110110;
assign LUT_3[15766] = 32'b00000000000000010100000100111101;
assign LUT_3[15767] = 32'b00000000000000011010110000011010;
assign LUT_3[15768] = 32'b00000000000000011010001000101001;
assign LUT_3[15769] = 32'b00000000000000100000110100000110;
assign LUT_3[15770] = 32'b00000000000000011100010000001101;
assign LUT_3[15771] = 32'b00000000000000100010111011101010;
assign LUT_3[15772] = 32'b00000000000000010111010110011111;
assign LUT_3[15773] = 32'b00000000000000011110000001111100;
assign LUT_3[15774] = 32'b00000000000000011001011110000011;
assign LUT_3[15775] = 32'b00000000000000100000001001100000;
assign LUT_3[15776] = 32'b00000000000000010010101011000000;
assign LUT_3[15777] = 32'b00000000000000011001010110011101;
assign LUT_3[15778] = 32'b00000000000000010100110010100100;
assign LUT_3[15779] = 32'b00000000000000011011011110000001;
assign LUT_3[15780] = 32'b00000000000000001111111000110110;
assign LUT_3[15781] = 32'b00000000000000010110100100010011;
assign LUT_3[15782] = 32'b00000000000000010010000000011010;
assign LUT_3[15783] = 32'b00000000000000011000101011110111;
assign LUT_3[15784] = 32'b00000000000000011000000100000110;
assign LUT_3[15785] = 32'b00000000000000011110101111100011;
assign LUT_3[15786] = 32'b00000000000000011010001011101010;
assign LUT_3[15787] = 32'b00000000000000100000110111000111;
assign LUT_3[15788] = 32'b00000000000000010101010001111100;
assign LUT_3[15789] = 32'b00000000000000011011111101011001;
assign LUT_3[15790] = 32'b00000000000000010111011001100000;
assign LUT_3[15791] = 32'b00000000000000011110000100111101;
assign LUT_3[15792] = 32'b00000000000000010101111110000011;
assign LUT_3[15793] = 32'b00000000000000011100101001100000;
assign LUT_3[15794] = 32'b00000000000000011000000101100111;
assign LUT_3[15795] = 32'b00000000000000011110110001000100;
assign LUT_3[15796] = 32'b00000000000000010011001011111001;
assign LUT_3[15797] = 32'b00000000000000011001110111010110;
assign LUT_3[15798] = 32'b00000000000000010101010011011101;
assign LUT_3[15799] = 32'b00000000000000011011111110111010;
assign LUT_3[15800] = 32'b00000000000000011011010111001001;
assign LUT_3[15801] = 32'b00000000000000100010000010100110;
assign LUT_3[15802] = 32'b00000000000000011101011110101101;
assign LUT_3[15803] = 32'b00000000000000100100001010001010;
assign LUT_3[15804] = 32'b00000000000000011000100100111111;
assign LUT_3[15805] = 32'b00000000000000011111010000011100;
assign LUT_3[15806] = 32'b00000000000000011010101100100011;
assign LUT_3[15807] = 32'b00000000000000100001011000000000;
assign LUT_3[15808] = 32'b00000000000000010001010101001011;
assign LUT_3[15809] = 32'b00000000000000011000000000101000;
assign LUT_3[15810] = 32'b00000000000000010011011100101111;
assign LUT_3[15811] = 32'b00000000000000011010001000001100;
assign LUT_3[15812] = 32'b00000000000000001110100011000001;
assign LUT_3[15813] = 32'b00000000000000010101001110011110;
assign LUT_3[15814] = 32'b00000000000000010000101010100101;
assign LUT_3[15815] = 32'b00000000000000010111010110000010;
assign LUT_3[15816] = 32'b00000000000000010110101110010001;
assign LUT_3[15817] = 32'b00000000000000011101011001101110;
assign LUT_3[15818] = 32'b00000000000000011000110101110101;
assign LUT_3[15819] = 32'b00000000000000011111100001010010;
assign LUT_3[15820] = 32'b00000000000000010011111100000111;
assign LUT_3[15821] = 32'b00000000000000011010100111100100;
assign LUT_3[15822] = 32'b00000000000000010110000011101011;
assign LUT_3[15823] = 32'b00000000000000011100101111001000;
assign LUT_3[15824] = 32'b00000000000000010100101000001110;
assign LUT_3[15825] = 32'b00000000000000011011010011101011;
assign LUT_3[15826] = 32'b00000000000000010110101111110010;
assign LUT_3[15827] = 32'b00000000000000011101011011001111;
assign LUT_3[15828] = 32'b00000000000000010001110110000100;
assign LUT_3[15829] = 32'b00000000000000011000100001100001;
assign LUT_3[15830] = 32'b00000000000000010011111101101000;
assign LUT_3[15831] = 32'b00000000000000011010101001000101;
assign LUT_3[15832] = 32'b00000000000000011010000001010100;
assign LUT_3[15833] = 32'b00000000000000100000101100110001;
assign LUT_3[15834] = 32'b00000000000000011100001000111000;
assign LUT_3[15835] = 32'b00000000000000100010110100010101;
assign LUT_3[15836] = 32'b00000000000000010111001111001010;
assign LUT_3[15837] = 32'b00000000000000011101111010100111;
assign LUT_3[15838] = 32'b00000000000000011001010110101110;
assign LUT_3[15839] = 32'b00000000000000100000000010001011;
assign LUT_3[15840] = 32'b00000000000000010010100011101011;
assign LUT_3[15841] = 32'b00000000000000011001001111001000;
assign LUT_3[15842] = 32'b00000000000000010100101011001111;
assign LUT_3[15843] = 32'b00000000000000011011010110101100;
assign LUT_3[15844] = 32'b00000000000000001111110001100001;
assign LUT_3[15845] = 32'b00000000000000010110011100111110;
assign LUT_3[15846] = 32'b00000000000000010001111001000101;
assign LUT_3[15847] = 32'b00000000000000011000100100100010;
assign LUT_3[15848] = 32'b00000000000000010111111100110001;
assign LUT_3[15849] = 32'b00000000000000011110101000001110;
assign LUT_3[15850] = 32'b00000000000000011010000100010101;
assign LUT_3[15851] = 32'b00000000000000100000101111110010;
assign LUT_3[15852] = 32'b00000000000000010101001010100111;
assign LUT_3[15853] = 32'b00000000000000011011110110000100;
assign LUT_3[15854] = 32'b00000000000000010111010010001011;
assign LUT_3[15855] = 32'b00000000000000011101111101101000;
assign LUT_3[15856] = 32'b00000000000000010101110110101110;
assign LUT_3[15857] = 32'b00000000000000011100100010001011;
assign LUT_3[15858] = 32'b00000000000000010111111110010010;
assign LUT_3[15859] = 32'b00000000000000011110101001101111;
assign LUT_3[15860] = 32'b00000000000000010011000100100100;
assign LUT_3[15861] = 32'b00000000000000011001110000000001;
assign LUT_3[15862] = 32'b00000000000000010101001100001000;
assign LUT_3[15863] = 32'b00000000000000011011110111100101;
assign LUT_3[15864] = 32'b00000000000000011011001111110100;
assign LUT_3[15865] = 32'b00000000000000100001111011010001;
assign LUT_3[15866] = 32'b00000000000000011101010111011000;
assign LUT_3[15867] = 32'b00000000000000100100000010110101;
assign LUT_3[15868] = 32'b00000000000000011000011101101010;
assign LUT_3[15869] = 32'b00000000000000011111001001000111;
assign LUT_3[15870] = 32'b00000000000000011010100101001110;
assign LUT_3[15871] = 32'b00000000000000100001010000101011;
assign LUT_3[15872] = 32'b00000000000000010110010111001101;
assign LUT_3[15873] = 32'b00000000000000011101000010101010;
assign LUT_3[15874] = 32'b00000000000000011000011110110001;
assign LUT_3[15875] = 32'b00000000000000011111001010001110;
assign LUT_3[15876] = 32'b00000000000000010011100101000011;
assign LUT_3[15877] = 32'b00000000000000011010010000100000;
assign LUT_3[15878] = 32'b00000000000000010101101100100111;
assign LUT_3[15879] = 32'b00000000000000011100011000000100;
assign LUT_3[15880] = 32'b00000000000000011011110000010011;
assign LUT_3[15881] = 32'b00000000000000100010011011110000;
assign LUT_3[15882] = 32'b00000000000000011101110111110111;
assign LUT_3[15883] = 32'b00000000000000100100100011010100;
assign LUT_3[15884] = 32'b00000000000000011000111110001001;
assign LUT_3[15885] = 32'b00000000000000011111101001100110;
assign LUT_3[15886] = 32'b00000000000000011011000101101101;
assign LUT_3[15887] = 32'b00000000000000100001110001001010;
assign LUT_3[15888] = 32'b00000000000000011001101010010000;
assign LUT_3[15889] = 32'b00000000000000100000010101101101;
assign LUT_3[15890] = 32'b00000000000000011011110001110100;
assign LUT_3[15891] = 32'b00000000000000100010011101010001;
assign LUT_3[15892] = 32'b00000000000000010110111000000110;
assign LUT_3[15893] = 32'b00000000000000011101100011100011;
assign LUT_3[15894] = 32'b00000000000000011000111111101010;
assign LUT_3[15895] = 32'b00000000000000011111101011000111;
assign LUT_3[15896] = 32'b00000000000000011111000011010110;
assign LUT_3[15897] = 32'b00000000000000100101101110110011;
assign LUT_3[15898] = 32'b00000000000000100001001010111010;
assign LUT_3[15899] = 32'b00000000000000100111110110010111;
assign LUT_3[15900] = 32'b00000000000000011100010001001100;
assign LUT_3[15901] = 32'b00000000000000100010111100101001;
assign LUT_3[15902] = 32'b00000000000000011110011000110000;
assign LUT_3[15903] = 32'b00000000000000100101000100001101;
assign LUT_3[15904] = 32'b00000000000000010111100101101101;
assign LUT_3[15905] = 32'b00000000000000011110010001001010;
assign LUT_3[15906] = 32'b00000000000000011001101101010001;
assign LUT_3[15907] = 32'b00000000000000100000011000101110;
assign LUT_3[15908] = 32'b00000000000000010100110011100011;
assign LUT_3[15909] = 32'b00000000000000011011011111000000;
assign LUT_3[15910] = 32'b00000000000000010110111011000111;
assign LUT_3[15911] = 32'b00000000000000011101100110100100;
assign LUT_3[15912] = 32'b00000000000000011100111110110011;
assign LUT_3[15913] = 32'b00000000000000100011101010010000;
assign LUT_3[15914] = 32'b00000000000000011111000110010111;
assign LUT_3[15915] = 32'b00000000000000100101110001110100;
assign LUT_3[15916] = 32'b00000000000000011010001100101001;
assign LUT_3[15917] = 32'b00000000000000100000111000000110;
assign LUT_3[15918] = 32'b00000000000000011100010100001101;
assign LUT_3[15919] = 32'b00000000000000100010111111101010;
assign LUT_3[15920] = 32'b00000000000000011010111000110000;
assign LUT_3[15921] = 32'b00000000000000100001100100001101;
assign LUT_3[15922] = 32'b00000000000000011101000000010100;
assign LUT_3[15923] = 32'b00000000000000100011101011110001;
assign LUT_3[15924] = 32'b00000000000000011000000110100110;
assign LUT_3[15925] = 32'b00000000000000011110110010000011;
assign LUT_3[15926] = 32'b00000000000000011010001110001010;
assign LUT_3[15927] = 32'b00000000000000100000111001100111;
assign LUT_3[15928] = 32'b00000000000000100000010001110110;
assign LUT_3[15929] = 32'b00000000000000100110111101010011;
assign LUT_3[15930] = 32'b00000000000000100010011001011010;
assign LUT_3[15931] = 32'b00000000000000101001000100110111;
assign LUT_3[15932] = 32'b00000000000000011101011111101100;
assign LUT_3[15933] = 32'b00000000000000100100001011001001;
assign LUT_3[15934] = 32'b00000000000000011111100111010000;
assign LUT_3[15935] = 32'b00000000000000100110010010101101;
assign LUT_3[15936] = 32'b00000000000000010110001111111000;
assign LUT_3[15937] = 32'b00000000000000011100111011010101;
assign LUT_3[15938] = 32'b00000000000000011000010111011100;
assign LUT_3[15939] = 32'b00000000000000011111000010111001;
assign LUT_3[15940] = 32'b00000000000000010011011101101110;
assign LUT_3[15941] = 32'b00000000000000011010001001001011;
assign LUT_3[15942] = 32'b00000000000000010101100101010010;
assign LUT_3[15943] = 32'b00000000000000011100010000101111;
assign LUT_3[15944] = 32'b00000000000000011011101000111110;
assign LUT_3[15945] = 32'b00000000000000100010010100011011;
assign LUT_3[15946] = 32'b00000000000000011101110000100010;
assign LUT_3[15947] = 32'b00000000000000100100011011111111;
assign LUT_3[15948] = 32'b00000000000000011000110110110100;
assign LUT_3[15949] = 32'b00000000000000011111100010010001;
assign LUT_3[15950] = 32'b00000000000000011010111110011000;
assign LUT_3[15951] = 32'b00000000000000100001101001110101;
assign LUT_3[15952] = 32'b00000000000000011001100010111011;
assign LUT_3[15953] = 32'b00000000000000100000001110011000;
assign LUT_3[15954] = 32'b00000000000000011011101010011111;
assign LUT_3[15955] = 32'b00000000000000100010010101111100;
assign LUT_3[15956] = 32'b00000000000000010110110000110001;
assign LUT_3[15957] = 32'b00000000000000011101011100001110;
assign LUT_3[15958] = 32'b00000000000000011000111000010101;
assign LUT_3[15959] = 32'b00000000000000011111100011110010;
assign LUT_3[15960] = 32'b00000000000000011110111100000001;
assign LUT_3[15961] = 32'b00000000000000100101100111011110;
assign LUT_3[15962] = 32'b00000000000000100001000011100101;
assign LUT_3[15963] = 32'b00000000000000100111101111000010;
assign LUT_3[15964] = 32'b00000000000000011100001001110111;
assign LUT_3[15965] = 32'b00000000000000100010110101010100;
assign LUT_3[15966] = 32'b00000000000000011110010001011011;
assign LUT_3[15967] = 32'b00000000000000100100111100111000;
assign LUT_3[15968] = 32'b00000000000000010111011110011000;
assign LUT_3[15969] = 32'b00000000000000011110001001110101;
assign LUT_3[15970] = 32'b00000000000000011001100101111100;
assign LUT_3[15971] = 32'b00000000000000100000010001011001;
assign LUT_3[15972] = 32'b00000000000000010100101100001110;
assign LUT_3[15973] = 32'b00000000000000011011010111101011;
assign LUT_3[15974] = 32'b00000000000000010110110011110010;
assign LUT_3[15975] = 32'b00000000000000011101011111001111;
assign LUT_3[15976] = 32'b00000000000000011100110111011110;
assign LUT_3[15977] = 32'b00000000000000100011100010111011;
assign LUT_3[15978] = 32'b00000000000000011110111111000010;
assign LUT_3[15979] = 32'b00000000000000100101101010011111;
assign LUT_3[15980] = 32'b00000000000000011010000101010100;
assign LUT_3[15981] = 32'b00000000000000100000110000110001;
assign LUT_3[15982] = 32'b00000000000000011100001100111000;
assign LUT_3[15983] = 32'b00000000000000100010111000010101;
assign LUT_3[15984] = 32'b00000000000000011010110001011011;
assign LUT_3[15985] = 32'b00000000000000100001011100111000;
assign LUT_3[15986] = 32'b00000000000000011100111000111111;
assign LUT_3[15987] = 32'b00000000000000100011100100011100;
assign LUT_3[15988] = 32'b00000000000000010111111111010001;
assign LUT_3[15989] = 32'b00000000000000011110101010101110;
assign LUT_3[15990] = 32'b00000000000000011010000110110101;
assign LUT_3[15991] = 32'b00000000000000100000110010010010;
assign LUT_3[15992] = 32'b00000000000000100000001010100001;
assign LUT_3[15993] = 32'b00000000000000100110110101111110;
assign LUT_3[15994] = 32'b00000000000000100010010010000101;
assign LUT_3[15995] = 32'b00000000000000101000111101100010;
assign LUT_3[15996] = 32'b00000000000000011101011000010111;
assign LUT_3[15997] = 32'b00000000000000100100000011110100;
assign LUT_3[15998] = 32'b00000000000000011111011111111011;
assign LUT_3[15999] = 32'b00000000000000100110001011011000;
assign LUT_3[16000] = 32'b00000000000000011000100010001011;
assign LUT_3[16001] = 32'b00000000000000011111001101101000;
assign LUT_3[16002] = 32'b00000000000000011010101001101111;
assign LUT_3[16003] = 32'b00000000000000100001010101001100;
assign LUT_3[16004] = 32'b00000000000000010101110000000001;
assign LUT_3[16005] = 32'b00000000000000011100011011011110;
assign LUT_3[16006] = 32'b00000000000000010111110111100101;
assign LUT_3[16007] = 32'b00000000000000011110100011000010;
assign LUT_3[16008] = 32'b00000000000000011101111011010001;
assign LUT_3[16009] = 32'b00000000000000100100100110101110;
assign LUT_3[16010] = 32'b00000000000000100000000010110101;
assign LUT_3[16011] = 32'b00000000000000100110101110010010;
assign LUT_3[16012] = 32'b00000000000000011011001001000111;
assign LUT_3[16013] = 32'b00000000000000100001110100100100;
assign LUT_3[16014] = 32'b00000000000000011101010000101011;
assign LUT_3[16015] = 32'b00000000000000100011111100001000;
assign LUT_3[16016] = 32'b00000000000000011011110101001110;
assign LUT_3[16017] = 32'b00000000000000100010100000101011;
assign LUT_3[16018] = 32'b00000000000000011101111100110010;
assign LUT_3[16019] = 32'b00000000000000100100101000001111;
assign LUT_3[16020] = 32'b00000000000000011001000011000100;
assign LUT_3[16021] = 32'b00000000000000011111101110100001;
assign LUT_3[16022] = 32'b00000000000000011011001010101000;
assign LUT_3[16023] = 32'b00000000000000100001110110000101;
assign LUT_3[16024] = 32'b00000000000000100001001110010100;
assign LUT_3[16025] = 32'b00000000000000100111111001110001;
assign LUT_3[16026] = 32'b00000000000000100011010101111000;
assign LUT_3[16027] = 32'b00000000000000101010000001010101;
assign LUT_3[16028] = 32'b00000000000000011110011100001010;
assign LUT_3[16029] = 32'b00000000000000100101000111100111;
assign LUT_3[16030] = 32'b00000000000000100000100011101110;
assign LUT_3[16031] = 32'b00000000000000100111001111001011;
assign LUT_3[16032] = 32'b00000000000000011001110000101011;
assign LUT_3[16033] = 32'b00000000000000100000011100001000;
assign LUT_3[16034] = 32'b00000000000000011011111000001111;
assign LUT_3[16035] = 32'b00000000000000100010100011101100;
assign LUT_3[16036] = 32'b00000000000000010110111110100001;
assign LUT_3[16037] = 32'b00000000000000011101101001111110;
assign LUT_3[16038] = 32'b00000000000000011001000110000101;
assign LUT_3[16039] = 32'b00000000000000011111110001100010;
assign LUT_3[16040] = 32'b00000000000000011111001001110001;
assign LUT_3[16041] = 32'b00000000000000100101110101001110;
assign LUT_3[16042] = 32'b00000000000000100001010001010101;
assign LUT_3[16043] = 32'b00000000000000100111111100110010;
assign LUT_3[16044] = 32'b00000000000000011100010111100111;
assign LUT_3[16045] = 32'b00000000000000100011000011000100;
assign LUT_3[16046] = 32'b00000000000000011110011111001011;
assign LUT_3[16047] = 32'b00000000000000100101001010101000;
assign LUT_3[16048] = 32'b00000000000000011101000011101110;
assign LUT_3[16049] = 32'b00000000000000100011101111001011;
assign LUT_3[16050] = 32'b00000000000000011111001011010010;
assign LUT_3[16051] = 32'b00000000000000100101110110101111;
assign LUT_3[16052] = 32'b00000000000000011010010001100100;
assign LUT_3[16053] = 32'b00000000000000100000111101000001;
assign LUT_3[16054] = 32'b00000000000000011100011001001000;
assign LUT_3[16055] = 32'b00000000000000100011000100100101;
assign LUT_3[16056] = 32'b00000000000000100010011100110100;
assign LUT_3[16057] = 32'b00000000000000101001001000010001;
assign LUT_3[16058] = 32'b00000000000000100100100100011000;
assign LUT_3[16059] = 32'b00000000000000101011001111110101;
assign LUT_3[16060] = 32'b00000000000000011111101010101010;
assign LUT_3[16061] = 32'b00000000000000100110010110000111;
assign LUT_3[16062] = 32'b00000000000000100001110010001110;
assign LUT_3[16063] = 32'b00000000000000101000011101101011;
assign LUT_3[16064] = 32'b00000000000000011000011010110110;
assign LUT_3[16065] = 32'b00000000000000011111000110010011;
assign LUT_3[16066] = 32'b00000000000000011010100010011010;
assign LUT_3[16067] = 32'b00000000000000100001001101110111;
assign LUT_3[16068] = 32'b00000000000000010101101000101100;
assign LUT_3[16069] = 32'b00000000000000011100010100001001;
assign LUT_3[16070] = 32'b00000000000000010111110000010000;
assign LUT_3[16071] = 32'b00000000000000011110011011101101;
assign LUT_3[16072] = 32'b00000000000000011101110011111100;
assign LUT_3[16073] = 32'b00000000000000100100011111011001;
assign LUT_3[16074] = 32'b00000000000000011111111011100000;
assign LUT_3[16075] = 32'b00000000000000100110100110111101;
assign LUT_3[16076] = 32'b00000000000000011011000001110010;
assign LUT_3[16077] = 32'b00000000000000100001101101001111;
assign LUT_3[16078] = 32'b00000000000000011101001001010110;
assign LUT_3[16079] = 32'b00000000000000100011110100110011;
assign LUT_3[16080] = 32'b00000000000000011011101101111001;
assign LUT_3[16081] = 32'b00000000000000100010011001010110;
assign LUT_3[16082] = 32'b00000000000000011101110101011101;
assign LUT_3[16083] = 32'b00000000000000100100100000111010;
assign LUT_3[16084] = 32'b00000000000000011000111011101111;
assign LUT_3[16085] = 32'b00000000000000011111100111001100;
assign LUT_3[16086] = 32'b00000000000000011011000011010011;
assign LUT_3[16087] = 32'b00000000000000100001101110110000;
assign LUT_3[16088] = 32'b00000000000000100001000110111111;
assign LUT_3[16089] = 32'b00000000000000100111110010011100;
assign LUT_3[16090] = 32'b00000000000000100011001110100011;
assign LUT_3[16091] = 32'b00000000000000101001111010000000;
assign LUT_3[16092] = 32'b00000000000000011110010100110101;
assign LUT_3[16093] = 32'b00000000000000100101000000010010;
assign LUT_3[16094] = 32'b00000000000000100000011100011001;
assign LUT_3[16095] = 32'b00000000000000100111000111110110;
assign LUT_3[16096] = 32'b00000000000000011001101001010110;
assign LUT_3[16097] = 32'b00000000000000100000010100110011;
assign LUT_3[16098] = 32'b00000000000000011011110000111010;
assign LUT_3[16099] = 32'b00000000000000100010011100010111;
assign LUT_3[16100] = 32'b00000000000000010110110111001100;
assign LUT_3[16101] = 32'b00000000000000011101100010101001;
assign LUT_3[16102] = 32'b00000000000000011000111110110000;
assign LUT_3[16103] = 32'b00000000000000011111101010001101;
assign LUT_3[16104] = 32'b00000000000000011111000010011100;
assign LUT_3[16105] = 32'b00000000000000100101101101111001;
assign LUT_3[16106] = 32'b00000000000000100001001010000000;
assign LUT_3[16107] = 32'b00000000000000100111110101011101;
assign LUT_3[16108] = 32'b00000000000000011100010000010010;
assign LUT_3[16109] = 32'b00000000000000100010111011101111;
assign LUT_3[16110] = 32'b00000000000000011110010111110110;
assign LUT_3[16111] = 32'b00000000000000100101000011010011;
assign LUT_3[16112] = 32'b00000000000000011100111100011001;
assign LUT_3[16113] = 32'b00000000000000100011100111110110;
assign LUT_3[16114] = 32'b00000000000000011111000011111101;
assign LUT_3[16115] = 32'b00000000000000100101101111011010;
assign LUT_3[16116] = 32'b00000000000000011010001010001111;
assign LUT_3[16117] = 32'b00000000000000100000110101101100;
assign LUT_3[16118] = 32'b00000000000000011100010001110011;
assign LUT_3[16119] = 32'b00000000000000100010111101010000;
assign LUT_3[16120] = 32'b00000000000000100010010101011111;
assign LUT_3[16121] = 32'b00000000000000101001000000111100;
assign LUT_3[16122] = 32'b00000000000000100100011101000011;
assign LUT_3[16123] = 32'b00000000000000101011001000100000;
assign LUT_3[16124] = 32'b00000000000000011111100011010101;
assign LUT_3[16125] = 32'b00000000000000100110001110110010;
assign LUT_3[16126] = 32'b00000000000000100001101010111001;
assign LUT_3[16127] = 32'b00000000000000101000010110010110;
assign LUT_3[16128] = 32'b00000000000000010010100110101110;
assign LUT_3[16129] = 32'b00000000000000011001010010001011;
assign LUT_3[16130] = 32'b00000000000000010100101110010010;
assign LUT_3[16131] = 32'b00000000000000011011011001101111;
assign LUT_3[16132] = 32'b00000000000000001111110100100100;
assign LUT_3[16133] = 32'b00000000000000010110100000000001;
assign LUT_3[16134] = 32'b00000000000000010001111100001000;
assign LUT_3[16135] = 32'b00000000000000011000100111100101;
assign LUT_3[16136] = 32'b00000000000000010111111111110100;
assign LUT_3[16137] = 32'b00000000000000011110101011010001;
assign LUT_3[16138] = 32'b00000000000000011010000111011000;
assign LUT_3[16139] = 32'b00000000000000100000110010110101;
assign LUT_3[16140] = 32'b00000000000000010101001101101010;
assign LUT_3[16141] = 32'b00000000000000011011111001000111;
assign LUT_3[16142] = 32'b00000000000000010111010101001110;
assign LUT_3[16143] = 32'b00000000000000011110000000101011;
assign LUT_3[16144] = 32'b00000000000000010101111001110001;
assign LUT_3[16145] = 32'b00000000000000011100100101001110;
assign LUT_3[16146] = 32'b00000000000000011000000001010101;
assign LUT_3[16147] = 32'b00000000000000011110101100110010;
assign LUT_3[16148] = 32'b00000000000000010011000111100111;
assign LUT_3[16149] = 32'b00000000000000011001110011000100;
assign LUT_3[16150] = 32'b00000000000000010101001111001011;
assign LUT_3[16151] = 32'b00000000000000011011111010101000;
assign LUT_3[16152] = 32'b00000000000000011011010010110111;
assign LUT_3[16153] = 32'b00000000000000100001111110010100;
assign LUT_3[16154] = 32'b00000000000000011101011010011011;
assign LUT_3[16155] = 32'b00000000000000100100000101111000;
assign LUT_3[16156] = 32'b00000000000000011000100000101101;
assign LUT_3[16157] = 32'b00000000000000011111001100001010;
assign LUT_3[16158] = 32'b00000000000000011010101000010001;
assign LUT_3[16159] = 32'b00000000000000100001010011101110;
assign LUT_3[16160] = 32'b00000000000000010011110101001110;
assign LUT_3[16161] = 32'b00000000000000011010100000101011;
assign LUT_3[16162] = 32'b00000000000000010101111100110010;
assign LUT_3[16163] = 32'b00000000000000011100101000001111;
assign LUT_3[16164] = 32'b00000000000000010001000011000100;
assign LUT_3[16165] = 32'b00000000000000010111101110100001;
assign LUT_3[16166] = 32'b00000000000000010011001010101000;
assign LUT_3[16167] = 32'b00000000000000011001110110000101;
assign LUT_3[16168] = 32'b00000000000000011001001110010100;
assign LUT_3[16169] = 32'b00000000000000011111111001110001;
assign LUT_3[16170] = 32'b00000000000000011011010101111000;
assign LUT_3[16171] = 32'b00000000000000100010000001010101;
assign LUT_3[16172] = 32'b00000000000000010110011100001010;
assign LUT_3[16173] = 32'b00000000000000011101000111100111;
assign LUT_3[16174] = 32'b00000000000000011000100011101110;
assign LUT_3[16175] = 32'b00000000000000011111001111001011;
assign LUT_3[16176] = 32'b00000000000000010111001000010001;
assign LUT_3[16177] = 32'b00000000000000011101110011101110;
assign LUT_3[16178] = 32'b00000000000000011001001111110101;
assign LUT_3[16179] = 32'b00000000000000011111111011010010;
assign LUT_3[16180] = 32'b00000000000000010100010110000111;
assign LUT_3[16181] = 32'b00000000000000011011000001100100;
assign LUT_3[16182] = 32'b00000000000000010110011101101011;
assign LUT_3[16183] = 32'b00000000000000011101001001001000;
assign LUT_3[16184] = 32'b00000000000000011100100001010111;
assign LUT_3[16185] = 32'b00000000000000100011001100110100;
assign LUT_3[16186] = 32'b00000000000000011110101000111011;
assign LUT_3[16187] = 32'b00000000000000100101010100011000;
assign LUT_3[16188] = 32'b00000000000000011001101111001101;
assign LUT_3[16189] = 32'b00000000000000100000011010101010;
assign LUT_3[16190] = 32'b00000000000000011011110110110001;
assign LUT_3[16191] = 32'b00000000000000100010100010001110;
assign LUT_3[16192] = 32'b00000000000000010010011111011001;
assign LUT_3[16193] = 32'b00000000000000011001001010110110;
assign LUT_3[16194] = 32'b00000000000000010100100110111101;
assign LUT_3[16195] = 32'b00000000000000011011010010011010;
assign LUT_3[16196] = 32'b00000000000000001111101101001111;
assign LUT_3[16197] = 32'b00000000000000010110011000101100;
assign LUT_3[16198] = 32'b00000000000000010001110100110011;
assign LUT_3[16199] = 32'b00000000000000011000100000010000;
assign LUT_3[16200] = 32'b00000000000000010111111000011111;
assign LUT_3[16201] = 32'b00000000000000011110100011111100;
assign LUT_3[16202] = 32'b00000000000000011010000000000011;
assign LUT_3[16203] = 32'b00000000000000100000101011100000;
assign LUT_3[16204] = 32'b00000000000000010101000110010101;
assign LUT_3[16205] = 32'b00000000000000011011110001110010;
assign LUT_3[16206] = 32'b00000000000000010111001101111001;
assign LUT_3[16207] = 32'b00000000000000011101111001010110;
assign LUT_3[16208] = 32'b00000000000000010101110010011100;
assign LUT_3[16209] = 32'b00000000000000011100011101111001;
assign LUT_3[16210] = 32'b00000000000000010111111010000000;
assign LUT_3[16211] = 32'b00000000000000011110100101011101;
assign LUT_3[16212] = 32'b00000000000000010011000000010010;
assign LUT_3[16213] = 32'b00000000000000011001101011101111;
assign LUT_3[16214] = 32'b00000000000000010101000111110110;
assign LUT_3[16215] = 32'b00000000000000011011110011010011;
assign LUT_3[16216] = 32'b00000000000000011011001011100010;
assign LUT_3[16217] = 32'b00000000000000100001110110111111;
assign LUT_3[16218] = 32'b00000000000000011101010011000110;
assign LUT_3[16219] = 32'b00000000000000100011111110100011;
assign LUT_3[16220] = 32'b00000000000000011000011001011000;
assign LUT_3[16221] = 32'b00000000000000011111000100110101;
assign LUT_3[16222] = 32'b00000000000000011010100000111100;
assign LUT_3[16223] = 32'b00000000000000100001001100011001;
assign LUT_3[16224] = 32'b00000000000000010011101101111001;
assign LUT_3[16225] = 32'b00000000000000011010011001010110;
assign LUT_3[16226] = 32'b00000000000000010101110101011101;
assign LUT_3[16227] = 32'b00000000000000011100100000111010;
assign LUT_3[16228] = 32'b00000000000000010000111011101111;
assign LUT_3[16229] = 32'b00000000000000010111100111001100;
assign LUT_3[16230] = 32'b00000000000000010011000011010011;
assign LUT_3[16231] = 32'b00000000000000011001101110110000;
assign LUT_3[16232] = 32'b00000000000000011001000110111111;
assign LUT_3[16233] = 32'b00000000000000011111110010011100;
assign LUT_3[16234] = 32'b00000000000000011011001110100011;
assign LUT_3[16235] = 32'b00000000000000100001111010000000;
assign LUT_3[16236] = 32'b00000000000000010110010100110101;
assign LUT_3[16237] = 32'b00000000000000011101000000010010;
assign LUT_3[16238] = 32'b00000000000000011000011100011001;
assign LUT_3[16239] = 32'b00000000000000011111000111110110;
assign LUT_3[16240] = 32'b00000000000000010111000000111100;
assign LUT_3[16241] = 32'b00000000000000011101101100011001;
assign LUT_3[16242] = 32'b00000000000000011001001000100000;
assign LUT_3[16243] = 32'b00000000000000011111110011111101;
assign LUT_3[16244] = 32'b00000000000000010100001110110010;
assign LUT_3[16245] = 32'b00000000000000011010111010001111;
assign LUT_3[16246] = 32'b00000000000000010110010110010110;
assign LUT_3[16247] = 32'b00000000000000011101000001110011;
assign LUT_3[16248] = 32'b00000000000000011100011010000010;
assign LUT_3[16249] = 32'b00000000000000100011000101011111;
assign LUT_3[16250] = 32'b00000000000000011110100001100110;
assign LUT_3[16251] = 32'b00000000000000100101001101000011;
assign LUT_3[16252] = 32'b00000000000000011001100111111000;
assign LUT_3[16253] = 32'b00000000000000100000010011010101;
assign LUT_3[16254] = 32'b00000000000000011011101111011100;
assign LUT_3[16255] = 32'b00000000000000100010011010111001;
assign LUT_3[16256] = 32'b00000000000000010100110001101100;
assign LUT_3[16257] = 32'b00000000000000011011011101001001;
assign LUT_3[16258] = 32'b00000000000000010110111001010000;
assign LUT_3[16259] = 32'b00000000000000011101100100101101;
assign LUT_3[16260] = 32'b00000000000000010001111111100010;
assign LUT_3[16261] = 32'b00000000000000011000101010111111;
assign LUT_3[16262] = 32'b00000000000000010100000111000110;
assign LUT_3[16263] = 32'b00000000000000011010110010100011;
assign LUT_3[16264] = 32'b00000000000000011010001010110010;
assign LUT_3[16265] = 32'b00000000000000100000110110001111;
assign LUT_3[16266] = 32'b00000000000000011100010010010110;
assign LUT_3[16267] = 32'b00000000000000100010111101110011;
assign LUT_3[16268] = 32'b00000000000000010111011000101000;
assign LUT_3[16269] = 32'b00000000000000011110000100000101;
assign LUT_3[16270] = 32'b00000000000000011001100000001100;
assign LUT_3[16271] = 32'b00000000000000100000001011101001;
assign LUT_3[16272] = 32'b00000000000000011000000100101111;
assign LUT_3[16273] = 32'b00000000000000011110110000001100;
assign LUT_3[16274] = 32'b00000000000000011010001100010011;
assign LUT_3[16275] = 32'b00000000000000100000110111110000;
assign LUT_3[16276] = 32'b00000000000000010101010010100101;
assign LUT_3[16277] = 32'b00000000000000011011111110000010;
assign LUT_3[16278] = 32'b00000000000000010111011010001001;
assign LUT_3[16279] = 32'b00000000000000011110000101100110;
assign LUT_3[16280] = 32'b00000000000000011101011101110101;
assign LUT_3[16281] = 32'b00000000000000100100001001010010;
assign LUT_3[16282] = 32'b00000000000000011111100101011001;
assign LUT_3[16283] = 32'b00000000000000100110010000110110;
assign LUT_3[16284] = 32'b00000000000000011010101011101011;
assign LUT_3[16285] = 32'b00000000000000100001010111001000;
assign LUT_3[16286] = 32'b00000000000000011100110011001111;
assign LUT_3[16287] = 32'b00000000000000100011011110101100;
assign LUT_3[16288] = 32'b00000000000000010110000000001100;
assign LUT_3[16289] = 32'b00000000000000011100101011101001;
assign LUT_3[16290] = 32'b00000000000000011000000111110000;
assign LUT_3[16291] = 32'b00000000000000011110110011001101;
assign LUT_3[16292] = 32'b00000000000000010011001110000010;
assign LUT_3[16293] = 32'b00000000000000011001111001011111;
assign LUT_3[16294] = 32'b00000000000000010101010101100110;
assign LUT_3[16295] = 32'b00000000000000011100000001000011;
assign LUT_3[16296] = 32'b00000000000000011011011001010010;
assign LUT_3[16297] = 32'b00000000000000100010000100101111;
assign LUT_3[16298] = 32'b00000000000000011101100000110110;
assign LUT_3[16299] = 32'b00000000000000100100001100010011;
assign LUT_3[16300] = 32'b00000000000000011000100111001000;
assign LUT_3[16301] = 32'b00000000000000011111010010100101;
assign LUT_3[16302] = 32'b00000000000000011010101110101100;
assign LUT_3[16303] = 32'b00000000000000100001011010001001;
assign LUT_3[16304] = 32'b00000000000000011001010011001111;
assign LUT_3[16305] = 32'b00000000000000011111111110101100;
assign LUT_3[16306] = 32'b00000000000000011011011010110011;
assign LUT_3[16307] = 32'b00000000000000100010000110010000;
assign LUT_3[16308] = 32'b00000000000000010110100001000101;
assign LUT_3[16309] = 32'b00000000000000011101001100100010;
assign LUT_3[16310] = 32'b00000000000000011000101000101001;
assign LUT_3[16311] = 32'b00000000000000011111010100000110;
assign LUT_3[16312] = 32'b00000000000000011110101100010101;
assign LUT_3[16313] = 32'b00000000000000100101010111110010;
assign LUT_3[16314] = 32'b00000000000000100000110011111001;
assign LUT_3[16315] = 32'b00000000000000100111011111010110;
assign LUT_3[16316] = 32'b00000000000000011011111010001011;
assign LUT_3[16317] = 32'b00000000000000100010100101101000;
assign LUT_3[16318] = 32'b00000000000000011110000001101111;
assign LUT_3[16319] = 32'b00000000000000100100101101001100;
assign LUT_3[16320] = 32'b00000000000000010100101010010111;
assign LUT_3[16321] = 32'b00000000000000011011010101110100;
assign LUT_3[16322] = 32'b00000000000000010110110001111011;
assign LUT_3[16323] = 32'b00000000000000011101011101011000;
assign LUT_3[16324] = 32'b00000000000000010001111000001101;
assign LUT_3[16325] = 32'b00000000000000011000100011101010;
assign LUT_3[16326] = 32'b00000000000000010011111111110001;
assign LUT_3[16327] = 32'b00000000000000011010101011001110;
assign LUT_3[16328] = 32'b00000000000000011010000011011101;
assign LUT_3[16329] = 32'b00000000000000100000101110111010;
assign LUT_3[16330] = 32'b00000000000000011100001011000001;
assign LUT_3[16331] = 32'b00000000000000100010110110011110;
assign LUT_3[16332] = 32'b00000000000000010111010001010011;
assign LUT_3[16333] = 32'b00000000000000011101111100110000;
assign LUT_3[16334] = 32'b00000000000000011001011000110111;
assign LUT_3[16335] = 32'b00000000000000100000000100010100;
assign LUT_3[16336] = 32'b00000000000000010111111101011010;
assign LUT_3[16337] = 32'b00000000000000011110101000110111;
assign LUT_3[16338] = 32'b00000000000000011010000100111110;
assign LUT_3[16339] = 32'b00000000000000100000110000011011;
assign LUT_3[16340] = 32'b00000000000000010101001011010000;
assign LUT_3[16341] = 32'b00000000000000011011110110101101;
assign LUT_3[16342] = 32'b00000000000000010111010010110100;
assign LUT_3[16343] = 32'b00000000000000011101111110010001;
assign LUT_3[16344] = 32'b00000000000000011101010110100000;
assign LUT_3[16345] = 32'b00000000000000100100000001111101;
assign LUT_3[16346] = 32'b00000000000000011111011110000100;
assign LUT_3[16347] = 32'b00000000000000100110001001100001;
assign LUT_3[16348] = 32'b00000000000000011010100100010110;
assign LUT_3[16349] = 32'b00000000000000100001001111110011;
assign LUT_3[16350] = 32'b00000000000000011100101011111010;
assign LUT_3[16351] = 32'b00000000000000100011010111010111;
assign LUT_3[16352] = 32'b00000000000000010101111000110111;
assign LUT_3[16353] = 32'b00000000000000011100100100010100;
assign LUT_3[16354] = 32'b00000000000000011000000000011011;
assign LUT_3[16355] = 32'b00000000000000011110101011111000;
assign LUT_3[16356] = 32'b00000000000000010011000110101101;
assign LUT_3[16357] = 32'b00000000000000011001110010001010;
assign LUT_3[16358] = 32'b00000000000000010101001110010001;
assign LUT_3[16359] = 32'b00000000000000011011111001101110;
assign LUT_3[16360] = 32'b00000000000000011011010001111101;
assign LUT_3[16361] = 32'b00000000000000100001111101011010;
assign LUT_3[16362] = 32'b00000000000000011101011001100001;
assign LUT_3[16363] = 32'b00000000000000100100000100111110;
assign LUT_3[16364] = 32'b00000000000000011000011111110011;
assign LUT_3[16365] = 32'b00000000000000011111001011010000;
assign LUT_3[16366] = 32'b00000000000000011010100111010111;
assign LUT_3[16367] = 32'b00000000000000100001010010110100;
assign LUT_3[16368] = 32'b00000000000000011001001011111010;
assign LUT_3[16369] = 32'b00000000000000011111110111010111;
assign LUT_3[16370] = 32'b00000000000000011011010011011110;
assign LUT_3[16371] = 32'b00000000000000100001111110111011;
assign LUT_3[16372] = 32'b00000000000000010110011001110000;
assign LUT_3[16373] = 32'b00000000000000011101000101001101;
assign LUT_3[16374] = 32'b00000000000000011000100001010100;
assign LUT_3[16375] = 32'b00000000000000011111001100110001;
assign LUT_3[16376] = 32'b00000000000000011110100101000000;
assign LUT_3[16377] = 32'b00000000000000100101010000011101;
assign LUT_3[16378] = 32'b00000000000000100000101100100100;
assign LUT_3[16379] = 32'b00000000000000100111011000000001;
assign LUT_3[16380] = 32'b00000000000000011011110010110110;
assign LUT_3[16381] = 32'b00000000000000100010011110010011;
assign LUT_3[16382] = 32'b00000000000000011101111010011010;
assign LUT_3[16383] = 32'b00000000000000100100100101110111;
assign LUT_3[16384] = 32'b00000000000000000100101110100111;
assign LUT_3[16385] = 32'b00000000000000001011011010000100;
assign LUT_3[16386] = 32'b00000000000000000110110110001011;
assign LUT_3[16387] = 32'b00000000000000001101100001101000;
assign LUT_3[16388] = 32'b00000000000000000001111100011101;
assign LUT_3[16389] = 32'b00000000000000001000100111111010;
assign LUT_3[16390] = 32'b00000000000000000100000100000001;
assign LUT_3[16391] = 32'b00000000000000001010101111011110;
assign LUT_3[16392] = 32'b00000000000000001010000111101101;
assign LUT_3[16393] = 32'b00000000000000010000110011001010;
assign LUT_3[16394] = 32'b00000000000000001100001111010001;
assign LUT_3[16395] = 32'b00000000000000010010111010101110;
assign LUT_3[16396] = 32'b00000000000000000111010101100011;
assign LUT_3[16397] = 32'b00000000000000001110000001000000;
assign LUT_3[16398] = 32'b00000000000000001001011101000111;
assign LUT_3[16399] = 32'b00000000000000010000001000100100;
assign LUT_3[16400] = 32'b00000000000000001000000001101010;
assign LUT_3[16401] = 32'b00000000000000001110101101000111;
assign LUT_3[16402] = 32'b00000000000000001010001001001110;
assign LUT_3[16403] = 32'b00000000000000010000110100101011;
assign LUT_3[16404] = 32'b00000000000000000101001111100000;
assign LUT_3[16405] = 32'b00000000000000001011111010111101;
assign LUT_3[16406] = 32'b00000000000000000111010111000100;
assign LUT_3[16407] = 32'b00000000000000001110000010100001;
assign LUT_3[16408] = 32'b00000000000000001101011010110000;
assign LUT_3[16409] = 32'b00000000000000010100000110001101;
assign LUT_3[16410] = 32'b00000000000000001111100010010100;
assign LUT_3[16411] = 32'b00000000000000010110001101110001;
assign LUT_3[16412] = 32'b00000000000000001010101000100110;
assign LUT_3[16413] = 32'b00000000000000010001010100000011;
assign LUT_3[16414] = 32'b00000000000000001100110000001010;
assign LUT_3[16415] = 32'b00000000000000010011011011100111;
assign LUT_3[16416] = 32'b00000000000000000101111101000111;
assign LUT_3[16417] = 32'b00000000000000001100101000100100;
assign LUT_3[16418] = 32'b00000000000000001000000100101011;
assign LUT_3[16419] = 32'b00000000000000001110110000001000;
assign LUT_3[16420] = 32'b00000000000000000011001010111101;
assign LUT_3[16421] = 32'b00000000000000001001110110011010;
assign LUT_3[16422] = 32'b00000000000000000101010010100001;
assign LUT_3[16423] = 32'b00000000000000001011111101111110;
assign LUT_3[16424] = 32'b00000000000000001011010110001101;
assign LUT_3[16425] = 32'b00000000000000010010000001101010;
assign LUT_3[16426] = 32'b00000000000000001101011101110001;
assign LUT_3[16427] = 32'b00000000000000010100001001001110;
assign LUT_3[16428] = 32'b00000000000000001000100100000011;
assign LUT_3[16429] = 32'b00000000000000001111001111100000;
assign LUT_3[16430] = 32'b00000000000000001010101011100111;
assign LUT_3[16431] = 32'b00000000000000010001010111000100;
assign LUT_3[16432] = 32'b00000000000000001001010000001010;
assign LUT_3[16433] = 32'b00000000000000001111111011100111;
assign LUT_3[16434] = 32'b00000000000000001011010111101110;
assign LUT_3[16435] = 32'b00000000000000010010000011001011;
assign LUT_3[16436] = 32'b00000000000000000110011110000000;
assign LUT_3[16437] = 32'b00000000000000001101001001011101;
assign LUT_3[16438] = 32'b00000000000000001000100101100100;
assign LUT_3[16439] = 32'b00000000000000001111010001000001;
assign LUT_3[16440] = 32'b00000000000000001110101001010000;
assign LUT_3[16441] = 32'b00000000000000010101010100101101;
assign LUT_3[16442] = 32'b00000000000000010000110000110100;
assign LUT_3[16443] = 32'b00000000000000010111011100010001;
assign LUT_3[16444] = 32'b00000000000000001011110111000110;
assign LUT_3[16445] = 32'b00000000000000010010100010100011;
assign LUT_3[16446] = 32'b00000000000000001101111110101010;
assign LUT_3[16447] = 32'b00000000000000010100101010000111;
assign LUT_3[16448] = 32'b00000000000000000100100111010010;
assign LUT_3[16449] = 32'b00000000000000001011010010101111;
assign LUT_3[16450] = 32'b00000000000000000110101110110110;
assign LUT_3[16451] = 32'b00000000000000001101011010010011;
assign LUT_3[16452] = 32'b00000000000000000001110101001000;
assign LUT_3[16453] = 32'b00000000000000001000100000100101;
assign LUT_3[16454] = 32'b00000000000000000011111100101100;
assign LUT_3[16455] = 32'b00000000000000001010101000001001;
assign LUT_3[16456] = 32'b00000000000000001010000000011000;
assign LUT_3[16457] = 32'b00000000000000010000101011110101;
assign LUT_3[16458] = 32'b00000000000000001100000111111100;
assign LUT_3[16459] = 32'b00000000000000010010110011011001;
assign LUT_3[16460] = 32'b00000000000000000111001110001110;
assign LUT_3[16461] = 32'b00000000000000001101111001101011;
assign LUT_3[16462] = 32'b00000000000000001001010101110010;
assign LUT_3[16463] = 32'b00000000000000010000000001001111;
assign LUT_3[16464] = 32'b00000000000000000111111010010101;
assign LUT_3[16465] = 32'b00000000000000001110100101110010;
assign LUT_3[16466] = 32'b00000000000000001010000001111001;
assign LUT_3[16467] = 32'b00000000000000010000101101010110;
assign LUT_3[16468] = 32'b00000000000000000101001000001011;
assign LUT_3[16469] = 32'b00000000000000001011110011101000;
assign LUT_3[16470] = 32'b00000000000000000111001111101111;
assign LUT_3[16471] = 32'b00000000000000001101111011001100;
assign LUT_3[16472] = 32'b00000000000000001101010011011011;
assign LUT_3[16473] = 32'b00000000000000010011111110111000;
assign LUT_3[16474] = 32'b00000000000000001111011010111111;
assign LUT_3[16475] = 32'b00000000000000010110000110011100;
assign LUT_3[16476] = 32'b00000000000000001010100001010001;
assign LUT_3[16477] = 32'b00000000000000010001001100101110;
assign LUT_3[16478] = 32'b00000000000000001100101000110101;
assign LUT_3[16479] = 32'b00000000000000010011010100010010;
assign LUT_3[16480] = 32'b00000000000000000101110101110010;
assign LUT_3[16481] = 32'b00000000000000001100100001001111;
assign LUT_3[16482] = 32'b00000000000000000111111101010110;
assign LUT_3[16483] = 32'b00000000000000001110101000110011;
assign LUT_3[16484] = 32'b00000000000000000011000011101000;
assign LUT_3[16485] = 32'b00000000000000001001101111000101;
assign LUT_3[16486] = 32'b00000000000000000101001011001100;
assign LUT_3[16487] = 32'b00000000000000001011110110101001;
assign LUT_3[16488] = 32'b00000000000000001011001110111000;
assign LUT_3[16489] = 32'b00000000000000010001111010010101;
assign LUT_3[16490] = 32'b00000000000000001101010110011100;
assign LUT_3[16491] = 32'b00000000000000010100000001111001;
assign LUT_3[16492] = 32'b00000000000000001000011100101110;
assign LUT_3[16493] = 32'b00000000000000001111001000001011;
assign LUT_3[16494] = 32'b00000000000000001010100100010010;
assign LUT_3[16495] = 32'b00000000000000010001001111101111;
assign LUT_3[16496] = 32'b00000000000000001001001000110101;
assign LUT_3[16497] = 32'b00000000000000001111110100010010;
assign LUT_3[16498] = 32'b00000000000000001011010000011001;
assign LUT_3[16499] = 32'b00000000000000010001111011110110;
assign LUT_3[16500] = 32'b00000000000000000110010110101011;
assign LUT_3[16501] = 32'b00000000000000001101000010001000;
assign LUT_3[16502] = 32'b00000000000000001000011110001111;
assign LUT_3[16503] = 32'b00000000000000001111001001101100;
assign LUT_3[16504] = 32'b00000000000000001110100001111011;
assign LUT_3[16505] = 32'b00000000000000010101001101011000;
assign LUT_3[16506] = 32'b00000000000000010000101001011111;
assign LUT_3[16507] = 32'b00000000000000010111010100111100;
assign LUT_3[16508] = 32'b00000000000000001011101111110001;
assign LUT_3[16509] = 32'b00000000000000010010011011001110;
assign LUT_3[16510] = 32'b00000000000000001101110111010101;
assign LUT_3[16511] = 32'b00000000000000010100100010110010;
assign LUT_3[16512] = 32'b00000000000000000110111001100101;
assign LUT_3[16513] = 32'b00000000000000001101100101000010;
assign LUT_3[16514] = 32'b00000000000000001001000001001001;
assign LUT_3[16515] = 32'b00000000000000001111101100100110;
assign LUT_3[16516] = 32'b00000000000000000100000111011011;
assign LUT_3[16517] = 32'b00000000000000001010110010111000;
assign LUT_3[16518] = 32'b00000000000000000110001110111111;
assign LUT_3[16519] = 32'b00000000000000001100111010011100;
assign LUT_3[16520] = 32'b00000000000000001100010010101011;
assign LUT_3[16521] = 32'b00000000000000010010111110001000;
assign LUT_3[16522] = 32'b00000000000000001110011010001111;
assign LUT_3[16523] = 32'b00000000000000010101000101101100;
assign LUT_3[16524] = 32'b00000000000000001001100000100001;
assign LUT_3[16525] = 32'b00000000000000010000001011111110;
assign LUT_3[16526] = 32'b00000000000000001011101000000101;
assign LUT_3[16527] = 32'b00000000000000010010010011100010;
assign LUT_3[16528] = 32'b00000000000000001010001100101000;
assign LUT_3[16529] = 32'b00000000000000010000111000000101;
assign LUT_3[16530] = 32'b00000000000000001100010100001100;
assign LUT_3[16531] = 32'b00000000000000010010111111101001;
assign LUT_3[16532] = 32'b00000000000000000111011010011110;
assign LUT_3[16533] = 32'b00000000000000001110000101111011;
assign LUT_3[16534] = 32'b00000000000000001001100010000010;
assign LUT_3[16535] = 32'b00000000000000010000001101011111;
assign LUT_3[16536] = 32'b00000000000000001111100101101110;
assign LUT_3[16537] = 32'b00000000000000010110010001001011;
assign LUT_3[16538] = 32'b00000000000000010001101101010010;
assign LUT_3[16539] = 32'b00000000000000011000011000101111;
assign LUT_3[16540] = 32'b00000000000000001100110011100100;
assign LUT_3[16541] = 32'b00000000000000010011011111000001;
assign LUT_3[16542] = 32'b00000000000000001110111011001000;
assign LUT_3[16543] = 32'b00000000000000010101100110100101;
assign LUT_3[16544] = 32'b00000000000000001000001000000101;
assign LUT_3[16545] = 32'b00000000000000001110110011100010;
assign LUT_3[16546] = 32'b00000000000000001010001111101001;
assign LUT_3[16547] = 32'b00000000000000010000111011000110;
assign LUT_3[16548] = 32'b00000000000000000101010101111011;
assign LUT_3[16549] = 32'b00000000000000001100000001011000;
assign LUT_3[16550] = 32'b00000000000000000111011101011111;
assign LUT_3[16551] = 32'b00000000000000001110001000111100;
assign LUT_3[16552] = 32'b00000000000000001101100001001011;
assign LUT_3[16553] = 32'b00000000000000010100001100101000;
assign LUT_3[16554] = 32'b00000000000000001111101000101111;
assign LUT_3[16555] = 32'b00000000000000010110010100001100;
assign LUT_3[16556] = 32'b00000000000000001010101111000001;
assign LUT_3[16557] = 32'b00000000000000010001011010011110;
assign LUT_3[16558] = 32'b00000000000000001100110110100101;
assign LUT_3[16559] = 32'b00000000000000010011100010000010;
assign LUT_3[16560] = 32'b00000000000000001011011011001000;
assign LUT_3[16561] = 32'b00000000000000010010000110100101;
assign LUT_3[16562] = 32'b00000000000000001101100010101100;
assign LUT_3[16563] = 32'b00000000000000010100001110001001;
assign LUT_3[16564] = 32'b00000000000000001000101000111110;
assign LUT_3[16565] = 32'b00000000000000001111010100011011;
assign LUT_3[16566] = 32'b00000000000000001010110000100010;
assign LUT_3[16567] = 32'b00000000000000010001011011111111;
assign LUT_3[16568] = 32'b00000000000000010000110100001110;
assign LUT_3[16569] = 32'b00000000000000010111011111101011;
assign LUT_3[16570] = 32'b00000000000000010010111011110010;
assign LUT_3[16571] = 32'b00000000000000011001100111001111;
assign LUT_3[16572] = 32'b00000000000000001110000010000100;
assign LUT_3[16573] = 32'b00000000000000010100101101100001;
assign LUT_3[16574] = 32'b00000000000000010000001001101000;
assign LUT_3[16575] = 32'b00000000000000010110110101000101;
assign LUT_3[16576] = 32'b00000000000000000110110010010000;
assign LUT_3[16577] = 32'b00000000000000001101011101101101;
assign LUT_3[16578] = 32'b00000000000000001000111001110100;
assign LUT_3[16579] = 32'b00000000000000001111100101010001;
assign LUT_3[16580] = 32'b00000000000000000100000000000110;
assign LUT_3[16581] = 32'b00000000000000001010101011100011;
assign LUT_3[16582] = 32'b00000000000000000110000111101010;
assign LUT_3[16583] = 32'b00000000000000001100110011000111;
assign LUT_3[16584] = 32'b00000000000000001100001011010110;
assign LUT_3[16585] = 32'b00000000000000010010110110110011;
assign LUT_3[16586] = 32'b00000000000000001110010010111010;
assign LUT_3[16587] = 32'b00000000000000010100111110010111;
assign LUT_3[16588] = 32'b00000000000000001001011001001100;
assign LUT_3[16589] = 32'b00000000000000010000000100101001;
assign LUT_3[16590] = 32'b00000000000000001011100000110000;
assign LUT_3[16591] = 32'b00000000000000010010001100001101;
assign LUT_3[16592] = 32'b00000000000000001010000101010011;
assign LUT_3[16593] = 32'b00000000000000010000110000110000;
assign LUT_3[16594] = 32'b00000000000000001100001100110111;
assign LUT_3[16595] = 32'b00000000000000010010111000010100;
assign LUT_3[16596] = 32'b00000000000000000111010011001001;
assign LUT_3[16597] = 32'b00000000000000001101111110100110;
assign LUT_3[16598] = 32'b00000000000000001001011010101101;
assign LUT_3[16599] = 32'b00000000000000010000000110001010;
assign LUT_3[16600] = 32'b00000000000000001111011110011001;
assign LUT_3[16601] = 32'b00000000000000010110001001110110;
assign LUT_3[16602] = 32'b00000000000000010001100101111101;
assign LUT_3[16603] = 32'b00000000000000011000010001011010;
assign LUT_3[16604] = 32'b00000000000000001100101100001111;
assign LUT_3[16605] = 32'b00000000000000010011010111101100;
assign LUT_3[16606] = 32'b00000000000000001110110011110011;
assign LUT_3[16607] = 32'b00000000000000010101011111010000;
assign LUT_3[16608] = 32'b00000000000000001000000000110000;
assign LUT_3[16609] = 32'b00000000000000001110101100001101;
assign LUT_3[16610] = 32'b00000000000000001010001000010100;
assign LUT_3[16611] = 32'b00000000000000010000110011110001;
assign LUT_3[16612] = 32'b00000000000000000101001110100110;
assign LUT_3[16613] = 32'b00000000000000001011111010000011;
assign LUT_3[16614] = 32'b00000000000000000111010110001010;
assign LUT_3[16615] = 32'b00000000000000001110000001100111;
assign LUT_3[16616] = 32'b00000000000000001101011001110110;
assign LUT_3[16617] = 32'b00000000000000010100000101010011;
assign LUT_3[16618] = 32'b00000000000000001111100001011010;
assign LUT_3[16619] = 32'b00000000000000010110001100110111;
assign LUT_3[16620] = 32'b00000000000000001010100111101100;
assign LUT_3[16621] = 32'b00000000000000010001010011001001;
assign LUT_3[16622] = 32'b00000000000000001100101111010000;
assign LUT_3[16623] = 32'b00000000000000010011011010101101;
assign LUT_3[16624] = 32'b00000000000000001011010011110011;
assign LUT_3[16625] = 32'b00000000000000010001111111010000;
assign LUT_3[16626] = 32'b00000000000000001101011011010111;
assign LUT_3[16627] = 32'b00000000000000010100000110110100;
assign LUT_3[16628] = 32'b00000000000000001000100001101001;
assign LUT_3[16629] = 32'b00000000000000001111001101000110;
assign LUT_3[16630] = 32'b00000000000000001010101001001101;
assign LUT_3[16631] = 32'b00000000000000010001010100101010;
assign LUT_3[16632] = 32'b00000000000000010000101100111001;
assign LUT_3[16633] = 32'b00000000000000010111011000010110;
assign LUT_3[16634] = 32'b00000000000000010010110100011101;
assign LUT_3[16635] = 32'b00000000000000011001011111111010;
assign LUT_3[16636] = 32'b00000000000000001101111010101111;
assign LUT_3[16637] = 32'b00000000000000010100100110001100;
assign LUT_3[16638] = 32'b00000000000000010000000010010011;
assign LUT_3[16639] = 32'b00000000000000010110101101110000;
assign LUT_3[16640] = 32'b00000000000000000000111110001000;
assign LUT_3[16641] = 32'b00000000000000000111101001100101;
assign LUT_3[16642] = 32'b00000000000000000011000101101100;
assign LUT_3[16643] = 32'b00000000000000001001110001001001;
assign LUT_3[16644] = 32'b11111111111111111110001011111110;
assign LUT_3[16645] = 32'b00000000000000000100110111011011;
assign LUT_3[16646] = 32'b00000000000000000000010011100010;
assign LUT_3[16647] = 32'b00000000000000000110111110111111;
assign LUT_3[16648] = 32'b00000000000000000110010111001110;
assign LUT_3[16649] = 32'b00000000000000001101000010101011;
assign LUT_3[16650] = 32'b00000000000000001000011110110010;
assign LUT_3[16651] = 32'b00000000000000001111001010001111;
assign LUT_3[16652] = 32'b00000000000000000011100101000100;
assign LUT_3[16653] = 32'b00000000000000001010010000100001;
assign LUT_3[16654] = 32'b00000000000000000101101100101000;
assign LUT_3[16655] = 32'b00000000000000001100011000000101;
assign LUT_3[16656] = 32'b00000000000000000100010001001011;
assign LUT_3[16657] = 32'b00000000000000001010111100101000;
assign LUT_3[16658] = 32'b00000000000000000110011000101111;
assign LUT_3[16659] = 32'b00000000000000001101000100001100;
assign LUT_3[16660] = 32'b00000000000000000001011111000001;
assign LUT_3[16661] = 32'b00000000000000001000001010011110;
assign LUT_3[16662] = 32'b00000000000000000011100110100101;
assign LUT_3[16663] = 32'b00000000000000001010010010000010;
assign LUT_3[16664] = 32'b00000000000000001001101010010001;
assign LUT_3[16665] = 32'b00000000000000010000010101101110;
assign LUT_3[16666] = 32'b00000000000000001011110001110101;
assign LUT_3[16667] = 32'b00000000000000010010011101010010;
assign LUT_3[16668] = 32'b00000000000000000110111000000111;
assign LUT_3[16669] = 32'b00000000000000001101100011100100;
assign LUT_3[16670] = 32'b00000000000000001000111111101011;
assign LUT_3[16671] = 32'b00000000000000001111101011001000;
assign LUT_3[16672] = 32'b00000000000000000010001100101000;
assign LUT_3[16673] = 32'b00000000000000001000111000000101;
assign LUT_3[16674] = 32'b00000000000000000100010100001100;
assign LUT_3[16675] = 32'b00000000000000001010111111101001;
assign LUT_3[16676] = 32'b11111111111111111111011010011110;
assign LUT_3[16677] = 32'b00000000000000000110000101111011;
assign LUT_3[16678] = 32'b00000000000000000001100010000010;
assign LUT_3[16679] = 32'b00000000000000001000001101011111;
assign LUT_3[16680] = 32'b00000000000000000111100101101110;
assign LUT_3[16681] = 32'b00000000000000001110010001001011;
assign LUT_3[16682] = 32'b00000000000000001001101101010010;
assign LUT_3[16683] = 32'b00000000000000010000011000101111;
assign LUT_3[16684] = 32'b00000000000000000100110011100100;
assign LUT_3[16685] = 32'b00000000000000001011011111000001;
assign LUT_3[16686] = 32'b00000000000000000110111011001000;
assign LUT_3[16687] = 32'b00000000000000001101100110100101;
assign LUT_3[16688] = 32'b00000000000000000101011111101011;
assign LUT_3[16689] = 32'b00000000000000001100001011001000;
assign LUT_3[16690] = 32'b00000000000000000111100111001111;
assign LUT_3[16691] = 32'b00000000000000001110010010101100;
assign LUT_3[16692] = 32'b00000000000000000010101101100001;
assign LUT_3[16693] = 32'b00000000000000001001011000111110;
assign LUT_3[16694] = 32'b00000000000000000100110101000101;
assign LUT_3[16695] = 32'b00000000000000001011100000100010;
assign LUT_3[16696] = 32'b00000000000000001010111000110001;
assign LUT_3[16697] = 32'b00000000000000010001100100001110;
assign LUT_3[16698] = 32'b00000000000000001101000000010101;
assign LUT_3[16699] = 32'b00000000000000010011101011110010;
assign LUT_3[16700] = 32'b00000000000000001000000110100111;
assign LUT_3[16701] = 32'b00000000000000001110110010000100;
assign LUT_3[16702] = 32'b00000000000000001010001110001011;
assign LUT_3[16703] = 32'b00000000000000010000111001101000;
assign LUT_3[16704] = 32'b00000000000000000000110110110011;
assign LUT_3[16705] = 32'b00000000000000000111100010010000;
assign LUT_3[16706] = 32'b00000000000000000010111110010111;
assign LUT_3[16707] = 32'b00000000000000001001101001110100;
assign LUT_3[16708] = 32'b11111111111111111110000100101001;
assign LUT_3[16709] = 32'b00000000000000000100110000000110;
assign LUT_3[16710] = 32'b00000000000000000000001100001101;
assign LUT_3[16711] = 32'b00000000000000000110110111101010;
assign LUT_3[16712] = 32'b00000000000000000110001111111001;
assign LUT_3[16713] = 32'b00000000000000001100111011010110;
assign LUT_3[16714] = 32'b00000000000000001000010111011101;
assign LUT_3[16715] = 32'b00000000000000001111000010111010;
assign LUT_3[16716] = 32'b00000000000000000011011101101111;
assign LUT_3[16717] = 32'b00000000000000001010001001001100;
assign LUT_3[16718] = 32'b00000000000000000101100101010011;
assign LUT_3[16719] = 32'b00000000000000001100010000110000;
assign LUT_3[16720] = 32'b00000000000000000100001001110110;
assign LUT_3[16721] = 32'b00000000000000001010110101010011;
assign LUT_3[16722] = 32'b00000000000000000110010001011010;
assign LUT_3[16723] = 32'b00000000000000001100111100110111;
assign LUT_3[16724] = 32'b00000000000000000001010111101100;
assign LUT_3[16725] = 32'b00000000000000001000000011001001;
assign LUT_3[16726] = 32'b00000000000000000011011111010000;
assign LUT_3[16727] = 32'b00000000000000001010001010101101;
assign LUT_3[16728] = 32'b00000000000000001001100010111100;
assign LUT_3[16729] = 32'b00000000000000010000001110011001;
assign LUT_3[16730] = 32'b00000000000000001011101010100000;
assign LUT_3[16731] = 32'b00000000000000010010010101111101;
assign LUT_3[16732] = 32'b00000000000000000110110000110010;
assign LUT_3[16733] = 32'b00000000000000001101011100001111;
assign LUT_3[16734] = 32'b00000000000000001000111000010110;
assign LUT_3[16735] = 32'b00000000000000001111100011110011;
assign LUT_3[16736] = 32'b00000000000000000010000101010011;
assign LUT_3[16737] = 32'b00000000000000001000110000110000;
assign LUT_3[16738] = 32'b00000000000000000100001100110111;
assign LUT_3[16739] = 32'b00000000000000001010111000010100;
assign LUT_3[16740] = 32'b11111111111111111111010011001001;
assign LUT_3[16741] = 32'b00000000000000000101111110100110;
assign LUT_3[16742] = 32'b00000000000000000001011010101101;
assign LUT_3[16743] = 32'b00000000000000001000000110001010;
assign LUT_3[16744] = 32'b00000000000000000111011110011001;
assign LUT_3[16745] = 32'b00000000000000001110001001110110;
assign LUT_3[16746] = 32'b00000000000000001001100101111101;
assign LUT_3[16747] = 32'b00000000000000010000010001011010;
assign LUT_3[16748] = 32'b00000000000000000100101100001111;
assign LUT_3[16749] = 32'b00000000000000001011010111101100;
assign LUT_3[16750] = 32'b00000000000000000110110011110011;
assign LUT_3[16751] = 32'b00000000000000001101011111010000;
assign LUT_3[16752] = 32'b00000000000000000101011000010110;
assign LUT_3[16753] = 32'b00000000000000001100000011110011;
assign LUT_3[16754] = 32'b00000000000000000111011111111010;
assign LUT_3[16755] = 32'b00000000000000001110001011010111;
assign LUT_3[16756] = 32'b00000000000000000010100110001100;
assign LUT_3[16757] = 32'b00000000000000001001010001101001;
assign LUT_3[16758] = 32'b00000000000000000100101101110000;
assign LUT_3[16759] = 32'b00000000000000001011011001001101;
assign LUT_3[16760] = 32'b00000000000000001010110001011100;
assign LUT_3[16761] = 32'b00000000000000010001011100111001;
assign LUT_3[16762] = 32'b00000000000000001100111001000000;
assign LUT_3[16763] = 32'b00000000000000010011100100011101;
assign LUT_3[16764] = 32'b00000000000000000111111111010010;
assign LUT_3[16765] = 32'b00000000000000001110101010101111;
assign LUT_3[16766] = 32'b00000000000000001010000110110110;
assign LUT_3[16767] = 32'b00000000000000010000110010010011;
assign LUT_3[16768] = 32'b00000000000000000011001001000110;
assign LUT_3[16769] = 32'b00000000000000001001110100100011;
assign LUT_3[16770] = 32'b00000000000000000101010000101010;
assign LUT_3[16771] = 32'b00000000000000001011111100000111;
assign LUT_3[16772] = 32'b00000000000000000000010110111100;
assign LUT_3[16773] = 32'b00000000000000000111000010011001;
assign LUT_3[16774] = 32'b00000000000000000010011110100000;
assign LUT_3[16775] = 32'b00000000000000001001001001111101;
assign LUT_3[16776] = 32'b00000000000000001000100010001100;
assign LUT_3[16777] = 32'b00000000000000001111001101101001;
assign LUT_3[16778] = 32'b00000000000000001010101001110000;
assign LUT_3[16779] = 32'b00000000000000010001010101001101;
assign LUT_3[16780] = 32'b00000000000000000101110000000010;
assign LUT_3[16781] = 32'b00000000000000001100011011011111;
assign LUT_3[16782] = 32'b00000000000000000111110111100110;
assign LUT_3[16783] = 32'b00000000000000001110100011000011;
assign LUT_3[16784] = 32'b00000000000000000110011100001001;
assign LUT_3[16785] = 32'b00000000000000001101000111100110;
assign LUT_3[16786] = 32'b00000000000000001000100011101101;
assign LUT_3[16787] = 32'b00000000000000001111001111001010;
assign LUT_3[16788] = 32'b00000000000000000011101001111111;
assign LUT_3[16789] = 32'b00000000000000001010010101011100;
assign LUT_3[16790] = 32'b00000000000000000101110001100011;
assign LUT_3[16791] = 32'b00000000000000001100011101000000;
assign LUT_3[16792] = 32'b00000000000000001011110101001111;
assign LUT_3[16793] = 32'b00000000000000010010100000101100;
assign LUT_3[16794] = 32'b00000000000000001101111100110011;
assign LUT_3[16795] = 32'b00000000000000010100101000010000;
assign LUT_3[16796] = 32'b00000000000000001001000011000101;
assign LUT_3[16797] = 32'b00000000000000001111101110100010;
assign LUT_3[16798] = 32'b00000000000000001011001010101001;
assign LUT_3[16799] = 32'b00000000000000010001110110000110;
assign LUT_3[16800] = 32'b00000000000000000100010111100110;
assign LUT_3[16801] = 32'b00000000000000001011000011000011;
assign LUT_3[16802] = 32'b00000000000000000110011111001010;
assign LUT_3[16803] = 32'b00000000000000001101001010100111;
assign LUT_3[16804] = 32'b00000000000000000001100101011100;
assign LUT_3[16805] = 32'b00000000000000001000010000111001;
assign LUT_3[16806] = 32'b00000000000000000011101101000000;
assign LUT_3[16807] = 32'b00000000000000001010011000011101;
assign LUT_3[16808] = 32'b00000000000000001001110000101100;
assign LUT_3[16809] = 32'b00000000000000010000011100001001;
assign LUT_3[16810] = 32'b00000000000000001011111000010000;
assign LUT_3[16811] = 32'b00000000000000010010100011101101;
assign LUT_3[16812] = 32'b00000000000000000110111110100010;
assign LUT_3[16813] = 32'b00000000000000001101101001111111;
assign LUT_3[16814] = 32'b00000000000000001001000110000110;
assign LUT_3[16815] = 32'b00000000000000001111110001100011;
assign LUT_3[16816] = 32'b00000000000000000111101010101001;
assign LUT_3[16817] = 32'b00000000000000001110010110000110;
assign LUT_3[16818] = 32'b00000000000000001001110010001101;
assign LUT_3[16819] = 32'b00000000000000010000011101101010;
assign LUT_3[16820] = 32'b00000000000000000100111000011111;
assign LUT_3[16821] = 32'b00000000000000001011100011111100;
assign LUT_3[16822] = 32'b00000000000000000111000000000011;
assign LUT_3[16823] = 32'b00000000000000001101101011100000;
assign LUT_3[16824] = 32'b00000000000000001101000011101111;
assign LUT_3[16825] = 32'b00000000000000010011101111001100;
assign LUT_3[16826] = 32'b00000000000000001111001011010011;
assign LUT_3[16827] = 32'b00000000000000010101110110110000;
assign LUT_3[16828] = 32'b00000000000000001010010001100101;
assign LUT_3[16829] = 32'b00000000000000010000111101000010;
assign LUT_3[16830] = 32'b00000000000000001100011001001001;
assign LUT_3[16831] = 32'b00000000000000010011000100100110;
assign LUT_3[16832] = 32'b00000000000000000011000001110001;
assign LUT_3[16833] = 32'b00000000000000001001101101001110;
assign LUT_3[16834] = 32'b00000000000000000101001001010101;
assign LUT_3[16835] = 32'b00000000000000001011110100110010;
assign LUT_3[16836] = 32'b00000000000000000000001111100111;
assign LUT_3[16837] = 32'b00000000000000000110111011000100;
assign LUT_3[16838] = 32'b00000000000000000010010111001011;
assign LUT_3[16839] = 32'b00000000000000001001000010101000;
assign LUT_3[16840] = 32'b00000000000000001000011010110111;
assign LUT_3[16841] = 32'b00000000000000001111000110010100;
assign LUT_3[16842] = 32'b00000000000000001010100010011011;
assign LUT_3[16843] = 32'b00000000000000010001001101111000;
assign LUT_3[16844] = 32'b00000000000000000101101000101101;
assign LUT_3[16845] = 32'b00000000000000001100010100001010;
assign LUT_3[16846] = 32'b00000000000000000111110000010001;
assign LUT_3[16847] = 32'b00000000000000001110011011101110;
assign LUT_3[16848] = 32'b00000000000000000110010100110100;
assign LUT_3[16849] = 32'b00000000000000001101000000010001;
assign LUT_3[16850] = 32'b00000000000000001000011100011000;
assign LUT_3[16851] = 32'b00000000000000001111000111110101;
assign LUT_3[16852] = 32'b00000000000000000011100010101010;
assign LUT_3[16853] = 32'b00000000000000001010001110000111;
assign LUT_3[16854] = 32'b00000000000000000101101010001110;
assign LUT_3[16855] = 32'b00000000000000001100010101101011;
assign LUT_3[16856] = 32'b00000000000000001011101101111010;
assign LUT_3[16857] = 32'b00000000000000010010011001010111;
assign LUT_3[16858] = 32'b00000000000000001101110101011110;
assign LUT_3[16859] = 32'b00000000000000010100100000111011;
assign LUT_3[16860] = 32'b00000000000000001000111011110000;
assign LUT_3[16861] = 32'b00000000000000001111100111001101;
assign LUT_3[16862] = 32'b00000000000000001011000011010100;
assign LUT_3[16863] = 32'b00000000000000010001101110110001;
assign LUT_3[16864] = 32'b00000000000000000100010000010001;
assign LUT_3[16865] = 32'b00000000000000001010111011101110;
assign LUT_3[16866] = 32'b00000000000000000110010111110101;
assign LUT_3[16867] = 32'b00000000000000001101000011010010;
assign LUT_3[16868] = 32'b00000000000000000001011110000111;
assign LUT_3[16869] = 32'b00000000000000001000001001100100;
assign LUT_3[16870] = 32'b00000000000000000011100101101011;
assign LUT_3[16871] = 32'b00000000000000001010010001001000;
assign LUT_3[16872] = 32'b00000000000000001001101001010111;
assign LUT_3[16873] = 32'b00000000000000010000010100110100;
assign LUT_3[16874] = 32'b00000000000000001011110000111011;
assign LUT_3[16875] = 32'b00000000000000010010011100011000;
assign LUT_3[16876] = 32'b00000000000000000110110111001101;
assign LUT_3[16877] = 32'b00000000000000001101100010101010;
assign LUT_3[16878] = 32'b00000000000000001000111110110001;
assign LUT_3[16879] = 32'b00000000000000001111101010001110;
assign LUT_3[16880] = 32'b00000000000000000111100011010100;
assign LUT_3[16881] = 32'b00000000000000001110001110110001;
assign LUT_3[16882] = 32'b00000000000000001001101010111000;
assign LUT_3[16883] = 32'b00000000000000010000010110010101;
assign LUT_3[16884] = 32'b00000000000000000100110001001010;
assign LUT_3[16885] = 32'b00000000000000001011011100100111;
assign LUT_3[16886] = 32'b00000000000000000110111000101110;
assign LUT_3[16887] = 32'b00000000000000001101100100001011;
assign LUT_3[16888] = 32'b00000000000000001100111100011010;
assign LUT_3[16889] = 32'b00000000000000010011100111110111;
assign LUT_3[16890] = 32'b00000000000000001111000011111110;
assign LUT_3[16891] = 32'b00000000000000010101101111011011;
assign LUT_3[16892] = 32'b00000000000000001010001010010000;
assign LUT_3[16893] = 32'b00000000000000010000110101101101;
assign LUT_3[16894] = 32'b00000000000000001100010001110100;
assign LUT_3[16895] = 32'b00000000000000010010111101010001;
assign LUT_3[16896] = 32'b00000000000000001000000011110011;
assign LUT_3[16897] = 32'b00000000000000001110101111010000;
assign LUT_3[16898] = 32'b00000000000000001010001011010111;
assign LUT_3[16899] = 32'b00000000000000010000110110110100;
assign LUT_3[16900] = 32'b00000000000000000101010001101001;
assign LUT_3[16901] = 32'b00000000000000001011111101000110;
assign LUT_3[16902] = 32'b00000000000000000111011001001101;
assign LUT_3[16903] = 32'b00000000000000001110000100101010;
assign LUT_3[16904] = 32'b00000000000000001101011100111001;
assign LUT_3[16905] = 32'b00000000000000010100001000010110;
assign LUT_3[16906] = 32'b00000000000000001111100100011101;
assign LUT_3[16907] = 32'b00000000000000010110001111111010;
assign LUT_3[16908] = 32'b00000000000000001010101010101111;
assign LUT_3[16909] = 32'b00000000000000010001010110001100;
assign LUT_3[16910] = 32'b00000000000000001100110010010011;
assign LUT_3[16911] = 32'b00000000000000010011011101110000;
assign LUT_3[16912] = 32'b00000000000000001011010110110110;
assign LUT_3[16913] = 32'b00000000000000010010000010010011;
assign LUT_3[16914] = 32'b00000000000000001101011110011010;
assign LUT_3[16915] = 32'b00000000000000010100001001110111;
assign LUT_3[16916] = 32'b00000000000000001000100100101100;
assign LUT_3[16917] = 32'b00000000000000001111010000001001;
assign LUT_3[16918] = 32'b00000000000000001010101100010000;
assign LUT_3[16919] = 32'b00000000000000010001010111101101;
assign LUT_3[16920] = 32'b00000000000000010000101111111100;
assign LUT_3[16921] = 32'b00000000000000010111011011011001;
assign LUT_3[16922] = 32'b00000000000000010010110111100000;
assign LUT_3[16923] = 32'b00000000000000011001100010111101;
assign LUT_3[16924] = 32'b00000000000000001101111101110010;
assign LUT_3[16925] = 32'b00000000000000010100101001001111;
assign LUT_3[16926] = 32'b00000000000000010000000101010110;
assign LUT_3[16927] = 32'b00000000000000010110110000110011;
assign LUT_3[16928] = 32'b00000000000000001001010010010011;
assign LUT_3[16929] = 32'b00000000000000001111111101110000;
assign LUT_3[16930] = 32'b00000000000000001011011001110111;
assign LUT_3[16931] = 32'b00000000000000010010000101010100;
assign LUT_3[16932] = 32'b00000000000000000110100000001001;
assign LUT_3[16933] = 32'b00000000000000001101001011100110;
assign LUT_3[16934] = 32'b00000000000000001000100111101101;
assign LUT_3[16935] = 32'b00000000000000001111010011001010;
assign LUT_3[16936] = 32'b00000000000000001110101011011001;
assign LUT_3[16937] = 32'b00000000000000010101010110110110;
assign LUT_3[16938] = 32'b00000000000000010000110010111101;
assign LUT_3[16939] = 32'b00000000000000010111011110011010;
assign LUT_3[16940] = 32'b00000000000000001011111001001111;
assign LUT_3[16941] = 32'b00000000000000010010100100101100;
assign LUT_3[16942] = 32'b00000000000000001110000000110011;
assign LUT_3[16943] = 32'b00000000000000010100101100010000;
assign LUT_3[16944] = 32'b00000000000000001100100101010110;
assign LUT_3[16945] = 32'b00000000000000010011010000110011;
assign LUT_3[16946] = 32'b00000000000000001110101100111010;
assign LUT_3[16947] = 32'b00000000000000010101011000010111;
assign LUT_3[16948] = 32'b00000000000000001001110011001100;
assign LUT_3[16949] = 32'b00000000000000010000011110101001;
assign LUT_3[16950] = 32'b00000000000000001011111010110000;
assign LUT_3[16951] = 32'b00000000000000010010100110001101;
assign LUT_3[16952] = 32'b00000000000000010001111110011100;
assign LUT_3[16953] = 32'b00000000000000011000101001111001;
assign LUT_3[16954] = 32'b00000000000000010100000110000000;
assign LUT_3[16955] = 32'b00000000000000011010110001011101;
assign LUT_3[16956] = 32'b00000000000000001111001100010010;
assign LUT_3[16957] = 32'b00000000000000010101110111101111;
assign LUT_3[16958] = 32'b00000000000000010001010011110110;
assign LUT_3[16959] = 32'b00000000000000010111111111010011;
assign LUT_3[16960] = 32'b00000000000000000111111100011110;
assign LUT_3[16961] = 32'b00000000000000001110100111111011;
assign LUT_3[16962] = 32'b00000000000000001010000100000010;
assign LUT_3[16963] = 32'b00000000000000010000101111011111;
assign LUT_3[16964] = 32'b00000000000000000101001010010100;
assign LUT_3[16965] = 32'b00000000000000001011110101110001;
assign LUT_3[16966] = 32'b00000000000000000111010001111000;
assign LUT_3[16967] = 32'b00000000000000001101111101010101;
assign LUT_3[16968] = 32'b00000000000000001101010101100100;
assign LUT_3[16969] = 32'b00000000000000010100000001000001;
assign LUT_3[16970] = 32'b00000000000000001111011101001000;
assign LUT_3[16971] = 32'b00000000000000010110001000100101;
assign LUT_3[16972] = 32'b00000000000000001010100011011010;
assign LUT_3[16973] = 32'b00000000000000010001001110110111;
assign LUT_3[16974] = 32'b00000000000000001100101010111110;
assign LUT_3[16975] = 32'b00000000000000010011010110011011;
assign LUT_3[16976] = 32'b00000000000000001011001111100001;
assign LUT_3[16977] = 32'b00000000000000010001111010111110;
assign LUT_3[16978] = 32'b00000000000000001101010111000101;
assign LUT_3[16979] = 32'b00000000000000010100000010100010;
assign LUT_3[16980] = 32'b00000000000000001000011101010111;
assign LUT_3[16981] = 32'b00000000000000001111001000110100;
assign LUT_3[16982] = 32'b00000000000000001010100100111011;
assign LUT_3[16983] = 32'b00000000000000010001010000011000;
assign LUT_3[16984] = 32'b00000000000000010000101000100111;
assign LUT_3[16985] = 32'b00000000000000010111010100000100;
assign LUT_3[16986] = 32'b00000000000000010010110000001011;
assign LUT_3[16987] = 32'b00000000000000011001011011101000;
assign LUT_3[16988] = 32'b00000000000000001101110110011101;
assign LUT_3[16989] = 32'b00000000000000010100100001111010;
assign LUT_3[16990] = 32'b00000000000000001111111110000001;
assign LUT_3[16991] = 32'b00000000000000010110101001011110;
assign LUT_3[16992] = 32'b00000000000000001001001010111110;
assign LUT_3[16993] = 32'b00000000000000001111110110011011;
assign LUT_3[16994] = 32'b00000000000000001011010010100010;
assign LUT_3[16995] = 32'b00000000000000010001111101111111;
assign LUT_3[16996] = 32'b00000000000000000110011000110100;
assign LUT_3[16997] = 32'b00000000000000001101000100010001;
assign LUT_3[16998] = 32'b00000000000000001000100000011000;
assign LUT_3[16999] = 32'b00000000000000001111001011110101;
assign LUT_3[17000] = 32'b00000000000000001110100100000100;
assign LUT_3[17001] = 32'b00000000000000010101001111100001;
assign LUT_3[17002] = 32'b00000000000000010000101011101000;
assign LUT_3[17003] = 32'b00000000000000010111010111000101;
assign LUT_3[17004] = 32'b00000000000000001011110001111010;
assign LUT_3[17005] = 32'b00000000000000010010011101010111;
assign LUT_3[17006] = 32'b00000000000000001101111001011110;
assign LUT_3[17007] = 32'b00000000000000010100100100111011;
assign LUT_3[17008] = 32'b00000000000000001100011110000001;
assign LUT_3[17009] = 32'b00000000000000010011001001011110;
assign LUT_3[17010] = 32'b00000000000000001110100101100101;
assign LUT_3[17011] = 32'b00000000000000010101010001000010;
assign LUT_3[17012] = 32'b00000000000000001001101011110111;
assign LUT_3[17013] = 32'b00000000000000010000010111010100;
assign LUT_3[17014] = 32'b00000000000000001011110011011011;
assign LUT_3[17015] = 32'b00000000000000010010011110111000;
assign LUT_3[17016] = 32'b00000000000000010001110111000111;
assign LUT_3[17017] = 32'b00000000000000011000100010100100;
assign LUT_3[17018] = 32'b00000000000000010011111110101011;
assign LUT_3[17019] = 32'b00000000000000011010101010001000;
assign LUT_3[17020] = 32'b00000000000000001111000100111101;
assign LUT_3[17021] = 32'b00000000000000010101110000011010;
assign LUT_3[17022] = 32'b00000000000000010001001100100001;
assign LUT_3[17023] = 32'b00000000000000010111110111111110;
assign LUT_3[17024] = 32'b00000000000000001010001110110001;
assign LUT_3[17025] = 32'b00000000000000010000111010001110;
assign LUT_3[17026] = 32'b00000000000000001100010110010101;
assign LUT_3[17027] = 32'b00000000000000010011000001110010;
assign LUT_3[17028] = 32'b00000000000000000111011100100111;
assign LUT_3[17029] = 32'b00000000000000001110001000000100;
assign LUT_3[17030] = 32'b00000000000000001001100100001011;
assign LUT_3[17031] = 32'b00000000000000010000001111101000;
assign LUT_3[17032] = 32'b00000000000000001111100111110111;
assign LUT_3[17033] = 32'b00000000000000010110010011010100;
assign LUT_3[17034] = 32'b00000000000000010001101111011011;
assign LUT_3[17035] = 32'b00000000000000011000011010111000;
assign LUT_3[17036] = 32'b00000000000000001100110101101101;
assign LUT_3[17037] = 32'b00000000000000010011100001001010;
assign LUT_3[17038] = 32'b00000000000000001110111101010001;
assign LUT_3[17039] = 32'b00000000000000010101101000101110;
assign LUT_3[17040] = 32'b00000000000000001101100001110100;
assign LUT_3[17041] = 32'b00000000000000010100001101010001;
assign LUT_3[17042] = 32'b00000000000000001111101001011000;
assign LUT_3[17043] = 32'b00000000000000010110010100110101;
assign LUT_3[17044] = 32'b00000000000000001010101111101010;
assign LUT_3[17045] = 32'b00000000000000010001011011000111;
assign LUT_3[17046] = 32'b00000000000000001100110111001110;
assign LUT_3[17047] = 32'b00000000000000010011100010101011;
assign LUT_3[17048] = 32'b00000000000000010010111010111010;
assign LUT_3[17049] = 32'b00000000000000011001100110010111;
assign LUT_3[17050] = 32'b00000000000000010101000010011110;
assign LUT_3[17051] = 32'b00000000000000011011101101111011;
assign LUT_3[17052] = 32'b00000000000000010000001000110000;
assign LUT_3[17053] = 32'b00000000000000010110110100001101;
assign LUT_3[17054] = 32'b00000000000000010010010000010100;
assign LUT_3[17055] = 32'b00000000000000011000111011110001;
assign LUT_3[17056] = 32'b00000000000000001011011101010001;
assign LUT_3[17057] = 32'b00000000000000010010001000101110;
assign LUT_3[17058] = 32'b00000000000000001101100100110101;
assign LUT_3[17059] = 32'b00000000000000010100010000010010;
assign LUT_3[17060] = 32'b00000000000000001000101011000111;
assign LUT_3[17061] = 32'b00000000000000001111010110100100;
assign LUT_3[17062] = 32'b00000000000000001010110010101011;
assign LUT_3[17063] = 32'b00000000000000010001011110001000;
assign LUT_3[17064] = 32'b00000000000000010000110110010111;
assign LUT_3[17065] = 32'b00000000000000010111100001110100;
assign LUT_3[17066] = 32'b00000000000000010010111101111011;
assign LUT_3[17067] = 32'b00000000000000011001101001011000;
assign LUT_3[17068] = 32'b00000000000000001110000100001101;
assign LUT_3[17069] = 32'b00000000000000010100101111101010;
assign LUT_3[17070] = 32'b00000000000000010000001011110001;
assign LUT_3[17071] = 32'b00000000000000010110110111001110;
assign LUT_3[17072] = 32'b00000000000000001110110000010100;
assign LUT_3[17073] = 32'b00000000000000010101011011110001;
assign LUT_3[17074] = 32'b00000000000000010000110111111000;
assign LUT_3[17075] = 32'b00000000000000010111100011010101;
assign LUT_3[17076] = 32'b00000000000000001011111110001010;
assign LUT_3[17077] = 32'b00000000000000010010101001100111;
assign LUT_3[17078] = 32'b00000000000000001110000101101110;
assign LUT_3[17079] = 32'b00000000000000010100110001001011;
assign LUT_3[17080] = 32'b00000000000000010100001001011010;
assign LUT_3[17081] = 32'b00000000000000011010110100110111;
assign LUT_3[17082] = 32'b00000000000000010110010000111110;
assign LUT_3[17083] = 32'b00000000000000011100111100011011;
assign LUT_3[17084] = 32'b00000000000000010001010111010000;
assign LUT_3[17085] = 32'b00000000000000011000000010101101;
assign LUT_3[17086] = 32'b00000000000000010011011110110100;
assign LUT_3[17087] = 32'b00000000000000011010001010010001;
assign LUT_3[17088] = 32'b00000000000000001010000111011100;
assign LUT_3[17089] = 32'b00000000000000010000110010111001;
assign LUT_3[17090] = 32'b00000000000000001100001111000000;
assign LUT_3[17091] = 32'b00000000000000010010111010011101;
assign LUT_3[17092] = 32'b00000000000000000111010101010010;
assign LUT_3[17093] = 32'b00000000000000001110000000101111;
assign LUT_3[17094] = 32'b00000000000000001001011100110110;
assign LUT_3[17095] = 32'b00000000000000010000001000010011;
assign LUT_3[17096] = 32'b00000000000000001111100000100010;
assign LUT_3[17097] = 32'b00000000000000010110001011111111;
assign LUT_3[17098] = 32'b00000000000000010001101000000110;
assign LUT_3[17099] = 32'b00000000000000011000010011100011;
assign LUT_3[17100] = 32'b00000000000000001100101110011000;
assign LUT_3[17101] = 32'b00000000000000010011011001110101;
assign LUT_3[17102] = 32'b00000000000000001110110101111100;
assign LUT_3[17103] = 32'b00000000000000010101100001011001;
assign LUT_3[17104] = 32'b00000000000000001101011010011111;
assign LUT_3[17105] = 32'b00000000000000010100000101111100;
assign LUT_3[17106] = 32'b00000000000000001111100010000011;
assign LUT_3[17107] = 32'b00000000000000010110001101100000;
assign LUT_3[17108] = 32'b00000000000000001010101000010101;
assign LUT_3[17109] = 32'b00000000000000010001010011110010;
assign LUT_3[17110] = 32'b00000000000000001100101111111001;
assign LUT_3[17111] = 32'b00000000000000010011011011010110;
assign LUT_3[17112] = 32'b00000000000000010010110011100101;
assign LUT_3[17113] = 32'b00000000000000011001011111000010;
assign LUT_3[17114] = 32'b00000000000000010100111011001001;
assign LUT_3[17115] = 32'b00000000000000011011100110100110;
assign LUT_3[17116] = 32'b00000000000000010000000001011011;
assign LUT_3[17117] = 32'b00000000000000010110101100111000;
assign LUT_3[17118] = 32'b00000000000000010010001000111111;
assign LUT_3[17119] = 32'b00000000000000011000110100011100;
assign LUT_3[17120] = 32'b00000000000000001011010101111100;
assign LUT_3[17121] = 32'b00000000000000010010000001011001;
assign LUT_3[17122] = 32'b00000000000000001101011101100000;
assign LUT_3[17123] = 32'b00000000000000010100001000111101;
assign LUT_3[17124] = 32'b00000000000000001000100011110010;
assign LUT_3[17125] = 32'b00000000000000001111001111001111;
assign LUT_3[17126] = 32'b00000000000000001010101011010110;
assign LUT_3[17127] = 32'b00000000000000010001010110110011;
assign LUT_3[17128] = 32'b00000000000000010000101111000010;
assign LUT_3[17129] = 32'b00000000000000010111011010011111;
assign LUT_3[17130] = 32'b00000000000000010010110110100110;
assign LUT_3[17131] = 32'b00000000000000011001100010000011;
assign LUT_3[17132] = 32'b00000000000000001101111100111000;
assign LUT_3[17133] = 32'b00000000000000010100101000010101;
assign LUT_3[17134] = 32'b00000000000000010000000100011100;
assign LUT_3[17135] = 32'b00000000000000010110101111111001;
assign LUT_3[17136] = 32'b00000000000000001110101000111111;
assign LUT_3[17137] = 32'b00000000000000010101010100011100;
assign LUT_3[17138] = 32'b00000000000000010000110000100011;
assign LUT_3[17139] = 32'b00000000000000010111011100000000;
assign LUT_3[17140] = 32'b00000000000000001011110110110101;
assign LUT_3[17141] = 32'b00000000000000010010100010010010;
assign LUT_3[17142] = 32'b00000000000000001101111110011001;
assign LUT_3[17143] = 32'b00000000000000010100101001110110;
assign LUT_3[17144] = 32'b00000000000000010100000010000101;
assign LUT_3[17145] = 32'b00000000000000011010101101100010;
assign LUT_3[17146] = 32'b00000000000000010110001001101001;
assign LUT_3[17147] = 32'b00000000000000011100110101000110;
assign LUT_3[17148] = 32'b00000000000000010001001111111011;
assign LUT_3[17149] = 32'b00000000000000010111111011011000;
assign LUT_3[17150] = 32'b00000000000000010011010111011111;
assign LUT_3[17151] = 32'b00000000000000011010000010111100;
assign LUT_3[17152] = 32'b00000000000000000100010011010100;
assign LUT_3[17153] = 32'b00000000000000001010111110110001;
assign LUT_3[17154] = 32'b00000000000000000110011010111000;
assign LUT_3[17155] = 32'b00000000000000001101000110010101;
assign LUT_3[17156] = 32'b00000000000000000001100001001010;
assign LUT_3[17157] = 32'b00000000000000001000001100100111;
assign LUT_3[17158] = 32'b00000000000000000011101000101110;
assign LUT_3[17159] = 32'b00000000000000001010010100001011;
assign LUT_3[17160] = 32'b00000000000000001001101100011010;
assign LUT_3[17161] = 32'b00000000000000010000010111110111;
assign LUT_3[17162] = 32'b00000000000000001011110011111110;
assign LUT_3[17163] = 32'b00000000000000010010011111011011;
assign LUT_3[17164] = 32'b00000000000000000110111010010000;
assign LUT_3[17165] = 32'b00000000000000001101100101101101;
assign LUT_3[17166] = 32'b00000000000000001001000001110100;
assign LUT_3[17167] = 32'b00000000000000001111101101010001;
assign LUT_3[17168] = 32'b00000000000000000111100110010111;
assign LUT_3[17169] = 32'b00000000000000001110010001110100;
assign LUT_3[17170] = 32'b00000000000000001001101101111011;
assign LUT_3[17171] = 32'b00000000000000010000011001011000;
assign LUT_3[17172] = 32'b00000000000000000100110100001101;
assign LUT_3[17173] = 32'b00000000000000001011011111101010;
assign LUT_3[17174] = 32'b00000000000000000110111011110001;
assign LUT_3[17175] = 32'b00000000000000001101100111001110;
assign LUT_3[17176] = 32'b00000000000000001100111111011101;
assign LUT_3[17177] = 32'b00000000000000010011101010111010;
assign LUT_3[17178] = 32'b00000000000000001111000111000001;
assign LUT_3[17179] = 32'b00000000000000010101110010011110;
assign LUT_3[17180] = 32'b00000000000000001010001101010011;
assign LUT_3[17181] = 32'b00000000000000010000111000110000;
assign LUT_3[17182] = 32'b00000000000000001100010100110111;
assign LUT_3[17183] = 32'b00000000000000010011000000010100;
assign LUT_3[17184] = 32'b00000000000000000101100001110100;
assign LUT_3[17185] = 32'b00000000000000001100001101010001;
assign LUT_3[17186] = 32'b00000000000000000111101001011000;
assign LUT_3[17187] = 32'b00000000000000001110010100110101;
assign LUT_3[17188] = 32'b00000000000000000010101111101010;
assign LUT_3[17189] = 32'b00000000000000001001011011000111;
assign LUT_3[17190] = 32'b00000000000000000100110111001110;
assign LUT_3[17191] = 32'b00000000000000001011100010101011;
assign LUT_3[17192] = 32'b00000000000000001010111010111010;
assign LUT_3[17193] = 32'b00000000000000010001100110010111;
assign LUT_3[17194] = 32'b00000000000000001101000010011110;
assign LUT_3[17195] = 32'b00000000000000010011101101111011;
assign LUT_3[17196] = 32'b00000000000000001000001000110000;
assign LUT_3[17197] = 32'b00000000000000001110110100001101;
assign LUT_3[17198] = 32'b00000000000000001010010000010100;
assign LUT_3[17199] = 32'b00000000000000010000111011110001;
assign LUT_3[17200] = 32'b00000000000000001000110100110111;
assign LUT_3[17201] = 32'b00000000000000001111100000010100;
assign LUT_3[17202] = 32'b00000000000000001010111100011011;
assign LUT_3[17203] = 32'b00000000000000010001100111111000;
assign LUT_3[17204] = 32'b00000000000000000110000010101101;
assign LUT_3[17205] = 32'b00000000000000001100101110001010;
assign LUT_3[17206] = 32'b00000000000000001000001010010001;
assign LUT_3[17207] = 32'b00000000000000001110110101101110;
assign LUT_3[17208] = 32'b00000000000000001110001101111101;
assign LUT_3[17209] = 32'b00000000000000010100111001011010;
assign LUT_3[17210] = 32'b00000000000000010000010101100001;
assign LUT_3[17211] = 32'b00000000000000010111000000111110;
assign LUT_3[17212] = 32'b00000000000000001011011011110011;
assign LUT_3[17213] = 32'b00000000000000010010000111010000;
assign LUT_3[17214] = 32'b00000000000000001101100011010111;
assign LUT_3[17215] = 32'b00000000000000010100001110110100;
assign LUT_3[17216] = 32'b00000000000000000100001011111111;
assign LUT_3[17217] = 32'b00000000000000001010110111011100;
assign LUT_3[17218] = 32'b00000000000000000110010011100011;
assign LUT_3[17219] = 32'b00000000000000001100111111000000;
assign LUT_3[17220] = 32'b00000000000000000001011001110101;
assign LUT_3[17221] = 32'b00000000000000001000000101010010;
assign LUT_3[17222] = 32'b00000000000000000011100001011001;
assign LUT_3[17223] = 32'b00000000000000001010001100110110;
assign LUT_3[17224] = 32'b00000000000000001001100101000101;
assign LUT_3[17225] = 32'b00000000000000010000010000100010;
assign LUT_3[17226] = 32'b00000000000000001011101100101001;
assign LUT_3[17227] = 32'b00000000000000010010011000000110;
assign LUT_3[17228] = 32'b00000000000000000110110010111011;
assign LUT_3[17229] = 32'b00000000000000001101011110011000;
assign LUT_3[17230] = 32'b00000000000000001000111010011111;
assign LUT_3[17231] = 32'b00000000000000001111100101111100;
assign LUT_3[17232] = 32'b00000000000000000111011111000010;
assign LUT_3[17233] = 32'b00000000000000001110001010011111;
assign LUT_3[17234] = 32'b00000000000000001001100110100110;
assign LUT_3[17235] = 32'b00000000000000010000010010000011;
assign LUT_3[17236] = 32'b00000000000000000100101100111000;
assign LUT_3[17237] = 32'b00000000000000001011011000010101;
assign LUT_3[17238] = 32'b00000000000000000110110100011100;
assign LUT_3[17239] = 32'b00000000000000001101011111111001;
assign LUT_3[17240] = 32'b00000000000000001100111000001000;
assign LUT_3[17241] = 32'b00000000000000010011100011100101;
assign LUT_3[17242] = 32'b00000000000000001110111111101100;
assign LUT_3[17243] = 32'b00000000000000010101101011001001;
assign LUT_3[17244] = 32'b00000000000000001010000101111110;
assign LUT_3[17245] = 32'b00000000000000010000110001011011;
assign LUT_3[17246] = 32'b00000000000000001100001101100010;
assign LUT_3[17247] = 32'b00000000000000010010111000111111;
assign LUT_3[17248] = 32'b00000000000000000101011010011111;
assign LUT_3[17249] = 32'b00000000000000001100000101111100;
assign LUT_3[17250] = 32'b00000000000000000111100010000011;
assign LUT_3[17251] = 32'b00000000000000001110001101100000;
assign LUT_3[17252] = 32'b00000000000000000010101000010101;
assign LUT_3[17253] = 32'b00000000000000001001010011110010;
assign LUT_3[17254] = 32'b00000000000000000100101111111001;
assign LUT_3[17255] = 32'b00000000000000001011011011010110;
assign LUT_3[17256] = 32'b00000000000000001010110011100101;
assign LUT_3[17257] = 32'b00000000000000010001011111000010;
assign LUT_3[17258] = 32'b00000000000000001100111011001001;
assign LUT_3[17259] = 32'b00000000000000010011100110100110;
assign LUT_3[17260] = 32'b00000000000000001000000001011011;
assign LUT_3[17261] = 32'b00000000000000001110101100111000;
assign LUT_3[17262] = 32'b00000000000000001010001000111111;
assign LUT_3[17263] = 32'b00000000000000010000110100011100;
assign LUT_3[17264] = 32'b00000000000000001000101101100010;
assign LUT_3[17265] = 32'b00000000000000001111011000111111;
assign LUT_3[17266] = 32'b00000000000000001010110101000110;
assign LUT_3[17267] = 32'b00000000000000010001100000100011;
assign LUT_3[17268] = 32'b00000000000000000101111011011000;
assign LUT_3[17269] = 32'b00000000000000001100100110110101;
assign LUT_3[17270] = 32'b00000000000000001000000010111100;
assign LUT_3[17271] = 32'b00000000000000001110101110011001;
assign LUT_3[17272] = 32'b00000000000000001110000110101000;
assign LUT_3[17273] = 32'b00000000000000010100110010000101;
assign LUT_3[17274] = 32'b00000000000000010000001110001100;
assign LUT_3[17275] = 32'b00000000000000010110111001101001;
assign LUT_3[17276] = 32'b00000000000000001011010100011110;
assign LUT_3[17277] = 32'b00000000000000010001111111111011;
assign LUT_3[17278] = 32'b00000000000000001101011100000010;
assign LUT_3[17279] = 32'b00000000000000010100000111011111;
assign LUT_3[17280] = 32'b00000000000000000110011110010010;
assign LUT_3[17281] = 32'b00000000000000001101001001101111;
assign LUT_3[17282] = 32'b00000000000000001000100101110110;
assign LUT_3[17283] = 32'b00000000000000001111010001010011;
assign LUT_3[17284] = 32'b00000000000000000011101100001000;
assign LUT_3[17285] = 32'b00000000000000001010010111100101;
assign LUT_3[17286] = 32'b00000000000000000101110011101100;
assign LUT_3[17287] = 32'b00000000000000001100011111001001;
assign LUT_3[17288] = 32'b00000000000000001011110111011000;
assign LUT_3[17289] = 32'b00000000000000010010100010110101;
assign LUT_3[17290] = 32'b00000000000000001101111110111100;
assign LUT_3[17291] = 32'b00000000000000010100101010011001;
assign LUT_3[17292] = 32'b00000000000000001001000101001110;
assign LUT_3[17293] = 32'b00000000000000001111110000101011;
assign LUT_3[17294] = 32'b00000000000000001011001100110010;
assign LUT_3[17295] = 32'b00000000000000010001111000001111;
assign LUT_3[17296] = 32'b00000000000000001001110001010101;
assign LUT_3[17297] = 32'b00000000000000010000011100110010;
assign LUT_3[17298] = 32'b00000000000000001011111000111001;
assign LUT_3[17299] = 32'b00000000000000010010100100010110;
assign LUT_3[17300] = 32'b00000000000000000110111111001011;
assign LUT_3[17301] = 32'b00000000000000001101101010101000;
assign LUT_3[17302] = 32'b00000000000000001001000110101111;
assign LUT_3[17303] = 32'b00000000000000001111110010001100;
assign LUT_3[17304] = 32'b00000000000000001111001010011011;
assign LUT_3[17305] = 32'b00000000000000010101110101111000;
assign LUT_3[17306] = 32'b00000000000000010001010001111111;
assign LUT_3[17307] = 32'b00000000000000010111111101011100;
assign LUT_3[17308] = 32'b00000000000000001100011000010001;
assign LUT_3[17309] = 32'b00000000000000010011000011101110;
assign LUT_3[17310] = 32'b00000000000000001110011111110101;
assign LUT_3[17311] = 32'b00000000000000010101001011010010;
assign LUT_3[17312] = 32'b00000000000000000111101100110010;
assign LUT_3[17313] = 32'b00000000000000001110011000001111;
assign LUT_3[17314] = 32'b00000000000000001001110100010110;
assign LUT_3[17315] = 32'b00000000000000010000011111110011;
assign LUT_3[17316] = 32'b00000000000000000100111010101000;
assign LUT_3[17317] = 32'b00000000000000001011100110000101;
assign LUT_3[17318] = 32'b00000000000000000111000010001100;
assign LUT_3[17319] = 32'b00000000000000001101101101101001;
assign LUT_3[17320] = 32'b00000000000000001101000101111000;
assign LUT_3[17321] = 32'b00000000000000010011110001010101;
assign LUT_3[17322] = 32'b00000000000000001111001101011100;
assign LUT_3[17323] = 32'b00000000000000010101111000111001;
assign LUT_3[17324] = 32'b00000000000000001010010011101110;
assign LUT_3[17325] = 32'b00000000000000010000111111001011;
assign LUT_3[17326] = 32'b00000000000000001100011011010010;
assign LUT_3[17327] = 32'b00000000000000010011000110101111;
assign LUT_3[17328] = 32'b00000000000000001010111111110101;
assign LUT_3[17329] = 32'b00000000000000010001101011010010;
assign LUT_3[17330] = 32'b00000000000000001101000111011001;
assign LUT_3[17331] = 32'b00000000000000010011110010110110;
assign LUT_3[17332] = 32'b00000000000000001000001101101011;
assign LUT_3[17333] = 32'b00000000000000001110111001001000;
assign LUT_3[17334] = 32'b00000000000000001010010101001111;
assign LUT_3[17335] = 32'b00000000000000010001000000101100;
assign LUT_3[17336] = 32'b00000000000000010000011000111011;
assign LUT_3[17337] = 32'b00000000000000010111000100011000;
assign LUT_3[17338] = 32'b00000000000000010010100000011111;
assign LUT_3[17339] = 32'b00000000000000011001001011111100;
assign LUT_3[17340] = 32'b00000000000000001101100110110001;
assign LUT_3[17341] = 32'b00000000000000010100010010001110;
assign LUT_3[17342] = 32'b00000000000000001111101110010101;
assign LUT_3[17343] = 32'b00000000000000010110011001110010;
assign LUT_3[17344] = 32'b00000000000000000110010110111101;
assign LUT_3[17345] = 32'b00000000000000001101000010011010;
assign LUT_3[17346] = 32'b00000000000000001000011110100001;
assign LUT_3[17347] = 32'b00000000000000001111001001111110;
assign LUT_3[17348] = 32'b00000000000000000011100100110011;
assign LUT_3[17349] = 32'b00000000000000001010010000010000;
assign LUT_3[17350] = 32'b00000000000000000101101100010111;
assign LUT_3[17351] = 32'b00000000000000001100010111110100;
assign LUT_3[17352] = 32'b00000000000000001011110000000011;
assign LUT_3[17353] = 32'b00000000000000010010011011100000;
assign LUT_3[17354] = 32'b00000000000000001101110111100111;
assign LUT_3[17355] = 32'b00000000000000010100100011000100;
assign LUT_3[17356] = 32'b00000000000000001000111101111001;
assign LUT_3[17357] = 32'b00000000000000001111101001010110;
assign LUT_3[17358] = 32'b00000000000000001011000101011101;
assign LUT_3[17359] = 32'b00000000000000010001110000111010;
assign LUT_3[17360] = 32'b00000000000000001001101010000000;
assign LUT_3[17361] = 32'b00000000000000010000010101011101;
assign LUT_3[17362] = 32'b00000000000000001011110001100100;
assign LUT_3[17363] = 32'b00000000000000010010011101000001;
assign LUT_3[17364] = 32'b00000000000000000110110111110110;
assign LUT_3[17365] = 32'b00000000000000001101100011010011;
assign LUT_3[17366] = 32'b00000000000000001000111111011010;
assign LUT_3[17367] = 32'b00000000000000001111101010110111;
assign LUT_3[17368] = 32'b00000000000000001111000011000110;
assign LUT_3[17369] = 32'b00000000000000010101101110100011;
assign LUT_3[17370] = 32'b00000000000000010001001010101010;
assign LUT_3[17371] = 32'b00000000000000010111110110000111;
assign LUT_3[17372] = 32'b00000000000000001100010000111100;
assign LUT_3[17373] = 32'b00000000000000010010111100011001;
assign LUT_3[17374] = 32'b00000000000000001110011000100000;
assign LUT_3[17375] = 32'b00000000000000010101000011111101;
assign LUT_3[17376] = 32'b00000000000000000111100101011101;
assign LUT_3[17377] = 32'b00000000000000001110010000111010;
assign LUT_3[17378] = 32'b00000000000000001001101101000001;
assign LUT_3[17379] = 32'b00000000000000010000011000011110;
assign LUT_3[17380] = 32'b00000000000000000100110011010011;
assign LUT_3[17381] = 32'b00000000000000001011011110110000;
assign LUT_3[17382] = 32'b00000000000000000110111010110111;
assign LUT_3[17383] = 32'b00000000000000001101100110010100;
assign LUT_3[17384] = 32'b00000000000000001100111110100011;
assign LUT_3[17385] = 32'b00000000000000010011101010000000;
assign LUT_3[17386] = 32'b00000000000000001111000110000111;
assign LUT_3[17387] = 32'b00000000000000010101110001100100;
assign LUT_3[17388] = 32'b00000000000000001010001100011001;
assign LUT_3[17389] = 32'b00000000000000010000110111110110;
assign LUT_3[17390] = 32'b00000000000000001100010011111101;
assign LUT_3[17391] = 32'b00000000000000010010111111011010;
assign LUT_3[17392] = 32'b00000000000000001010111000100000;
assign LUT_3[17393] = 32'b00000000000000010001100011111101;
assign LUT_3[17394] = 32'b00000000000000001101000000000100;
assign LUT_3[17395] = 32'b00000000000000010011101011100001;
assign LUT_3[17396] = 32'b00000000000000001000000110010110;
assign LUT_3[17397] = 32'b00000000000000001110110001110011;
assign LUT_3[17398] = 32'b00000000000000001010001101111010;
assign LUT_3[17399] = 32'b00000000000000010000111001010111;
assign LUT_3[17400] = 32'b00000000000000010000010001100110;
assign LUT_3[17401] = 32'b00000000000000010110111101000011;
assign LUT_3[17402] = 32'b00000000000000010010011001001010;
assign LUT_3[17403] = 32'b00000000000000011001000100100111;
assign LUT_3[17404] = 32'b00000000000000001101011111011100;
assign LUT_3[17405] = 32'b00000000000000010100001010111001;
assign LUT_3[17406] = 32'b00000000000000001111100111000000;
assign LUT_3[17407] = 32'b00000000000000010110010010011101;
assign LUT_3[17408] = 32'b00000000000000001011010011100100;
assign LUT_3[17409] = 32'b00000000000000010001111111000001;
assign LUT_3[17410] = 32'b00000000000000001101011011001000;
assign LUT_3[17411] = 32'b00000000000000010100000110100101;
assign LUT_3[17412] = 32'b00000000000000001000100001011010;
assign LUT_3[17413] = 32'b00000000000000001111001100110111;
assign LUT_3[17414] = 32'b00000000000000001010101000111110;
assign LUT_3[17415] = 32'b00000000000000010001010100011011;
assign LUT_3[17416] = 32'b00000000000000010000101100101010;
assign LUT_3[17417] = 32'b00000000000000010111011000000111;
assign LUT_3[17418] = 32'b00000000000000010010110100001110;
assign LUT_3[17419] = 32'b00000000000000011001011111101011;
assign LUT_3[17420] = 32'b00000000000000001101111010100000;
assign LUT_3[17421] = 32'b00000000000000010100100101111101;
assign LUT_3[17422] = 32'b00000000000000010000000010000100;
assign LUT_3[17423] = 32'b00000000000000010110101101100001;
assign LUT_3[17424] = 32'b00000000000000001110100110100111;
assign LUT_3[17425] = 32'b00000000000000010101010010000100;
assign LUT_3[17426] = 32'b00000000000000010000101110001011;
assign LUT_3[17427] = 32'b00000000000000010111011001101000;
assign LUT_3[17428] = 32'b00000000000000001011110100011101;
assign LUT_3[17429] = 32'b00000000000000010010011111111010;
assign LUT_3[17430] = 32'b00000000000000001101111100000001;
assign LUT_3[17431] = 32'b00000000000000010100100111011110;
assign LUT_3[17432] = 32'b00000000000000010011111111101101;
assign LUT_3[17433] = 32'b00000000000000011010101011001010;
assign LUT_3[17434] = 32'b00000000000000010110000111010001;
assign LUT_3[17435] = 32'b00000000000000011100110010101110;
assign LUT_3[17436] = 32'b00000000000000010001001101100011;
assign LUT_3[17437] = 32'b00000000000000010111111001000000;
assign LUT_3[17438] = 32'b00000000000000010011010101000111;
assign LUT_3[17439] = 32'b00000000000000011010000000100100;
assign LUT_3[17440] = 32'b00000000000000001100100010000100;
assign LUT_3[17441] = 32'b00000000000000010011001101100001;
assign LUT_3[17442] = 32'b00000000000000001110101001101000;
assign LUT_3[17443] = 32'b00000000000000010101010101000101;
assign LUT_3[17444] = 32'b00000000000000001001101111111010;
assign LUT_3[17445] = 32'b00000000000000010000011011010111;
assign LUT_3[17446] = 32'b00000000000000001011110111011110;
assign LUT_3[17447] = 32'b00000000000000010010100010111011;
assign LUT_3[17448] = 32'b00000000000000010001111011001010;
assign LUT_3[17449] = 32'b00000000000000011000100110100111;
assign LUT_3[17450] = 32'b00000000000000010100000010101110;
assign LUT_3[17451] = 32'b00000000000000011010101110001011;
assign LUT_3[17452] = 32'b00000000000000001111001001000000;
assign LUT_3[17453] = 32'b00000000000000010101110100011101;
assign LUT_3[17454] = 32'b00000000000000010001010000100100;
assign LUT_3[17455] = 32'b00000000000000010111111100000001;
assign LUT_3[17456] = 32'b00000000000000001111110101000111;
assign LUT_3[17457] = 32'b00000000000000010110100000100100;
assign LUT_3[17458] = 32'b00000000000000010001111100101011;
assign LUT_3[17459] = 32'b00000000000000011000101000001000;
assign LUT_3[17460] = 32'b00000000000000001101000010111101;
assign LUT_3[17461] = 32'b00000000000000010011101110011010;
assign LUT_3[17462] = 32'b00000000000000001111001010100001;
assign LUT_3[17463] = 32'b00000000000000010101110101111110;
assign LUT_3[17464] = 32'b00000000000000010101001110001101;
assign LUT_3[17465] = 32'b00000000000000011011111001101010;
assign LUT_3[17466] = 32'b00000000000000010111010101110001;
assign LUT_3[17467] = 32'b00000000000000011110000001001110;
assign LUT_3[17468] = 32'b00000000000000010010011100000011;
assign LUT_3[17469] = 32'b00000000000000011001000111100000;
assign LUT_3[17470] = 32'b00000000000000010100100011100111;
assign LUT_3[17471] = 32'b00000000000000011011001111000100;
assign LUT_3[17472] = 32'b00000000000000001011001100001111;
assign LUT_3[17473] = 32'b00000000000000010001110111101100;
assign LUT_3[17474] = 32'b00000000000000001101010011110011;
assign LUT_3[17475] = 32'b00000000000000010011111111010000;
assign LUT_3[17476] = 32'b00000000000000001000011010000101;
assign LUT_3[17477] = 32'b00000000000000001111000101100010;
assign LUT_3[17478] = 32'b00000000000000001010100001101001;
assign LUT_3[17479] = 32'b00000000000000010001001101000110;
assign LUT_3[17480] = 32'b00000000000000010000100101010101;
assign LUT_3[17481] = 32'b00000000000000010111010000110010;
assign LUT_3[17482] = 32'b00000000000000010010101100111001;
assign LUT_3[17483] = 32'b00000000000000011001011000010110;
assign LUT_3[17484] = 32'b00000000000000001101110011001011;
assign LUT_3[17485] = 32'b00000000000000010100011110101000;
assign LUT_3[17486] = 32'b00000000000000001111111010101111;
assign LUT_3[17487] = 32'b00000000000000010110100110001100;
assign LUT_3[17488] = 32'b00000000000000001110011111010010;
assign LUT_3[17489] = 32'b00000000000000010101001010101111;
assign LUT_3[17490] = 32'b00000000000000010000100110110110;
assign LUT_3[17491] = 32'b00000000000000010111010010010011;
assign LUT_3[17492] = 32'b00000000000000001011101101001000;
assign LUT_3[17493] = 32'b00000000000000010010011000100101;
assign LUT_3[17494] = 32'b00000000000000001101110100101100;
assign LUT_3[17495] = 32'b00000000000000010100100000001001;
assign LUT_3[17496] = 32'b00000000000000010011111000011000;
assign LUT_3[17497] = 32'b00000000000000011010100011110101;
assign LUT_3[17498] = 32'b00000000000000010101111111111100;
assign LUT_3[17499] = 32'b00000000000000011100101011011001;
assign LUT_3[17500] = 32'b00000000000000010001000110001110;
assign LUT_3[17501] = 32'b00000000000000010111110001101011;
assign LUT_3[17502] = 32'b00000000000000010011001101110010;
assign LUT_3[17503] = 32'b00000000000000011001111001001111;
assign LUT_3[17504] = 32'b00000000000000001100011010101111;
assign LUT_3[17505] = 32'b00000000000000010011000110001100;
assign LUT_3[17506] = 32'b00000000000000001110100010010011;
assign LUT_3[17507] = 32'b00000000000000010101001101110000;
assign LUT_3[17508] = 32'b00000000000000001001101000100101;
assign LUT_3[17509] = 32'b00000000000000010000010100000010;
assign LUT_3[17510] = 32'b00000000000000001011110000001001;
assign LUT_3[17511] = 32'b00000000000000010010011011100110;
assign LUT_3[17512] = 32'b00000000000000010001110011110101;
assign LUT_3[17513] = 32'b00000000000000011000011111010010;
assign LUT_3[17514] = 32'b00000000000000010011111011011001;
assign LUT_3[17515] = 32'b00000000000000011010100110110110;
assign LUT_3[17516] = 32'b00000000000000001111000001101011;
assign LUT_3[17517] = 32'b00000000000000010101101101001000;
assign LUT_3[17518] = 32'b00000000000000010001001001001111;
assign LUT_3[17519] = 32'b00000000000000010111110100101100;
assign LUT_3[17520] = 32'b00000000000000001111101101110010;
assign LUT_3[17521] = 32'b00000000000000010110011001001111;
assign LUT_3[17522] = 32'b00000000000000010001110101010110;
assign LUT_3[17523] = 32'b00000000000000011000100000110011;
assign LUT_3[17524] = 32'b00000000000000001100111011101000;
assign LUT_3[17525] = 32'b00000000000000010011100111000101;
assign LUT_3[17526] = 32'b00000000000000001111000011001100;
assign LUT_3[17527] = 32'b00000000000000010101101110101001;
assign LUT_3[17528] = 32'b00000000000000010101000110111000;
assign LUT_3[17529] = 32'b00000000000000011011110010010101;
assign LUT_3[17530] = 32'b00000000000000010111001110011100;
assign LUT_3[17531] = 32'b00000000000000011101111001111001;
assign LUT_3[17532] = 32'b00000000000000010010010100101110;
assign LUT_3[17533] = 32'b00000000000000011001000000001011;
assign LUT_3[17534] = 32'b00000000000000010100011100010010;
assign LUT_3[17535] = 32'b00000000000000011011000111101111;
assign LUT_3[17536] = 32'b00000000000000001101011110100010;
assign LUT_3[17537] = 32'b00000000000000010100001001111111;
assign LUT_3[17538] = 32'b00000000000000001111100110000110;
assign LUT_3[17539] = 32'b00000000000000010110010001100011;
assign LUT_3[17540] = 32'b00000000000000001010101100011000;
assign LUT_3[17541] = 32'b00000000000000010001010111110101;
assign LUT_3[17542] = 32'b00000000000000001100110011111100;
assign LUT_3[17543] = 32'b00000000000000010011011111011001;
assign LUT_3[17544] = 32'b00000000000000010010110111101000;
assign LUT_3[17545] = 32'b00000000000000011001100011000101;
assign LUT_3[17546] = 32'b00000000000000010100111111001100;
assign LUT_3[17547] = 32'b00000000000000011011101010101001;
assign LUT_3[17548] = 32'b00000000000000010000000101011110;
assign LUT_3[17549] = 32'b00000000000000010110110000111011;
assign LUT_3[17550] = 32'b00000000000000010010001101000010;
assign LUT_3[17551] = 32'b00000000000000011000111000011111;
assign LUT_3[17552] = 32'b00000000000000010000110001100101;
assign LUT_3[17553] = 32'b00000000000000010111011101000010;
assign LUT_3[17554] = 32'b00000000000000010010111001001001;
assign LUT_3[17555] = 32'b00000000000000011001100100100110;
assign LUT_3[17556] = 32'b00000000000000001101111111011011;
assign LUT_3[17557] = 32'b00000000000000010100101010111000;
assign LUT_3[17558] = 32'b00000000000000010000000110111111;
assign LUT_3[17559] = 32'b00000000000000010110110010011100;
assign LUT_3[17560] = 32'b00000000000000010110001010101011;
assign LUT_3[17561] = 32'b00000000000000011100110110001000;
assign LUT_3[17562] = 32'b00000000000000011000010010001111;
assign LUT_3[17563] = 32'b00000000000000011110111101101100;
assign LUT_3[17564] = 32'b00000000000000010011011000100001;
assign LUT_3[17565] = 32'b00000000000000011010000011111110;
assign LUT_3[17566] = 32'b00000000000000010101100000000101;
assign LUT_3[17567] = 32'b00000000000000011100001011100010;
assign LUT_3[17568] = 32'b00000000000000001110101101000010;
assign LUT_3[17569] = 32'b00000000000000010101011000011111;
assign LUT_3[17570] = 32'b00000000000000010000110100100110;
assign LUT_3[17571] = 32'b00000000000000010111100000000011;
assign LUT_3[17572] = 32'b00000000000000001011111010111000;
assign LUT_3[17573] = 32'b00000000000000010010100110010101;
assign LUT_3[17574] = 32'b00000000000000001110000010011100;
assign LUT_3[17575] = 32'b00000000000000010100101101111001;
assign LUT_3[17576] = 32'b00000000000000010100000110001000;
assign LUT_3[17577] = 32'b00000000000000011010110001100101;
assign LUT_3[17578] = 32'b00000000000000010110001101101100;
assign LUT_3[17579] = 32'b00000000000000011100111001001001;
assign LUT_3[17580] = 32'b00000000000000010001010011111110;
assign LUT_3[17581] = 32'b00000000000000010111111111011011;
assign LUT_3[17582] = 32'b00000000000000010011011011100010;
assign LUT_3[17583] = 32'b00000000000000011010000110111111;
assign LUT_3[17584] = 32'b00000000000000010010000000000101;
assign LUT_3[17585] = 32'b00000000000000011000101011100010;
assign LUT_3[17586] = 32'b00000000000000010100000111101001;
assign LUT_3[17587] = 32'b00000000000000011010110011000110;
assign LUT_3[17588] = 32'b00000000000000001111001101111011;
assign LUT_3[17589] = 32'b00000000000000010101111001011000;
assign LUT_3[17590] = 32'b00000000000000010001010101011111;
assign LUT_3[17591] = 32'b00000000000000011000000000111100;
assign LUT_3[17592] = 32'b00000000000000010111011001001011;
assign LUT_3[17593] = 32'b00000000000000011110000100101000;
assign LUT_3[17594] = 32'b00000000000000011001100000101111;
assign LUT_3[17595] = 32'b00000000000000100000001100001100;
assign LUT_3[17596] = 32'b00000000000000010100100111000001;
assign LUT_3[17597] = 32'b00000000000000011011010010011110;
assign LUT_3[17598] = 32'b00000000000000010110101110100101;
assign LUT_3[17599] = 32'b00000000000000011101011010000010;
assign LUT_3[17600] = 32'b00000000000000001101010111001101;
assign LUT_3[17601] = 32'b00000000000000010100000010101010;
assign LUT_3[17602] = 32'b00000000000000001111011110110001;
assign LUT_3[17603] = 32'b00000000000000010110001010001110;
assign LUT_3[17604] = 32'b00000000000000001010100101000011;
assign LUT_3[17605] = 32'b00000000000000010001010000100000;
assign LUT_3[17606] = 32'b00000000000000001100101100100111;
assign LUT_3[17607] = 32'b00000000000000010011011000000100;
assign LUT_3[17608] = 32'b00000000000000010010110000010011;
assign LUT_3[17609] = 32'b00000000000000011001011011110000;
assign LUT_3[17610] = 32'b00000000000000010100110111110111;
assign LUT_3[17611] = 32'b00000000000000011011100011010100;
assign LUT_3[17612] = 32'b00000000000000001111111110001001;
assign LUT_3[17613] = 32'b00000000000000010110101001100110;
assign LUT_3[17614] = 32'b00000000000000010010000101101101;
assign LUT_3[17615] = 32'b00000000000000011000110001001010;
assign LUT_3[17616] = 32'b00000000000000010000101010010000;
assign LUT_3[17617] = 32'b00000000000000010111010101101101;
assign LUT_3[17618] = 32'b00000000000000010010110001110100;
assign LUT_3[17619] = 32'b00000000000000011001011101010001;
assign LUT_3[17620] = 32'b00000000000000001101111000000110;
assign LUT_3[17621] = 32'b00000000000000010100100011100011;
assign LUT_3[17622] = 32'b00000000000000001111111111101010;
assign LUT_3[17623] = 32'b00000000000000010110101011000111;
assign LUT_3[17624] = 32'b00000000000000010110000011010110;
assign LUT_3[17625] = 32'b00000000000000011100101110110011;
assign LUT_3[17626] = 32'b00000000000000011000001010111010;
assign LUT_3[17627] = 32'b00000000000000011110110110010111;
assign LUT_3[17628] = 32'b00000000000000010011010001001100;
assign LUT_3[17629] = 32'b00000000000000011001111100101001;
assign LUT_3[17630] = 32'b00000000000000010101011000110000;
assign LUT_3[17631] = 32'b00000000000000011100000100001101;
assign LUT_3[17632] = 32'b00000000000000001110100101101101;
assign LUT_3[17633] = 32'b00000000000000010101010001001010;
assign LUT_3[17634] = 32'b00000000000000010000101101010001;
assign LUT_3[17635] = 32'b00000000000000010111011000101110;
assign LUT_3[17636] = 32'b00000000000000001011110011100011;
assign LUT_3[17637] = 32'b00000000000000010010011111000000;
assign LUT_3[17638] = 32'b00000000000000001101111011000111;
assign LUT_3[17639] = 32'b00000000000000010100100110100100;
assign LUT_3[17640] = 32'b00000000000000010011111110110011;
assign LUT_3[17641] = 32'b00000000000000011010101010010000;
assign LUT_3[17642] = 32'b00000000000000010110000110010111;
assign LUT_3[17643] = 32'b00000000000000011100110001110100;
assign LUT_3[17644] = 32'b00000000000000010001001100101001;
assign LUT_3[17645] = 32'b00000000000000010111111000000110;
assign LUT_3[17646] = 32'b00000000000000010011010100001101;
assign LUT_3[17647] = 32'b00000000000000011001111111101010;
assign LUT_3[17648] = 32'b00000000000000010001111000110000;
assign LUT_3[17649] = 32'b00000000000000011000100100001101;
assign LUT_3[17650] = 32'b00000000000000010100000000010100;
assign LUT_3[17651] = 32'b00000000000000011010101011110001;
assign LUT_3[17652] = 32'b00000000000000001111000110100110;
assign LUT_3[17653] = 32'b00000000000000010101110010000011;
assign LUT_3[17654] = 32'b00000000000000010001001110001010;
assign LUT_3[17655] = 32'b00000000000000010111111001100111;
assign LUT_3[17656] = 32'b00000000000000010111010001110110;
assign LUT_3[17657] = 32'b00000000000000011101111101010011;
assign LUT_3[17658] = 32'b00000000000000011001011001011010;
assign LUT_3[17659] = 32'b00000000000000100000000100110111;
assign LUT_3[17660] = 32'b00000000000000010100011111101100;
assign LUT_3[17661] = 32'b00000000000000011011001011001001;
assign LUT_3[17662] = 32'b00000000000000010110100111010000;
assign LUT_3[17663] = 32'b00000000000000011101010010101101;
assign LUT_3[17664] = 32'b00000000000000000111100011000101;
assign LUT_3[17665] = 32'b00000000000000001110001110100010;
assign LUT_3[17666] = 32'b00000000000000001001101010101001;
assign LUT_3[17667] = 32'b00000000000000010000010110000110;
assign LUT_3[17668] = 32'b00000000000000000100110000111011;
assign LUT_3[17669] = 32'b00000000000000001011011100011000;
assign LUT_3[17670] = 32'b00000000000000000110111000011111;
assign LUT_3[17671] = 32'b00000000000000001101100011111100;
assign LUT_3[17672] = 32'b00000000000000001100111100001011;
assign LUT_3[17673] = 32'b00000000000000010011100111101000;
assign LUT_3[17674] = 32'b00000000000000001111000011101111;
assign LUT_3[17675] = 32'b00000000000000010101101111001100;
assign LUT_3[17676] = 32'b00000000000000001010001010000001;
assign LUT_3[17677] = 32'b00000000000000010000110101011110;
assign LUT_3[17678] = 32'b00000000000000001100010001100101;
assign LUT_3[17679] = 32'b00000000000000010010111101000010;
assign LUT_3[17680] = 32'b00000000000000001010110110001000;
assign LUT_3[17681] = 32'b00000000000000010001100001100101;
assign LUT_3[17682] = 32'b00000000000000001100111101101100;
assign LUT_3[17683] = 32'b00000000000000010011101001001001;
assign LUT_3[17684] = 32'b00000000000000001000000011111110;
assign LUT_3[17685] = 32'b00000000000000001110101111011011;
assign LUT_3[17686] = 32'b00000000000000001010001011100010;
assign LUT_3[17687] = 32'b00000000000000010000110110111111;
assign LUT_3[17688] = 32'b00000000000000010000001111001110;
assign LUT_3[17689] = 32'b00000000000000010110111010101011;
assign LUT_3[17690] = 32'b00000000000000010010010110110010;
assign LUT_3[17691] = 32'b00000000000000011001000010001111;
assign LUT_3[17692] = 32'b00000000000000001101011101000100;
assign LUT_3[17693] = 32'b00000000000000010100001000100001;
assign LUT_3[17694] = 32'b00000000000000001111100100101000;
assign LUT_3[17695] = 32'b00000000000000010110010000000101;
assign LUT_3[17696] = 32'b00000000000000001000110001100101;
assign LUT_3[17697] = 32'b00000000000000001111011101000010;
assign LUT_3[17698] = 32'b00000000000000001010111001001001;
assign LUT_3[17699] = 32'b00000000000000010001100100100110;
assign LUT_3[17700] = 32'b00000000000000000101111111011011;
assign LUT_3[17701] = 32'b00000000000000001100101010111000;
assign LUT_3[17702] = 32'b00000000000000001000000110111111;
assign LUT_3[17703] = 32'b00000000000000001110110010011100;
assign LUT_3[17704] = 32'b00000000000000001110001010101011;
assign LUT_3[17705] = 32'b00000000000000010100110110001000;
assign LUT_3[17706] = 32'b00000000000000010000010010001111;
assign LUT_3[17707] = 32'b00000000000000010110111101101100;
assign LUT_3[17708] = 32'b00000000000000001011011000100001;
assign LUT_3[17709] = 32'b00000000000000010010000011111110;
assign LUT_3[17710] = 32'b00000000000000001101100000000101;
assign LUT_3[17711] = 32'b00000000000000010100001011100010;
assign LUT_3[17712] = 32'b00000000000000001100000100101000;
assign LUT_3[17713] = 32'b00000000000000010010110000000101;
assign LUT_3[17714] = 32'b00000000000000001110001100001100;
assign LUT_3[17715] = 32'b00000000000000010100110111101001;
assign LUT_3[17716] = 32'b00000000000000001001010010011110;
assign LUT_3[17717] = 32'b00000000000000001111111101111011;
assign LUT_3[17718] = 32'b00000000000000001011011010000010;
assign LUT_3[17719] = 32'b00000000000000010010000101011111;
assign LUT_3[17720] = 32'b00000000000000010001011101101110;
assign LUT_3[17721] = 32'b00000000000000011000001001001011;
assign LUT_3[17722] = 32'b00000000000000010011100101010010;
assign LUT_3[17723] = 32'b00000000000000011010010000101111;
assign LUT_3[17724] = 32'b00000000000000001110101011100100;
assign LUT_3[17725] = 32'b00000000000000010101010111000001;
assign LUT_3[17726] = 32'b00000000000000010000110011001000;
assign LUT_3[17727] = 32'b00000000000000010111011110100101;
assign LUT_3[17728] = 32'b00000000000000000111011011110000;
assign LUT_3[17729] = 32'b00000000000000001110000111001101;
assign LUT_3[17730] = 32'b00000000000000001001100011010100;
assign LUT_3[17731] = 32'b00000000000000010000001110110001;
assign LUT_3[17732] = 32'b00000000000000000100101001100110;
assign LUT_3[17733] = 32'b00000000000000001011010101000011;
assign LUT_3[17734] = 32'b00000000000000000110110001001010;
assign LUT_3[17735] = 32'b00000000000000001101011100100111;
assign LUT_3[17736] = 32'b00000000000000001100110100110110;
assign LUT_3[17737] = 32'b00000000000000010011100000010011;
assign LUT_3[17738] = 32'b00000000000000001110111100011010;
assign LUT_3[17739] = 32'b00000000000000010101100111110111;
assign LUT_3[17740] = 32'b00000000000000001010000010101100;
assign LUT_3[17741] = 32'b00000000000000010000101110001001;
assign LUT_3[17742] = 32'b00000000000000001100001010010000;
assign LUT_3[17743] = 32'b00000000000000010010110101101101;
assign LUT_3[17744] = 32'b00000000000000001010101110110011;
assign LUT_3[17745] = 32'b00000000000000010001011010010000;
assign LUT_3[17746] = 32'b00000000000000001100110110010111;
assign LUT_3[17747] = 32'b00000000000000010011100001110100;
assign LUT_3[17748] = 32'b00000000000000000111111100101001;
assign LUT_3[17749] = 32'b00000000000000001110101000000110;
assign LUT_3[17750] = 32'b00000000000000001010000100001101;
assign LUT_3[17751] = 32'b00000000000000010000101111101010;
assign LUT_3[17752] = 32'b00000000000000010000000111111001;
assign LUT_3[17753] = 32'b00000000000000010110110011010110;
assign LUT_3[17754] = 32'b00000000000000010010001111011101;
assign LUT_3[17755] = 32'b00000000000000011000111010111010;
assign LUT_3[17756] = 32'b00000000000000001101010101101111;
assign LUT_3[17757] = 32'b00000000000000010100000001001100;
assign LUT_3[17758] = 32'b00000000000000001111011101010011;
assign LUT_3[17759] = 32'b00000000000000010110001000110000;
assign LUT_3[17760] = 32'b00000000000000001000101010010000;
assign LUT_3[17761] = 32'b00000000000000001111010101101101;
assign LUT_3[17762] = 32'b00000000000000001010110001110100;
assign LUT_3[17763] = 32'b00000000000000010001011101010001;
assign LUT_3[17764] = 32'b00000000000000000101111000000110;
assign LUT_3[17765] = 32'b00000000000000001100100011100011;
assign LUT_3[17766] = 32'b00000000000000000111111111101010;
assign LUT_3[17767] = 32'b00000000000000001110101011000111;
assign LUT_3[17768] = 32'b00000000000000001110000011010110;
assign LUT_3[17769] = 32'b00000000000000010100101110110011;
assign LUT_3[17770] = 32'b00000000000000010000001010111010;
assign LUT_3[17771] = 32'b00000000000000010110110110010111;
assign LUT_3[17772] = 32'b00000000000000001011010001001100;
assign LUT_3[17773] = 32'b00000000000000010001111100101001;
assign LUT_3[17774] = 32'b00000000000000001101011000110000;
assign LUT_3[17775] = 32'b00000000000000010100000100001101;
assign LUT_3[17776] = 32'b00000000000000001011111101010011;
assign LUT_3[17777] = 32'b00000000000000010010101000110000;
assign LUT_3[17778] = 32'b00000000000000001110000100110111;
assign LUT_3[17779] = 32'b00000000000000010100110000010100;
assign LUT_3[17780] = 32'b00000000000000001001001011001001;
assign LUT_3[17781] = 32'b00000000000000001111110110100110;
assign LUT_3[17782] = 32'b00000000000000001011010010101101;
assign LUT_3[17783] = 32'b00000000000000010001111110001010;
assign LUT_3[17784] = 32'b00000000000000010001010110011001;
assign LUT_3[17785] = 32'b00000000000000011000000001110110;
assign LUT_3[17786] = 32'b00000000000000010011011101111101;
assign LUT_3[17787] = 32'b00000000000000011010001001011010;
assign LUT_3[17788] = 32'b00000000000000001110100100001111;
assign LUT_3[17789] = 32'b00000000000000010101001111101100;
assign LUT_3[17790] = 32'b00000000000000010000101011110011;
assign LUT_3[17791] = 32'b00000000000000010111010111010000;
assign LUT_3[17792] = 32'b00000000000000001001101110000011;
assign LUT_3[17793] = 32'b00000000000000010000011001100000;
assign LUT_3[17794] = 32'b00000000000000001011110101100111;
assign LUT_3[17795] = 32'b00000000000000010010100001000100;
assign LUT_3[17796] = 32'b00000000000000000110111011111001;
assign LUT_3[17797] = 32'b00000000000000001101100111010110;
assign LUT_3[17798] = 32'b00000000000000001001000011011101;
assign LUT_3[17799] = 32'b00000000000000001111101110111010;
assign LUT_3[17800] = 32'b00000000000000001111000111001001;
assign LUT_3[17801] = 32'b00000000000000010101110010100110;
assign LUT_3[17802] = 32'b00000000000000010001001110101101;
assign LUT_3[17803] = 32'b00000000000000010111111010001010;
assign LUT_3[17804] = 32'b00000000000000001100010100111111;
assign LUT_3[17805] = 32'b00000000000000010011000000011100;
assign LUT_3[17806] = 32'b00000000000000001110011100100011;
assign LUT_3[17807] = 32'b00000000000000010101001000000000;
assign LUT_3[17808] = 32'b00000000000000001101000001000110;
assign LUT_3[17809] = 32'b00000000000000010011101100100011;
assign LUT_3[17810] = 32'b00000000000000001111001000101010;
assign LUT_3[17811] = 32'b00000000000000010101110100000111;
assign LUT_3[17812] = 32'b00000000000000001010001110111100;
assign LUT_3[17813] = 32'b00000000000000010000111010011001;
assign LUT_3[17814] = 32'b00000000000000001100010110100000;
assign LUT_3[17815] = 32'b00000000000000010011000001111101;
assign LUT_3[17816] = 32'b00000000000000010010011010001100;
assign LUT_3[17817] = 32'b00000000000000011001000101101001;
assign LUT_3[17818] = 32'b00000000000000010100100001110000;
assign LUT_3[17819] = 32'b00000000000000011011001101001101;
assign LUT_3[17820] = 32'b00000000000000001111101000000010;
assign LUT_3[17821] = 32'b00000000000000010110010011011111;
assign LUT_3[17822] = 32'b00000000000000010001101111100110;
assign LUT_3[17823] = 32'b00000000000000011000011011000011;
assign LUT_3[17824] = 32'b00000000000000001010111100100011;
assign LUT_3[17825] = 32'b00000000000000010001101000000000;
assign LUT_3[17826] = 32'b00000000000000001101000100000111;
assign LUT_3[17827] = 32'b00000000000000010011101111100100;
assign LUT_3[17828] = 32'b00000000000000001000001010011001;
assign LUT_3[17829] = 32'b00000000000000001110110101110110;
assign LUT_3[17830] = 32'b00000000000000001010010001111101;
assign LUT_3[17831] = 32'b00000000000000010000111101011010;
assign LUT_3[17832] = 32'b00000000000000010000010101101001;
assign LUT_3[17833] = 32'b00000000000000010111000001000110;
assign LUT_3[17834] = 32'b00000000000000010010011101001101;
assign LUT_3[17835] = 32'b00000000000000011001001000101010;
assign LUT_3[17836] = 32'b00000000000000001101100011011111;
assign LUT_3[17837] = 32'b00000000000000010100001110111100;
assign LUT_3[17838] = 32'b00000000000000001111101011000011;
assign LUT_3[17839] = 32'b00000000000000010110010110100000;
assign LUT_3[17840] = 32'b00000000000000001110001111100110;
assign LUT_3[17841] = 32'b00000000000000010100111011000011;
assign LUT_3[17842] = 32'b00000000000000010000010111001010;
assign LUT_3[17843] = 32'b00000000000000010111000010100111;
assign LUT_3[17844] = 32'b00000000000000001011011101011100;
assign LUT_3[17845] = 32'b00000000000000010010001000111001;
assign LUT_3[17846] = 32'b00000000000000001101100101000000;
assign LUT_3[17847] = 32'b00000000000000010100010000011101;
assign LUT_3[17848] = 32'b00000000000000010011101000101100;
assign LUT_3[17849] = 32'b00000000000000011010010100001001;
assign LUT_3[17850] = 32'b00000000000000010101110000010000;
assign LUT_3[17851] = 32'b00000000000000011100011011101101;
assign LUT_3[17852] = 32'b00000000000000010000110110100010;
assign LUT_3[17853] = 32'b00000000000000010111100001111111;
assign LUT_3[17854] = 32'b00000000000000010010111110000110;
assign LUT_3[17855] = 32'b00000000000000011001101001100011;
assign LUT_3[17856] = 32'b00000000000000001001100110101110;
assign LUT_3[17857] = 32'b00000000000000010000010010001011;
assign LUT_3[17858] = 32'b00000000000000001011101110010010;
assign LUT_3[17859] = 32'b00000000000000010010011001101111;
assign LUT_3[17860] = 32'b00000000000000000110110100100100;
assign LUT_3[17861] = 32'b00000000000000001101100000000001;
assign LUT_3[17862] = 32'b00000000000000001000111100001000;
assign LUT_3[17863] = 32'b00000000000000001111100111100101;
assign LUT_3[17864] = 32'b00000000000000001110111111110100;
assign LUT_3[17865] = 32'b00000000000000010101101011010001;
assign LUT_3[17866] = 32'b00000000000000010001000111011000;
assign LUT_3[17867] = 32'b00000000000000010111110010110101;
assign LUT_3[17868] = 32'b00000000000000001100001101101010;
assign LUT_3[17869] = 32'b00000000000000010010111001000111;
assign LUT_3[17870] = 32'b00000000000000001110010101001110;
assign LUT_3[17871] = 32'b00000000000000010101000000101011;
assign LUT_3[17872] = 32'b00000000000000001100111001110001;
assign LUT_3[17873] = 32'b00000000000000010011100101001110;
assign LUT_3[17874] = 32'b00000000000000001111000001010101;
assign LUT_3[17875] = 32'b00000000000000010101101100110010;
assign LUT_3[17876] = 32'b00000000000000001010000111100111;
assign LUT_3[17877] = 32'b00000000000000010000110011000100;
assign LUT_3[17878] = 32'b00000000000000001100001111001011;
assign LUT_3[17879] = 32'b00000000000000010010111010101000;
assign LUT_3[17880] = 32'b00000000000000010010010010110111;
assign LUT_3[17881] = 32'b00000000000000011000111110010100;
assign LUT_3[17882] = 32'b00000000000000010100011010011011;
assign LUT_3[17883] = 32'b00000000000000011011000101111000;
assign LUT_3[17884] = 32'b00000000000000001111100000101101;
assign LUT_3[17885] = 32'b00000000000000010110001100001010;
assign LUT_3[17886] = 32'b00000000000000010001101000010001;
assign LUT_3[17887] = 32'b00000000000000011000010011101110;
assign LUT_3[17888] = 32'b00000000000000001010110101001110;
assign LUT_3[17889] = 32'b00000000000000010001100000101011;
assign LUT_3[17890] = 32'b00000000000000001100111100110010;
assign LUT_3[17891] = 32'b00000000000000010011101000001111;
assign LUT_3[17892] = 32'b00000000000000001000000011000100;
assign LUT_3[17893] = 32'b00000000000000001110101110100001;
assign LUT_3[17894] = 32'b00000000000000001010001010101000;
assign LUT_3[17895] = 32'b00000000000000010000110110000101;
assign LUT_3[17896] = 32'b00000000000000010000001110010100;
assign LUT_3[17897] = 32'b00000000000000010110111001110001;
assign LUT_3[17898] = 32'b00000000000000010010010101111000;
assign LUT_3[17899] = 32'b00000000000000011001000001010101;
assign LUT_3[17900] = 32'b00000000000000001101011100001010;
assign LUT_3[17901] = 32'b00000000000000010100000111100111;
assign LUT_3[17902] = 32'b00000000000000001111100011101110;
assign LUT_3[17903] = 32'b00000000000000010110001111001011;
assign LUT_3[17904] = 32'b00000000000000001110001000010001;
assign LUT_3[17905] = 32'b00000000000000010100110011101110;
assign LUT_3[17906] = 32'b00000000000000010000001111110101;
assign LUT_3[17907] = 32'b00000000000000010110111011010010;
assign LUT_3[17908] = 32'b00000000000000001011010110000111;
assign LUT_3[17909] = 32'b00000000000000010010000001100100;
assign LUT_3[17910] = 32'b00000000000000001101011101101011;
assign LUT_3[17911] = 32'b00000000000000010100001001001000;
assign LUT_3[17912] = 32'b00000000000000010011100001010111;
assign LUT_3[17913] = 32'b00000000000000011010001100110100;
assign LUT_3[17914] = 32'b00000000000000010101101000111011;
assign LUT_3[17915] = 32'b00000000000000011100010100011000;
assign LUT_3[17916] = 32'b00000000000000010000101111001101;
assign LUT_3[17917] = 32'b00000000000000010111011010101010;
assign LUT_3[17918] = 32'b00000000000000010010110110110001;
assign LUT_3[17919] = 32'b00000000000000011001100010001110;
assign LUT_3[17920] = 32'b00000000000000001110101000110000;
assign LUT_3[17921] = 32'b00000000000000010101010100001101;
assign LUT_3[17922] = 32'b00000000000000010000110000010100;
assign LUT_3[17923] = 32'b00000000000000010111011011110001;
assign LUT_3[17924] = 32'b00000000000000001011110110100110;
assign LUT_3[17925] = 32'b00000000000000010010100010000011;
assign LUT_3[17926] = 32'b00000000000000001101111110001010;
assign LUT_3[17927] = 32'b00000000000000010100101001100111;
assign LUT_3[17928] = 32'b00000000000000010100000001110110;
assign LUT_3[17929] = 32'b00000000000000011010101101010011;
assign LUT_3[17930] = 32'b00000000000000010110001001011010;
assign LUT_3[17931] = 32'b00000000000000011100110100110111;
assign LUT_3[17932] = 32'b00000000000000010001001111101100;
assign LUT_3[17933] = 32'b00000000000000010111111011001001;
assign LUT_3[17934] = 32'b00000000000000010011010111010000;
assign LUT_3[17935] = 32'b00000000000000011010000010101101;
assign LUT_3[17936] = 32'b00000000000000010001111011110011;
assign LUT_3[17937] = 32'b00000000000000011000100111010000;
assign LUT_3[17938] = 32'b00000000000000010100000011010111;
assign LUT_3[17939] = 32'b00000000000000011010101110110100;
assign LUT_3[17940] = 32'b00000000000000001111001001101001;
assign LUT_3[17941] = 32'b00000000000000010101110101000110;
assign LUT_3[17942] = 32'b00000000000000010001010001001101;
assign LUT_3[17943] = 32'b00000000000000010111111100101010;
assign LUT_3[17944] = 32'b00000000000000010111010100111001;
assign LUT_3[17945] = 32'b00000000000000011110000000010110;
assign LUT_3[17946] = 32'b00000000000000011001011100011101;
assign LUT_3[17947] = 32'b00000000000000100000000111111010;
assign LUT_3[17948] = 32'b00000000000000010100100010101111;
assign LUT_3[17949] = 32'b00000000000000011011001110001100;
assign LUT_3[17950] = 32'b00000000000000010110101010010011;
assign LUT_3[17951] = 32'b00000000000000011101010101110000;
assign LUT_3[17952] = 32'b00000000000000001111110111010000;
assign LUT_3[17953] = 32'b00000000000000010110100010101101;
assign LUT_3[17954] = 32'b00000000000000010001111110110100;
assign LUT_3[17955] = 32'b00000000000000011000101010010001;
assign LUT_3[17956] = 32'b00000000000000001101000101000110;
assign LUT_3[17957] = 32'b00000000000000010011110000100011;
assign LUT_3[17958] = 32'b00000000000000001111001100101010;
assign LUT_3[17959] = 32'b00000000000000010101111000000111;
assign LUT_3[17960] = 32'b00000000000000010101010000010110;
assign LUT_3[17961] = 32'b00000000000000011011111011110011;
assign LUT_3[17962] = 32'b00000000000000010111010111111010;
assign LUT_3[17963] = 32'b00000000000000011110000011010111;
assign LUT_3[17964] = 32'b00000000000000010010011110001100;
assign LUT_3[17965] = 32'b00000000000000011001001001101001;
assign LUT_3[17966] = 32'b00000000000000010100100101110000;
assign LUT_3[17967] = 32'b00000000000000011011010001001101;
assign LUT_3[17968] = 32'b00000000000000010011001010010011;
assign LUT_3[17969] = 32'b00000000000000011001110101110000;
assign LUT_3[17970] = 32'b00000000000000010101010001110111;
assign LUT_3[17971] = 32'b00000000000000011011111101010100;
assign LUT_3[17972] = 32'b00000000000000010000011000001001;
assign LUT_3[17973] = 32'b00000000000000010111000011100110;
assign LUT_3[17974] = 32'b00000000000000010010011111101101;
assign LUT_3[17975] = 32'b00000000000000011001001011001010;
assign LUT_3[17976] = 32'b00000000000000011000100011011001;
assign LUT_3[17977] = 32'b00000000000000011111001110110110;
assign LUT_3[17978] = 32'b00000000000000011010101010111101;
assign LUT_3[17979] = 32'b00000000000000100001010110011010;
assign LUT_3[17980] = 32'b00000000000000010101110001001111;
assign LUT_3[17981] = 32'b00000000000000011100011100101100;
assign LUT_3[17982] = 32'b00000000000000010111111000110011;
assign LUT_3[17983] = 32'b00000000000000011110100100010000;
assign LUT_3[17984] = 32'b00000000000000001110100001011011;
assign LUT_3[17985] = 32'b00000000000000010101001100111000;
assign LUT_3[17986] = 32'b00000000000000010000101000111111;
assign LUT_3[17987] = 32'b00000000000000010111010100011100;
assign LUT_3[17988] = 32'b00000000000000001011101111010001;
assign LUT_3[17989] = 32'b00000000000000010010011010101110;
assign LUT_3[17990] = 32'b00000000000000001101110110110101;
assign LUT_3[17991] = 32'b00000000000000010100100010010010;
assign LUT_3[17992] = 32'b00000000000000010011111010100001;
assign LUT_3[17993] = 32'b00000000000000011010100101111110;
assign LUT_3[17994] = 32'b00000000000000010110000010000101;
assign LUT_3[17995] = 32'b00000000000000011100101101100010;
assign LUT_3[17996] = 32'b00000000000000010001001000010111;
assign LUT_3[17997] = 32'b00000000000000010111110011110100;
assign LUT_3[17998] = 32'b00000000000000010011001111111011;
assign LUT_3[17999] = 32'b00000000000000011001111011011000;
assign LUT_3[18000] = 32'b00000000000000010001110100011110;
assign LUT_3[18001] = 32'b00000000000000011000011111111011;
assign LUT_3[18002] = 32'b00000000000000010011111100000010;
assign LUT_3[18003] = 32'b00000000000000011010100111011111;
assign LUT_3[18004] = 32'b00000000000000001111000010010100;
assign LUT_3[18005] = 32'b00000000000000010101101101110001;
assign LUT_3[18006] = 32'b00000000000000010001001001111000;
assign LUT_3[18007] = 32'b00000000000000010111110101010101;
assign LUT_3[18008] = 32'b00000000000000010111001101100100;
assign LUT_3[18009] = 32'b00000000000000011101111001000001;
assign LUT_3[18010] = 32'b00000000000000011001010101001000;
assign LUT_3[18011] = 32'b00000000000000100000000000100101;
assign LUT_3[18012] = 32'b00000000000000010100011011011010;
assign LUT_3[18013] = 32'b00000000000000011011000110110111;
assign LUT_3[18014] = 32'b00000000000000010110100010111110;
assign LUT_3[18015] = 32'b00000000000000011101001110011011;
assign LUT_3[18016] = 32'b00000000000000001111101111111011;
assign LUT_3[18017] = 32'b00000000000000010110011011011000;
assign LUT_3[18018] = 32'b00000000000000010001110111011111;
assign LUT_3[18019] = 32'b00000000000000011000100010111100;
assign LUT_3[18020] = 32'b00000000000000001100111101110001;
assign LUT_3[18021] = 32'b00000000000000010011101001001110;
assign LUT_3[18022] = 32'b00000000000000001111000101010101;
assign LUT_3[18023] = 32'b00000000000000010101110000110010;
assign LUT_3[18024] = 32'b00000000000000010101001001000001;
assign LUT_3[18025] = 32'b00000000000000011011110100011110;
assign LUT_3[18026] = 32'b00000000000000010111010000100101;
assign LUT_3[18027] = 32'b00000000000000011101111100000010;
assign LUT_3[18028] = 32'b00000000000000010010010110110111;
assign LUT_3[18029] = 32'b00000000000000011001000010010100;
assign LUT_3[18030] = 32'b00000000000000010100011110011011;
assign LUT_3[18031] = 32'b00000000000000011011001001111000;
assign LUT_3[18032] = 32'b00000000000000010011000010111110;
assign LUT_3[18033] = 32'b00000000000000011001101110011011;
assign LUT_3[18034] = 32'b00000000000000010101001010100010;
assign LUT_3[18035] = 32'b00000000000000011011110101111111;
assign LUT_3[18036] = 32'b00000000000000010000010000110100;
assign LUT_3[18037] = 32'b00000000000000010110111100010001;
assign LUT_3[18038] = 32'b00000000000000010010011000011000;
assign LUT_3[18039] = 32'b00000000000000011001000011110101;
assign LUT_3[18040] = 32'b00000000000000011000011100000100;
assign LUT_3[18041] = 32'b00000000000000011111000111100001;
assign LUT_3[18042] = 32'b00000000000000011010100011101000;
assign LUT_3[18043] = 32'b00000000000000100001001111000101;
assign LUT_3[18044] = 32'b00000000000000010101101001111010;
assign LUT_3[18045] = 32'b00000000000000011100010101010111;
assign LUT_3[18046] = 32'b00000000000000010111110001011110;
assign LUT_3[18047] = 32'b00000000000000011110011100111011;
assign LUT_3[18048] = 32'b00000000000000010000110011101110;
assign LUT_3[18049] = 32'b00000000000000010111011111001011;
assign LUT_3[18050] = 32'b00000000000000010010111011010010;
assign LUT_3[18051] = 32'b00000000000000011001100110101111;
assign LUT_3[18052] = 32'b00000000000000001110000001100100;
assign LUT_3[18053] = 32'b00000000000000010100101101000001;
assign LUT_3[18054] = 32'b00000000000000010000001001001000;
assign LUT_3[18055] = 32'b00000000000000010110110100100101;
assign LUT_3[18056] = 32'b00000000000000010110001100110100;
assign LUT_3[18057] = 32'b00000000000000011100111000010001;
assign LUT_3[18058] = 32'b00000000000000011000010100011000;
assign LUT_3[18059] = 32'b00000000000000011110111111110101;
assign LUT_3[18060] = 32'b00000000000000010011011010101010;
assign LUT_3[18061] = 32'b00000000000000011010000110000111;
assign LUT_3[18062] = 32'b00000000000000010101100010001110;
assign LUT_3[18063] = 32'b00000000000000011100001101101011;
assign LUT_3[18064] = 32'b00000000000000010100000110110001;
assign LUT_3[18065] = 32'b00000000000000011010110010001110;
assign LUT_3[18066] = 32'b00000000000000010110001110010101;
assign LUT_3[18067] = 32'b00000000000000011100111001110010;
assign LUT_3[18068] = 32'b00000000000000010001010100100111;
assign LUT_3[18069] = 32'b00000000000000011000000000000100;
assign LUT_3[18070] = 32'b00000000000000010011011100001011;
assign LUT_3[18071] = 32'b00000000000000011010000111101000;
assign LUT_3[18072] = 32'b00000000000000011001011111110111;
assign LUT_3[18073] = 32'b00000000000000100000001011010100;
assign LUT_3[18074] = 32'b00000000000000011011100111011011;
assign LUT_3[18075] = 32'b00000000000000100010010010111000;
assign LUT_3[18076] = 32'b00000000000000010110101101101101;
assign LUT_3[18077] = 32'b00000000000000011101011001001010;
assign LUT_3[18078] = 32'b00000000000000011000110101010001;
assign LUT_3[18079] = 32'b00000000000000011111100000101110;
assign LUT_3[18080] = 32'b00000000000000010010000010001110;
assign LUT_3[18081] = 32'b00000000000000011000101101101011;
assign LUT_3[18082] = 32'b00000000000000010100001001110010;
assign LUT_3[18083] = 32'b00000000000000011010110101001111;
assign LUT_3[18084] = 32'b00000000000000001111010000000100;
assign LUT_3[18085] = 32'b00000000000000010101111011100001;
assign LUT_3[18086] = 32'b00000000000000010001010111101000;
assign LUT_3[18087] = 32'b00000000000000011000000011000101;
assign LUT_3[18088] = 32'b00000000000000010111011011010100;
assign LUT_3[18089] = 32'b00000000000000011110000110110001;
assign LUT_3[18090] = 32'b00000000000000011001100010111000;
assign LUT_3[18091] = 32'b00000000000000100000001110010101;
assign LUT_3[18092] = 32'b00000000000000010100101001001010;
assign LUT_3[18093] = 32'b00000000000000011011010100100111;
assign LUT_3[18094] = 32'b00000000000000010110110000101110;
assign LUT_3[18095] = 32'b00000000000000011101011100001011;
assign LUT_3[18096] = 32'b00000000000000010101010101010001;
assign LUT_3[18097] = 32'b00000000000000011100000000101110;
assign LUT_3[18098] = 32'b00000000000000010111011100110101;
assign LUT_3[18099] = 32'b00000000000000011110001000010010;
assign LUT_3[18100] = 32'b00000000000000010010100011000111;
assign LUT_3[18101] = 32'b00000000000000011001001110100100;
assign LUT_3[18102] = 32'b00000000000000010100101010101011;
assign LUT_3[18103] = 32'b00000000000000011011010110001000;
assign LUT_3[18104] = 32'b00000000000000011010101110010111;
assign LUT_3[18105] = 32'b00000000000000100001011001110100;
assign LUT_3[18106] = 32'b00000000000000011100110101111011;
assign LUT_3[18107] = 32'b00000000000000100011100001011000;
assign LUT_3[18108] = 32'b00000000000000010111111100001101;
assign LUT_3[18109] = 32'b00000000000000011110100111101010;
assign LUT_3[18110] = 32'b00000000000000011010000011110001;
assign LUT_3[18111] = 32'b00000000000000100000101111001110;
assign LUT_3[18112] = 32'b00000000000000010000101100011001;
assign LUT_3[18113] = 32'b00000000000000010111010111110110;
assign LUT_3[18114] = 32'b00000000000000010010110011111101;
assign LUT_3[18115] = 32'b00000000000000011001011111011010;
assign LUT_3[18116] = 32'b00000000000000001101111010001111;
assign LUT_3[18117] = 32'b00000000000000010100100101101100;
assign LUT_3[18118] = 32'b00000000000000010000000001110011;
assign LUT_3[18119] = 32'b00000000000000010110101101010000;
assign LUT_3[18120] = 32'b00000000000000010110000101011111;
assign LUT_3[18121] = 32'b00000000000000011100110000111100;
assign LUT_3[18122] = 32'b00000000000000011000001101000011;
assign LUT_3[18123] = 32'b00000000000000011110111000100000;
assign LUT_3[18124] = 32'b00000000000000010011010011010101;
assign LUT_3[18125] = 32'b00000000000000011001111110110010;
assign LUT_3[18126] = 32'b00000000000000010101011010111001;
assign LUT_3[18127] = 32'b00000000000000011100000110010110;
assign LUT_3[18128] = 32'b00000000000000010011111111011100;
assign LUT_3[18129] = 32'b00000000000000011010101010111001;
assign LUT_3[18130] = 32'b00000000000000010110000111000000;
assign LUT_3[18131] = 32'b00000000000000011100110010011101;
assign LUT_3[18132] = 32'b00000000000000010001001101010010;
assign LUT_3[18133] = 32'b00000000000000010111111000101111;
assign LUT_3[18134] = 32'b00000000000000010011010100110110;
assign LUT_3[18135] = 32'b00000000000000011010000000010011;
assign LUT_3[18136] = 32'b00000000000000011001011000100010;
assign LUT_3[18137] = 32'b00000000000000100000000011111111;
assign LUT_3[18138] = 32'b00000000000000011011100000000110;
assign LUT_3[18139] = 32'b00000000000000100010001011100011;
assign LUT_3[18140] = 32'b00000000000000010110100110011000;
assign LUT_3[18141] = 32'b00000000000000011101010001110101;
assign LUT_3[18142] = 32'b00000000000000011000101101111100;
assign LUT_3[18143] = 32'b00000000000000011111011001011001;
assign LUT_3[18144] = 32'b00000000000000010001111010111001;
assign LUT_3[18145] = 32'b00000000000000011000100110010110;
assign LUT_3[18146] = 32'b00000000000000010100000010011101;
assign LUT_3[18147] = 32'b00000000000000011010101101111010;
assign LUT_3[18148] = 32'b00000000000000001111001000101111;
assign LUT_3[18149] = 32'b00000000000000010101110100001100;
assign LUT_3[18150] = 32'b00000000000000010001010000010011;
assign LUT_3[18151] = 32'b00000000000000010111111011110000;
assign LUT_3[18152] = 32'b00000000000000010111010011111111;
assign LUT_3[18153] = 32'b00000000000000011101111111011100;
assign LUT_3[18154] = 32'b00000000000000011001011011100011;
assign LUT_3[18155] = 32'b00000000000000100000000111000000;
assign LUT_3[18156] = 32'b00000000000000010100100001110101;
assign LUT_3[18157] = 32'b00000000000000011011001101010010;
assign LUT_3[18158] = 32'b00000000000000010110101001011001;
assign LUT_3[18159] = 32'b00000000000000011101010100110110;
assign LUT_3[18160] = 32'b00000000000000010101001101111100;
assign LUT_3[18161] = 32'b00000000000000011011111001011001;
assign LUT_3[18162] = 32'b00000000000000010111010101100000;
assign LUT_3[18163] = 32'b00000000000000011110000000111101;
assign LUT_3[18164] = 32'b00000000000000010010011011110010;
assign LUT_3[18165] = 32'b00000000000000011001000111001111;
assign LUT_3[18166] = 32'b00000000000000010100100011010110;
assign LUT_3[18167] = 32'b00000000000000011011001110110011;
assign LUT_3[18168] = 32'b00000000000000011010100111000010;
assign LUT_3[18169] = 32'b00000000000000100001010010011111;
assign LUT_3[18170] = 32'b00000000000000011100101110100110;
assign LUT_3[18171] = 32'b00000000000000100011011010000011;
assign LUT_3[18172] = 32'b00000000000000010111110100111000;
assign LUT_3[18173] = 32'b00000000000000011110100000010101;
assign LUT_3[18174] = 32'b00000000000000011001111100011100;
assign LUT_3[18175] = 32'b00000000000000100000100111111001;
assign LUT_3[18176] = 32'b00000000000000001010111000010001;
assign LUT_3[18177] = 32'b00000000000000010001100011101110;
assign LUT_3[18178] = 32'b00000000000000001100111111110101;
assign LUT_3[18179] = 32'b00000000000000010011101011010010;
assign LUT_3[18180] = 32'b00000000000000001000000110000111;
assign LUT_3[18181] = 32'b00000000000000001110110001100100;
assign LUT_3[18182] = 32'b00000000000000001010001101101011;
assign LUT_3[18183] = 32'b00000000000000010000111001001000;
assign LUT_3[18184] = 32'b00000000000000010000010001010111;
assign LUT_3[18185] = 32'b00000000000000010110111100110100;
assign LUT_3[18186] = 32'b00000000000000010010011000111011;
assign LUT_3[18187] = 32'b00000000000000011001000100011000;
assign LUT_3[18188] = 32'b00000000000000001101011111001101;
assign LUT_3[18189] = 32'b00000000000000010100001010101010;
assign LUT_3[18190] = 32'b00000000000000001111100110110001;
assign LUT_3[18191] = 32'b00000000000000010110010010001110;
assign LUT_3[18192] = 32'b00000000000000001110001011010100;
assign LUT_3[18193] = 32'b00000000000000010100110110110001;
assign LUT_3[18194] = 32'b00000000000000010000010010111000;
assign LUT_3[18195] = 32'b00000000000000010110111110010101;
assign LUT_3[18196] = 32'b00000000000000001011011001001010;
assign LUT_3[18197] = 32'b00000000000000010010000100100111;
assign LUT_3[18198] = 32'b00000000000000001101100000101110;
assign LUT_3[18199] = 32'b00000000000000010100001100001011;
assign LUT_3[18200] = 32'b00000000000000010011100100011010;
assign LUT_3[18201] = 32'b00000000000000011010001111110111;
assign LUT_3[18202] = 32'b00000000000000010101101011111110;
assign LUT_3[18203] = 32'b00000000000000011100010111011011;
assign LUT_3[18204] = 32'b00000000000000010000110010010000;
assign LUT_3[18205] = 32'b00000000000000010111011101101101;
assign LUT_3[18206] = 32'b00000000000000010010111001110100;
assign LUT_3[18207] = 32'b00000000000000011001100101010001;
assign LUT_3[18208] = 32'b00000000000000001100000110110001;
assign LUT_3[18209] = 32'b00000000000000010010110010001110;
assign LUT_3[18210] = 32'b00000000000000001110001110010101;
assign LUT_3[18211] = 32'b00000000000000010100111001110010;
assign LUT_3[18212] = 32'b00000000000000001001010100100111;
assign LUT_3[18213] = 32'b00000000000000010000000000000100;
assign LUT_3[18214] = 32'b00000000000000001011011100001011;
assign LUT_3[18215] = 32'b00000000000000010010000111101000;
assign LUT_3[18216] = 32'b00000000000000010001011111110111;
assign LUT_3[18217] = 32'b00000000000000011000001011010100;
assign LUT_3[18218] = 32'b00000000000000010011100111011011;
assign LUT_3[18219] = 32'b00000000000000011010010010111000;
assign LUT_3[18220] = 32'b00000000000000001110101101101101;
assign LUT_3[18221] = 32'b00000000000000010101011001001010;
assign LUT_3[18222] = 32'b00000000000000010000110101010001;
assign LUT_3[18223] = 32'b00000000000000010111100000101110;
assign LUT_3[18224] = 32'b00000000000000001111011001110100;
assign LUT_3[18225] = 32'b00000000000000010110000101010001;
assign LUT_3[18226] = 32'b00000000000000010001100001011000;
assign LUT_3[18227] = 32'b00000000000000011000001100110101;
assign LUT_3[18228] = 32'b00000000000000001100100111101010;
assign LUT_3[18229] = 32'b00000000000000010011010011000111;
assign LUT_3[18230] = 32'b00000000000000001110101111001110;
assign LUT_3[18231] = 32'b00000000000000010101011010101011;
assign LUT_3[18232] = 32'b00000000000000010100110010111010;
assign LUT_3[18233] = 32'b00000000000000011011011110010111;
assign LUT_3[18234] = 32'b00000000000000010110111010011110;
assign LUT_3[18235] = 32'b00000000000000011101100101111011;
assign LUT_3[18236] = 32'b00000000000000010010000000110000;
assign LUT_3[18237] = 32'b00000000000000011000101100001101;
assign LUT_3[18238] = 32'b00000000000000010100001000010100;
assign LUT_3[18239] = 32'b00000000000000011010110011110001;
assign LUT_3[18240] = 32'b00000000000000001010110000111100;
assign LUT_3[18241] = 32'b00000000000000010001011100011001;
assign LUT_3[18242] = 32'b00000000000000001100111000100000;
assign LUT_3[18243] = 32'b00000000000000010011100011111101;
assign LUT_3[18244] = 32'b00000000000000000111111110110010;
assign LUT_3[18245] = 32'b00000000000000001110101010001111;
assign LUT_3[18246] = 32'b00000000000000001010000110010110;
assign LUT_3[18247] = 32'b00000000000000010000110001110011;
assign LUT_3[18248] = 32'b00000000000000010000001010000010;
assign LUT_3[18249] = 32'b00000000000000010110110101011111;
assign LUT_3[18250] = 32'b00000000000000010010010001100110;
assign LUT_3[18251] = 32'b00000000000000011000111101000011;
assign LUT_3[18252] = 32'b00000000000000001101010111111000;
assign LUT_3[18253] = 32'b00000000000000010100000011010101;
assign LUT_3[18254] = 32'b00000000000000001111011111011100;
assign LUT_3[18255] = 32'b00000000000000010110001010111001;
assign LUT_3[18256] = 32'b00000000000000001110000011111111;
assign LUT_3[18257] = 32'b00000000000000010100101111011100;
assign LUT_3[18258] = 32'b00000000000000010000001011100011;
assign LUT_3[18259] = 32'b00000000000000010110110111000000;
assign LUT_3[18260] = 32'b00000000000000001011010001110101;
assign LUT_3[18261] = 32'b00000000000000010001111101010010;
assign LUT_3[18262] = 32'b00000000000000001101011001011001;
assign LUT_3[18263] = 32'b00000000000000010100000100110110;
assign LUT_3[18264] = 32'b00000000000000010011011101000101;
assign LUT_3[18265] = 32'b00000000000000011010001000100010;
assign LUT_3[18266] = 32'b00000000000000010101100100101001;
assign LUT_3[18267] = 32'b00000000000000011100010000000110;
assign LUT_3[18268] = 32'b00000000000000010000101010111011;
assign LUT_3[18269] = 32'b00000000000000010111010110011000;
assign LUT_3[18270] = 32'b00000000000000010010110010011111;
assign LUT_3[18271] = 32'b00000000000000011001011101111100;
assign LUT_3[18272] = 32'b00000000000000001011111111011100;
assign LUT_3[18273] = 32'b00000000000000010010101010111001;
assign LUT_3[18274] = 32'b00000000000000001110000111000000;
assign LUT_3[18275] = 32'b00000000000000010100110010011101;
assign LUT_3[18276] = 32'b00000000000000001001001101010010;
assign LUT_3[18277] = 32'b00000000000000001111111000101111;
assign LUT_3[18278] = 32'b00000000000000001011010100110110;
assign LUT_3[18279] = 32'b00000000000000010010000000010011;
assign LUT_3[18280] = 32'b00000000000000010001011000100010;
assign LUT_3[18281] = 32'b00000000000000011000000011111111;
assign LUT_3[18282] = 32'b00000000000000010011100000000110;
assign LUT_3[18283] = 32'b00000000000000011010001011100011;
assign LUT_3[18284] = 32'b00000000000000001110100110011000;
assign LUT_3[18285] = 32'b00000000000000010101010001110101;
assign LUT_3[18286] = 32'b00000000000000010000101101111100;
assign LUT_3[18287] = 32'b00000000000000010111011001011001;
assign LUT_3[18288] = 32'b00000000000000001111010010011111;
assign LUT_3[18289] = 32'b00000000000000010101111101111100;
assign LUT_3[18290] = 32'b00000000000000010001011010000011;
assign LUT_3[18291] = 32'b00000000000000011000000101100000;
assign LUT_3[18292] = 32'b00000000000000001100100000010101;
assign LUT_3[18293] = 32'b00000000000000010011001011110010;
assign LUT_3[18294] = 32'b00000000000000001110100111111001;
assign LUT_3[18295] = 32'b00000000000000010101010011010110;
assign LUT_3[18296] = 32'b00000000000000010100101011100101;
assign LUT_3[18297] = 32'b00000000000000011011010111000010;
assign LUT_3[18298] = 32'b00000000000000010110110011001001;
assign LUT_3[18299] = 32'b00000000000000011101011110100110;
assign LUT_3[18300] = 32'b00000000000000010001111001011011;
assign LUT_3[18301] = 32'b00000000000000011000100100111000;
assign LUT_3[18302] = 32'b00000000000000010100000000111111;
assign LUT_3[18303] = 32'b00000000000000011010101100011100;
assign LUT_3[18304] = 32'b00000000000000001101000011001111;
assign LUT_3[18305] = 32'b00000000000000010011101110101100;
assign LUT_3[18306] = 32'b00000000000000001111001010110011;
assign LUT_3[18307] = 32'b00000000000000010101110110010000;
assign LUT_3[18308] = 32'b00000000000000001010010001000101;
assign LUT_3[18309] = 32'b00000000000000010000111100100010;
assign LUT_3[18310] = 32'b00000000000000001100011000101001;
assign LUT_3[18311] = 32'b00000000000000010011000100000110;
assign LUT_3[18312] = 32'b00000000000000010010011100010101;
assign LUT_3[18313] = 32'b00000000000000011001000111110010;
assign LUT_3[18314] = 32'b00000000000000010100100011111001;
assign LUT_3[18315] = 32'b00000000000000011011001111010110;
assign LUT_3[18316] = 32'b00000000000000001111101010001011;
assign LUT_3[18317] = 32'b00000000000000010110010101101000;
assign LUT_3[18318] = 32'b00000000000000010001110001101111;
assign LUT_3[18319] = 32'b00000000000000011000011101001100;
assign LUT_3[18320] = 32'b00000000000000010000010110010010;
assign LUT_3[18321] = 32'b00000000000000010111000001101111;
assign LUT_3[18322] = 32'b00000000000000010010011101110110;
assign LUT_3[18323] = 32'b00000000000000011001001001010011;
assign LUT_3[18324] = 32'b00000000000000001101100100001000;
assign LUT_3[18325] = 32'b00000000000000010100001111100101;
assign LUT_3[18326] = 32'b00000000000000001111101011101100;
assign LUT_3[18327] = 32'b00000000000000010110010111001001;
assign LUT_3[18328] = 32'b00000000000000010101101111011000;
assign LUT_3[18329] = 32'b00000000000000011100011010110101;
assign LUT_3[18330] = 32'b00000000000000010111110110111100;
assign LUT_3[18331] = 32'b00000000000000011110100010011001;
assign LUT_3[18332] = 32'b00000000000000010010111101001110;
assign LUT_3[18333] = 32'b00000000000000011001101000101011;
assign LUT_3[18334] = 32'b00000000000000010101000100110010;
assign LUT_3[18335] = 32'b00000000000000011011110000001111;
assign LUT_3[18336] = 32'b00000000000000001110010001101111;
assign LUT_3[18337] = 32'b00000000000000010100111101001100;
assign LUT_3[18338] = 32'b00000000000000010000011001010011;
assign LUT_3[18339] = 32'b00000000000000010111000100110000;
assign LUT_3[18340] = 32'b00000000000000001011011111100101;
assign LUT_3[18341] = 32'b00000000000000010010001011000010;
assign LUT_3[18342] = 32'b00000000000000001101100111001001;
assign LUT_3[18343] = 32'b00000000000000010100010010100110;
assign LUT_3[18344] = 32'b00000000000000010011101010110101;
assign LUT_3[18345] = 32'b00000000000000011010010110010010;
assign LUT_3[18346] = 32'b00000000000000010101110010011001;
assign LUT_3[18347] = 32'b00000000000000011100011101110110;
assign LUT_3[18348] = 32'b00000000000000010000111000101011;
assign LUT_3[18349] = 32'b00000000000000010111100100001000;
assign LUT_3[18350] = 32'b00000000000000010011000000001111;
assign LUT_3[18351] = 32'b00000000000000011001101011101100;
assign LUT_3[18352] = 32'b00000000000000010001100100110010;
assign LUT_3[18353] = 32'b00000000000000011000010000001111;
assign LUT_3[18354] = 32'b00000000000000010011101100010110;
assign LUT_3[18355] = 32'b00000000000000011010010111110011;
assign LUT_3[18356] = 32'b00000000000000001110110010101000;
assign LUT_3[18357] = 32'b00000000000000010101011110000101;
assign LUT_3[18358] = 32'b00000000000000010000111010001100;
assign LUT_3[18359] = 32'b00000000000000010111100101101001;
assign LUT_3[18360] = 32'b00000000000000010110111101111000;
assign LUT_3[18361] = 32'b00000000000000011101101001010101;
assign LUT_3[18362] = 32'b00000000000000011001000101011100;
assign LUT_3[18363] = 32'b00000000000000011111110000111001;
assign LUT_3[18364] = 32'b00000000000000010100001011101110;
assign LUT_3[18365] = 32'b00000000000000011010110111001011;
assign LUT_3[18366] = 32'b00000000000000010110010011010010;
assign LUT_3[18367] = 32'b00000000000000011100111110101111;
assign LUT_3[18368] = 32'b00000000000000001100111011111010;
assign LUT_3[18369] = 32'b00000000000000010011100111010111;
assign LUT_3[18370] = 32'b00000000000000001111000011011110;
assign LUT_3[18371] = 32'b00000000000000010101101110111011;
assign LUT_3[18372] = 32'b00000000000000001010001001110000;
assign LUT_3[18373] = 32'b00000000000000010000110101001101;
assign LUT_3[18374] = 32'b00000000000000001100010001010100;
assign LUT_3[18375] = 32'b00000000000000010010111100110001;
assign LUT_3[18376] = 32'b00000000000000010010010101000000;
assign LUT_3[18377] = 32'b00000000000000011001000000011101;
assign LUT_3[18378] = 32'b00000000000000010100011100100100;
assign LUT_3[18379] = 32'b00000000000000011011001000000001;
assign LUT_3[18380] = 32'b00000000000000001111100010110110;
assign LUT_3[18381] = 32'b00000000000000010110001110010011;
assign LUT_3[18382] = 32'b00000000000000010001101010011010;
assign LUT_3[18383] = 32'b00000000000000011000010101110111;
assign LUT_3[18384] = 32'b00000000000000010000001110111101;
assign LUT_3[18385] = 32'b00000000000000010110111010011010;
assign LUT_3[18386] = 32'b00000000000000010010010110100001;
assign LUT_3[18387] = 32'b00000000000000011001000001111110;
assign LUT_3[18388] = 32'b00000000000000001101011100110011;
assign LUT_3[18389] = 32'b00000000000000010100001000010000;
assign LUT_3[18390] = 32'b00000000000000001111100100010111;
assign LUT_3[18391] = 32'b00000000000000010110001111110100;
assign LUT_3[18392] = 32'b00000000000000010101101000000011;
assign LUT_3[18393] = 32'b00000000000000011100010011100000;
assign LUT_3[18394] = 32'b00000000000000010111101111100111;
assign LUT_3[18395] = 32'b00000000000000011110011011000100;
assign LUT_3[18396] = 32'b00000000000000010010110101111001;
assign LUT_3[18397] = 32'b00000000000000011001100001010110;
assign LUT_3[18398] = 32'b00000000000000010100111101011101;
assign LUT_3[18399] = 32'b00000000000000011011101000111010;
assign LUT_3[18400] = 32'b00000000000000001110001010011010;
assign LUT_3[18401] = 32'b00000000000000010100110101110111;
assign LUT_3[18402] = 32'b00000000000000010000010001111110;
assign LUT_3[18403] = 32'b00000000000000010110111101011011;
assign LUT_3[18404] = 32'b00000000000000001011011000010000;
assign LUT_3[18405] = 32'b00000000000000010010000011101101;
assign LUT_3[18406] = 32'b00000000000000001101011111110100;
assign LUT_3[18407] = 32'b00000000000000010100001011010001;
assign LUT_3[18408] = 32'b00000000000000010011100011100000;
assign LUT_3[18409] = 32'b00000000000000011010001110111101;
assign LUT_3[18410] = 32'b00000000000000010101101011000100;
assign LUT_3[18411] = 32'b00000000000000011100010110100001;
assign LUT_3[18412] = 32'b00000000000000010000110001010110;
assign LUT_3[18413] = 32'b00000000000000010111011100110011;
assign LUT_3[18414] = 32'b00000000000000010010111000111010;
assign LUT_3[18415] = 32'b00000000000000011001100100010111;
assign LUT_3[18416] = 32'b00000000000000010001011101011101;
assign LUT_3[18417] = 32'b00000000000000011000001000111010;
assign LUT_3[18418] = 32'b00000000000000010011100101000001;
assign LUT_3[18419] = 32'b00000000000000011010010000011110;
assign LUT_3[18420] = 32'b00000000000000001110101011010011;
assign LUT_3[18421] = 32'b00000000000000010101010110110000;
assign LUT_3[18422] = 32'b00000000000000010000110010110111;
assign LUT_3[18423] = 32'b00000000000000010111011110010100;
assign LUT_3[18424] = 32'b00000000000000010110110110100011;
assign LUT_3[18425] = 32'b00000000000000011101100010000000;
assign LUT_3[18426] = 32'b00000000000000011000111110000111;
assign LUT_3[18427] = 32'b00000000000000011111101001100100;
assign LUT_3[18428] = 32'b00000000000000010100000100011001;
assign LUT_3[18429] = 32'b00000000000000011010101111110110;
assign LUT_3[18430] = 32'b00000000000000010110001011111101;
assign LUT_3[18431] = 32'b00000000000000011100110111011010;
assign LUT_3[18432] = 32'b00000000000000000110100100110101;
assign LUT_3[18433] = 32'b00000000000000001101010000010010;
assign LUT_3[18434] = 32'b00000000000000001000101100011001;
assign LUT_3[18435] = 32'b00000000000000001111010111110110;
assign LUT_3[18436] = 32'b00000000000000000011110010101011;
assign LUT_3[18437] = 32'b00000000000000001010011110001000;
assign LUT_3[18438] = 32'b00000000000000000101111010001111;
assign LUT_3[18439] = 32'b00000000000000001100100101101100;
assign LUT_3[18440] = 32'b00000000000000001011111101111011;
assign LUT_3[18441] = 32'b00000000000000010010101001011000;
assign LUT_3[18442] = 32'b00000000000000001110000101011111;
assign LUT_3[18443] = 32'b00000000000000010100110000111100;
assign LUT_3[18444] = 32'b00000000000000001001001011110001;
assign LUT_3[18445] = 32'b00000000000000001111110111001110;
assign LUT_3[18446] = 32'b00000000000000001011010011010101;
assign LUT_3[18447] = 32'b00000000000000010001111110110010;
assign LUT_3[18448] = 32'b00000000000000001001110111111000;
assign LUT_3[18449] = 32'b00000000000000010000100011010101;
assign LUT_3[18450] = 32'b00000000000000001011111111011100;
assign LUT_3[18451] = 32'b00000000000000010010101010111001;
assign LUT_3[18452] = 32'b00000000000000000111000101101110;
assign LUT_3[18453] = 32'b00000000000000001101110001001011;
assign LUT_3[18454] = 32'b00000000000000001001001101010010;
assign LUT_3[18455] = 32'b00000000000000001111111000101111;
assign LUT_3[18456] = 32'b00000000000000001111010000111110;
assign LUT_3[18457] = 32'b00000000000000010101111100011011;
assign LUT_3[18458] = 32'b00000000000000010001011000100010;
assign LUT_3[18459] = 32'b00000000000000011000000011111111;
assign LUT_3[18460] = 32'b00000000000000001100011110110100;
assign LUT_3[18461] = 32'b00000000000000010011001010010001;
assign LUT_3[18462] = 32'b00000000000000001110100110011000;
assign LUT_3[18463] = 32'b00000000000000010101010001110101;
assign LUT_3[18464] = 32'b00000000000000000111110011010101;
assign LUT_3[18465] = 32'b00000000000000001110011110110010;
assign LUT_3[18466] = 32'b00000000000000001001111010111001;
assign LUT_3[18467] = 32'b00000000000000010000100110010110;
assign LUT_3[18468] = 32'b00000000000000000101000001001011;
assign LUT_3[18469] = 32'b00000000000000001011101100101000;
assign LUT_3[18470] = 32'b00000000000000000111001000101111;
assign LUT_3[18471] = 32'b00000000000000001101110100001100;
assign LUT_3[18472] = 32'b00000000000000001101001100011011;
assign LUT_3[18473] = 32'b00000000000000010011110111111000;
assign LUT_3[18474] = 32'b00000000000000001111010011111111;
assign LUT_3[18475] = 32'b00000000000000010101111111011100;
assign LUT_3[18476] = 32'b00000000000000001010011010010001;
assign LUT_3[18477] = 32'b00000000000000010001000101101110;
assign LUT_3[18478] = 32'b00000000000000001100100001110101;
assign LUT_3[18479] = 32'b00000000000000010011001101010010;
assign LUT_3[18480] = 32'b00000000000000001011000110011000;
assign LUT_3[18481] = 32'b00000000000000010001110001110101;
assign LUT_3[18482] = 32'b00000000000000001101001101111100;
assign LUT_3[18483] = 32'b00000000000000010011111001011001;
assign LUT_3[18484] = 32'b00000000000000001000010100001110;
assign LUT_3[18485] = 32'b00000000000000001110111111101011;
assign LUT_3[18486] = 32'b00000000000000001010011011110010;
assign LUT_3[18487] = 32'b00000000000000010001000111001111;
assign LUT_3[18488] = 32'b00000000000000010000011111011110;
assign LUT_3[18489] = 32'b00000000000000010111001010111011;
assign LUT_3[18490] = 32'b00000000000000010010100111000010;
assign LUT_3[18491] = 32'b00000000000000011001010010011111;
assign LUT_3[18492] = 32'b00000000000000001101101101010100;
assign LUT_3[18493] = 32'b00000000000000010100011000110001;
assign LUT_3[18494] = 32'b00000000000000001111110100111000;
assign LUT_3[18495] = 32'b00000000000000010110100000010101;
assign LUT_3[18496] = 32'b00000000000000000110011101100000;
assign LUT_3[18497] = 32'b00000000000000001101001000111101;
assign LUT_3[18498] = 32'b00000000000000001000100101000100;
assign LUT_3[18499] = 32'b00000000000000001111010000100001;
assign LUT_3[18500] = 32'b00000000000000000011101011010110;
assign LUT_3[18501] = 32'b00000000000000001010010110110011;
assign LUT_3[18502] = 32'b00000000000000000101110010111010;
assign LUT_3[18503] = 32'b00000000000000001100011110010111;
assign LUT_3[18504] = 32'b00000000000000001011110110100110;
assign LUT_3[18505] = 32'b00000000000000010010100010000011;
assign LUT_3[18506] = 32'b00000000000000001101111110001010;
assign LUT_3[18507] = 32'b00000000000000010100101001100111;
assign LUT_3[18508] = 32'b00000000000000001001000100011100;
assign LUT_3[18509] = 32'b00000000000000001111101111111001;
assign LUT_3[18510] = 32'b00000000000000001011001100000000;
assign LUT_3[18511] = 32'b00000000000000010001110111011101;
assign LUT_3[18512] = 32'b00000000000000001001110000100011;
assign LUT_3[18513] = 32'b00000000000000010000011100000000;
assign LUT_3[18514] = 32'b00000000000000001011111000000111;
assign LUT_3[18515] = 32'b00000000000000010010100011100100;
assign LUT_3[18516] = 32'b00000000000000000110111110011001;
assign LUT_3[18517] = 32'b00000000000000001101101001110110;
assign LUT_3[18518] = 32'b00000000000000001001000101111101;
assign LUT_3[18519] = 32'b00000000000000001111110001011010;
assign LUT_3[18520] = 32'b00000000000000001111001001101001;
assign LUT_3[18521] = 32'b00000000000000010101110101000110;
assign LUT_3[18522] = 32'b00000000000000010001010001001101;
assign LUT_3[18523] = 32'b00000000000000010111111100101010;
assign LUT_3[18524] = 32'b00000000000000001100010111011111;
assign LUT_3[18525] = 32'b00000000000000010011000010111100;
assign LUT_3[18526] = 32'b00000000000000001110011111000011;
assign LUT_3[18527] = 32'b00000000000000010101001010100000;
assign LUT_3[18528] = 32'b00000000000000000111101100000000;
assign LUT_3[18529] = 32'b00000000000000001110010111011101;
assign LUT_3[18530] = 32'b00000000000000001001110011100100;
assign LUT_3[18531] = 32'b00000000000000010000011111000001;
assign LUT_3[18532] = 32'b00000000000000000100111001110110;
assign LUT_3[18533] = 32'b00000000000000001011100101010011;
assign LUT_3[18534] = 32'b00000000000000000111000001011010;
assign LUT_3[18535] = 32'b00000000000000001101101100110111;
assign LUT_3[18536] = 32'b00000000000000001101000101000110;
assign LUT_3[18537] = 32'b00000000000000010011110000100011;
assign LUT_3[18538] = 32'b00000000000000001111001100101010;
assign LUT_3[18539] = 32'b00000000000000010101111000000111;
assign LUT_3[18540] = 32'b00000000000000001010010010111100;
assign LUT_3[18541] = 32'b00000000000000010000111110011001;
assign LUT_3[18542] = 32'b00000000000000001100011010100000;
assign LUT_3[18543] = 32'b00000000000000010011000101111101;
assign LUT_3[18544] = 32'b00000000000000001010111111000011;
assign LUT_3[18545] = 32'b00000000000000010001101010100000;
assign LUT_3[18546] = 32'b00000000000000001101000110100111;
assign LUT_3[18547] = 32'b00000000000000010011110010000100;
assign LUT_3[18548] = 32'b00000000000000001000001100111001;
assign LUT_3[18549] = 32'b00000000000000001110111000010110;
assign LUT_3[18550] = 32'b00000000000000001010010100011101;
assign LUT_3[18551] = 32'b00000000000000010000111111111010;
assign LUT_3[18552] = 32'b00000000000000010000011000001001;
assign LUT_3[18553] = 32'b00000000000000010111000011100110;
assign LUT_3[18554] = 32'b00000000000000010010011111101101;
assign LUT_3[18555] = 32'b00000000000000011001001011001010;
assign LUT_3[18556] = 32'b00000000000000001101100101111111;
assign LUT_3[18557] = 32'b00000000000000010100010001011100;
assign LUT_3[18558] = 32'b00000000000000001111101101100011;
assign LUT_3[18559] = 32'b00000000000000010110011001000000;
assign LUT_3[18560] = 32'b00000000000000001000101111110011;
assign LUT_3[18561] = 32'b00000000000000001111011011010000;
assign LUT_3[18562] = 32'b00000000000000001010110111010111;
assign LUT_3[18563] = 32'b00000000000000010001100010110100;
assign LUT_3[18564] = 32'b00000000000000000101111101101001;
assign LUT_3[18565] = 32'b00000000000000001100101001000110;
assign LUT_3[18566] = 32'b00000000000000001000000101001101;
assign LUT_3[18567] = 32'b00000000000000001110110000101010;
assign LUT_3[18568] = 32'b00000000000000001110001000111001;
assign LUT_3[18569] = 32'b00000000000000010100110100010110;
assign LUT_3[18570] = 32'b00000000000000010000010000011101;
assign LUT_3[18571] = 32'b00000000000000010110111011111010;
assign LUT_3[18572] = 32'b00000000000000001011010110101111;
assign LUT_3[18573] = 32'b00000000000000010010000010001100;
assign LUT_3[18574] = 32'b00000000000000001101011110010011;
assign LUT_3[18575] = 32'b00000000000000010100001001110000;
assign LUT_3[18576] = 32'b00000000000000001100000010110110;
assign LUT_3[18577] = 32'b00000000000000010010101110010011;
assign LUT_3[18578] = 32'b00000000000000001110001010011010;
assign LUT_3[18579] = 32'b00000000000000010100110101110111;
assign LUT_3[18580] = 32'b00000000000000001001010000101100;
assign LUT_3[18581] = 32'b00000000000000001111111100001001;
assign LUT_3[18582] = 32'b00000000000000001011011000010000;
assign LUT_3[18583] = 32'b00000000000000010010000011101101;
assign LUT_3[18584] = 32'b00000000000000010001011011111100;
assign LUT_3[18585] = 32'b00000000000000011000000111011001;
assign LUT_3[18586] = 32'b00000000000000010011100011100000;
assign LUT_3[18587] = 32'b00000000000000011010001110111101;
assign LUT_3[18588] = 32'b00000000000000001110101001110010;
assign LUT_3[18589] = 32'b00000000000000010101010101001111;
assign LUT_3[18590] = 32'b00000000000000010000110001010110;
assign LUT_3[18591] = 32'b00000000000000010111011100110011;
assign LUT_3[18592] = 32'b00000000000000001001111110010011;
assign LUT_3[18593] = 32'b00000000000000010000101001110000;
assign LUT_3[18594] = 32'b00000000000000001100000101110111;
assign LUT_3[18595] = 32'b00000000000000010010110001010100;
assign LUT_3[18596] = 32'b00000000000000000111001100001001;
assign LUT_3[18597] = 32'b00000000000000001101110111100110;
assign LUT_3[18598] = 32'b00000000000000001001010011101101;
assign LUT_3[18599] = 32'b00000000000000001111111111001010;
assign LUT_3[18600] = 32'b00000000000000001111010111011001;
assign LUT_3[18601] = 32'b00000000000000010110000010110110;
assign LUT_3[18602] = 32'b00000000000000010001011110111101;
assign LUT_3[18603] = 32'b00000000000000011000001010011010;
assign LUT_3[18604] = 32'b00000000000000001100100101001111;
assign LUT_3[18605] = 32'b00000000000000010011010000101100;
assign LUT_3[18606] = 32'b00000000000000001110101100110011;
assign LUT_3[18607] = 32'b00000000000000010101011000010000;
assign LUT_3[18608] = 32'b00000000000000001101010001010110;
assign LUT_3[18609] = 32'b00000000000000010011111100110011;
assign LUT_3[18610] = 32'b00000000000000001111011000111010;
assign LUT_3[18611] = 32'b00000000000000010110000100010111;
assign LUT_3[18612] = 32'b00000000000000001010011111001100;
assign LUT_3[18613] = 32'b00000000000000010001001010101001;
assign LUT_3[18614] = 32'b00000000000000001100100110110000;
assign LUT_3[18615] = 32'b00000000000000010011010010001101;
assign LUT_3[18616] = 32'b00000000000000010010101010011100;
assign LUT_3[18617] = 32'b00000000000000011001010101111001;
assign LUT_3[18618] = 32'b00000000000000010100110010000000;
assign LUT_3[18619] = 32'b00000000000000011011011101011101;
assign LUT_3[18620] = 32'b00000000000000001111111000010010;
assign LUT_3[18621] = 32'b00000000000000010110100011101111;
assign LUT_3[18622] = 32'b00000000000000010001111111110110;
assign LUT_3[18623] = 32'b00000000000000011000101011010011;
assign LUT_3[18624] = 32'b00000000000000001000101000011110;
assign LUT_3[18625] = 32'b00000000000000001111010011111011;
assign LUT_3[18626] = 32'b00000000000000001010110000000010;
assign LUT_3[18627] = 32'b00000000000000010001011011011111;
assign LUT_3[18628] = 32'b00000000000000000101110110010100;
assign LUT_3[18629] = 32'b00000000000000001100100001110001;
assign LUT_3[18630] = 32'b00000000000000000111111101111000;
assign LUT_3[18631] = 32'b00000000000000001110101001010101;
assign LUT_3[18632] = 32'b00000000000000001110000001100100;
assign LUT_3[18633] = 32'b00000000000000010100101101000001;
assign LUT_3[18634] = 32'b00000000000000010000001001001000;
assign LUT_3[18635] = 32'b00000000000000010110110100100101;
assign LUT_3[18636] = 32'b00000000000000001011001111011010;
assign LUT_3[18637] = 32'b00000000000000010001111010110111;
assign LUT_3[18638] = 32'b00000000000000001101010110111110;
assign LUT_3[18639] = 32'b00000000000000010100000010011011;
assign LUT_3[18640] = 32'b00000000000000001011111011100001;
assign LUT_3[18641] = 32'b00000000000000010010100110111110;
assign LUT_3[18642] = 32'b00000000000000001110000011000101;
assign LUT_3[18643] = 32'b00000000000000010100101110100010;
assign LUT_3[18644] = 32'b00000000000000001001001001010111;
assign LUT_3[18645] = 32'b00000000000000001111110100110100;
assign LUT_3[18646] = 32'b00000000000000001011010000111011;
assign LUT_3[18647] = 32'b00000000000000010001111100011000;
assign LUT_3[18648] = 32'b00000000000000010001010100100111;
assign LUT_3[18649] = 32'b00000000000000011000000000000100;
assign LUT_3[18650] = 32'b00000000000000010011011100001011;
assign LUT_3[18651] = 32'b00000000000000011010000111101000;
assign LUT_3[18652] = 32'b00000000000000001110100010011101;
assign LUT_3[18653] = 32'b00000000000000010101001101111010;
assign LUT_3[18654] = 32'b00000000000000010000101010000001;
assign LUT_3[18655] = 32'b00000000000000010111010101011110;
assign LUT_3[18656] = 32'b00000000000000001001110110111110;
assign LUT_3[18657] = 32'b00000000000000010000100010011011;
assign LUT_3[18658] = 32'b00000000000000001011111110100010;
assign LUT_3[18659] = 32'b00000000000000010010101001111111;
assign LUT_3[18660] = 32'b00000000000000000111000100110100;
assign LUT_3[18661] = 32'b00000000000000001101110000010001;
assign LUT_3[18662] = 32'b00000000000000001001001100011000;
assign LUT_3[18663] = 32'b00000000000000001111110111110101;
assign LUT_3[18664] = 32'b00000000000000001111010000000100;
assign LUT_3[18665] = 32'b00000000000000010101111011100001;
assign LUT_3[18666] = 32'b00000000000000010001010111101000;
assign LUT_3[18667] = 32'b00000000000000011000000011000101;
assign LUT_3[18668] = 32'b00000000000000001100011101111010;
assign LUT_3[18669] = 32'b00000000000000010011001001010111;
assign LUT_3[18670] = 32'b00000000000000001110100101011110;
assign LUT_3[18671] = 32'b00000000000000010101010000111011;
assign LUT_3[18672] = 32'b00000000000000001101001010000001;
assign LUT_3[18673] = 32'b00000000000000010011110101011110;
assign LUT_3[18674] = 32'b00000000000000001111010001100101;
assign LUT_3[18675] = 32'b00000000000000010101111101000010;
assign LUT_3[18676] = 32'b00000000000000001010010111110111;
assign LUT_3[18677] = 32'b00000000000000010001000011010100;
assign LUT_3[18678] = 32'b00000000000000001100011111011011;
assign LUT_3[18679] = 32'b00000000000000010011001010111000;
assign LUT_3[18680] = 32'b00000000000000010010100011000111;
assign LUT_3[18681] = 32'b00000000000000011001001110100100;
assign LUT_3[18682] = 32'b00000000000000010100101010101011;
assign LUT_3[18683] = 32'b00000000000000011011010110001000;
assign LUT_3[18684] = 32'b00000000000000001111110000111101;
assign LUT_3[18685] = 32'b00000000000000010110011100011010;
assign LUT_3[18686] = 32'b00000000000000010001111000100001;
assign LUT_3[18687] = 32'b00000000000000011000100011111110;
assign LUT_3[18688] = 32'b00000000000000000010110100010110;
assign LUT_3[18689] = 32'b00000000000000001001011111110011;
assign LUT_3[18690] = 32'b00000000000000000100111011111010;
assign LUT_3[18691] = 32'b00000000000000001011100111010111;
assign LUT_3[18692] = 32'b00000000000000000000000010001100;
assign LUT_3[18693] = 32'b00000000000000000110101101101001;
assign LUT_3[18694] = 32'b00000000000000000010001001110000;
assign LUT_3[18695] = 32'b00000000000000001000110101001101;
assign LUT_3[18696] = 32'b00000000000000001000001101011100;
assign LUT_3[18697] = 32'b00000000000000001110111000111001;
assign LUT_3[18698] = 32'b00000000000000001010010101000000;
assign LUT_3[18699] = 32'b00000000000000010001000000011101;
assign LUT_3[18700] = 32'b00000000000000000101011011010010;
assign LUT_3[18701] = 32'b00000000000000001100000110101111;
assign LUT_3[18702] = 32'b00000000000000000111100010110110;
assign LUT_3[18703] = 32'b00000000000000001110001110010011;
assign LUT_3[18704] = 32'b00000000000000000110000111011001;
assign LUT_3[18705] = 32'b00000000000000001100110010110110;
assign LUT_3[18706] = 32'b00000000000000001000001110111101;
assign LUT_3[18707] = 32'b00000000000000001110111010011010;
assign LUT_3[18708] = 32'b00000000000000000011010101001111;
assign LUT_3[18709] = 32'b00000000000000001010000000101100;
assign LUT_3[18710] = 32'b00000000000000000101011100110011;
assign LUT_3[18711] = 32'b00000000000000001100001000010000;
assign LUT_3[18712] = 32'b00000000000000001011100000011111;
assign LUT_3[18713] = 32'b00000000000000010010001011111100;
assign LUT_3[18714] = 32'b00000000000000001101101000000011;
assign LUT_3[18715] = 32'b00000000000000010100010011100000;
assign LUT_3[18716] = 32'b00000000000000001000101110010101;
assign LUT_3[18717] = 32'b00000000000000001111011001110010;
assign LUT_3[18718] = 32'b00000000000000001010110101111001;
assign LUT_3[18719] = 32'b00000000000000010001100001010110;
assign LUT_3[18720] = 32'b00000000000000000100000010110110;
assign LUT_3[18721] = 32'b00000000000000001010101110010011;
assign LUT_3[18722] = 32'b00000000000000000110001010011010;
assign LUT_3[18723] = 32'b00000000000000001100110101110111;
assign LUT_3[18724] = 32'b00000000000000000001010000101100;
assign LUT_3[18725] = 32'b00000000000000000111111100001001;
assign LUT_3[18726] = 32'b00000000000000000011011000010000;
assign LUT_3[18727] = 32'b00000000000000001010000011101101;
assign LUT_3[18728] = 32'b00000000000000001001011011111100;
assign LUT_3[18729] = 32'b00000000000000010000000111011001;
assign LUT_3[18730] = 32'b00000000000000001011100011100000;
assign LUT_3[18731] = 32'b00000000000000010010001110111101;
assign LUT_3[18732] = 32'b00000000000000000110101001110010;
assign LUT_3[18733] = 32'b00000000000000001101010101001111;
assign LUT_3[18734] = 32'b00000000000000001000110001010110;
assign LUT_3[18735] = 32'b00000000000000001111011100110011;
assign LUT_3[18736] = 32'b00000000000000000111010101111001;
assign LUT_3[18737] = 32'b00000000000000001110000001010110;
assign LUT_3[18738] = 32'b00000000000000001001011101011101;
assign LUT_3[18739] = 32'b00000000000000010000001000111010;
assign LUT_3[18740] = 32'b00000000000000000100100011101111;
assign LUT_3[18741] = 32'b00000000000000001011001111001100;
assign LUT_3[18742] = 32'b00000000000000000110101011010011;
assign LUT_3[18743] = 32'b00000000000000001101010110110000;
assign LUT_3[18744] = 32'b00000000000000001100101110111111;
assign LUT_3[18745] = 32'b00000000000000010011011010011100;
assign LUT_3[18746] = 32'b00000000000000001110110110100011;
assign LUT_3[18747] = 32'b00000000000000010101100010000000;
assign LUT_3[18748] = 32'b00000000000000001001111100110101;
assign LUT_3[18749] = 32'b00000000000000010000101000010010;
assign LUT_3[18750] = 32'b00000000000000001100000100011001;
assign LUT_3[18751] = 32'b00000000000000010010101111110110;
assign LUT_3[18752] = 32'b00000000000000000010101101000001;
assign LUT_3[18753] = 32'b00000000000000001001011000011110;
assign LUT_3[18754] = 32'b00000000000000000100110100100101;
assign LUT_3[18755] = 32'b00000000000000001011100000000010;
assign LUT_3[18756] = 32'b11111111111111111111111010110111;
assign LUT_3[18757] = 32'b00000000000000000110100110010100;
assign LUT_3[18758] = 32'b00000000000000000010000010011011;
assign LUT_3[18759] = 32'b00000000000000001000101101111000;
assign LUT_3[18760] = 32'b00000000000000001000000110000111;
assign LUT_3[18761] = 32'b00000000000000001110110001100100;
assign LUT_3[18762] = 32'b00000000000000001010001101101011;
assign LUT_3[18763] = 32'b00000000000000010000111001001000;
assign LUT_3[18764] = 32'b00000000000000000101010011111101;
assign LUT_3[18765] = 32'b00000000000000001011111111011010;
assign LUT_3[18766] = 32'b00000000000000000111011011100001;
assign LUT_3[18767] = 32'b00000000000000001110000110111110;
assign LUT_3[18768] = 32'b00000000000000000110000000000100;
assign LUT_3[18769] = 32'b00000000000000001100101011100001;
assign LUT_3[18770] = 32'b00000000000000001000000111101000;
assign LUT_3[18771] = 32'b00000000000000001110110011000101;
assign LUT_3[18772] = 32'b00000000000000000011001101111010;
assign LUT_3[18773] = 32'b00000000000000001001111001010111;
assign LUT_3[18774] = 32'b00000000000000000101010101011110;
assign LUT_3[18775] = 32'b00000000000000001100000000111011;
assign LUT_3[18776] = 32'b00000000000000001011011001001010;
assign LUT_3[18777] = 32'b00000000000000010010000100100111;
assign LUT_3[18778] = 32'b00000000000000001101100000101110;
assign LUT_3[18779] = 32'b00000000000000010100001100001011;
assign LUT_3[18780] = 32'b00000000000000001000100111000000;
assign LUT_3[18781] = 32'b00000000000000001111010010011101;
assign LUT_3[18782] = 32'b00000000000000001010101110100100;
assign LUT_3[18783] = 32'b00000000000000010001011010000001;
assign LUT_3[18784] = 32'b00000000000000000011111011100001;
assign LUT_3[18785] = 32'b00000000000000001010100110111110;
assign LUT_3[18786] = 32'b00000000000000000110000011000101;
assign LUT_3[18787] = 32'b00000000000000001100101110100010;
assign LUT_3[18788] = 32'b00000000000000000001001001010111;
assign LUT_3[18789] = 32'b00000000000000000111110100110100;
assign LUT_3[18790] = 32'b00000000000000000011010000111011;
assign LUT_3[18791] = 32'b00000000000000001001111100011000;
assign LUT_3[18792] = 32'b00000000000000001001010100100111;
assign LUT_3[18793] = 32'b00000000000000010000000000000100;
assign LUT_3[18794] = 32'b00000000000000001011011100001011;
assign LUT_3[18795] = 32'b00000000000000010010000111101000;
assign LUT_3[18796] = 32'b00000000000000000110100010011101;
assign LUT_3[18797] = 32'b00000000000000001101001101111010;
assign LUT_3[18798] = 32'b00000000000000001000101010000001;
assign LUT_3[18799] = 32'b00000000000000001111010101011110;
assign LUT_3[18800] = 32'b00000000000000000111001110100100;
assign LUT_3[18801] = 32'b00000000000000001101111010000001;
assign LUT_3[18802] = 32'b00000000000000001001010110001000;
assign LUT_3[18803] = 32'b00000000000000010000000001100101;
assign LUT_3[18804] = 32'b00000000000000000100011100011010;
assign LUT_3[18805] = 32'b00000000000000001011000111110111;
assign LUT_3[18806] = 32'b00000000000000000110100011111110;
assign LUT_3[18807] = 32'b00000000000000001101001111011011;
assign LUT_3[18808] = 32'b00000000000000001100100111101010;
assign LUT_3[18809] = 32'b00000000000000010011010011000111;
assign LUT_3[18810] = 32'b00000000000000001110101111001110;
assign LUT_3[18811] = 32'b00000000000000010101011010101011;
assign LUT_3[18812] = 32'b00000000000000001001110101100000;
assign LUT_3[18813] = 32'b00000000000000010000100000111101;
assign LUT_3[18814] = 32'b00000000000000001011111101000100;
assign LUT_3[18815] = 32'b00000000000000010010101000100001;
assign LUT_3[18816] = 32'b00000000000000000100111111010100;
assign LUT_3[18817] = 32'b00000000000000001011101010110001;
assign LUT_3[18818] = 32'b00000000000000000111000110111000;
assign LUT_3[18819] = 32'b00000000000000001101110010010101;
assign LUT_3[18820] = 32'b00000000000000000010001101001010;
assign LUT_3[18821] = 32'b00000000000000001000111000100111;
assign LUT_3[18822] = 32'b00000000000000000100010100101110;
assign LUT_3[18823] = 32'b00000000000000001011000000001011;
assign LUT_3[18824] = 32'b00000000000000001010011000011010;
assign LUT_3[18825] = 32'b00000000000000010001000011110111;
assign LUT_3[18826] = 32'b00000000000000001100011111111110;
assign LUT_3[18827] = 32'b00000000000000010011001011011011;
assign LUT_3[18828] = 32'b00000000000000000111100110010000;
assign LUT_3[18829] = 32'b00000000000000001110010001101101;
assign LUT_3[18830] = 32'b00000000000000001001101101110100;
assign LUT_3[18831] = 32'b00000000000000010000011001010001;
assign LUT_3[18832] = 32'b00000000000000001000010010010111;
assign LUT_3[18833] = 32'b00000000000000001110111101110100;
assign LUT_3[18834] = 32'b00000000000000001010011001111011;
assign LUT_3[18835] = 32'b00000000000000010001000101011000;
assign LUT_3[18836] = 32'b00000000000000000101100000001101;
assign LUT_3[18837] = 32'b00000000000000001100001011101010;
assign LUT_3[18838] = 32'b00000000000000000111100111110001;
assign LUT_3[18839] = 32'b00000000000000001110010011001110;
assign LUT_3[18840] = 32'b00000000000000001101101011011101;
assign LUT_3[18841] = 32'b00000000000000010100010110111010;
assign LUT_3[18842] = 32'b00000000000000001111110011000001;
assign LUT_3[18843] = 32'b00000000000000010110011110011110;
assign LUT_3[18844] = 32'b00000000000000001010111001010011;
assign LUT_3[18845] = 32'b00000000000000010001100100110000;
assign LUT_3[18846] = 32'b00000000000000001101000000110111;
assign LUT_3[18847] = 32'b00000000000000010011101100010100;
assign LUT_3[18848] = 32'b00000000000000000110001101110100;
assign LUT_3[18849] = 32'b00000000000000001100111001010001;
assign LUT_3[18850] = 32'b00000000000000001000010101011000;
assign LUT_3[18851] = 32'b00000000000000001111000000110101;
assign LUT_3[18852] = 32'b00000000000000000011011011101010;
assign LUT_3[18853] = 32'b00000000000000001010000111000111;
assign LUT_3[18854] = 32'b00000000000000000101100011001110;
assign LUT_3[18855] = 32'b00000000000000001100001110101011;
assign LUT_3[18856] = 32'b00000000000000001011100110111010;
assign LUT_3[18857] = 32'b00000000000000010010010010010111;
assign LUT_3[18858] = 32'b00000000000000001101101110011110;
assign LUT_3[18859] = 32'b00000000000000010100011001111011;
assign LUT_3[18860] = 32'b00000000000000001000110100110000;
assign LUT_3[18861] = 32'b00000000000000001111100000001101;
assign LUT_3[18862] = 32'b00000000000000001010111100010100;
assign LUT_3[18863] = 32'b00000000000000010001100111110001;
assign LUT_3[18864] = 32'b00000000000000001001100000110111;
assign LUT_3[18865] = 32'b00000000000000010000001100010100;
assign LUT_3[18866] = 32'b00000000000000001011101000011011;
assign LUT_3[18867] = 32'b00000000000000010010010011111000;
assign LUT_3[18868] = 32'b00000000000000000110101110101101;
assign LUT_3[18869] = 32'b00000000000000001101011010001010;
assign LUT_3[18870] = 32'b00000000000000001000110110010001;
assign LUT_3[18871] = 32'b00000000000000001111100001101110;
assign LUT_3[18872] = 32'b00000000000000001110111001111101;
assign LUT_3[18873] = 32'b00000000000000010101100101011010;
assign LUT_3[18874] = 32'b00000000000000010001000001100001;
assign LUT_3[18875] = 32'b00000000000000010111101100111110;
assign LUT_3[18876] = 32'b00000000000000001100000111110011;
assign LUT_3[18877] = 32'b00000000000000010010110011010000;
assign LUT_3[18878] = 32'b00000000000000001110001111010111;
assign LUT_3[18879] = 32'b00000000000000010100111010110100;
assign LUT_3[18880] = 32'b00000000000000000100110111111111;
assign LUT_3[18881] = 32'b00000000000000001011100011011100;
assign LUT_3[18882] = 32'b00000000000000000110111111100011;
assign LUT_3[18883] = 32'b00000000000000001101101011000000;
assign LUT_3[18884] = 32'b00000000000000000010000101110101;
assign LUT_3[18885] = 32'b00000000000000001000110001010010;
assign LUT_3[18886] = 32'b00000000000000000100001101011001;
assign LUT_3[18887] = 32'b00000000000000001010111000110110;
assign LUT_3[18888] = 32'b00000000000000001010010001000101;
assign LUT_3[18889] = 32'b00000000000000010000111100100010;
assign LUT_3[18890] = 32'b00000000000000001100011000101001;
assign LUT_3[18891] = 32'b00000000000000010011000100000110;
assign LUT_3[18892] = 32'b00000000000000000111011110111011;
assign LUT_3[18893] = 32'b00000000000000001110001010011000;
assign LUT_3[18894] = 32'b00000000000000001001100110011111;
assign LUT_3[18895] = 32'b00000000000000010000010001111100;
assign LUT_3[18896] = 32'b00000000000000001000001011000010;
assign LUT_3[18897] = 32'b00000000000000001110110110011111;
assign LUT_3[18898] = 32'b00000000000000001010010010100110;
assign LUT_3[18899] = 32'b00000000000000010000111110000011;
assign LUT_3[18900] = 32'b00000000000000000101011000111000;
assign LUT_3[18901] = 32'b00000000000000001100000100010101;
assign LUT_3[18902] = 32'b00000000000000000111100000011100;
assign LUT_3[18903] = 32'b00000000000000001110001011111001;
assign LUT_3[18904] = 32'b00000000000000001101100100001000;
assign LUT_3[18905] = 32'b00000000000000010100001111100101;
assign LUT_3[18906] = 32'b00000000000000001111101011101100;
assign LUT_3[18907] = 32'b00000000000000010110010111001001;
assign LUT_3[18908] = 32'b00000000000000001010110001111110;
assign LUT_3[18909] = 32'b00000000000000010001011101011011;
assign LUT_3[18910] = 32'b00000000000000001100111001100010;
assign LUT_3[18911] = 32'b00000000000000010011100100111111;
assign LUT_3[18912] = 32'b00000000000000000110000110011111;
assign LUT_3[18913] = 32'b00000000000000001100110001111100;
assign LUT_3[18914] = 32'b00000000000000001000001110000011;
assign LUT_3[18915] = 32'b00000000000000001110111001100000;
assign LUT_3[18916] = 32'b00000000000000000011010100010101;
assign LUT_3[18917] = 32'b00000000000000001001111111110010;
assign LUT_3[18918] = 32'b00000000000000000101011011111001;
assign LUT_3[18919] = 32'b00000000000000001100000111010110;
assign LUT_3[18920] = 32'b00000000000000001011011111100101;
assign LUT_3[18921] = 32'b00000000000000010010001011000010;
assign LUT_3[18922] = 32'b00000000000000001101100111001001;
assign LUT_3[18923] = 32'b00000000000000010100010010100110;
assign LUT_3[18924] = 32'b00000000000000001000101101011011;
assign LUT_3[18925] = 32'b00000000000000001111011000111000;
assign LUT_3[18926] = 32'b00000000000000001010110100111111;
assign LUT_3[18927] = 32'b00000000000000010001100000011100;
assign LUT_3[18928] = 32'b00000000000000001001011001100010;
assign LUT_3[18929] = 32'b00000000000000010000000100111111;
assign LUT_3[18930] = 32'b00000000000000001011100001000110;
assign LUT_3[18931] = 32'b00000000000000010010001100100011;
assign LUT_3[18932] = 32'b00000000000000000110100111011000;
assign LUT_3[18933] = 32'b00000000000000001101010010110101;
assign LUT_3[18934] = 32'b00000000000000001000101110111100;
assign LUT_3[18935] = 32'b00000000000000001111011010011001;
assign LUT_3[18936] = 32'b00000000000000001110110010101000;
assign LUT_3[18937] = 32'b00000000000000010101011110000101;
assign LUT_3[18938] = 32'b00000000000000010000111010001100;
assign LUT_3[18939] = 32'b00000000000000010111100101101001;
assign LUT_3[18940] = 32'b00000000000000001100000000011110;
assign LUT_3[18941] = 32'b00000000000000010010101011111011;
assign LUT_3[18942] = 32'b00000000000000001110001000000010;
assign LUT_3[18943] = 32'b00000000000000010100110011011111;
assign LUT_3[18944] = 32'b00000000000000001001111010000001;
assign LUT_3[18945] = 32'b00000000000000010000100101011110;
assign LUT_3[18946] = 32'b00000000000000001100000001100101;
assign LUT_3[18947] = 32'b00000000000000010010101101000010;
assign LUT_3[18948] = 32'b00000000000000000111000111110111;
assign LUT_3[18949] = 32'b00000000000000001101110011010100;
assign LUT_3[18950] = 32'b00000000000000001001001111011011;
assign LUT_3[18951] = 32'b00000000000000001111111010111000;
assign LUT_3[18952] = 32'b00000000000000001111010011000111;
assign LUT_3[18953] = 32'b00000000000000010101111110100100;
assign LUT_3[18954] = 32'b00000000000000010001011010101011;
assign LUT_3[18955] = 32'b00000000000000011000000110001000;
assign LUT_3[18956] = 32'b00000000000000001100100000111101;
assign LUT_3[18957] = 32'b00000000000000010011001100011010;
assign LUT_3[18958] = 32'b00000000000000001110101000100001;
assign LUT_3[18959] = 32'b00000000000000010101010011111110;
assign LUT_3[18960] = 32'b00000000000000001101001101000100;
assign LUT_3[18961] = 32'b00000000000000010011111000100001;
assign LUT_3[18962] = 32'b00000000000000001111010100101000;
assign LUT_3[18963] = 32'b00000000000000010110000000000101;
assign LUT_3[18964] = 32'b00000000000000001010011010111010;
assign LUT_3[18965] = 32'b00000000000000010001000110010111;
assign LUT_3[18966] = 32'b00000000000000001100100010011110;
assign LUT_3[18967] = 32'b00000000000000010011001101111011;
assign LUT_3[18968] = 32'b00000000000000010010100110001010;
assign LUT_3[18969] = 32'b00000000000000011001010001100111;
assign LUT_3[18970] = 32'b00000000000000010100101101101110;
assign LUT_3[18971] = 32'b00000000000000011011011001001011;
assign LUT_3[18972] = 32'b00000000000000001111110100000000;
assign LUT_3[18973] = 32'b00000000000000010110011111011101;
assign LUT_3[18974] = 32'b00000000000000010001111011100100;
assign LUT_3[18975] = 32'b00000000000000011000100111000001;
assign LUT_3[18976] = 32'b00000000000000001011001000100001;
assign LUT_3[18977] = 32'b00000000000000010001110011111110;
assign LUT_3[18978] = 32'b00000000000000001101010000000101;
assign LUT_3[18979] = 32'b00000000000000010011111011100010;
assign LUT_3[18980] = 32'b00000000000000001000010110010111;
assign LUT_3[18981] = 32'b00000000000000001111000001110100;
assign LUT_3[18982] = 32'b00000000000000001010011101111011;
assign LUT_3[18983] = 32'b00000000000000010001001001011000;
assign LUT_3[18984] = 32'b00000000000000010000100001100111;
assign LUT_3[18985] = 32'b00000000000000010111001101000100;
assign LUT_3[18986] = 32'b00000000000000010010101001001011;
assign LUT_3[18987] = 32'b00000000000000011001010100101000;
assign LUT_3[18988] = 32'b00000000000000001101101111011101;
assign LUT_3[18989] = 32'b00000000000000010100011010111010;
assign LUT_3[18990] = 32'b00000000000000001111110111000001;
assign LUT_3[18991] = 32'b00000000000000010110100010011110;
assign LUT_3[18992] = 32'b00000000000000001110011011100100;
assign LUT_3[18993] = 32'b00000000000000010101000111000001;
assign LUT_3[18994] = 32'b00000000000000010000100011001000;
assign LUT_3[18995] = 32'b00000000000000010111001110100101;
assign LUT_3[18996] = 32'b00000000000000001011101001011010;
assign LUT_3[18997] = 32'b00000000000000010010010100110111;
assign LUT_3[18998] = 32'b00000000000000001101110000111110;
assign LUT_3[18999] = 32'b00000000000000010100011100011011;
assign LUT_3[19000] = 32'b00000000000000010011110100101010;
assign LUT_3[19001] = 32'b00000000000000011010100000000111;
assign LUT_3[19002] = 32'b00000000000000010101111100001110;
assign LUT_3[19003] = 32'b00000000000000011100100111101011;
assign LUT_3[19004] = 32'b00000000000000010001000010100000;
assign LUT_3[19005] = 32'b00000000000000010111101101111101;
assign LUT_3[19006] = 32'b00000000000000010011001010000100;
assign LUT_3[19007] = 32'b00000000000000011001110101100001;
assign LUT_3[19008] = 32'b00000000000000001001110010101100;
assign LUT_3[19009] = 32'b00000000000000010000011110001001;
assign LUT_3[19010] = 32'b00000000000000001011111010010000;
assign LUT_3[19011] = 32'b00000000000000010010100101101101;
assign LUT_3[19012] = 32'b00000000000000000111000000100010;
assign LUT_3[19013] = 32'b00000000000000001101101011111111;
assign LUT_3[19014] = 32'b00000000000000001001001000000110;
assign LUT_3[19015] = 32'b00000000000000001111110011100011;
assign LUT_3[19016] = 32'b00000000000000001111001011110010;
assign LUT_3[19017] = 32'b00000000000000010101110111001111;
assign LUT_3[19018] = 32'b00000000000000010001010011010110;
assign LUT_3[19019] = 32'b00000000000000010111111110110011;
assign LUT_3[19020] = 32'b00000000000000001100011001101000;
assign LUT_3[19021] = 32'b00000000000000010011000101000101;
assign LUT_3[19022] = 32'b00000000000000001110100001001100;
assign LUT_3[19023] = 32'b00000000000000010101001100101001;
assign LUT_3[19024] = 32'b00000000000000001101000101101111;
assign LUT_3[19025] = 32'b00000000000000010011110001001100;
assign LUT_3[19026] = 32'b00000000000000001111001101010011;
assign LUT_3[19027] = 32'b00000000000000010101111000110000;
assign LUT_3[19028] = 32'b00000000000000001010010011100101;
assign LUT_3[19029] = 32'b00000000000000010000111111000010;
assign LUT_3[19030] = 32'b00000000000000001100011011001001;
assign LUT_3[19031] = 32'b00000000000000010011000110100110;
assign LUT_3[19032] = 32'b00000000000000010010011110110101;
assign LUT_3[19033] = 32'b00000000000000011001001010010010;
assign LUT_3[19034] = 32'b00000000000000010100100110011001;
assign LUT_3[19035] = 32'b00000000000000011011010001110110;
assign LUT_3[19036] = 32'b00000000000000001111101100101011;
assign LUT_3[19037] = 32'b00000000000000010110011000001000;
assign LUT_3[19038] = 32'b00000000000000010001110100001111;
assign LUT_3[19039] = 32'b00000000000000011000011111101100;
assign LUT_3[19040] = 32'b00000000000000001011000001001100;
assign LUT_3[19041] = 32'b00000000000000010001101100101001;
assign LUT_3[19042] = 32'b00000000000000001101001000110000;
assign LUT_3[19043] = 32'b00000000000000010011110100001101;
assign LUT_3[19044] = 32'b00000000000000001000001111000010;
assign LUT_3[19045] = 32'b00000000000000001110111010011111;
assign LUT_3[19046] = 32'b00000000000000001010010110100110;
assign LUT_3[19047] = 32'b00000000000000010001000010000011;
assign LUT_3[19048] = 32'b00000000000000010000011010010010;
assign LUT_3[19049] = 32'b00000000000000010111000101101111;
assign LUT_3[19050] = 32'b00000000000000010010100001110110;
assign LUT_3[19051] = 32'b00000000000000011001001101010011;
assign LUT_3[19052] = 32'b00000000000000001101101000001000;
assign LUT_3[19053] = 32'b00000000000000010100010011100101;
assign LUT_3[19054] = 32'b00000000000000001111101111101100;
assign LUT_3[19055] = 32'b00000000000000010110011011001001;
assign LUT_3[19056] = 32'b00000000000000001110010100001111;
assign LUT_3[19057] = 32'b00000000000000010100111111101100;
assign LUT_3[19058] = 32'b00000000000000010000011011110011;
assign LUT_3[19059] = 32'b00000000000000010111000111010000;
assign LUT_3[19060] = 32'b00000000000000001011100010000101;
assign LUT_3[19061] = 32'b00000000000000010010001101100010;
assign LUT_3[19062] = 32'b00000000000000001101101001101001;
assign LUT_3[19063] = 32'b00000000000000010100010101000110;
assign LUT_3[19064] = 32'b00000000000000010011101101010101;
assign LUT_3[19065] = 32'b00000000000000011010011000110010;
assign LUT_3[19066] = 32'b00000000000000010101110100111001;
assign LUT_3[19067] = 32'b00000000000000011100100000010110;
assign LUT_3[19068] = 32'b00000000000000010000111011001011;
assign LUT_3[19069] = 32'b00000000000000010111100110101000;
assign LUT_3[19070] = 32'b00000000000000010011000010101111;
assign LUT_3[19071] = 32'b00000000000000011001101110001100;
assign LUT_3[19072] = 32'b00000000000000001100000100111111;
assign LUT_3[19073] = 32'b00000000000000010010110000011100;
assign LUT_3[19074] = 32'b00000000000000001110001100100011;
assign LUT_3[19075] = 32'b00000000000000010100111000000000;
assign LUT_3[19076] = 32'b00000000000000001001010010110101;
assign LUT_3[19077] = 32'b00000000000000001111111110010010;
assign LUT_3[19078] = 32'b00000000000000001011011010011001;
assign LUT_3[19079] = 32'b00000000000000010010000101110110;
assign LUT_3[19080] = 32'b00000000000000010001011110000101;
assign LUT_3[19081] = 32'b00000000000000011000001001100010;
assign LUT_3[19082] = 32'b00000000000000010011100101101001;
assign LUT_3[19083] = 32'b00000000000000011010010001000110;
assign LUT_3[19084] = 32'b00000000000000001110101011111011;
assign LUT_3[19085] = 32'b00000000000000010101010111011000;
assign LUT_3[19086] = 32'b00000000000000010000110011011111;
assign LUT_3[19087] = 32'b00000000000000010111011110111100;
assign LUT_3[19088] = 32'b00000000000000001111011000000010;
assign LUT_3[19089] = 32'b00000000000000010110000011011111;
assign LUT_3[19090] = 32'b00000000000000010001011111100110;
assign LUT_3[19091] = 32'b00000000000000011000001011000011;
assign LUT_3[19092] = 32'b00000000000000001100100101111000;
assign LUT_3[19093] = 32'b00000000000000010011010001010101;
assign LUT_3[19094] = 32'b00000000000000001110101101011100;
assign LUT_3[19095] = 32'b00000000000000010101011000111001;
assign LUT_3[19096] = 32'b00000000000000010100110001001000;
assign LUT_3[19097] = 32'b00000000000000011011011100100101;
assign LUT_3[19098] = 32'b00000000000000010110111000101100;
assign LUT_3[19099] = 32'b00000000000000011101100100001001;
assign LUT_3[19100] = 32'b00000000000000010001111110111110;
assign LUT_3[19101] = 32'b00000000000000011000101010011011;
assign LUT_3[19102] = 32'b00000000000000010100000110100010;
assign LUT_3[19103] = 32'b00000000000000011010110001111111;
assign LUT_3[19104] = 32'b00000000000000001101010011011111;
assign LUT_3[19105] = 32'b00000000000000010011111110111100;
assign LUT_3[19106] = 32'b00000000000000001111011011000011;
assign LUT_3[19107] = 32'b00000000000000010110000110100000;
assign LUT_3[19108] = 32'b00000000000000001010100001010101;
assign LUT_3[19109] = 32'b00000000000000010001001100110010;
assign LUT_3[19110] = 32'b00000000000000001100101000111001;
assign LUT_3[19111] = 32'b00000000000000010011010100010110;
assign LUT_3[19112] = 32'b00000000000000010010101100100101;
assign LUT_3[19113] = 32'b00000000000000011001011000000010;
assign LUT_3[19114] = 32'b00000000000000010100110100001001;
assign LUT_3[19115] = 32'b00000000000000011011011111100110;
assign LUT_3[19116] = 32'b00000000000000001111111010011011;
assign LUT_3[19117] = 32'b00000000000000010110100101111000;
assign LUT_3[19118] = 32'b00000000000000010010000001111111;
assign LUT_3[19119] = 32'b00000000000000011000101101011100;
assign LUT_3[19120] = 32'b00000000000000010000100110100010;
assign LUT_3[19121] = 32'b00000000000000010111010001111111;
assign LUT_3[19122] = 32'b00000000000000010010101110000110;
assign LUT_3[19123] = 32'b00000000000000011001011001100011;
assign LUT_3[19124] = 32'b00000000000000001101110100011000;
assign LUT_3[19125] = 32'b00000000000000010100011111110101;
assign LUT_3[19126] = 32'b00000000000000001111111011111100;
assign LUT_3[19127] = 32'b00000000000000010110100111011001;
assign LUT_3[19128] = 32'b00000000000000010101111111101000;
assign LUT_3[19129] = 32'b00000000000000011100101011000101;
assign LUT_3[19130] = 32'b00000000000000011000000111001100;
assign LUT_3[19131] = 32'b00000000000000011110110010101001;
assign LUT_3[19132] = 32'b00000000000000010011001101011110;
assign LUT_3[19133] = 32'b00000000000000011001111000111011;
assign LUT_3[19134] = 32'b00000000000000010101010101000010;
assign LUT_3[19135] = 32'b00000000000000011100000000011111;
assign LUT_3[19136] = 32'b00000000000000001011111101101010;
assign LUT_3[19137] = 32'b00000000000000010010101001000111;
assign LUT_3[19138] = 32'b00000000000000001110000101001110;
assign LUT_3[19139] = 32'b00000000000000010100110000101011;
assign LUT_3[19140] = 32'b00000000000000001001001011100000;
assign LUT_3[19141] = 32'b00000000000000001111110110111101;
assign LUT_3[19142] = 32'b00000000000000001011010011000100;
assign LUT_3[19143] = 32'b00000000000000010001111110100001;
assign LUT_3[19144] = 32'b00000000000000010001010110110000;
assign LUT_3[19145] = 32'b00000000000000011000000010001101;
assign LUT_3[19146] = 32'b00000000000000010011011110010100;
assign LUT_3[19147] = 32'b00000000000000011010001001110001;
assign LUT_3[19148] = 32'b00000000000000001110100100100110;
assign LUT_3[19149] = 32'b00000000000000010101010000000011;
assign LUT_3[19150] = 32'b00000000000000010000101100001010;
assign LUT_3[19151] = 32'b00000000000000010111010111100111;
assign LUT_3[19152] = 32'b00000000000000001111010000101101;
assign LUT_3[19153] = 32'b00000000000000010101111100001010;
assign LUT_3[19154] = 32'b00000000000000010001011000010001;
assign LUT_3[19155] = 32'b00000000000000011000000011101110;
assign LUT_3[19156] = 32'b00000000000000001100011110100011;
assign LUT_3[19157] = 32'b00000000000000010011001010000000;
assign LUT_3[19158] = 32'b00000000000000001110100110000111;
assign LUT_3[19159] = 32'b00000000000000010101010001100100;
assign LUT_3[19160] = 32'b00000000000000010100101001110011;
assign LUT_3[19161] = 32'b00000000000000011011010101010000;
assign LUT_3[19162] = 32'b00000000000000010110110001010111;
assign LUT_3[19163] = 32'b00000000000000011101011100110100;
assign LUT_3[19164] = 32'b00000000000000010001110111101001;
assign LUT_3[19165] = 32'b00000000000000011000100011000110;
assign LUT_3[19166] = 32'b00000000000000010011111111001101;
assign LUT_3[19167] = 32'b00000000000000011010101010101010;
assign LUT_3[19168] = 32'b00000000000000001101001100001010;
assign LUT_3[19169] = 32'b00000000000000010011110111100111;
assign LUT_3[19170] = 32'b00000000000000001111010011101110;
assign LUT_3[19171] = 32'b00000000000000010101111111001011;
assign LUT_3[19172] = 32'b00000000000000001010011010000000;
assign LUT_3[19173] = 32'b00000000000000010001000101011101;
assign LUT_3[19174] = 32'b00000000000000001100100001100100;
assign LUT_3[19175] = 32'b00000000000000010011001101000001;
assign LUT_3[19176] = 32'b00000000000000010010100101010000;
assign LUT_3[19177] = 32'b00000000000000011001010000101101;
assign LUT_3[19178] = 32'b00000000000000010100101100110100;
assign LUT_3[19179] = 32'b00000000000000011011011000010001;
assign LUT_3[19180] = 32'b00000000000000001111110011000110;
assign LUT_3[19181] = 32'b00000000000000010110011110100011;
assign LUT_3[19182] = 32'b00000000000000010001111010101010;
assign LUT_3[19183] = 32'b00000000000000011000100110000111;
assign LUT_3[19184] = 32'b00000000000000010000011111001101;
assign LUT_3[19185] = 32'b00000000000000010111001010101010;
assign LUT_3[19186] = 32'b00000000000000010010100110110001;
assign LUT_3[19187] = 32'b00000000000000011001010010001110;
assign LUT_3[19188] = 32'b00000000000000001101101101000011;
assign LUT_3[19189] = 32'b00000000000000010100011000100000;
assign LUT_3[19190] = 32'b00000000000000001111110100100111;
assign LUT_3[19191] = 32'b00000000000000010110100000000100;
assign LUT_3[19192] = 32'b00000000000000010101111000010011;
assign LUT_3[19193] = 32'b00000000000000011100100011110000;
assign LUT_3[19194] = 32'b00000000000000010111111111110111;
assign LUT_3[19195] = 32'b00000000000000011110101011010100;
assign LUT_3[19196] = 32'b00000000000000010011000110001001;
assign LUT_3[19197] = 32'b00000000000000011001110001100110;
assign LUT_3[19198] = 32'b00000000000000010101001101101101;
assign LUT_3[19199] = 32'b00000000000000011011111001001010;
assign LUT_3[19200] = 32'b00000000000000000110001001100010;
assign LUT_3[19201] = 32'b00000000000000001100110100111111;
assign LUT_3[19202] = 32'b00000000000000001000010001000110;
assign LUT_3[19203] = 32'b00000000000000001110111100100011;
assign LUT_3[19204] = 32'b00000000000000000011010111011000;
assign LUT_3[19205] = 32'b00000000000000001010000010110101;
assign LUT_3[19206] = 32'b00000000000000000101011110111100;
assign LUT_3[19207] = 32'b00000000000000001100001010011001;
assign LUT_3[19208] = 32'b00000000000000001011100010101000;
assign LUT_3[19209] = 32'b00000000000000010010001110000101;
assign LUT_3[19210] = 32'b00000000000000001101101010001100;
assign LUT_3[19211] = 32'b00000000000000010100010101101001;
assign LUT_3[19212] = 32'b00000000000000001000110000011110;
assign LUT_3[19213] = 32'b00000000000000001111011011111011;
assign LUT_3[19214] = 32'b00000000000000001010111000000010;
assign LUT_3[19215] = 32'b00000000000000010001100011011111;
assign LUT_3[19216] = 32'b00000000000000001001011100100101;
assign LUT_3[19217] = 32'b00000000000000010000001000000010;
assign LUT_3[19218] = 32'b00000000000000001011100100001001;
assign LUT_3[19219] = 32'b00000000000000010010001111100110;
assign LUT_3[19220] = 32'b00000000000000000110101010011011;
assign LUT_3[19221] = 32'b00000000000000001101010101111000;
assign LUT_3[19222] = 32'b00000000000000001000110001111111;
assign LUT_3[19223] = 32'b00000000000000001111011101011100;
assign LUT_3[19224] = 32'b00000000000000001110110101101011;
assign LUT_3[19225] = 32'b00000000000000010101100001001000;
assign LUT_3[19226] = 32'b00000000000000010000111101001111;
assign LUT_3[19227] = 32'b00000000000000010111101000101100;
assign LUT_3[19228] = 32'b00000000000000001100000011100001;
assign LUT_3[19229] = 32'b00000000000000010010101110111110;
assign LUT_3[19230] = 32'b00000000000000001110001011000101;
assign LUT_3[19231] = 32'b00000000000000010100110110100010;
assign LUT_3[19232] = 32'b00000000000000000111011000000010;
assign LUT_3[19233] = 32'b00000000000000001110000011011111;
assign LUT_3[19234] = 32'b00000000000000001001011111100110;
assign LUT_3[19235] = 32'b00000000000000010000001011000011;
assign LUT_3[19236] = 32'b00000000000000000100100101111000;
assign LUT_3[19237] = 32'b00000000000000001011010001010101;
assign LUT_3[19238] = 32'b00000000000000000110101101011100;
assign LUT_3[19239] = 32'b00000000000000001101011000111001;
assign LUT_3[19240] = 32'b00000000000000001100110001001000;
assign LUT_3[19241] = 32'b00000000000000010011011100100101;
assign LUT_3[19242] = 32'b00000000000000001110111000101100;
assign LUT_3[19243] = 32'b00000000000000010101100100001001;
assign LUT_3[19244] = 32'b00000000000000001001111110111110;
assign LUT_3[19245] = 32'b00000000000000010000101010011011;
assign LUT_3[19246] = 32'b00000000000000001100000110100010;
assign LUT_3[19247] = 32'b00000000000000010010110001111111;
assign LUT_3[19248] = 32'b00000000000000001010101011000101;
assign LUT_3[19249] = 32'b00000000000000010001010110100010;
assign LUT_3[19250] = 32'b00000000000000001100110010101001;
assign LUT_3[19251] = 32'b00000000000000010011011110000110;
assign LUT_3[19252] = 32'b00000000000000000111111000111011;
assign LUT_3[19253] = 32'b00000000000000001110100100011000;
assign LUT_3[19254] = 32'b00000000000000001010000000011111;
assign LUT_3[19255] = 32'b00000000000000010000101011111100;
assign LUT_3[19256] = 32'b00000000000000010000000100001011;
assign LUT_3[19257] = 32'b00000000000000010110101111101000;
assign LUT_3[19258] = 32'b00000000000000010010001011101111;
assign LUT_3[19259] = 32'b00000000000000011000110111001100;
assign LUT_3[19260] = 32'b00000000000000001101010010000001;
assign LUT_3[19261] = 32'b00000000000000010011111101011110;
assign LUT_3[19262] = 32'b00000000000000001111011001100101;
assign LUT_3[19263] = 32'b00000000000000010110000101000010;
assign LUT_3[19264] = 32'b00000000000000000110000010001101;
assign LUT_3[19265] = 32'b00000000000000001100101101101010;
assign LUT_3[19266] = 32'b00000000000000001000001001110001;
assign LUT_3[19267] = 32'b00000000000000001110110101001110;
assign LUT_3[19268] = 32'b00000000000000000011010000000011;
assign LUT_3[19269] = 32'b00000000000000001001111011100000;
assign LUT_3[19270] = 32'b00000000000000000101010111100111;
assign LUT_3[19271] = 32'b00000000000000001100000011000100;
assign LUT_3[19272] = 32'b00000000000000001011011011010011;
assign LUT_3[19273] = 32'b00000000000000010010000110110000;
assign LUT_3[19274] = 32'b00000000000000001101100010110111;
assign LUT_3[19275] = 32'b00000000000000010100001110010100;
assign LUT_3[19276] = 32'b00000000000000001000101001001001;
assign LUT_3[19277] = 32'b00000000000000001111010100100110;
assign LUT_3[19278] = 32'b00000000000000001010110000101101;
assign LUT_3[19279] = 32'b00000000000000010001011100001010;
assign LUT_3[19280] = 32'b00000000000000001001010101010000;
assign LUT_3[19281] = 32'b00000000000000010000000000101101;
assign LUT_3[19282] = 32'b00000000000000001011011100110100;
assign LUT_3[19283] = 32'b00000000000000010010001000010001;
assign LUT_3[19284] = 32'b00000000000000000110100011000110;
assign LUT_3[19285] = 32'b00000000000000001101001110100011;
assign LUT_3[19286] = 32'b00000000000000001000101010101010;
assign LUT_3[19287] = 32'b00000000000000001111010110000111;
assign LUT_3[19288] = 32'b00000000000000001110101110010110;
assign LUT_3[19289] = 32'b00000000000000010101011001110011;
assign LUT_3[19290] = 32'b00000000000000010000110101111010;
assign LUT_3[19291] = 32'b00000000000000010111100001010111;
assign LUT_3[19292] = 32'b00000000000000001011111100001100;
assign LUT_3[19293] = 32'b00000000000000010010100111101001;
assign LUT_3[19294] = 32'b00000000000000001110000011110000;
assign LUT_3[19295] = 32'b00000000000000010100101111001101;
assign LUT_3[19296] = 32'b00000000000000000111010000101101;
assign LUT_3[19297] = 32'b00000000000000001101111100001010;
assign LUT_3[19298] = 32'b00000000000000001001011000010001;
assign LUT_3[19299] = 32'b00000000000000010000000011101110;
assign LUT_3[19300] = 32'b00000000000000000100011110100011;
assign LUT_3[19301] = 32'b00000000000000001011001010000000;
assign LUT_3[19302] = 32'b00000000000000000110100110000111;
assign LUT_3[19303] = 32'b00000000000000001101010001100100;
assign LUT_3[19304] = 32'b00000000000000001100101001110011;
assign LUT_3[19305] = 32'b00000000000000010011010101010000;
assign LUT_3[19306] = 32'b00000000000000001110110001010111;
assign LUT_3[19307] = 32'b00000000000000010101011100110100;
assign LUT_3[19308] = 32'b00000000000000001001110111101001;
assign LUT_3[19309] = 32'b00000000000000010000100011000110;
assign LUT_3[19310] = 32'b00000000000000001011111111001101;
assign LUT_3[19311] = 32'b00000000000000010010101010101010;
assign LUT_3[19312] = 32'b00000000000000001010100011110000;
assign LUT_3[19313] = 32'b00000000000000010001001111001101;
assign LUT_3[19314] = 32'b00000000000000001100101011010100;
assign LUT_3[19315] = 32'b00000000000000010011010110110001;
assign LUT_3[19316] = 32'b00000000000000000111110001100110;
assign LUT_3[19317] = 32'b00000000000000001110011101000011;
assign LUT_3[19318] = 32'b00000000000000001001111001001010;
assign LUT_3[19319] = 32'b00000000000000010000100100100111;
assign LUT_3[19320] = 32'b00000000000000001111111100110110;
assign LUT_3[19321] = 32'b00000000000000010110101000010011;
assign LUT_3[19322] = 32'b00000000000000010010000100011010;
assign LUT_3[19323] = 32'b00000000000000011000101111110111;
assign LUT_3[19324] = 32'b00000000000000001101001010101100;
assign LUT_3[19325] = 32'b00000000000000010011110110001001;
assign LUT_3[19326] = 32'b00000000000000001111010010010000;
assign LUT_3[19327] = 32'b00000000000000010101111101101101;
assign LUT_3[19328] = 32'b00000000000000001000010100100000;
assign LUT_3[19329] = 32'b00000000000000001110111111111101;
assign LUT_3[19330] = 32'b00000000000000001010011100000100;
assign LUT_3[19331] = 32'b00000000000000010001000111100001;
assign LUT_3[19332] = 32'b00000000000000000101100010010110;
assign LUT_3[19333] = 32'b00000000000000001100001101110011;
assign LUT_3[19334] = 32'b00000000000000000111101001111010;
assign LUT_3[19335] = 32'b00000000000000001110010101010111;
assign LUT_3[19336] = 32'b00000000000000001101101101100110;
assign LUT_3[19337] = 32'b00000000000000010100011001000011;
assign LUT_3[19338] = 32'b00000000000000001111110101001010;
assign LUT_3[19339] = 32'b00000000000000010110100000100111;
assign LUT_3[19340] = 32'b00000000000000001010111011011100;
assign LUT_3[19341] = 32'b00000000000000010001100110111001;
assign LUT_3[19342] = 32'b00000000000000001101000011000000;
assign LUT_3[19343] = 32'b00000000000000010011101110011101;
assign LUT_3[19344] = 32'b00000000000000001011100111100011;
assign LUT_3[19345] = 32'b00000000000000010010010011000000;
assign LUT_3[19346] = 32'b00000000000000001101101111000111;
assign LUT_3[19347] = 32'b00000000000000010100011010100100;
assign LUT_3[19348] = 32'b00000000000000001000110101011001;
assign LUT_3[19349] = 32'b00000000000000001111100000110110;
assign LUT_3[19350] = 32'b00000000000000001010111100111101;
assign LUT_3[19351] = 32'b00000000000000010001101000011010;
assign LUT_3[19352] = 32'b00000000000000010001000000101001;
assign LUT_3[19353] = 32'b00000000000000010111101100000110;
assign LUT_3[19354] = 32'b00000000000000010011001000001101;
assign LUT_3[19355] = 32'b00000000000000011001110011101010;
assign LUT_3[19356] = 32'b00000000000000001110001110011111;
assign LUT_3[19357] = 32'b00000000000000010100111001111100;
assign LUT_3[19358] = 32'b00000000000000010000010110000011;
assign LUT_3[19359] = 32'b00000000000000010111000001100000;
assign LUT_3[19360] = 32'b00000000000000001001100011000000;
assign LUT_3[19361] = 32'b00000000000000010000001110011101;
assign LUT_3[19362] = 32'b00000000000000001011101010100100;
assign LUT_3[19363] = 32'b00000000000000010010010110000001;
assign LUT_3[19364] = 32'b00000000000000000110110000110110;
assign LUT_3[19365] = 32'b00000000000000001101011100010011;
assign LUT_3[19366] = 32'b00000000000000001000111000011010;
assign LUT_3[19367] = 32'b00000000000000001111100011110111;
assign LUT_3[19368] = 32'b00000000000000001110111100000110;
assign LUT_3[19369] = 32'b00000000000000010101100111100011;
assign LUT_3[19370] = 32'b00000000000000010001000011101010;
assign LUT_3[19371] = 32'b00000000000000010111101111000111;
assign LUT_3[19372] = 32'b00000000000000001100001001111100;
assign LUT_3[19373] = 32'b00000000000000010010110101011001;
assign LUT_3[19374] = 32'b00000000000000001110010001100000;
assign LUT_3[19375] = 32'b00000000000000010100111100111101;
assign LUT_3[19376] = 32'b00000000000000001100110110000011;
assign LUT_3[19377] = 32'b00000000000000010011100001100000;
assign LUT_3[19378] = 32'b00000000000000001110111101100111;
assign LUT_3[19379] = 32'b00000000000000010101101001000100;
assign LUT_3[19380] = 32'b00000000000000001010000011111001;
assign LUT_3[19381] = 32'b00000000000000010000101111010110;
assign LUT_3[19382] = 32'b00000000000000001100001011011101;
assign LUT_3[19383] = 32'b00000000000000010010110110111010;
assign LUT_3[19384] = 32'b00000000000000010010001111001001;
assign LUT_3[19385] = 32'b00000000000000011000111010100110;
assign LUT_3[19386] = 32'b00000000000000010100010110101101;
assign LUT_3[19387] = 32'b00000000000000011011000010001010;
assign LUT_3[19388] = 32'b00000000000000001111011100111111;
assign LUT_3[19389] = 32'b00000000000000010110001000011100;
assign LUT_3[19390] = 32'b00000000000000010001100100100011;
assign LUT_3[19391] = 32'b00000000000000011000010000000000;
assign LUT_3[19392] = 32'b00000000000000001000001101001011;
assign LUT_3[19393] = 32'b00000000000000001110111000101000;
assign LUT_3[19394] = 32'b00000000000000001010010100101111;
assign LUT_3[19395] = 32'b00000000000000010001000000001100;
assign LUT_3[19396] = 32'b00000000000000000101011011000001;
assign LUT_3[19397] = 32'b00000000000000001100000110011110;
assign LUT_3[19398] = 32'b00000000000000000111100010100101;
assign LUT_3[19399] = 32'b00000000000000001110001110000010;
assign LUT_3[19400] = 32'b00000000000000001101100110010001;
assign LUT_3[19401] = 32'b00000000000000010100010001101110;
assign LUT_3[19402] = 32'b00000000000000001111101101110101;
assign LUT_3[19403] = 32'b00000000000000010110011001010010;
assign LUT_3[19404] = 32'b00000000000000001010110100000111;
assign LUT_3[19405] = 32'b00000000000000010001011111100100;
assign LUT_3[19406] = 32'b00000000000000001100111011101011;
assign LUT_3[19407] = 32'b00000000000000010011100111001000;
assign LUT_3[19408] = 32'b00000000000000001011100000001110;
assign LUT_3[19409] = 32'b00000000000000010010001011101011;
assign LUT_3[19410] = 32'b00000000000000001101100111110010;
assign LUT_3[19411] = 32'b00000000000000010100010011001111;
assign LUT_3[19412] = 32'b00000000000000001000101110000100;
assign LUT_3[19413] = 32'b00000000000000001111011001100001;
assign LUT_3[19414] = 32'b00000000000000001010110101101000;
assign LUT_3[19415] = 32'b00000000000000010001100001000101;
assign LUT_3[19416] = 32'b00000000000000010000111001010100;
assign LUT_3[19417] = 32'b00000000000000010111100100110001;
assign LUT_3[19418] = 32'b00000000000000010011000000111000;
assign LUT_3[19419] = 32'b00000000000000011001101100010101;
assign LUT_3[19420] = 32'b00000000000000001110000111001010;
assign LUT_3[19421] = 32'b00000000000000010100110010100111;
assign LUT_3[19422] = 32'b00000000000000010000001110101110;
assign LUT_3[19423] = 32'b00000000000000010110111010001011;
assign LUT_3[19424] = 32'b00000000000000001001011011101011;
assign LUT_3[19425] = 32'b00000000000000010000000111001000;
assign LUT_3[19426] = 32'b00000000000000001011100011001111;
assign LUT_3[19427] = 32'b00000000000000010010001110101100;
assign LUT_3[19428] = 32'b00000000000000000110101001100001;
assign LUT_3[19429] = 32'b00000000000000001101010100111110;
assign LUT_3[19430] = 32'b00000000000000001000110001000101;
assign LUT_3[19431] = 32'b00000000000000001111011100100010;
assign LUT_3[19432] = 32'b00000000000000001110110100110001;
assign LUT_3[19433] = 32'b00000000000000010101100000001110;
assign LUT_3[19434] = 32'b00000000000000010000111100010101;
assign LUT_3[19435] = 32'b00000000000000010111100111110010;
assign LUT_3[19436] = 32'b00000000000000001100000010100111;
assign LUT_3[19437] = 32'b00000000000000010010101110000100;
assign LUT_3[19438] = 32'b00000000000000001110001010001011;
assign LUT_3[19439] = 32'b00000000000000010100110101101000;
assign LUT_3[19440] = 32'b00000000000000001100101110101110;
assign LUT_3[19441] = 32'b00000000000000010011011010001011;
assign LUT_3[19442] = 32'b00000000000000001110110110010010;
assign LUT_3[19443] = 32'b00000000000000010101100001101111;
assign LUT_3[19444] = 32'b00000000000000001001111100100100;
assign LUT_3[19445] = 32'b00000000000000010000101000000001;
assign LUT_3[19446] = 32'b00000000000000001100000100001000;
assign LUT_3[19447] = 32'b00000000000000010010101111100101;
assign LUT_3[19448] = 32'b00000000000000010010000111110100;
assign LUT_3[19449] = 32'b00000000000000011000110011010001;
assign LUT_3[19450] = 32'b00000000000000010100001111011000;
assign LUT_3[19451] = 32'b00000000000000011010111010110101;
assign LUT_3[19452] = 32'b00000000000000001111010101101010;
assign LUT_3[19453] = 32'b00000000000000010110000001000111;
assign LUT_3[19454] = 32'b00000000000000010001011101001110;
assign LUT_3[19455] = 32'b00000000000000011000001000101011;
assign LUT_3[19456] = 32'b00000000000000001101001001110010;
assign LUT_3[19457] = 32'b00000000000000010011110101001111;
assign LUT_3[19458] = 32'b00000000000000001111010001010110;
assign LUT_3[19459] = 32'b00000000000000010101111100110011;
assign LUT_3[19460] = 32'b00000000000000001010010111101000;
assign LUT_3[19461] = 32'b00000000000000010001000011000101;
assign LUT_3[19462] = 32'b00000000000000001100011111001100;
assign LUT_3[19463] = 32'b00000000000000010011001010101001;
assign LUT_3[19464] = 32'b00000000000000010010100010111000;
assign LUT_3[19465] = 32'b00000000000000011001001110010101;
assign LUT_3[19466] = 32'b00000000000000010100101010011100;
assign LUT_3[19467] = 32'b00000000000000011011010101111001;
assign LUT_3[19468] = 32'b00000000000000001111110000101110;
assign LUT_3[19469] = 32'b00000000000000010110011100001011;
assign LUT_3[19470] = 32'b00000000000000010001111000010010;
assign LUT_3[19471] = 32'b00000000000000011000100011101111;
assign LUT_3[19472] = 32'b00000000000000010000011100110101;
assign LUT_3[19473] = 32'b00000000000000010111001000010010;
assign LUT_3[19474] = 32'b00000000000000010010100100011001;
assign LUT_3[19475] = 32'b00000000000000011001001111110110;
assign LUT_3[19476] = 32'b00000000000000001101101010101011;
assign LUT_3[19477] = 32'b00000000000000010100010110001000;
assign LUT_3[19478] = 32'b00000000000000001111110010001111;
assign LUT_3[19479] = 32'b00000000000000010110011101101100;
assign LUT_3[19480] = 32'b00000000000000010101110101111011;
assign LUT_3[19481] = 32'b00000000000000011100100001011000;
assign LUT_3[19482] = 32'b00000000000000010111111101011111;
assign LUT_3[19483] = 32'b00000000000000011110101000111100;
assign LUT_3[19484] = 32'b00000000000000010011000011110001;
assign LUT_3[19485] = 32'b00000000000000011001101111001110;
assign LUT_3[19486] = 32'b00000000000000010101001011010101;
assign LUT_3[19487] = 32'b00000000000000011011110110110010;
assign LUT_3[19488] = 32'b00000000000000001110011000010010;
assign LUT_3[19489] = 32'b00000000000000010101000011101111;
assign LUT_3[19490] = 32'b00000000000000010000011111110110;
assign LUT_3[19491] = 32'b00000000000000010111001011010011;
assign LUT_3[19492] = 32'b00000000000000001011100110001000;
assign LUT_3[19493] = 32'b00000000000000010010010001100101;
assign LUT_3[19494] = 32'b00000000000000001101101101101100;
assign LUT_3[19495] = 32'b00000000000000010100011001001001;
assign LUT_3[19496] = 32'b00000000000000010011110001011000;
assign LUT_3[19497] = 32'b00000000000000011010011100110101;
assign LUT_3[19498] = 32'b00000000000000010101111000111100;
assign LUT_3[19499] = 32'b00000000000000011100100100011001;
assign LUT_3[19500] = 32'b00000000000000010000111111001110;
assign LUT_3[19501] = 32'b00000000000000010111101010101011;
assign LUT_3[19502] = 32'b00000000000000010011000110110010;
assign LUT_3[19503] = 32'b00000000000000011001110010001111;
assign LUT_3[19504] = 32'b00000000000000010001101011010101;
assign LUT_3[19505] = 32'b00000000000000011000010110110010;
assign LUT_3[19506] = 32'b00000000000000010011110010111001;
assign LUT_3[19507] = 32'b00000000000000011010011110010110;
assign LUT_3[19508] = 32'b00000000000000001110111001001011;
assign LUT_3[19509] = 32'b00000000000000010101100100101000;
assign LUT_3[19510] = 32'b00000000000000010001000000101111;
assign LUT_3[19511] = 32'b00000000000000010111101100001100;
assign LUT_3[19512] = 32'b00000000000000010111000100011011;
assign LUT_3[19513] = 32'b00000000000000011101101111111000;
assign LUT_3[19514] = 32'b00000000000000011001001011111111;
assign LUT_3[19515] = 32'b00000000000000011111110111011100;
assign LUT_3[19516] = 32'b00000000000000010100010010010001;
assign LUT_3[19517] = 32'b00000000000000011010111101101110;
assign LUT_3[19518] = 32'b00000000000000010110011001110101;
assign LUT_3[19519] = 32'b00000000000000011101000101010010;
assign LUT_3[19520] = 32'b00000000000000001101000010011101;
assign LUT_3[19521] = 32'b00000000000000010011101101111010;
assign LUT_3[19522] = 32'b00000000000000001111001010000001;
assign LUT_3[19523] = 32'b00000000000000010101110101011110;
assign LUT_3[19524] = 32'b00000000000000001010010000010011;
assign LUT_3[19525] = 32'b00000000000000010000111011110000;
assign LUT_3[19526] = 32'b00000000000000001100010111110111;
assign LUT_3[19527] = 32'b00000000000000010011000011010100;
assign LUT_3[19528] = 32'b00000000000000010010011011100011;
assign LUT_3[19529] = 32'b00000000000000011001000111000000;
assign LUT_3[19530] = 32'b00000000000000010100100011000111;
assign LUT_3[19531] = 32'b00000000000000011011001110100100;
assign LUT_3[19532] = 32'b00000000000000001111101001011001;
assign LUT_3[19533] = 32'b00000000000000010110010100110110;
assign LUT_3[19534] = 32'b00000000000000010001110000111101;
assign LUT_3[19535] = 32'b00000000000000011000011100011010;
assign LUT_3[19536] = 32'b00000000000000010000010101100000;
assign LUT_3[19537] = 32'b00000000000000010111000000111101;
assign LUT_3[19538] = 32'b00000000000000010010011101000100;
assign LUT_3[19539] = 32'b00000000000000011001001000100001;
assign LUT_3[19540] = 32'b00000000000000001101100011010110;
assign LUT_3[19541] = 32'b00000000000000010100001110110011;
assign LUT_3[19542] = 32'b00000000000000001111101010111010;
assign LUT_3[19543] = 32'b00000000000000010110010110010111;
assign LUT_3[19544] = 32'b00000000000000010101101110100110;
assign LUT_3[19545] = 32'b00000000000000011100011010000011;
assign LUT_3[19546] = 32'b00000000000000010111110110001010;
assign LUT_3[19547] = 32'b00000000000000011110100001100111;
assign LUT_3[19548] = 32'b00000000000000010010111100011100;
assign LUT_3[19549] = 32'b00000000000000011001100111111001;
assign LUT_3[19550] = 32'b00000000000000010101000100000000;
assign LUT_3[19551] = 32'b00000000000000011011101111011101;
assign LUT_3[19552] = 32'b00000000000000001110010000111101;
assign LUT_3[19553] = 32'b00000000000000010100111100011010;
assign LUT_3[19554] = 32'b00000000000000010000011000100001;
assign LUT_3[19555] = 32'b00000000000000010111000011111110;
assign LUT_3[19556] = 32'b00000000000000001011011110110011;
assign LUT_3[19557] = 32'b00000000000000010010001010010000;
assign LUT_3[19558] = 32'b00000000000000001101100110010111;
assign LUT_3[19559] = 32'b00000000000000010100010001110100;
assign LUT_3[19560] = 32'b00000000000000010011101010000011;
assign LUT_3[19561] = 32'b00000000000000011010010101100000;
assign LUT_3[19562] = 32'b00000000000000010101110001100111;
assign LUT_3[19563] = 32'b00000000000000011100011101000100;
assign LUT_3[19564] = 32'b00000000000000010000110111111001;
assign LUT_3[19565] = 32'b00000000000000010111100011010110;
assign LUT_3[19566] = 32'b00000000000000010010111111011101;
assign LUT_3[19567] = 32'b00000000000000011001101010111010;
assign LUT_3[19568] = 32'b00000000000000010001100100000000;
assign LUT_3[19569] = 32'b00000000000000011000001111011101;
assign LUT_3[19570] = 32'b00000000000000010011101011100100;
assign LUT_3[19571] = 32'b00000000000000011010010111000001;
assign LUT_3[19572] = 32'b00000000000000001110110001110110;
assign LUT_3[19573] = 32'b00000000000000010101011101010011;
assign LUT_3[19574] = 32'b00000000000000010000111001011010;
assign LUT_3[19575] = 32'b00000000000000010111100100110111;
assign LUT_3[19576] = 32'b00000000000000010110111101000110;
assign LUT_3[19577] = 32'b00000000000000011101101000100011;
assign LUT_3[19578] = 32'b00000000000000011001000100101010;
assign LUT_3[19579] = 32'b00000000000000011111110000000111;
assign LUT_3[19580] = 32'b00000000000000010100001010111100;
assign LUT_3[19581] = 32'b00000000000000011010110110011001;
assign LUT_3[19582] = 32'b00000000000000010110010010100000;
assign LUT_3[19583] = 32'b00000000000000011100111101111101;
assign LUT_3[19584] = 32'b00000000000000001111010100110000;
assign LUT_3[19585] = 32'b00000000000000010110000000001101;
assign LUT_3[19586] = 32'b00000000000000010001011100010100;
assign LUT_3[19587] = 32'b00000000000000011000000111110001;
assign LUT_3[19588] = 32'b00000000000000001100100010100110;
assign LUT_3[19589] = 32'b00000000000000010011001110000011;
assign LUT_3[19590] = 32'b00000000000000001110101010001010;
assign LUT_3[19591] = 32'b00000000000000010101010101100111;
assign LUT_3[19592] = 32'b00000000000000010100101101110110;
assign LUT_3[19593] = 32'b00000000000000011011011001010011;
assign LUT_3[19594] = 32'b00000000000000010110110101011010;
assign LUT_3[19595] = 32'b00000000000000011101100000110111;
assign LUT_3[19596] = 32'b00000000000000010001111011101100;
assign LUT_3[19597] = 32'b00000000000000011000100111001001;
assign LUT_3[19598] = 32'b00000000000000010100000011010000;
assign LUT_3[19599] = 32'b00000000000000011010101110101101;
assign LUT_3[19600] = 32'b00000000000000010010100111110011;
assign LUT_3[19601] = 32'b00000000000000011001010011010000;
assign LUT_3[19602] = 32'b00000000000000010100101111010111;
assign LUT_3[19603] = 32'b00000000000000011011011010110100;
assign LUT_3[19604] = 32'b00000000000000001111110101101001;
assign LUT_3[19605] = 32'b00000000000000010110100001000110;
assign LUT_3[19606] = 32'b00000000000000010001111101001101;
assign LUT_3[19607] = 32'b00000000000000011000101000101010;
assign LUT_3[19608] = 32'b00000000000000011000000000111001;
assign LUT_3[19609] = 32'b00000000000000011110101100010110;
assign LUT_3[19610] = 32'b00000000000000011010001000011101;
assign LUT_3[19611] = 32'b00000000000000100000110011111010;
assign LUT_3[19612] = 32'b00000000000000010101001110101111;
assign LUT_3[19613] = 32'b00000000000000011011111010001100;
assign LUT_3[19614] = 32'b00000000000000010111010110010011;
assign LUT_3[19615] = 32'b00000000000000011110000001110000;
assign LUT_3[19616] = 32'b00000000000000010000100011010000;
assign LUT_3[19617] = 32'b00000000000000010111001110101101;
assign LUT_3[19618] = 32'b00000000000000010010101010110100;
assign LUT_3[19619] = 32'b00000000000000011001010110010001;
assign LUT_3[19620] = 32'b00000000000000001101110001000110;
assign LUT_3[19621] = 32'b00000000000000010100011100100011;
assign LUT_3[19622] = 32'b00000000000000001111111000101010;
assign LUT_3[19623] = 32'b00000000000000010110100100000111;
assign LUT_3[19624] = 32'b00000000000000010101111100010110;
assign LUT_3[19625] = 32'b00000000000000011100100111110011;
assign LUT_3[19626] = 32'b00000000000000011000000011111010;
assign LUT_3[19627] = 32'b00000000000000011110101111010111;
assign LUT_3[19628] = 32'b00000000000000010011001010001100;
assign LUT_3[19629] = 32'b00000000000000011001110101101001;
assign LUT_3[19630] = 32'b00000000000000010101010001110000;
assign LUT_3[19631] = 32'b00000000000000011011111101001101;
assign LUT_3[19632] = 32'b00000000000000010011110110010011;
assign LUT_3[19633] = 32'b00000000000000011010100001110000;
assign LUT_3[19634] = 32'b00000000000000010101111101110111;
assign LUT_3[19635] = 32'b00000000000000011100101001010100;
assign LUT_3[19636] = 32'b00000000000000010001000100001001;
assign LUT_3[19637] = 32'b00000000000000010111101111100110;
assign LUT_3[19638] = 32'b00000000000000010011001011101101;
assign LUT_3[19639] = 32'b00000000000000011001110111001010;
assign LUT_3[19640] = 32'b00000000000000011001001111011001;
assign LUT_3[19641] = 32'b00000000000000011111111010110110;
assign LUT_3[19642] = 32'b00000000000000011011010110111101;
assign LUT_3[19643] = 32'b00000000000000100010000010011010;
assign LUT_3[19644] = 32'b00000000000000010110011101001111;
assign LUT_3[19645] = 32'b00000000000000011101001000101100;
assign LUT_3[19646] = 32'b00000000000000011000100100110011;
assign LUT_3[19647] = 32'b00000000000000011111010000010000;
assign LUT_3[19648] = 32'b00000000000000001111001101011011;
assign LUT_3[19649] = 32'b00000000000000010101111000111000;
assign LUT_3[19650] = 32'b00000000000000010001010100111111;
assign LUT_3[19651] = 32'b00000000000000011000000000011100;
assign LUT_3[19652] = 32'b00000000000000001100011011010001;
assign LUT_3[19653] = 32'b00000000000000010011000110101110;
assign LUT_3[19654] = 32'b00000000000000001110100010110101;
assign LUT_3[19655] = 32'b00000000000000010101001110010010;
assign LUT_3[19656] = 32'b00000000000000010100100110100001;
assign LUT_3[19657] = 32'b00000000000000011011010001111110;
assign LUT_3[19658] = 32'b00000000000000010110101110000101;
assign LUT_3[19659] = 32'b00000000000000011101011001100010;
assign LUT_3[19660] = 32'b00000000000000010001110100010111;
assign LUT_3[19661] = 32'b00000000000000011000011111110100;
assign LUT_3[19662] = 32'b00000000000000010011111011111011;
assign LUT_3[19663] = 32'b00000000000000011010100111011000;
assign LUT_3[19664] = 32'b00000000000000010010100000011110;
assign LUT_3[19665] = 32'b00000000000000011001001011111011;
assign LUT_3[19666] = 32'b00000000000000010100101000000010;
assign LUT_3[19667] = 32'b00000000000000011011010011011111;
assign LUT_3[19668] = 32'b00000000000000001111101110010100;
assign LUT_3[19669] = 32'b00000000000000010110011001110001;
assign LUT_3[19670] = 32'b00000000000000010001110101111000;
assign LUT_3[19671] = 32'b00000000000000011000100001010101;
assign LUT_3[19672] = 32'b00000000000000010111111001100100;
assign LUT_3[19673] = 32'b00000000000000011110100101000001;
assign LUT_3[19674] = 32'b00000000000000011010000001001000;
assign LUT_3[19675] = 32'b00000000000000100000101100100101;
assign LUT_3[19676] = 32'b00000000000000010101000111011010;
assign LUT_3[19677] = 32'b00000000000000011011110010110111;
assign LUT_3[19678] = 32'b00000000000000010111001110111110;
assign LUT_3[19679] = 32'b00000000000000011101111010011011;
assign LUT_3[19680] = 32'b00000000000000010000011011111011;
assign LUT_3[19681] = 32'b00000000000000010111000111011000;
assign LUT_3[19682] = 32'b00000000000000010010100011011111;
assign LUT_3[19683] = 32'b00000000000000011001001110111100;
assign LUT_3[19684] = 32'b00000000000000001101101001110001;
assign LUT_3[19685] = 32'b00000000000000010100010101001110;
assign LUT_3[19686] = 32'b00000000000000001111110001010101;
assign LUT_3[19687] = 32'b00000000000000010110011100110010;
assign LUT_3[19688] = 32'b00000000000000010101110101000001;
assign LUT_3[19689] = 32'b00000000000000011100100000011110;
assign LUT_3[19690] = 32'b00000000000000010111111100100101;
assign LUT_3[19691] = 32'b00000000000000011110101000000010;
assign LUT_3[19692] = 32'b00000000000000010011000010110111;
assign LUT_3[19693] = 32'b00000000000000011001101110010100;
assign LUT_3[19694] = 32'b00000000000000010101001010011011;
assign LUT_3[19695] = 32'b00000000000000011011110101111000;
assign LUT_3[19696] = 32'b00000000000000010011101110111110;
assign LUT_3[19697] = 32'b00000000000000011010011010011011;
assign LUT_3[19698] = 32'b00000000000000010101110110100010;
assign LUT_3[19699] = 32'b00000000000000011100100001111111;
assign LUT_3[19700] = 32'b00000000000000010000111100110100;
assign LUT_3[19701] = 32'b00000000000000010111101000010001;
assign LUT_3[19702] = 32'b00000000000000010011000100011000;
assign LUT_3[19703] = 32'b00000000000000011001101111110101;
assign LUT_3[19704] = 32'b00000000000000011001001000000100;
assign LUT_3[19705] = 32'b00000000000000011111110011100001;
assign LUT_3[19706] = 32'b00000000000000011011001111101000;
assign LUT_3[19707] = 32'b00000000000000100001111011000101;
assign LUT_3[19708] = 32'b00000000000000010110010101111010;
assign LUT_3[19709] = 32'b00000000000000011101000001010111;
assign LUT_3[19710] = 32'b00000000000000011000011101011110;
assign LUT_3[19711] = 32'b00000000000000011111001000111011;
assign LUT_3[19712] = 32'b00000000000000001001011001010011;
assign LUT_3[19713] = 32'b00000000000000010000000100110000;
assign LUT_3[19714] = 32'b00000000000000001011100000110111;
assign LUT_3[19715] = 32'b00000000000000010010001100010100;
assign LUT_3[19716] = 32'b00000000000000000110100111001001;
assign LUT_3[19717] = 32'b00000000000000001101010010100110;
assign LUT_3[19718] = 32'b00000000000000001000101110101101;
assign LUT_3[19719] = 32'b00000000000000001111011010001010;
assign LUT_3[19720] = 32'b00000000000000001110110010011001;
assign LUT_3[19721] = 32'b00000000000000010101011101110110;
assign LUT_3[19722] = 32'b00000000000000010000111001111101;
assign LUT_3[19723] = 32'b00000000000000010111100101011010;
assign LUT_3[19724] = 32'b00000000000000001100000000001111;
assign LUT_3[19725] = 32'b00000000000000010010101011101100;
assign LUT_3[19726] = 32'b00000000000000001110000111110011;
assign LUT_3[19727] = 32'b00000000000000010100110011010000;
assign LUT_3[19728] = 32'b00000000000000001100101100010110;
assign LUT_3[19729] = 32'b00000000000000010011010111110011;
assign LUT_3[19730] = 32'b00000000000000001110110011111010;
assign LUT_3[19731] = 32'b00000000000000010101011111010111;
assign LUT_3[19732] = 32'b00000000000000001001111010001100;
assign LUT_3[19733] = 32'b00000000000000010000100101101001;
assign LUT_3[19734] = 32'b00000000000000001100000001110000;
assign LUT_3[19735] = 32'b00000000000000010010101101001101;
assign LUT_3[19736] = 32'b00000000000000010010000101011100;
assign LUT_3[19737] = 32'b00000000000000011000110000111001;
assign LUT_3[19738] = 32'b00000000000000010100001101000000;
assign LUT_3[19739] = 32'b00000000000000011010111000011101;
assign LUT_3[19740] = 32'b00000000000000001111010011010010;
assign LUT_3[19741] = 32'b00000000000000010101111110101111;
assign LUT_3[19742] = 32'b00000000000000010001011010110110;
assign LUT_3[19743] = 32'b00000000000000011000000110010011;
assign LUT_3[19744] = 32'b00000000000000001010100111110011;
assign LUT_3[19745] = 32'b00000000000000010001010011010000;
assign LUT_3[19746] = 32'b00000000000000001100101111010111;
assign LUT_3[19747] = 32'b00000000000000010011011010110100;
assign LUT_3[19748] = 32'b00000000000000000111110101101001;
assign LUT_3[19749] = 32'b00000000000000001110100001000110;
assign LUT_3[19750] = 32'b00000000000000001001111101001101;
assign LUT_3[19751] = 32'b00000000000000010000101000101010;
assign LUT_3[19752] = 32'b00000000000000010000000000111001;
assign LUT_3[19753] = 32'b00000000000000010110101100010110;
assign LUT_3[19754] = 32'b00000000000000010010001000011101;
assign LUT_3[19755] = 32'b00000000000000011000110011111010;
assign LUT_3[19756] = 32'b00000000000000001101001110101111;
assign LUT_3[19757] = 32'b00000000000000010011111010001100;
assign LUT_3[19758] = 32'b00000000000000001111010110010011;
assign LUT_3[19759] = 32'b00000000000000010110000001110000;
assign LUT_3[19760] = 32'b00000000000000001101111010110110;
assign LUT_3[19761] = 32'b00000000000000010100100110010011;
assign LUT_3[19762] = 32'b00000000000000010000000010011010;
assign LUT_3[19763] = 32'b00000000000000010110101101110111;
assign LUT_3[19764] = 32'b00000000000000001011001000101100;
assign LUT_3[19765] = 32'b00000000000000010001110100001001;
assign LUT_3[19766] = 32'b00000000000000001101010000010000;
assign LUT_3[19767] = 32'b00000000000000010011111011101101;
assign LUT_3[19768] = 32'b00000000000000010011010011111100;
assign LUT_3[19769] = 32'b00000000000000011001111111011001;
assign LUT_3[19770] = 32'b00000000000000010101011011100000;
assign LUT_3[19771] = 32'b00000000000000011100000110111101;
assign LUT_3[19772] = 32'b00000000000000010000100001110010;
assign LUT_3[19773] = 32'b00000000000000010111001101001111;
assign LUT_3[19774] = 32'b00000000000000010010101001010110;
assign LUT_3[19775] = 32'b00000000000000011001010100110011;
assign LUT_3[19776] = 32'b00000000000000001001010001111110;
assign LUT_3[19777] = 32'b00000000000000001111111101011011;
assign LUT_3[19778] = 32'b00000000000000001011011001100010;
assign LUT_3[19779] = 32'b00000000000000010010000100111111;
assign LUT_3[19780] = 32'b00000000000000000110011111110100;
assign LUT_3[19781] = 32'b00000000000000001101001011010001;
assign LUT_3[19782] = 32'b00000000000000001000100111011000;
assign LUT_3[19783] = 32'b00000000000000001111010010110101;
assign LUT_3[19784] = 32'b00000000000000001110101011000100;
assign LUT_3[19785] = 32'b00000000000000010101010110100001;
assign LUT_3[19786] = 32'b00000000000000010000110010101000;
assign LUT_3[19787] = 32'b00000000000000010111011110000101;
assign LUT_3[19788] = 32'b00000000000000001011111000111010;
assign LUT_3[19789] = 32'b00000000000000010010100100010111;
assign LUT_3[19790] = 32'b00000000000000001110000000011110;
assign LUT_3[19791] = 32'b00000000000000010100101011111011;
assign LUT_3[19792] = 32'b00000000000000001100100101000001;
assign LUT_3[19793] = 32'b00000000000000010011010000011110;
assign LUT_3[19794] = 32'b00000000000000001110101100100101;
assign LUT_3[19795] = 32'b00000000000000010101011000000010;
assign LUT_3[19796] = 32'b00000000000000001001110010110111;
assign LUT_3[19797] = 32'b00000000000000010000011110010100;
assign LUT_3[19798] = 32'b00000000000000001011111010011011;
assign LUT_3[19799] = 32'b00000000000000010010100101111000;
assign LUT_3[19800] = 32'b00000000000000010001111110000111;
assign LUT_3[19801] = 32'b00000000000000011000101001100100;
assign LUT_3[19802] = 32'b00000000000000010100000101101011;
assign LUT_3[19803] = 32'b00000000000000011010110001001000;
assign LUT_3[19804] = 32'b00000000000000001111001011111101;
assign LUT_3[19805] = 32'b00000000000000010101110111011010;
assign LUT_3[19806] = 32'b00000000000000010001010011100001;
assign LUT_3[19807] = 32'b00000000000000010111111110111110;
assign LUT_3[19808] = 32'b00000000000000001010100000011110;
assign LUT_3[19809] = 32'b00000000000000010001001011111011;
assign LUT_3[19810] = 32'b00000000000000001100101000000010;
assign LUT_3[19811] = 32'b00000000000000010011010011011111;
assign LUT_3[19812] = 32'b00000000000000000111101110010100;
assign LUT_3[19813] = 32'b00000000000000001110011001110001;
assign LUT_3[19814] = 32'b00000000000000001001110101111000;
assign LUT_3[19815] = 32'b00000000000000010000100001010101;
assign LUT_3[19816] = 32'b00000000000000001111111001100100;
assign LUT_3[19817] = 32'b00000000000000010110100101000001;
assign LUT_3[19818] = 32'b00000000000000010010000001001000;
assign LUT_3[19819] = 32'b00000000000000011000101100100101;
assign LUT_3[19820] = 32'b00000000000000001101000111011010;
assign LUT_3[19821] = 32'b00000000000000010011110010110111;
assign LUT_3[19822] = 32'b00000000000000001111001110111110;
assign LUT_3[19823] = 32'b00000000000000010101111010011011;
assign LUT_3[19824] = 32'b00000000000000001101110011100001;
assign LUT_3[19825] = 32'b00000000000000010100011110111110;
assign LUT_3[19826] = 32'b00000000000000001111111011000101;
assign LUT_3[19827] = 32'b00000000000000010110100110100010;
assign LUT_3[19828] = 32'b00000000000000001011000001010111;
assign LUT_3[19829] = 32'b00000000000000010001101100110100;
assign LUT_3[19830] = 32'b00000000000000001101001000111011;
assign LUT_3[19831] = 32'b00000000000000010011110100011000;
assign LUT_3[19832] = 32'b00000000000000010011001100100111;
assign LUT_3[19833] = 32'b00000000000000011001111000000100;
assign LUT_3[19834] = 32'b00000000000000010101010100001011;
assign LUT_3[19835] = 32'b00000000000000011011111111101000;
assign LUT_3[19836] = 32'b00000000000000010000011010011101;
assign LUT_3[19837] = 32'b00000000000000010111000101111010;
assign LUT_3[19838] = 32'b00000000000000010010100010000001;
assign LUT_3[19839] = 32'b00000000000000011001001101011110;
assign LUT_3[19840] = 32'b00000000000000001011100100010001;
assign LUT_3[19841] = 32'b00000000000000010010001111101110;
assign LUT_3[19842] = 32'b00000000000000001101101011110101;
assign LUT_3[19843] = 32'b00000000000000010100010111010010;
assign LUT_3[19844] = 32'b00000000000000001000110010000111;
assign LUT_3[19845] = 32'b00000000000000001111011101100100;
assign LUT_3[19846] = 32'b00000000000000001010111001101011;
assign LUT_3[19847] = 32'b00000000000000010001100101001000;
assign LUT_3[19848] = 32'b00000000000000010000111101010111;
assign LUT_3[19849] = 32'b00000000000000010111101000110100;
assign LUT_3[19850] = 32'b00000000000000010011000100111011;
assign LUT_3[19851] = 32'b00000000000000011001110000011000;
assign LUT_3[19852] = 32'b00000000000000001110001011001101;
assign LUT_3[19853] = 32'b00000000000000010100110110101010;
assign LUT_3[19854] = 32'b00000000000000010000010010110001;
assign LUT_3[19855] = 32'b00000000000000010110111110001110;
assign LUT_3[19856] = 32'b00000000000000001110110111010100;
assign LUT_3[19857] = 32'b00000000000000010101100010110001;
assign LUT_3[19858] = 32'b00000000000000010000111110111000;
assign LUT_3[19859] = 32'b00000000000000010111101010010101;
assign LUT_3[19860] = 32'b00000000000000001100000101001010;
assign LUT_3[19861] = 32'b00000000000000010010110000100111;
assign LUT_3[19862] = 32'b00000000000000001110001100101110;
assign LUT_3[19863] = 32'b00000000000000010100111000001011;
assign LUT_3[19864] = 32'b00000000000000010100010000011010;
assign LUT_3[19865] = 32'b00000000000000011010111011110111;
assign LUT_3[19866] = 32'b00000000000000010110010111111110;
assign LUT_3[19867] = 32'b00000000000000011101000011011011;
assign LUT_3[19868] = 32'b00000000000000010001011110010000;
assign LUT_3[19869] = 32'b00000000000000011000001001101101;
assign LUT_3[19870] = 32'b00000000000000010011100101110100;
assign LUT_3[19871] = 32'b00000000000000011010010001010001;
assign LUT_3[19872] = 32'b00000000000000001100110010110001;
assign LUT_3[19873] = 32'b00000000000000010011011110001110;
assign LUT_3[19874] = 32'b00000000000000001110111010010101;
assign LUT_3[19875] = 32'b00000000000000010101100101110010;
assign LUT_3[19876] = 32'b00000000000000001010000000100111;
assign LUT_3[19877] = 32'b00000000000000010000101100000100;
assign LUT_3[19878] = 32'b00000000000000001100001000001011;
assign LUT_3[19879] = 32'b00000000000000010010110011101000;
assign LUT_3[19880] = 32'b00000000000000010010001011110111;
assign LUT_3[19881] = 32'b00000000000000011000110111010100;
assign LUT_3[19882] = 32'b00000000000000010100010011011011;
assign LUT_3[19883] = 32'b00000000000000011010111110111000;
assign LUT_3[19884] = 32'b00000000000000001111011001101101;
assign LUT_3[19885] = 32'b00000000000000010110000101001010;
assign LUT_3[19886] = 32'b00000000000000010001100001010001;
assign LUT_3[19887] = 32'b00000000000000011000001100101110;
assign LUT_3[19888] = 32'b00000000000000010000000101110100;
assign LUT_3[19889] = 32'b00000000000000010110110001010001;
assign LUT_3[19890] = 32'b00000000000000010010001101011000;
assign LUT_3[19891] = 32'b00000000000000011000111000110101;
assign LUT_3[19892] = 32'b00000000000000001101010011101010;
assign LUT_3[19893] = 32'b00000000000000010011111111000111;
assign LUT_3[19894] = 32'b00000000000000001111011011001110;
assign LUT_3[19895] = 32'b00000000000000010110000110101011;
assign LUT_3[19896] = 32'b00000000000000010101011110111010;
assign LUT_3[19897] = 32'b00000000000000011100001010010111;
assign LUT_3[19898] = 32'b00000000000000010111100110011110;
assign LUT_3[19899] = 32'b00000000000000011110010001111011;
assign LUT_3[19900] = 32'b00000000000000010010101100110000;
assign LUT_3[19901] = 32'b00000000000000011001011000001101;
assign LUT_3[19902] = 32'b00000000000000010100110100010100;
assign LUT_3[19903] = 32'b00000000000000011011011111110001;
assign LUT_3[19904] = 32'b00000000000000001011011100111100;
assign LUT_3[19905] = 32'b00000000000000010010001000011001;
assign LUT_3[19906] = 32'b00000000000000001101100100100000;
assign LUT_3[19907] = 32'b00000000000000010100001111111101;
assign LUT_3[19908] = 32'b00000000000000001000101010110010;
assign LUT_3[19909] = 32'b00000000000000001111010110001111;
assign LUT_3[19910] = 32'b00000000000000001010110010010110;
assign LUT_3[19911] = 32'b00000000000000010001011101110011;
assign LUT_3[19912] = 32'b00000000000000010000110110000010;
assign LUT_3[19913] = 32'b00000000000000010111100001011111;
assign LUT_3[19914] = 32'b00000000000000010010111101100110;
assign LUT_3[19915] = 32'b00000000000000011001101001000011;
assign LUT_3[19916] = 32'b00000000000000001110000011111000;
assign LUT_3[19917] = 32'b00000000000000010100101111010101;
assign LUT_3[19918] = 32'b00000000000000010000001011011100;
assign LUT_3[19919] = 32'b00000000000000010110110110111001;
assign LUT_3[19920] = 32'b00000000000000001110101111111111;
assign LUT_3[19921] = 32'b00000000000000010101011011011100;
assign LUT_3[19922] = 32'b00000000000000010000110111100011;
assign LUT_3[19923] = 32'b00000000000000010111100011000000;
assign LUT_3[19924] = 32'b00000000000000001011111101110101;
assign LUT_3[19925] = 32'b00000000000000010010101001010010;
assign LUT_3[19926] = 32'b00000000000000001110000101011001;
assign LUT_3[19927] = 32'b00000000000000010100110000110110;
assign LUT_3[19928] = 32'b00000000000000010100001001000101;
assign LUT_3[19929] = 32'b00000000000000011010110100100010;
assign LUT_3[19930] = 32'b00000000000000010110010000101001;
assign LUT_3[19931] = 32'b00000000000000011100111100000110;
assign LUT_3[19932] = 32'b00000000000000010001010110111011;
assign LUT_3[19933] = 32'b00000000000000011000000010011000;
assign LUT_3[19934] = 32'b00000000000000010011011110011111;
assign LUT_3[19935] = 32'b00000000000000011010001001111100;
assign LUT_3[19936] = 32'b00000000000000001100101011011100;
assign LUT_3[19937] = 32'b00000000000000010011010110111001;
assign LUT_3[19938] = 32'b00000000000000001110110011000000;
assign LUT_3[19939] = 32'b00000000000000010101011110011101;
assign LUT_3[19940] = 32'b00000000000000001001111001010010;
assign LUT_3[19941] = 32'b00000000000000010000100100101111;
assign LUT_3[19942] = 32'b00000000000000001100000000110110;
assign LUT_3[19943] = 32'b00000000000000010010101100010011;
assign LUT_3[19944] = 32'b00000000000000010010000100100010;
assign LUT_3[19945] = 32'b00000000000000011000101111111111;
assign LUT_3[19946] = 32'b00000000000000010100001100000110;
assign LUT_3[19947] = 32'b00000000000000011010110111100011;
assign LUT_3[19948] = 32'b00000000000000001111010010011000;
assign LUT_3[19949] = 32'b00000000000000010101111101110101;
assign LUT_3[19950] = 32'b00000000000000010001011001111100;
assign LUT_3[19951] = 32'b00000000000000011000000101011001;
assign LUT_3[19952] = 32'b00000000000000001111111110011111;
assign LUT_3[19953] = 32'b00000000000000010110101001111100;
assign LUT_3[19954] = 32'b00000000000000010010000110000011;
assign LUT_3[19955] = 32'b00000000000000011000110001100000;
assign LUT_3[19956] = 32'b00000000000000001101001100010101;
assign LUT_3[19957] = 32'b00000000000000010011110111110010;
assign LUT_3[19958] = 32'b00000000000000001111010011111001;
assign LUT_3[19959] = 32'b00000000000000010101111111010110;
assign LUT_3[19960] = 32'b00000000000000010101010111100101;
assign LUT_3[19961] = 32'b00000000000000011100000011000010;
assign LUT_3[19962] = 32'b00000000000000010111011111001001;
assign LUT_3[19963] = 32'b00000000000000011110001010100110;
assign LUT_3[19964] = 32'b00000000000000010010100101011011;
assign LUT_3[19965] = 32'b00000000000000011001010000111000;
assign LUT_3[19966] = 32'b00000000000000010100101100111111;
assign LUT_3[19967] = 32'b00000000000000011011011000011100;
assign LUT_3[19968] = 32'b00000000000000010000011110111110;
assign LUT_3[19969] = 32'b00000000000000010111001010011011;
assign LUT_3[19970] = 32'b00000000000000010010100110100010;
assign LUT_3[19971] = 32'b00000000000000011001010001111111;
assign LUT_3[19972] = 32'b00000000000000001101101100110100;
assign LUT_3[19973] = 32'b00000000000000010100011000010001;
assign LUT_3[19974] = 32'b00000000000000001111110100011000;
assign LUT_3[19975] = 32'b00000000000000010110011111110101;
assign LUT_3[19976] = 32'b00000000000000010101111000000100;
assign LUT_3[19977] = 32'b00000000000000011100100011100001;
assign LUT_3[19978] = 32'b00000000000000010111111111101000;
assign LUT_3[19979] = 32'b00000000000000011110101011000101;
assign LUT_3[19980] = 32'b00000000000000010011000101111010;
assign LUT_3[19981] = 32'b00000000000000011001110001010111;
assign LUT_3[19982] = 32'b00000000000000010101001101011110;
assign LUT_3[19983] = 32'b00000000000000011011111000111011;
assign LUT_3[19984] = 32'b00000000000000010011110010000001;
assign LUT_3[19985] = 32'b00000000000000011010011101011110;
assign LUT_3[19986] = 32'b00000000000000010101111001100101;
assign LUT_3[19987] = 32'b00000000000000011100100101000010;
assign LUT_3[19988] = 32'b00000000000000010000111111110111;
assign LUT_3[19989] = 32'b00000000000000010111101011010100;
assign LUT_3[19990] = 32'b00000000000000010011000111011011;
assign LUT_3[19991] = 32'b00000000000000011001110010111000;
assign LUT_3[19992] = 32'b00000000000000011001001011000111;
assign LUT_3[19993] = 32'b00000000000000011111110110100100;
assign LUT_3[19994] = 32'b00000000000000011011010010101011;
assign LUT_3[19995] = 32'b00000000000000100001111110001000;
assign LUT_3[19996] = 32'b00000000000000010110011000111101;
assign LUT_3[19997] = 32'b00000000000000011101000100011010;
assign LUT_3[19998] = 32'b00000000000000011000100000100001;
assign LUT_3[19999] = 32'b00000000000000011111001011111110;
assign LUT_3[20000] = 32'b00000000000000010001101101011110;
assign LUT_3[20001] = 32'b00000000000000011000011000111011;
assign LUT_3[20002] = 32'b00000000000000010011110101000010;
assign LUT_3[20003] = 32'b00000000000000011010100000011111;
assign LUT_3[20004] = 32'b00000000000000001110111011010100;
assign LUT_3[20005] = 32'b00000000000000010101100110110001;
assign LUT_3[20006] = 32'b00000000000000010001000010111000;
assign LUT_3[20007] = 32'b00000000000000010111101110010101;
assign LUT_3[20008] = 32'b00000000000000010111000110100100;
assign LUT_3[20009] = 32'b00000000000000011101110010000001;
assign LUT_3[20010] = 32'b00000000000000011001001110001000;
assign LUT_3[20011] = 32'b00000000000000011111111001100101;
assign LUT_3[20012] = 32'b00000000000000010100010100011010;
assign LUT_3[20013] = 32'b00000000000000011010111111110111;
assign LUT_3[20014] = 32'b00000000000000010110011011111110;
assign LUT_3[20015] = 32'b00000000000000011101000111011011;
assign LUT_3[20016] = 32'b00000000000000010101000000100001;
assign LUT_3[20017] = 32'b00000000000000011011101011111110;
assign LUT_3[20018] = 32'b00000000000000010111001000000101;
assign LUT_3[20019] = 32'b00000000000000011101110011100010;
assign LUT_3[20020] = 32'b00000000000000010010001110010111;
assign LUT_3[20021] = 32'b00000000000000011000111001110100;
assign LUT_3[20022] = 32'b00000000000000010100010101111011;
assign LUT_3[20023] = 32'b00000000000000011011000001011000;
assign LUT_3[20024] = 32'b00000000000000011010011001100111;
assign LUT_3[20025] = 32'b00000000000000100001000101000100;
assign LUT_3[20026] = 32'b00000000000000011100100001001011;
assign LUT_3[20027] = 32'b00000000000000100011001100101000;
assign LUT_3[20028] = 32'b00000000000000010111100111011101;
assign LUT_3[20029] = 32'b00000000000000011110010010111010;
assign LUT_3[20030] = 32'b00000000000000011001101111000001;
assign LUT_3[20031] = 32'b00000000000000100000011010011110;
assign LUT_3[20032] = 32'b00000000000000010000010111101001;
assign LUT_3[20033] = 32'b00000000000000010111000011000110;
assign LUT_3[20034] = 32'b00000000000000010010011111001101;
assign LUT_3[20035] = 32'b00000000000000011001001010101010;
assign LUT_3[20036] = 32'b00000000000000001101100101011111;
assign LUT_3[20037] = 32'b00000000000000010100010000111100;
assign LUT_3[20038] = 32'b00000000000000001111101101000011;
assign LUT_3[20039] = 32'b00000000000000010110011000100000;
assign LUT_3[20040] = 32'b00000000000000010101110000101111;
assign LUT_3[20041] = 32'b00000000000000011100011100001100;
assign LUT_3[20042] = 32'b00000000000000010111111000010011;
assign LUT_3[20043] = 32'b00000000000000011110100011110000;
assign LUT_3[20044] = 32'b00000000000000010010111110100101;
assign LUT_3[20045] = 32'b00000000000000011001101010000010;
assign LUT_3[20046] = 32'b00000000000000010101000110001001;
assign LUT_3[20047] = 32'b00000000000000011011110001100110;
assign LUT_3[20048] = 32'b00000000000000010011101010101100;
assign LUT_3[20049] = 32'b00000000000000011010010110001001;
assign LUT_3[20050] = 32'b00000000000000010101110010010000;
assign LUT_3[20051] = 32'b00000000000000011100011101101101;
assign LUT_3[20052] = 32'b00000000000000010000111000100010;
assign LUT_3[20053] = 32'b00000000000000010111100011111111;
assign LUT_3[20054] = 32'b00000000000000010011000000000110;
assign LUT_3[20055] = 32'b00000000000000011001101011100011;
assign LUT_3[20056] = 32'b00000000000000011001000011110010;
assign LUT_3[20057] = 32'b00000000000000011111101111001111;
assign LUT_3[20058] = 32'b00000000000000011011001011010110;
assign LUT_3[20059] = 32'b00000000000000100001110110110011;
assign LUT_3[20060] = 32'b00000000000000010110010001101000;
assign LUT_3[20061] = 32'b00000000000000011100111101000101;
assign LUT_3[20062] = 32'b00000000000000011000011001001100;
assign LUT_3[20063] = 32'b00000000000000011111000100101001;
assign LUT_3[20064] = 32'b00000000000000010001100110001001;
assign LUT_3[20065] = 32'b00000000000000011000010001100110;
assign LUT_3[20066] = 32'b00000000000000010011101101101101;
assign LUT_3[20067] = 32'b00000000000000011010011001001010;
assign LUT_3[20068] = 32'b00000000000000001110110011111111;
assign LUT_3[20069] = 32'b00000000000000010101011111011100;
assign LUT_3[20070] = 32'b00000000000000010000111011100011;
assign LUT_3[20071] = 32'b00000000000000010111100111000000;
assign LUT_3[20072] = 32'b00000000000000010110111111001111;
assign LUT_3[20073] = 32'b00000000000000011101101010101100;
assign LUT_3[20074] = 32'b00000000000000011001000110110011;
assign LUT_3[20075] = 32'b00000000000000011111110010010000;
assign LUT_3[20076] = 32'b00000000000000010100001101000101;
assign LUT_3[20077] = 32'b00000000000000011010111000100010;
assign LUT_3[20078] = 32'b00000000000000010110010100101001;
assign LUT_3[20079] = 32'b00000000000000011101000000000110;
assign LUT_3[20080] = 32'b00000000000000010100111001001100;
assign LUT_3[20081] = 32'b00000000000000011011100100101001;
assign LUT_3[20082] = 32'b00000000000000010111000000110000;
assign LUT_3[20083] = 32'b00000000000000011101101100001101;
assign LUT_3[20084] = 32'b00000000000000010010000111000010;
assign LUT_3[20085] = 32'b00000000000000011000110010011111;
assign LUT_3[20086] = 32'b00000000000000010100001110100110;
assign LUT_3[20087] = 32'b00000000000000011010111010000011;
assign LUT_3[20088] = 32'b00000000000000011010010010010010;
assign LUT_3[20089] = 32'b00000000000000100000111101101111;
assign LUT_3[20090] = 32'b00000000000000011100011001110110;
assign LUT_3[20091] = 32'b00000000000000100011000101010011;
assign LUT_3[20092] = 32'b00000000000000010111100000001000;
assign LUT_3[20093] = 32'b00000000000000011110001011100101;
assign LUT_3[20094] = 32'b00000000000000011001100111101100;
assign LUT_3[20095] = 32'b00000000000000100000010011001001;
assign LUT_3[20096] = 32'b00000000000000010010101001111100;
assign LUT_3[20097] = 32'b00000000000000011001010101011001;
assign LUT_3[20098] = 32'b00000000000000010100110001100000;
assign LUT_3[20099] = 32'b00000000000000011011011100111101;
assign LUT_3[20100] = 32'b00000000000000001111110111110010;
assign LUT_3[20101] = 32'b00000000000000010110100011001111;
assign LUT_3[20102] = 32'b00000000000000010001111111010110;
assign LUT_3[20103] = 32'b00000000000000011000101010110011;
assign LUT_3[20104] = 32'b00000000000000011000000011000010;
assign LUT_3[20105] = 32'b00000000000000011110101110011111;
assign LUT_3[20106] = 32'b00000000000000011010001010100110;
assign LUT_3[20107] = 32'b00000000000000100000110110000011;
assign LUT_3[20108] = 32'b00000000000000010101010000111000;
assign LUT_3[20109] = 32'b00000000000000011011111100010101;
assign LUT_3[20110] = 32'b00000000000000010111011000011100;
assign LUT_3[20111] = 32'b00000000000000011110000011111001;
assign LUT_3[20112] = 32'b00000000000000010101111100111111;
assign LUT_3[20113] = 32'b00000000000000011100101000011100;
assign LUT_3[20114] = 32'b00000000000000011000000100100011;
assign LUT_3[20115] = 32'b00000000000000011110110000000000;
assign LUT_3[20116] = 32'b00000000000000010011001010110101;
assign LUT_3[20117] = 32'b00000000000000011001110110010010;
assign LUT_3[20118] = 32'b00000000000000010101010010011001;
assign LUT_3[20119] = 32'b00000000000000011011111101110110;
assign LUT_3[20120] = 32'b00000000000000011011010110000101;
assign LUT_3[20121] = 32'b00000000000000100010000001100010;
assign LUT_3[20122] = 32'b00000000000000011101011101101001;
assign LUT_3[20123] = 32'b00000000000000100100001001000110;
assign LUT_3[20124] = 32'b00000000000000011000100011111011;
assign LUT_3[20125] = 32'b00000000000000011111001111011000;
assign LUT_3[20126] = 32'b00000000000000011010101011011111;
assign LUT_3[20127] = 32'b00000000000000100001010110111100;
assign LUT_3[20128] = 32'b00000000000000010011111000011100;
assign LUT_3[20129] = 32'b00000000000000011010100011111001;
assign LUT_3[20130] = 32'b00000000000000010110000000000000;
assign LUT_3[20131] = 32'b00000000000000011100101011011101;
assign LUT_3[20132] = 32'b00000000000000010001000110010010;
assign LUT_3[20133] = 32'b00000000000000010111110001101111;
assign LUT_3[20134] = 32'b00000000000000010011001101110110;
assign LUT_3[20135] = 32'b00000000000000011001111001010011;
assign LUT_3[20136] = 32'b00000000000000011001010001100010;
assign LUT_3[20137] = 32'b00000000000000011111111100111111;
assign LUT_3[20138] = 32'b00000000000000011011011001000110;
assign LUT_3[20139] = 32'b00000000000000100010000100100011;
assign LUT_3[20140] = 32'b00000000000000010110011111011000;
assign LUT_3[20141] = 32'b00000000000000011101001010110101;
assign LUT_3[20142] = 32'b00000000000000011000100110111100;
assign LUT_3[20143] = 32'b00000000000000011111010010011001;
assign LUT_3[20144] = 32'b00000000000000010111001011011111;
assign LUT_3[20145] = 32'b00000000000000011101110110111100;
assign LUT_3[20146] = 32'b00000000000000011001010011000011;
assign LUT_3[20147] = 32'b00000000000000011111111110100000;
assign LUT_3[20148] = 32'b00000000000000010100011001010101;
assign LUT_3[20149] = 32'b00000000000000011011000100110010;
assign LUT_3[20150] = 32'b00000000000000010110100000111001;
assign LUT_3[20151] = 32'b00000000000000011101001100010110;
assign LUT_3[20152] = 32'b00000000000000011100100100100101;
assign LUT_3[20153] = 32'b00000000000000100011010000000010;
assign LUT_3[20154] = 32'b00000000000000011110101100001001;
assign LUT_3[20155] = 32'b00000000000000100101010111100110;
assign LUT_3[20156] = 32'b00000000000000011001110010011011;
assign LUT_3[20157] = 32'b00000000000000100000011101111000;
assign LUT_3[20158] = 32'b00000000000000011011111001111111;
assign LUT_3[20159] = 32'b00000000000000100010100101011100;
assign LUT_3[20160] = 32'b00000000000000010010100010100111;
assign LUT_3[20161] = 32'b00000000000000011001001110000100;
assign LUT_3[20162] = 32'b00000000000000010100101010001011;
assign LUT_3[20163] = 32'b00000000000000011011010101101000;
assign LUT_3[20164] = 32'b00000000000000001111110000011101;
assign LUT_3[20165] = 32'b00000000000000010110011011111010;
assign LUT_3[20166] = 32'b00000000000000010001111000000001;
assign LUT_3[20167] = 32'b00000000000000011000100011011110;
assign LUT_3[20168] = 32'b00000000000000010111111011101101;
assign LUT_3[20169] = 32'b00000000000000011110100111001010;
assign LUT_3[20170] = 32'b00000000000000011010000011010001;
assign LUT_3[20171] = 32'b00000000000000100000101110101110;
assign LUT_3[20172] = 32'b00000000000000010101001001100011;
assign LUT_3[20173] = 32'b00000000000000011011110101000000;
assign LUT_3[20174] = 32'b00000000000000010111010001000111;
assign LUT_3[20175] = 32'b00000000000000011101111100100100;
assign LUT_3[20176] = 32'b00000000000000010101110101101010;
assign LUT_3[20177] = 32'b00000000000000011100100001000111;
assign LUT_3[20178] = 32'b00000000000000010111111101001110;
assign LUT_3[20179] = 32'b00000000000000011110101000101011;
assign LUT_3[20180] = 32'b00000000000000010011000011100000;
assign LUT_3[20181] = 32'b00000000000000011001101110111101;
assign LUT_3[20182] = 32'b00000000000000010101001011000100;
assign LUT_3[20183] = 32'b00000000000000011011110110100001;
assign LUT_3[20184] = 32'b00000000000000011011001110110000;
assign LUT_3[20185] = 32'b00000000000000100001111010001101;
assign LUT_3[20186] = 32'b00000000000000011101010110010100;
assign LUT_3[20187] = 32'b00000000000000100100000001110001;
assign LUT_3[20188] = 32'b00000000000000011000011100100110;
assign LUT_3[20189] = 32'b00000000000000011111001000000011;
assign LUT_3[20190] = 32'b00000000000000011010100100001010;
assign LUT_3[20191] = 32'b00000000000000100001001111100111;
assign LUT_3[20192] = 32'b00000000000000010011110001000111;
assign LUT_3[20193] = 32'b00000000000000011010011100100100;
assign LUT_3[20194] = 32'b00000000000000010101111000101011;
assign LUT_3[20195] = 32'b00000000000000011100100100001000;
assign LUT_3[20196] = 32'b00000000000000010000111110111101;
assign LUT_3[20197] = 32'b00000000000000010111101010011010;
assign LUT_3[20198] = 32'b00000000000000010011000110100001;
assign LUT_3[20199] = 32'b00000000000000011001110001111110;
assign LUT_3[20200] = 32'b00000000000000011001001010001101;
assign LUT_3[20201] = 32'b00000000000000011111110101101010;
assign LUT_3[20202] = 32'b00000000000000011011010001110001;
assign LUT_3[20203] = 32'b00000000000000100001111101001110;
assign LUT_3[20204] = 32'b00000000000000010110011000000011;
assign LUT_3[20205] = 32'b00000000000000011101000011100000;
assign LUT_3[20206] = 32'b00000000000000011000011111100111;
assign LUT_3[20207] = 32'b00000000000000011111001011000100;
assign LUT_3[20208] = 32'b00000000000000010111000100001010;
assign LUT_3[20209] = 32'b00000000000000011101101111100111;
assign LUT_3[20210] = 32'b00000000000000011001001011101110;
assign LUT_3[20211] = 32'b00000000000000011111110111001011;
assign LUT_3[20212] = 32'b00000000000000010100010010000000;
assign LUT_3[20213] = 32'b00000000000000011010111101011101;
assign LUT_3[20214] = 32'b00000000000000010110011001100100;
assign LUT_3[20215] = 32'b00000000000000011101000101000001;
assign LUT_3[20216] = 32'b00000000000000011100011101010000;
assign LUT_3[20217] = 32'b00000000000000100011001000101101;
assign LUT_3[20218] = 32'b00000000000000011110100100110100;
assign LUT_3[20219] = 32'b00000000000000100101010000010001;
assign LUT_3[20220] = 32'b00000000000000011001101011000110;
assign LUT_3[20221] = 32'b00000000000000100000010110100011;
assign LUT_3[20222] = 32'b00000000000000011011110010101010;
assign LUT_3[20223] = 32'b00000000000000100010011110000111;
assign LUT_3[20224] = 32'b00000000000000001100101110011111;
assign LUT_3[20225] = 32'b00000000000000010011011001111100;
assign LUT_3[20226] = 32'b00000000000000001110110110000011;
assign LUT_3[20227] = 32'b00000000000000010101100001100000;
assign LUT_3[20228] = 32'b00000000000000001001111100010101;
assign LUT_3[20229] = 32'b00000000000000010000100111110010;
assign LUT_3[20230] = 32'b00000000000000001100000011111001;
assign LUT_3[20231] = 32'b00000000000000010010101111010110;
assign LUT_3[20232] = 32'b00000000000000010010000111100101;
assign LUT_3[20233] = 32'b00000000000000011000110011000010;
assign LUT_3[20234] = 32'b00000000000000010100001111001001;
assign LUT_3[20235] = 32'b00000000000000011010111010100110;
assign LUT_3[20236] = 32'b00000000000000001111010101011011;
assign LUT_3[20237] = 32'b00000000000000010110000000111000;
assign LUT_3[20238] = 32'b00000000000000010001011100111111;
assign LUT_3[20239] = 32'b00000000000000011000001000011100;
assign LUT_3[20240] = 32'b00000000000000010000000001100010;
assign LUT_3[20241] = 32'b00000000000000010110101100111111;
assign LUT_3[20242] = 32'b00000000000000010010001001000110;
assign LUT_3[20243] = 32'b00000000000000011000110100100011;
assign LUT_3[20244] = 32'b00000000000000001101001111011000;
assign LUT_3[20245] = 32'b00000000000000010011111010110101;
assign LUT_3[20246] = 32'b00000000000000001111010110111100;
assign LUT_3[20247] = 32'b00000000000000010110000010011001;
assign LUT_3[20248] = 32'b00000000000000010101011010101000;
assign LUT_3[20249] = 32'b00000000000000011100000110000101;
assign LUT_3[20250] = 32'b00000000000000010111100010001100;
assign LUT_3[20251] = 32'b00000000000000011110001101101001;
assign LUT_3[20252] = 32'b00000000000000010010101000011110;
assign LUT_3[20253] = 32'b00000000000000011001010011111011;
assign LUT_3[20254] = 32'b00000000000000010100110000000010;
assign LUT_3[20255] = 32'b00000000000000011011011011011111;
assign LUT_3[20256] = 32'b00000000000000001101111100111111;
assign LUT_3[20257] = 32'b00000000000000010100101000011100;
assign LUT_3[20258] = 32'b00000000000000010000000100100011;
assign LUT_3[20259] = 32'b00000000000000010110110000000000;
assign LUT_3[20260] = 32'b00000000000000001011001010110101;
assign LUT_3[20261] = 32'b00000000000000010001110110010010;
assign LUT_3[20262] = 32'b00000000000000001101010010011001;
assign LUT_3[20263] = 32'b00000000000000010011111101110110;
assign LUT_3[20264] = 32'b00000000000000010011010110000101;
assign LUT_3[20265] = 32'b00000000000000011010000001100010;
assign LUT_3[20266] = 32'b00000000000000010101011101101001;
assign LUT_3[20267] = 32'b00000000000000011100001001000110;
assign LUT_3[20268] = 32'b00000000000000010000100011111011;
assign LUT_3[20269] = 32'b00000000000000010111001111011000;
assign LUT_3[20270] = 32'b00000000000000010010101011011111;
assign LUT_3[20271] = 32'b00000000000000011001010110111100;
assign LUT_3[20272] = 32'b00000000000000010001010000000010;
assign LUT_3[20273] = 32'b00000000000000010111111011011111;
assign LUT_3[20274] = 32'b00000000000000010011010111100110;
assign LUT_3[20275] = 32'b00000000000000011010000011000011;
assign LUT_3[20276] = 32'b00000000000000001110011101111000;
assign LUT_3[20277] = 32'b00000000000000010101001001010101;
assign LUT_3[20278] = 32'b00000000000000010000100101011100;
assign LUT_3[20279] = 32'b00000000000000010111010000111001;
assign LUT_3[20280] = 32'b00000000000000010110101001001000;
assign LUT_3[20281] = 32'b00000000000000011101010100100101;
assign LUT_3[20282] = 32'b00000000000000011000110000101100;
assign LUT_3[20283] = 32'b00000000000000011111011100001001;
assign LUT_3[20284] = 32'b00000000000000010011110110111110;
assign LUT_3[20285] = 32'b00000000000000011010100010011011;
assign LUT_3[20286] = 32'b00000000000000010101111110100010;
assign LUT_3[20287] = 32'b00000000000000011100101001111111;
assign LUT_3[20288] = 32'b00000000000000001100100111001010;
assign LUT_3[20289] = 32'b00000000000000010011010010100111;
assign LUT_3[20290] = 32'b00000000000000001110101110101110;
assign LUT_3[20291] = 32'b00000000000000010101011010001011;
assign LUT_3[20292] = 32'b00000000000000001001110101000000;
assign LUT_3[20293] = 32'b00000000000000010000100000011101;
assign LUT_3[20294] = 32'b00000000000000001011111100100100;
assign LUT_3[20295] = 32'b00000000000000010010101000000001;
assign LUT_3[20296] = 32'b00000000000000010010000000010000;
assign LUT_3[20297] = 32'b00000000000000011000101011101101;
assign LUT_3[20298] = 32'b00000000000000010100000111110100;
assign LUT_3[20299] = 32'b00000000000000011010110011010001;
assign LUT_3[20300] = 32'b00000000000000001111001110000110;
assign LUT_3[20301] = 32'b00000000000000010101111001100011;
assign LUT_3[20302] = 32'b00000000000000010001010101101010;
assign LUT_3[20303] = 32'b00000000000000011000000001000111;
assign LUT_3[20304] = 32'b00000000000000001111111010001101;
assign LUT_3[20305] = 32'b00000000000000010110100101101010;
assign LUT_3[20306] = 32'b00000000000000010010000001110001;
assign LUT_3[20307] = 32'b00000000000000011000101101001110;
assign LUT_3[20308] = 32'b00000000000000001101001000000011;
assign LUT_3[20309] = 32'b00000000000000010011110011100000;
assign LUT_3[20310] = 32'b00000000000000001111001111100111;
assign LUT_3[20311] = 32'b00000000000000010101111011000100;
assign LUT_3[20312] = 32'b00000000000000010101010011010011;
assign LUT_3[20313] = 32'b00000000000000011011111110110000;
assign LUT_3[20314] = 32'b00000000000000010111011010110111;
assign LUT_3[20315] = 32'b00000000000000011110000110010100;
assign LUT_3[20316] = 32'b00000000000000010010100001001001;
assign LUT_3[20317] = 32'b00000000000000011001001100100110;
assign LUT_3[20318] = 32'b00000000000000010100101000101101;
assign LUT_3[20319] = 32'b00000000000000011011010100001010;
assign LUT_3[20320] = 32'b00000000000000001101110101101010;
assign LUT_3[20321] = 32'b00000000000000010100100001000111;
assign LUT_3[20322] = 32'b00000000000000001111111101001110;
assign LUT_3[20323] = 32'b00000000000000010110101000101011;
assign LUT_3[20324] = 32'b00000000000000001011000011100000;
assign LUT_3[20325] = 32'b00000000000000010001101110111101;
assign LUT_3[20326] = 32'b00000000000000001101001011000100;
assign LUT_3[20327] = 32'b00000000000000010011110110100001;
assign LUT_3[20328] = 32'b00000000000000010011001110110000;
assign LUT_3[20329] = 32'b00000000000000011001111010001101;
assign LUT_3[20330] = 32'b00000000000000010101010110010100;
assign LUT_3[20331] = 32'b00000000000000011100000001110001;
assign LUT_3[20332] = 32'b00000000000000010000011100100110;
assign LUT_3[20333] = 32'b00000000000000010111001000000011;
assign LUT_3[20334] = 32'b00000000000000010010100100001010;
assign LUT_3[20335] = 32'b00000000000000011001001111100111;
assign LUT_3[20336] = 32'b00000000000000010001001000101101;
assign LUT_3[20337] = 32'b00000000000000010111110100001010;
assign LUT_3[20338] = 32'b00000000000000010011010000010001;
assign LUT_3[20339] = 32'b00000000000000011001111011101110;
assign LUT_3[20340] = 32'b00000000000000001110010110100011;
assign LUT_3[20341] = 32'b00000000000000010101000010000000;
assign LUT_3[20342] = 32'b00000000000000010000011110000111;
assign LUT_3[20343] = 32'b00000000000000010111001001100100;
assign LUT_3[20344] = 32'b00000000000000010110100001110011;
assign LUT_3[20345] = 32'b00000000000000011101001101010000;
assign LUT_3[20346] = 32'b00000000000000011000101001010111;
assign LUT_3[20347] = 32'b00000000000000011111010100110100;
assign LUT_3[20348] = 32'b00000000000000010011101111101001;
assign LUT_3[20349] = 32'b00000000000000011010011011000110;
assign LUT_3[20350] = 32'b00000000000000010101110111001101;
assign LUT_3[20351] = 32'b00000000000000011100100010101010;
assign LUT_3[20352] = 32'b00000000000000001110111001011101;
assign LUT_3[20353] = 32'b00000000000000010101100100111010;
assign LUT_3[20354] = 32'b00000000000000010001000001000001;
assign LUT_3[20355] = 32'b00000000000000010111101100011110;
assign LUT_3[20356] = 32'b00000000000000001100000111010011;
assign LUT_3[20357] = 32'b00000000000000010010110010110000;
assign LUT_3[20358] = 32'b00000000000000001110001110110111;
assign LUT_3[20359] = 32'b00000000000000010100111010010100;
assign LUT_3[20360] = 32'b00000000000000010100010010100011;
assign LUT_3[20361] = 32'b00000000000000011010111110000000;
assign LUT_3[20362] = 32'b00000000000000010110011010000111;
assign LUT_3[20363] = 32'b00000000000000011101000101100100;
assign LUT_3[20364] = 32'b00000000000000010001100000011001;
assign LUT_3[20365] = 32'b00000000000000011000001011110110;
assign LUT_3[20366] = 32'b00000000000000010011100111111101;
assign LUT_3[20367] = 32'b00000000000000011010010011011010;
assign LUT_3[20368] = 32'b00000000000000010010001100100000;
assign LUT_3[20369] = 32'b00000000000000011000110111111101;
assign LUT_3[20370] = 32'b00000000000000010100010100000100;
assign LUT_3[20371] = 32'b00000000000000011010111111100001;
assign LUT_3[20372] = 32'b00000000000000001111011010010110;
assign LUT_3[20373] = 32'b00000000000000010110000101110011;
assign LUT_3[20374] = 32'b00000000000000010001100001111010;
assign LUT_3[20375] = 32'b00000000000000011000001101010111;
assign LUT_3[20376] = 32'b00000000000000010111100101100110;
assign LUT_3[20377] = 32'b00000000000000011110010001000011;
assign LUT_3[20378] = 32'b00000000000000011001101101001010;
assign LUT_3[20379] = 32'b00000000000000100000011000100111;
assign LUT_3[20380] = 32'b00000000000000010100110011011100;
assign LUT_3[20381] = 32'b00000000000000011011011110111001;
assign LUT_3[20382] = 32'b00000000000000010110111011000000;
assign LUT_3[20383] = 32'b00000000000000011101100110011101;
assign LUT_3[20384] = 32'b00000000000000010000000111111101;
assign LUT_3[20385] = 32'b00000000000000010110110011011010;
assign LUT_3[20386] = 32'b00000000000000010010001111100001;
assign LUT_3[20387] = 32'b00000000000000011000111010111110;
assign LUT_3[20388] = 32'b00000000000000001101010101110011;
assign LUT_3[20389] = 32'b00000000000000010100000001010000;
assign LUT_3[20390] = 32'b00000000000000001111011101010111;
assign LUT_3[20391] = 32'b00000000000000010110001000110100;
assign LUT_3[20392] = 32'b00000000000000010101100001000011;
assign LUT_3[20393] = 32'b00000000000000011100001100100000;
assign LUT_3[20394] = 32'b00000000000000010111101000100111;
assign LUT_3[20395] = 32'b00000000000000011110010100000100;
assign LUT_3[20396] = 32'b00000000000000010010101110111001;
assign LUT_3[20397] = 32'b00000000000000011001011010010110;
assign LUT_3[20398] = 32'b00000000000000010100110110011101;
assign LUT_3[20399] = 32'b00000000000000011011100001111010;
assign LUT_3[20400] = 32'b00000000000000010011011011000000;
assign LUT_3[20401] = 32'b00000000000000011010000110011101;
assign LUT_3[20402] = 32'b00000000000000010101100010100100;
assign LUT_3[20403] = 32'b00000000000000011100001110000001;
assign LUT_3[20404] = 32'b00000000000000010000101000110110;
assign LUT_3[20405] = 32'b00000000000000010111010100010011;
assign LUT_3[20406] = 32'b00000000000000010010110000011010;
assign LUT_3[20407] = 32'b00000000000000011001011011110111;
assign LUT_3[20408] = 32'b00000000000000011000110100000110;
assign LUT_3[20409] = 32'b00000000000000011111011111100011;
assign LUT_3[20410] = 32'b00000000000000011010111011101010;
assign LUT_3[20411] = 32'b00000000000000100001100111000111;
assign LUT_3[20412] = 32'b00000000000000010110000001111100;
assign LUT_3[20413] = 32'b00000000000000011100101101011001;
assign LUT_3[20414] = 32'b00000000000000011000001001100000;
assign LUT_3[20415] = 32'b00000000000000011110110100111101;
assign LUT_3[20416] = 32'b00000000000000001110110010001000;
assign LUT_3[20417] = 32'b00000000000000010101011101100101;
assign LUT_3[20418] = 32'b00000000000000010000111001101100;
assign LUT_3[20419] = 32'b00000000000000010111100101001001;
assign LUT_3[20420] = 32'b00000000000000001011111111111110;
assign LUT_3[20421] = 32'b00000000000000010010101011011011;
assign LUT_3[20422] = 32'b00000000000000001110000111100010;
assign LUT_3[20423] = 32'b00000000000000010100110010111111;
assign LUT_3[20424] = 32'b00000000000000010100001011001110;
assign LUT_3[20425] = 32'b00000000000000011010110110101011;
assign LUT_3[20426] = 32'b00000000000000010110010010110010;
assign LUT_3[20427] = 32'b00000000000000011100111110001111;
assign LUT_3[20428] = 32'b00000000000000010001011001000100;
assign LUT_3[20429] = 32'b00000000000000011000000100100001;
assign LUT_3[20430] = 32'b00000000000000010011100000101000;
assign LUT_3[20431] = 32'b00000000000000011010001100000101;
assign LUT_3[20432] = 32'b00000000000000010010000101001011;
assign LUT_3[20433] = 32'b00000000000000011000110000101000;
assign LUT_3[20434] = 32'b00000000000000010100001100101111;
assign LUT_3[20435] = 32'b00000000000000011010111000001100;
assign LUT_3[20436] = 32'b00000000000000001111010011000001;
assign LUT_3[20437] = 32'b00000000000000010101111110011110;
assign LUT_3[20438] = 32'b00000000000000010001011010100101;
assign LUT_3[20439] = 32'b00000000000000011000000110000010;
assign LUT_3[20440] = 32'b00000000000000010111011110010001;
assign LUT_3[20441] = 32'b00000000000000011110001001101110;
assign LUT_3[20442] = 32'b00000000000000011001100101110101;
assign LUT_3[20443] = 32'b00000000000000100000010001010010;
assign LUT_3[20444] = 32'b00000000000000010100101100000111;
assign LUT_3[20445] = 32'b00000000000000011011010111100100;
assign LUT_3[20446] = 32'b00000000000000010110110011101011;
assign LUT_3[20447] = 32'b00000000000000011101011111001000;
assign LUT_3[20448] = 32'b00000000000000010000000000101000;
assign LUT_3[20449] = 32'b00000000000000010110101100000101;
assign LUT_3[20450] = 32'b00000000000000010010001000001100;
assign LUT_3[20451] = 32'b00000000000000011000110011101001;
assign LUT_3[20452] = 32'b00000000000000001101001110011110;
assign LUT_3[20453] = 32'b00000000000000010011111001111011;
assign LUT_3[20454] = 32'b00000000000000001111010110000010;
assign LUT_3[20455] = 32'b00000000000000010110000001011111;
assign LUT_3[20456] = 32'b00000000000000010101011001101110;
assign LUT_3[20457] = 32'b00000000000000011100000101001011;
assign LUT_3[20458] = 32'b00000000000000010111100001010010;
assign LUT_3[20459] = 32'b00000000000000011110001100101111;
assign LUT_3[20460] = 32'b00000000000000010010100111100100;
assign LUT_3[20461] = 32'b00000000000000011001010011000001;
assign LUT_3[20462] = 32'b00000000000000010100101111001000;
assign LUT_3[20463] = 32'b00000000000000011011011010100101;
assign LUT_3[20464] = 32'b00000000000000010011010011101011;
assign LUT_3[20465] = 32'b00000000000000011001111111001000;
assign LUT_3[20466] = 32'b00000000000000010101011011001111;
assign LUT_3[20467] = 32'b00000000000000011100000110101100;
assign LUT_3[20468] = 32'b00000000000000010000100001100001;
assign LUT_3[20469] = 32'b00000000000000010111001100111110;
assign LUT_3[20470] = 32'b00000000000000010010101001000101;
assign LUT_3[20471] = 32'b00000000000000011001010100100010;
assign LUT_3[20472] = 32'b00000000000000011000101100110001;
assign LUT_3[20473] = 32'b00000000000000011111011000001110;
assign LUT_3[20474] = 32'b00000000000000011010110100010101;
assign LUT_3[20475] = 32'b00000000000000100001011111110010;
assign LUT_3[20476] = 32'b00000000000000010101111010100111;
assign LUT_3[20477] = 32'b00000000000000011100100110000100;
assign LUT_3[20478] = 32'b00000000000000011000000010001011;
assign LUT_3[20479] = 32'b00000000000000011110101101101000;
assign LUT_3[20480] = 32'b00000000000000001001000000000010;
assign LUT_3[20481] = 32'b00000000000000001111101011011111;
assign LUT_3[20482] = 32'b00000000000000001011000111100110;
assign LUT_3[20483] = 32'b00000000000000010001110011000011;
assign LUT_3[20484] = 32'b00000000000000000110001101111000;
assign LUT_3[20485] = 32'b00000000000000001100111001010101;
assign LUT_3[20486] = 32'b00000000000000001000010101011100;
assign LUT_3[20487] = 32'b00000000000000001111000000111001;
assign LUT_3[20488] = 32'b00000000000000001110011001001000;
assign LUT_3[20489] = 32'b00000000000000010101000100100101;
assign LUT_3[20490] = 32'b00000000000000010000100000101100;
assign LUT_3[20491] = 32'b00000000000000010111001100001001;
assign LUT_3[20492] = 32'b00000000000000001011100110111110;
assign LUT_3[20493] = 32'b00000000000000010010010010011011;
assign LUT_3[20494] = 32'b00000000000000001101101110100010;
assign LUT_3[20495] = 32'b00000000000000010100011001111111;
assign LUT_3[20496] = 32'b00000000000000001100010011000101;
assign LUT_3[20497] = 32'b00000000000000010010111110100010;
assign LUT_3[20498] = 32'b00000000000000001110011010101001;
assign LUT_3[20499] = 32'b00000000000000010101000110000110;
assign LUT_3[20500] = 32'b00000000000000001001100000111011;
assign LUT_3[20501] = 32'b00000000000000010000001100011000;
assign LUT_3[20502] = 32'b00000000000000001011101000011111;
assign LUT_3[20503] = 32'b00000000000000010010010011111100;
assign LUT_3[20504] = 32'b00000000000000010001101100001011;
assign LUT_3[20505] = 32'b00000000000000011000010111101000;
assign LUT_3[20506] = 32'b00000000000000010011110011101111;
assign LUT_3[20507] = 32'b00000000000000011010011111001100;
assign LUT_3[20508] = 32'b00000000000000001110111010000001;
assign LUT_3[20509] = 32'b00000000000000010101100101011110;
assign LUT_3[20510] = 32'b00000000000000010001000001100101;
assign LUT_3[20511] = 32'b00000000000000010111101101000010;
assign LUT_3[20512] = 32'b00000000000000001010001110100010;
assign LUT_3[20513] = 32'b00000000000000010000111001111111;
assign LUT_3[20514] = 32'b00000000000000001100010110000110;
assign LUT_3[20515] = 32'b00000000000000010011000001100011;
assign LUT_3[20516] = 32'b00000000000000000111011100011000;
assign LUT_3[20517] = 32'b00000000000000001110000111110101;
assign LUT_3[20518] = 32'b00000000000000001001100011111100;
assign LUT_3[20519] = 32'b00000000000000010000001111011001;
assign LUT_3[20520] = 32'b00000000000000001111100111101000;
assign LUT_3[20521] = 32'b00000000000000010110010011000101;
assign LUT_3[20522] = 32'b00000000000000010001101111001100;
assign LUT_3[20523] = 32'b00000000000000011000011010101001;
assign LUT_3[20524] = 32'b00000000000000001100110101011110;
assign LUT_3[20525] = 32'b00000000000000010011100000111011;
assign LUT_3[20526] = 32'b00000000000000001110111101000010;
assign LUT_3[20527] = 32'b00000000000000010101101000011111;
assign LUT_3[20528] = 32'b00000000000000001101100001100101;
assign LUT_3[20529] = 32'b00000000000000010100001101000010;
assign LUT_3[20530] = 32'b00000000000000001111101001001001;
assign LUT_3[20531] = 32'b00000000000000010110010100100110;
assign LUT_3[20532] = 32'b00000000000000001010101111011011;
assign LUT_3[20533] = 32'b00000000000000010001011010111000;
assign LUT_3[20534] = 32'b00000000000000001100110110111111;
assign LUT_3[20535] = 32'b00000000000000010011100010011100;
assign LUT_3[20536] = 32'b00000000000000010010111010101011;
assign LUT_3[20537] = 32'b00000000000000011001100110001000;
assign LUT_3[20538] = 32'b00000000000000010101000010001111;
assign LUT_3[20539] = 32'b00000000000000011011101101101100;
assign LUT_3[20540] = 32'b00000000000000010000001000100001;
assign LUT_3[20541] = 32'b00000000000000010110110011111110;
assign LUT_3[20542] = 32'b00000000000000010010010000000101;
assign LUT_3[20543] = 32'b00000000000000011000111011100010;
assign LUT_3[20544] = 32'b00000000000000001000111000101101;
assign LUT_3[20545] = 32'b00000000000000001111100100001010;
assign LUT_3[20546] = 32'b00000000000000001011000000010001;
assign LUT_3[20547] = 32'b00000000000000010001101011101110;
assign LUT_3[20548] = 32'b00000000000000000110000110100011;
assign LUT_3[20549] = 32'b00000000000000001100110010000000;
assign LUT_3[20550] = 32'b00000000000000001000001110000111;
assign LUT_3[20551] = 32'b00000000000000001110111001100100;
assign LUT_3[20552] = 32'b00000000000000001110010001110011;
assign LUT_3[20553] = 32'b00000000000000010100111101010000;
assign LUT_3[20554] = 32'b00000000000000010000011001010111;
assign LUT_3[20555] = 32'b00000000000000010111000100110100;
assign LUT_3[20556] = 32'b00000000000000001011011111101001;
assign LUT_3[20557] = 32'b00000000000000010010001011000110;
assign LUT_3[20558] = 32'b00000000000000001101100111001101;
assign LUT_3[20559] = 32'b00000000000000010100010010101010;
assign LUT_3[20560] = 32'b00000000000000001100001011110000;
assign LUT_3[20561] = 32'b00000000000000010010110111001101;
assign LUT_3[20562] = 32'b00000000000000001110010011010100;
assign LUT_3[20563] = 32'b00000000000000010100111110110001;
assign LUT_3[20564] = 32'b00000000000000001001011001100110;
assign LUT_3[20565] = 32'b00000000000000010000000101000011;
assign LUT_3[20566] = 32'b00000000000000001011100001001010;
assign LUT_3[20567] = 32'b00000000000000010010001100100111;
assign LUT_3[20568] = 32'b00000000000000010001100100110110;
assign LUT_3[20569] = 32'b00000000000000011000010000010011;
assign LUT_3[20570] = 32'b00000000000000010011101100011010;
assign LUT_3[20571] = 32'b00000000000000011010010111110111;
assign LUT_3[20572] = 32'b00000000000000001110110010101100;
assign LUT_3[20573] = 32'b00000000000000010101011110001001;
assign LUT_3[20574] = 32'b00000000000000010000111010010000;
assign LUT_3[20575] = 32'b00000000000000010111100101101101;
assign LUT_3[20576] = 32'b00000000000000001010000111001101;
assign LUT_3[20577] = 32'b00000000000000010000110010101010;
assign LUT_3[20578] = 32'b00000000000000001100001110110001;
assign LUT_3[20579] = 32'b00000000000000010010111010001110;
assign LUT_3[20580] = 32'b00000000000000000111010101000011;
assign LUT_3[20581] = 32'b00000000000000001110000000100000;
assign LUT_3[20582] = 32'b00000000000000001001011100100111;
assign LUT_3[20583] = 32'b00000000000000010000001000000100;
assign LUT_3[20584] = 32'b00000000000000001111100000010011;
assign LUT_3[20585] = 32'b00000000000000010110001011110000;
assign LUT_3[20586] = 32'b00000000000000010001100111110111;
assign LUT_3[20587] = 32'b00000000000000011000010011010100;
assign LUT_3[20588] = 32'b00000000000000001100101110001001;
assign LUT_3[20589] = 32'b00000000000000010011011001100110;
assign LUT_3[20590] = 32'b00000000000000001110110101101101;
assign LUT_3[20591] = 32'b00000000000000010101100001001010;
assign LUT_3[20592] = 32'b00000000000000001101011010010000;
assign LUT_3[20593] = 32'b00000000000000010100000101101101;
assign LUT_3[20594] = 32'b00000000000000001111100001110100;
assign LUT_3[20595] = 32'b00000000000000010110001101010001;
assign LUT_3[20596] = 32'b00000000000000001010101000000110;
assign LUT_3[20597] = 32'b00000000000000010001010011100011;
assign LUT_3[20598] = 32'b00000000000000001100101111101010;
assign LUT_3[20599] = 32'b00000000000000010011011011000111;
assign LUT_3[20600] = 32'b00000000000000010010110011010110;
assign LUT_3[20601] = 32'b00000000000000011001011110110011;
assign LUT_3[20602] = 32'b00000000000000010100111010111010;
assign LUT_3[20603] = 32'b00000000000000011011100110010111;
assign LUT_3[20604] = 32'b00000000000000010000000001001100;
assign LUT_3[20605] = 32'b00000000000000010110101100101001;
assign LUT_3[20606] = 32'b00000000000000010010001000110000;
assign LUT_3[20607] = 32'b00000000000000011000110100001101;
assign LUT_3[20608] = 32'b00000000000000001011001011000000;
assign LUT_3[20609] = 32'b00000000000000010001110110011101;
assign LUT_3[20610] = 32'b00000000000000001101010010100100;
assign LUT_3[20611] = 32'b00000000000000010011111110000001;
assign LUT_3[20612] = 32'b00000000000000001000011000110110;
assign LUT_3[20613] = 32'b00000000000000001111000100010011;
assign LUT_3[20614] = 32'b00000000000000001010100000011010;
assign LUT_3[20615] = 32'b00000000000000010001001011110111;
assign LUT_3[20616] = 32'b00000000000000010000100100000110;
assign LUT_3[20617] = 32'b00000000000000010111001111100011;
assign LUT_3[20618] = 32'b00000000000000010010101011101010;
assign LUT_3[20619] = 32'b00000000000000011001010111000111;
assign LUT_3[20620] = 32'b00000000000000001101110001111100;
assign LUT_3[20621] = 32'b00000000000000010100011101011001;
assign LUT_3[20622] = 32'b00000000000000001111111001100000;
assign LUT_3[20623] = 32'b00000000000000010110100100111101;
assign LUT_3[20624] = 32'b00000000000000001110011110000011;
assign LUT_3[20625] = 32'b00000000000000010101001001100000;
assign LUT_3[20626] = 32'b00000000000000010000100101100111;
assign LUT_3[20627] = 32'b00000000000000010111010001000100;
assign LUT_3[20628] = 32'b00000000000000001011101011111001;
assign LUT_3[20629] = 32'b00000000000000010010010111010110;
assign LUT_3[20630] = 32'b00000000000000001101110011011101;
assign LUT_3[20631] = 32'b00000000000000010100011110111010;
assign LUT_3[20632] = 32'b00000000000000010011110111001001;
assign LUT_3[20633] = 32'b00000000000000011010100010100110;
assign LUT_3[20634] = 32'b00000000000000010101111110101101;
assign LUT_3[20635] = 32'b00000000000000011100101010001010;
assign LUT_3[20636] = 32'b00000000000000010001000100111111;
assign LUT_3[20637] = 32'b00000000000000010111110000011100;
assign LUT_3[20638] = 32'b00000000000000010011001100100011;
assign LUT_3[20639] = 32'b00000000000000011001111000000000;
assign LUT_3[20640] = 32'b00000000000000001100011001100000;
assign LUT_3[20641] = 32'b00000000000000010011000100111101;
assign LUT_3[20642] = 32'b00000000000000001110100001000100;
assign LUT_3[20643] = 32'b00000000000000010101001100100001;
assign LUT_3[20644] = 32'b00000000000000001001100111010110;
assign LUT_3[20645] = 32'b00000000000000010000010010110011;
assign LUT_3[20646] = 32'b00000000000000001011101110111010;
assign LUT_3[20647] = 32'b00000000000000010010011010010111;
assign LUT_3[20648] = 32'b00000000000000010001110010100110;
assign LUT_3[20649] = 32'b00000000000000011000011110000011;
assign LUT_3[20650] = 32'b00000000000000010011111010001010;
assign LUT_3[20651] = 32'b00000000000000011010100101100111;
assign LUT_3[20652] = 32'b00000000000000001111000000011100;
assign LUT_3[20653] = 32'b00000000000000010101101011111001;
assign LUT_3[20654] = 32'b00000000000000010001001000000000;
assign LUT_3[20655] = 32'b00000000000000010111110011011101;
assign LUT_3[20656] = 32'b00000000000000001111101100100011;
assign LUT_3[20657] = 32'b00000000000000010110011000000000;
assign LUT_3[20658] = 32'b00000000000000010001110100000111;
assign LUT_3[20659] = 32'b00000000000000011000011111100100;
assign LUT_3[20660] = 32'b00000000000000001100111010011001;
assign LUT_3[20661] = 32'b00000000000000010011100101110110;
assign LUT_3[20662] = 32'b00000000000000001111000001111101;
assign LUT_3[20663] = 32'b00000000000000010101101101011010;
assign LUT_3[20664] = 32'b00000000000000010101000101101001;
assign LUT_3[20665] = 32'b00000000000000011011110001000110;
assign LUT_3[20666] = 32'b00000000000000010111001101001101;
assign LUT_3[20667] = 32'b00000000000000011101111000101010;
assign LUT_3[20668] = 32'b00000000000000010010010011011111;
assign LUT_3[20669] = 32'b00000000000000011000111110111100;
assign LUT_3[20670] = 32'b00000000000000010100011011000011;
assign LUT_3[20671] = 32'b00000000000000011011000110100000;
assign LUT_3[20672] = 32'b00000000000000001011000011101011;
assign LUT_3[20673] = 32'b00000000000000010001101111001000;
assign LUT_3[20674] = 32'b00000000000000001101001011001111;
assign LUT_3[20675] = 32'b00000000000000010011110110101100;
assign LUT_3[20676] = 32'b00000000000000001000010001100001;
assign LUT_3[20677] = 32'b00000000000000001110111100111110;
assign LUT_3[20678] = 32'b00000000000000001010011001000101;
assign LUT_3[20679] = 32'b00000000000000010001000100100010;
assign LUT_3[20680] = 32'b00000000000000010000011100110001;
assign LUT_3[20681] = 32'b00000000000000010111001000001110;
assign LUT_3[20682] = 32'b00000000000000010010100100010101;
assign LUT_3[20683] = 32'b00000000000000011001001111110010;
assign LUT_3[20684] = 32'b00000000000000001101101010100111;
assign LUT_3[20685] = 32'b00000000000000010100010110000100;
assign LUT_3[20686] = 32'b00000000000000001111110010001011;
assign LUT_3[20687] = 32'b00000000000000010110011101101000;
assign LUT_3[20688] = 32'b00000000000000001110010110101110;
assign LUT_3[20689] = 32'b00000000000000010101000010001011;
assign LUT_3[20690] = 32'b00000000000000010000011110010010;
assign LUT_3[20691] = 32'b00000000000000010111001001101111;
assign LUT_3[20692] = 32'b00000000000000001011100100100100;
assign LUT_3[20693] = 32'b00000000000000010010010000000001;
assign LUT_3[20694] = 32'b00000000000000001101101100001000;
assign LUT_3[20695] = 32'b00000000000000010100010111100101;
assign LUT_3[20696] = 32'b00000000000000010011101111110100;
assign LUT_3[20697] = 32'b00000000000000011010011011010001;
assign LUT_3[20698] = 32'b00000000000000010101110111011000;
assign LUT_3[20699] = 32'b00000000000000011100100010110101;
assign LUT_3[20700] = 32'b00000000000000010000111101101010;
assign LUT_3[20701] = 32'b00000000000000010111101001000111;
assign LUT_3[20702] = 32'b00000000000000010011000101001110;
assign LUT_3[20703] = 32'b00000000000000011001110000101011;
assign LUT_3[20704] = 32'b00000000000000001100010010001011;
assign LUT_3[20705] = 32'b00000000000000010010111101101000;
assign LUT_3[20706] = 32'b00000000000000001110011001101111;
assign LUT_3[20707] = 32'b00000000000000010101000101001100;
assign LUT_3[20708] = 32'b00000000000000001001100000000001;
assign LUT_3[20709] = 32'b00000000000000010000001011011110;
assign LUT_3[20710] = 32'b00000000000000001011100111100101;
assign LUT_3[20711] = 32'b00000000000000010010010011000010;
assign LUT_3[20712] = 32'b00000000000000010001101011010001;
assign LUT_3[20713] = 32'b00000000000000011000010110101110;
assign LUT_3[20714] = 32'b00000000000000010011110010110101;
assign LUT_3[20715] = 32'b00000000000000011010011110010010;
assign LUT_3[20716] = 32'b00000000000000001110111001000111;
assign LUT_3[20717] = 32'b00000000000000010101100100100100;
assign LUT_3[20718] = 32'b00000000000000010001000000101011;
assign LUT_3[20719] = 32'b00000000000000010111101100001000;
assign LUT_3[20720] = 32'b00000000000000001111100101001110;
assign LUT_3[20721] = 32'b00000000000000010110010000101011;
assign LUT_3[20722] = 32'b00000000000000010001101100110010;
assign LUT_3[20723] = 32'b00000000000000011000011000001111;
assign LUT_3[20724] = 32'b00000000000000001100110011000100;
assign LUT_3[20725] = 32'b00000000000000010011011110100001;
assign LUT_3[20726] = 32'b00000000000000001110111010101000;
assign LUT_3[20727] = 32'b00000000000000010101100110000101;
assign LUT_3[20728] = 32'b00000000000000010100111110010100;
assign LUT_3[20729] = 32'b00000000000000011011101001110001;
assign LUT_3[20730] = 32'b00000000000000010111000101111000;
assign LUT_3[20731] = 32'b00000000000000011101110001010101;
assign LUT_3[20732] = 32'b00000000000000010010001100001010;
assign LUT_3[20733] = 32'b00000000000000011000110111100111;
assign LUT_3[20734] = 32'b00000000000000010100010011101110;
assign LUT_3[20735] = 32'b00000000000000011010111111001011;
assign LUT_3[20736] = 32'b00000000000000000101001111100011;
assign LUT_3[20737] = 32'b00000000000000001011111011000000;
assign LUT_3[20738] = 32'b00000000000000000111010111000111;
assign LUT_3[20739] = 32'b00000000000000001110000010100100;
assign LUT_3[20740] = 32'b00000000000000000010011101011001;
assign LUT_3[20741] = 32'b00000000000000001001001000110110;
assign LUT_3[20742] = 32'b00000000000000000100100100111101;
assign LUT_3[20743] = 32'b00000000000000001011010000011010;
assign LUT_3[20744] = 32'b00000000000000001010101000101001;
assign LUT_3[20745] = 32'b00000000000000010001010100000110;
assign LUT_3[20746] = 32'b00000000000000001100110000001101;
assign LUT_3[20747] = 32'b00000000000000010011011011101010;
assign LUT_3[20748] = 32'b00000000000000000111110110011111;
assign LUT_3[20749] = 32'b00000000000000001110100001111100;
assign LUT_3[20750] = 32'b00000000000000001001111110000011;
assign LUT_3[20751] = 32'b00000000000000010000101001100000;
assign LUT_3[20752] = 32'b00000000000000001000100010100110;
assign LUT_3[20753] = 32'b00000000000000001111001110000011;
assign LUT_3[20754] = 32'b00000000000000001010101010001010;
assign LUT_3[20755] = 32'b00000000000000010001010101100111;
assign LUT_3[20756] = 32'b00000000000000000101110000011100;
assign LUT_3[20757] = 32'b00000000000000001100011011111001;
assign LUT_3[20758] = 32'b00000000000000000111111000000000;
assign LUT_3[20759] = 32'b00000000000000001110100011011101;
assign LUT_3[20760] = 32'b00000000000000001101111011101100;
assign LUT_3[20761] = 32'b00000000000000010100100111001001;
assign LUT_3[20762] = 32'b00000000000000010000000011010000;
assign LUT_3[20763] = 32'b00000000000000010110101110101101;
assign LUT_3[20764] = 32'b00000000000000001011001001100010;
assign LUT_3[20765] = 32'b00000000000000010001110100111111;
assign LUT_3[20766] = 32'b00000000000000001101010001000110;
assign LUT_3[20767] = 32'b00000000000000010011111100100011;
assign LUT_3[20768] = 32'b00000000000000000110011110000011;
assign LUT_3[20769] = 32'b00000000000000001101001001100000;
assign LUT_3[20770] = 32'b00000000000000001000100101100111;
assign LUT_3[20771] = 32'b00000000000000001111010001000100;
assign LUT_3[20772] = 32'b00000000000000000011101011111001;
assign LUT_3[20773] = 32'b00000000000000001010010111010110;
assign LUT_3[20774] = 32'b00000000000000000101110011011101;
assign LUT_3[20775] = 32'b00000000000000001100011110111010;
assign LUT_3[20776] = 32'b00000000000000001011110111001001;
assign LUT_3[20777] = 32'b00000000000000010010100010100110;
assign LUT_3[20778] = 32'b00000000000000001101111110101101;
assign LUT_3[20779] = 32'b00000000000000010100101010001010;
assign LUT_3[20780] = 32'b00000000000000001001000100111111;
assign LUT_3[20781] = 32'b00000000000000001111110000011100;
assign LUT_3[20782] = 32'b00000000000000001011001100100011;
assign LUT_3[20783] = 32'b00000000000000010001111000000000;
assign LUT_3[20784] = 32'b00000000000000001001110001000110;
assign LUT_3[20785] = 32'b00000000000000010000011100100011;
assign LUT_3[20786] = 32'b00000000000000001011111000101010;
assign LUT_3[20787] = 32'b00000000000000010010100100000111;
assign LUT_3[20788] = 32'b00000000000000000110111110111100;
assign LUT_3[20789] = 32'b00000000000000001101101010011001;
assign LUT_3[20790] = 32'b00000000000000001001000110100000;
assign LUT_3[20791] = 32'b00000000000000001111110001111101;
assign LUT_3[20792] = 32'b00000000000000001111001010001100;
assign LUT_3[20793] = 32'b00000000000000010101110101101001;
assign LUT_3[20794] = 32'b00000000000000010001010001110000;
assign LUT_3[20795] = 32'b00000000000000010111111101001101;
assign LUT_3[20796] = 32'b00000000000000001100011000000010;
assign LUT_3[20797] = 32'b00000000000000010011000011011111;
assign LUT_3[20798] = 32'b00000000000000001110011111100110;
assign LUT_3[20799] = 32'b00000000000000010101001011000011;
assign LUT_3[20800] = 32'b00000000000000000101001000001110;
assign LUT_3[20801] = 32'b00000000000000001011110011101011;
assign LUT_3[20802] = 32'b00000000000000000111001111110010;
assign LUT_3[20803] = 32'b00000000000000001101111011001111;
assign LUT_3[20804] = 32'b00000000000000000010010110000100;
assign LUT_3[20805] = 32'b00000000000000001001000001100001;
assign LUT_3[20806] = 32'b00000000000000000100011101101000;
assign LUT_3[20807] = 32'b00000000000000001011001001000101;
assign LUT_3[20808] = 32'b00000000000000001010100001010100;
assign LUT_3[20809] = 32'b00000000000000010001001100110001;
assign LUT_3[20810] = 32'b00000000000000001100101000111000;
assign LUT_3[20811] = 32'b00000000000000010011010100010101;
assign LUT_3[20812] = 32'b00000000000000000111101111001010;
assign LUT_3[20813] = 32'b00000000000000001110011010100111;
assign LUT_3[20814] = 32'b00000000000000001001110110101110;
assign LUT_3[20815] = 32'b00000000000000010000100010001011;
assign LUT_3[20816] = 32'b00000000000000001000011011010001;
assign LUT_3[20817] = 32'b00000000000000001111000110101110;
assign LUT_3[20818] = 32'b00000000000000001010100010110101;
assign LUT_3[20819] = 32'b00000000000000010001001110010010;
assign LUT_3[20820] = 32'b00000000000000000101101001000111;
assign LUT_3[20821] = 32'b00000000000000001100010100100100;
assign LUT_3[20822] = 32'b00000000000000000111110000101011;
assign LUT_3[20823] = 32'b00000000000000001110011100001000;
assign LUT_3[20824] = 32'b00000000000000001101110100010111;
assign LUT_3[20825] = 32'b00000000000000010100011111110100;
assign LUT_3[20826] = 32'b00000000000000001111111011111011;
assign LUT_3[20827] = 32'b00000000000000010110100111011000;
assign LUT_3[20828] = 32'b00000000000000001011000010001101;
assign LUT_3[20829] = 32'b00000000000000010001101101101010;
assign LUT_3[20830] = 32'b00000000000000001101001001110001;
assign LUT_3[20831] = 32'b00000000000000010011110101001110;
assign LUT_3[20832] = 32'b00000000000000000110010110101110;
assign LUT_3[20833] = 32'b00000000000000001101000010001011;
assign LUT_3[20834] = 32'b00000000000000001000011110010010;
assign LUT_3[20835] = 32'b00000000000000001111001001101111;
assign LUT_3[20836] = 32'b00000000000000000011100100100100;
assign LUT_3[20837] = 32'b00000000000000001010010000000001;
assign LUT_3[20838] = 32'b00000000000000000101101100001000;
assign LUT_3[20839] = 32'b00000000000000001100010111100101;
assign LUT_3[20840] = 32'b00000000000000001011101111110100;
assign LUT_3[20841] = 32'b00000000000000010010011011010001;
assign LUT_3[20842] = 32'b00000000000000001101110111011000;
assign LUT_3[20843] = 32'b00000000000000010100100010110101;
assign LUT_3[20844] = 32'b00000000000000001000111101101010;
assign LUT_3[20845] = 32'b00000000000000001111101001000111;
assign LUT_3[20846] = 32'b00000000000000001011000101001110;
assign LUT_3[20847] = 32'b00000000000000010001110000101011;
assign LUT_3[20848] = 32'b00000000000000001001101001110001;
assign LUT_3[20849] = 32'b00000000000000010000010101001110;
assign LUT_3[20850] = 32'b00000000000000001011110001010101;
assign LUT_3[20851] = 32'b00000000000000010010011100110010;
assign LUT_3[20852] = 32'b00000000000000000110110111100111;
assign LUT_3[20853] = 32'b00000000000000001101100011000100;
assign LUT_3[20854] = 32'b00000000000000001000111111001011;
assign LUT_3[20855] = 32'b00000000000000001111101010101000;
assign LUT_3[20856] = 32'b00000000000000001111000010110111;
assign LUT_3[20857] = 32'b00000000000000010101101110010100;
assign LUT_3[20858] = 32'b00000000000000010001001010011011;
assign LUT_3[20859] = 32'b00000000000000010111110101111000;
assign LUT_3[20860] = 32'b00000000000000001100010000101101;
assign LUT_3[20861] = 32'b00000000000000010010111100001010;
assign LUT_3[20862] = 32'b00000000000000001110011000010001;
assign LUT_3[20863] = 32'b00000000000000010101000011101110;
assign LUT_3[20864] = 32'b00000000000000000111011010100001;
assign LUT_3[20865] = 32'b00000000000000001110000101111110;
assign LUT_3[20866] = 32'b00000000000000001001100010000101;
assign LUT_3[20867] = 32'b00000000000000010000001101100010;
assign LUT_3[20868] = 32'b00000000000000000100101000010111;
assign LUT_3[20869] = 32'b00000000000000001011010011110100;
assign LUT_3[20870] = 32'b00000000000000000110101111111011;
assign LUT_3[20871] = 32'b00000000000000001101011011011000;
assign LUT_3[20872] = 32'b00000000000000001100110011100111;
assign LUT_3[20873] = 32'b00000000000000010011011111000100;
assign LUT_3[20874] = 32'b00000000000000001110111011001011;
assign LUT_3[20875] = 32'b00000000000000010101100110101000;
assign LUT_3[20876] = 32'b00000000000000001010000001011101;
assign LUT_3[20877] = 32'b00000000000000010000101100111010;
assign LUT_3[20878] = 32'b00000000000000001100001001000001;
assign LUT_3[20879] = 32'b00000000000000010010110100011110;
assign LUT_3[20880] = 32'b00000000000000001010101101100100;
assign LUT_3[20881] = 32'b00000000000000010001011001000001;
assign LUT_3[20882] = 32'b00000000000000001100110101001000;
assign LUT_3[20883] = 32'b00000000000000010011100000100101;
assign LUT_3[20884] = 32'b00000000000000000111111011011010;
assign LUT_3[20885] = 32'b00000000000000001110100110110111;
assign LUT_3[20886] = 32'b00000000000000001010000010111110;
assign LUT_3[20887] = 32'b00000000000000010000101110011011;
assign LUT_3[20888] = 32'b00000000000000010000000110101010;
assign LUT_3[20889] = 32'b00000000000000010110110010000111;
assign LUT_3[20890] = 32'b00000000000000010010001110001110;
assign LUT_3[20891] = 32'b00000000000000011000111001101011;
assign LUT_3[20892] = 32'b00000000000000001101010100100000;
assign LUT_3[20893] = 32'b00000000000000010011111111111101;
assign LUT_3[20894] = 32'b00000000000000001111011100000100;
assign LUT_3[20895] = 32'b00000000000000010110000111100001;
assign LUT_3[20896] = 32'b00000000000000001000101001000001;
assign LUT_3[20897] = 32'b00000000000000001111010100011110;
assign LUT_3[20898] = 32'b00000000000000001010110000100101;
assign LUT_3[20899] = 32'b00000000000000010001011100000010;
assign LUT_3[20900] = 32'b00000000000000000101110110110111;
assign LUT_3[20901] = 32'b00000000000000001100100010010100;
assign LUT_3[20902] = 32'b00000000000000000111111110011011;
assign LUT_3[20903] = 32'b00000000000000001110101001111000;
assign LUT_3[20904] = 32'b00000000000000001110000010000111;
assign LUT_3[20905] = 32'b00000000000000010100101101100100;
assign LUT_3[20906] = 32'b00000000000000010000001001101011;
assign LUT_3[20907] = 32'b00000000000000010110110101001000;
assign LUT_3[20908] = 32'b00000000000000001011001111111101;
assign LUT_3[20909] = 32'b00000000000000010001111011011010;
assign LUT_3[20910] = 32'b00000000000000001101010111100001;
assign LUT_3[20911] = 32'b00000000000000010100000010111110;
assign LUT_3[20912] = 32'b00000000000000001011111100000100;
assign LUT_3[20913] = 32'b00000000000000010010100111100001;
assign LUT_3[20914] = 32'b00000000000000001110000011101000;
assign LUT_3[20915] = 32'b00000000000000010100101111000101;
assign LUT_3[20916] = 32'b00000000000000001001001001111010;
assign LUT_3[20917] = 32'b00000000000000001111110101010111;
assign LUT_3[20918] = 32'b00000000000000001011010001011110;
assign LUT_3[20919] = 32'b00000000000000010001111100111011;
assign LUT_3[20920] = 32'b00000000000000010001010101001010;
assign LUT_3[20921] = 32'b00000000000000011000000000100111;
assign LUT_3[20922] = 32'b00000000000000010011011100101110;
assign LUT_3[20923] = 32'b00000000000000011010001000001011;
assign LUT_3[20924] = 32'b00000000000000001110100011000000;
assign LUT_3[20925] = 32'b00000000000000010101001110011101;
assign LUT_3[20926] = 32'b00000000000000010000101010100100;
assign LUT_3[20927] = 32'b00000000000000010111010110000001;
assign LUT_3[20928] = 32'b00000000000000000111010011001100;
assign LUT_3[20929] = 32'b00000000000000001101111110101001;
assign LUT_3[20930] = 32'b00000000000000001001011010110000;
assign LUT_3[20931] = 32'b00000000000000010000000110001101;
assign LUT_3[20932] = 32'b00000000000000000100100001000010;
assign LUT_3[20933] = 32'b00000000000000001011001100011111;
assign LUT_3[20934] = 32'b00000000000000000110101000100110;
assign LUT_3[20935] = 32'b00000000000000001101010100000011;
assign LUT_3[20936] = 32'b00000000000000001100101100010010;
assign LUT_3[20937] = 32'b00000000000000010011010111101111;
assign LUT_3[20938] = 32'b00000000000000001110110011110110;
assign LUT_3[20939] = 32'b00000000000000010101011111010011;
assign LUT_3[20940] = 32'b00000000000000001001111010001000;
assign LUT_3[20941] = 32'b00000000000000010000100101100101;
assign LUT_3[20942] = 32'b00000000000000001100000001101100;
assign LUT_3[20943] = 32'b00000000000000010010101101001001;
assign LUT_3[20944] = 32'b00000000000000001010100110001111;
assign LUT_3[20945] = 32'b00000000000000010001010001101100;
assign LUT_3[20946] = 32'b00000000000000001100101101110011;
assign LUT_3[20947] = 32'b00000000000000010011011001010000;
assign LUT_3[20948] = 32'b00000000000000000111110100000101;
assign LUT_3[20949] = 32'b00000000000000001110011111100010;
assign LUT_3[20950] = 32'b00000000000000001001111011101001;
assign LUT_3[20951] = 32'b00000000000000010000100111000110;
assign LUT_3[20952] = 32'b00000000000000001111111111010101;
assign LUT_3[20953] = 32'b00000000000000010110101010110010;
assign LUT_3[20954] = 32'b00000000000000010010000110111001;
assign LUT_3[20955] = 32'b00000000000000011000110010010110;
assign LUT_3[20956] = 32'b00000000000000001101001101001011;
assign LUT_3[20957] = 32'b00000000000000010011111000101000;
assign LUT_3[20958] = 32'b00000000000000001111010100101111;
assign LUT_3[20959] = 32'b00000000000000010110000000001100;
assign LUT_3[20960] = 32'b00000000000000001000100001101100;
assign LUT_3[20961] = 32'b00000000000000001111001101001001;
assign LUT_3[20962] = 32'b00000000000000001010101001010000;
assign LUT_3[20963] = 32'b00000000000000010001010100101101;
assign LUT_3[20964] = 32'b00000000000000000101101111100010;
assign LUT_3[20965] = 32'b00000000000000001100011010111111;
assign LUT_3[20966] = 32'b00000000000000000111110111000110;
assign LUT_3[20967] = 32'b00000000000000001110100010100011;
assign LUT_3[20968] = 32'b00000000000000001101111010110010;
assign LUT_3[20969] = 32'b00000000000000010100100110001111;
assign LUT_3[20970] = 32'b00000000000000010000000010010110;
assign LUT_3[20971] = 32'b00000000000000010110101101110011;
assign LUT_3[20972] = 32'b00000000000000001011001000101000;
assign LUT_3[20973] = 32'b00000000000000010001110100000101;
assign LUT_3[20974] = 32'b00000000000000001101010000001100;
assign LUT_3[20975] = 32'b00000000000000010011111011101001;
assign LUT_3[20976] = 32'b00000000000000001011110100101111;
assign LUT_3[20977] = 32'b00000000000000010010100000001100;
assign LUT_3[20978] = 32'b00000000000000001101111100010011;
assign LUT_3[20979] = 32'b00000000000000010100100111110000;
assign LUT_3[20980] = 32'b00000000000000001001000010100101;
assign LUT_3[20981] = 32'b00000000000000001111101110000010;
assign LUT_3[20982] = 32'b00000000000000001011001010001001;
assign LUT_3[20983] = 32'b00000000000000010001110101100110;
assign LUT_3[20984] = 32'b00000000000000010001001101110101;
assign LUT_3[20985] = 32'b00000000000000010111111001010010;
assign LUT_3[20986] = 32'b00000000000000010011010101011001;
assign LUT_3[20987] = 32'b00000000000000011010000000110110;
assign LUT_3[20988] = 32'b00000000000000001110011011101011;
assign LUT_3[20989] = 32'b00000000000000010101000111001000;
assign LUT_3[20990] = 32'b00000000000000010000100011001111;
assign LUT_3[20991] = 32'b00000000000000010111001110101100;
assign LUT_3[20992] = 32'b00000000000000001100010101001110;
assign LUT_3[20993] = 32'b00000000000000010011000000101011;
assign LUT_3[20994] = 32'b00000000000000001110011100110010;
assign LUT_3[20995] = 32'b00000000000000010101001000001111;
assign LUT_3[20996] = 32'b00000000000000001001100011000100;
assign LUT_3[20997] = 32'b00000000000000010000001110100001;
assign LUT_3[20998] = 32'b00000000000000001011101010101000;
assign LUT_3[20999] = 32'b00000000000000010010010110000101;
assign LUT_3[21000] = 32'b00000000000000010001101110010100;
assign LUT_3[21001] = 32'b00000000000000011000011001110001;
assign LUT_3[21002] = 32'b00000000000000010011110101111000;
assign LUT_3[21003] = 32'b00000000000000011010100001010101;
assign LUT_3[21004] = 32'b00000000000000001110111100001010;
assign LUT_3[21005] = 32'b00000000000000010101100111100111;
assign LUT_3[21006] = 32'b00000000000000010001000011101110;
assign LUT_3[21007] = 32'b00000000000000010111101111001011;
assign LUT_3[21008] = 32'b00000000000000001111101000010001;
assign LUT_3[21009] = 32'b00000000000000010110010011101110;
assign LUT_3[21010] = 32'b00000000000000010001101111110101;
assign LUT_3[21011] = 32'b00000000000000011000011011010010;
assign LUT_3[21012] = 32'b00000000000000001100110110000111;
assign LUT_3[21013] = 32'b00000000000000010011100001100100;
assign LUT_3[21014] = 32'b00000000000000001110111101101011;
assign LUT_3[21015] = 32'b00000000000000010101101001001000;
assign LUT_3[21016] = 32'b00000000000000010101000001010111;
assign LUT_3[21017] = 32'b00000000000000011011101100110100;
assign LUT_3[21018] = 32'b00000000000000010111001000111011;
assign LUT_3[21019] = 32'b00000000000000011101110100011000;
assign LUT_3[21020] = 32'b00000000000000010010001111001101;
assign LUT_3[21021] = 32'b00000000000000011000111010101010;
assign LUT_3[21022] = 32'b00000000000000010100010110110001;
assign LUT_3[21023] = 32'b00000000000000011011000010001110;
assign LUT_3[21024] = 32'b00000000000000001101100011101110;
assign LUT_3[21025] = 32'b00000000000000010100001111001011;
assign LUT_3[21026] = 32'b00000000000000001111101011010010;
assign LUT_3[21027] = 32'b00000000000000010110010110101111;
assign LUT_3[21028] = 32'b00000000000000001010110001100100;
assign LUT_3[21029] = 32'b00000000000000010001011101000001;
assign LUT_3[21030] = 32'b00000000000000001100111001001000;
assign LUT_3[21031] = 32'b00000000000000010011100100100101;
assign LUT_3[21032] = 32'b00000000000000010010111100110100;
assign LUT_3[21033] = 32'b00000000000000011001101000010001;
assign LUT_3[21034] = 32'b00000000000000010101000100011000;
assign LUT_3[21035] = 32'b00000000000000011011101111110101;
assign LUT_3[21036] = 32'b00000000000000010000001010101010;
assign LUT_3[21037] = 32'b00000000000000010110110110000111;
assign LUT_3[21038] = 32'b00000000000000010010010010001110;
assign LUT_3[21039] = 32'b00000000000000011000111101101011;
assign LUT_3[21040] = 32'b00000000000000010000110110110001;
assign LUT_3[21041] = 32'b00000000000000010111100010001110;
assign LUT_3[21042] = 32'b00000000000000010010111110010101;
assign LUT_3[21043] = 32'b00000000000000011001101001110010;
assign LUT_3[21044] = 32'b00000000000000001110000100100111;
assign LUT_3[21045] = 32'b00000000000000010100110000000100;
assign LUT_3[21046] = 32'b00000000000000010000001100001011;
assign LUT_3[21047] = 32'b00000000000000010110110111101000;
assign LUT_3[21048] = 32'b00000000000000010110001111110111;
assign LUT_3[21049] = 32'b00000000000000011100111011010100;
assign LUT_3[21050] = 32'b00000000000000011000010111011011;
assign LUT_3[21051] = 32'b00000000000000011111000010111000;
assign LUT_3[21052] = 32'b00000000000000010011011101101101;
assign LUT_3[21053] = 32'b00000000000000011010001001001010;
assign LUT_3[21054] = 32'b00000000000000010101100101010001;
assign LUT_3[21055] = 32'b00000000000000011100010000101110;
assign LUT_3[21056] = 32'b00000000000000001100001101111001;
assign LUT_3[21057] = 32'b00000000000000010010111001010110;
assign LUT_3[21058] = 32'b00000000000000001110010101011101;
assign LUT_3[21059] = 32'b00000000000000010101000000111010;
assign LUT_3[21060] = 32'b00000000000000001001011011101111;
assign LUT_3[21061] = 32'b00000000000000010000000111001100;
assign LUT_3[21062] = 32'b00000000000000001011100011010011;
assign LUT_3[21063] = 32'b00000000000000010010001110110000;
assign LUT_3[21064] = 32'b00000000000000010001100110111111;
assign LUT_3[21065] = 32'b00000000000000011000010010011100;
assign LUT_3[21066] = 32'b00000000000000010011101110100011;
assign LUT_3[21067] = 32'b00000000000000011010011010000000;
assign LUT_3[21068] = 32'b00000000000000001110110100110101;
assign LUT_3[21069] = 32'b00000000000000010101100000010010;
assign LUT_3[21070] = 32'b00000000000000010000111100011001;
assign LUT_3[21071] = 32'b00000000000000010111100111110110;
assign LUT_3[21072] = 32'b00000000000000001111100000111100;
assign LUT_3[21073] = 32'b00000000000000010110001100011001;
assign LUT_3[21074] = 32'b00000000000000010001101000100000;
assign LUT_3[21075] = 32'b00000000000000011000010011111101;
assign LUT_3[21076] = 32'b00000000000000001100101110110010;
assign LUT_3[21077] = 32'b00000000000000010011011010001111;
assign LUT_3[21078] = 32'b00000000000000001110110110010110;
assign LUT_3[21079] = 32'b00000000000000010101100001110011;
assign LUT_3[21080] = 32'b00000000000000010100111010000010;
assign LUT_3[21081] = 32'b00000000000000011011100101011111;
assign LUT_3[21082] = 32'b00000000000000010111000001100110;
assign LUT_3[21083] = 32'b00000000000000011101101101000011;
assign LUT_3[21084] = 32'b00000000000000010010000111111000;
assign LUT_3[21085] = 32'b00000000000000011000110011010101;
assign LUT_3[21086] = 32'b00000000000000010100001111011100;
assign LUT_3[21087] = 32'b00000000000000011010111010111001;
assign LUT_3[21088] = 32'b00000000000000001101011100011001;
assign LUT_3[21089] = 32'b00000000000000010100000111110110;
assign LUT_3[21090] = 32'b00000000000000001111100011111101;
assign LUT_3[21091] = 32'b00000000000000010110001111011010;
assign LUT_3[21092] = 32'b00000000000000001010101010001111;
assign LUT_3[21093] = 32'b00000000000000010001010101101100;
assign LUT_3[21094] = 32'b00000000000000001100110001110011;
assign LUT_3[21095] = 32'b00000000000000010011011101010000;
assign LUT_3[21096] = 32'b00000000000000010010110101011111;
assign LUT_3[21097] = 32'b00000000000000011001100000111100;
assign LUT_3[21098] = 32'b00000000000000010100111101000011;
assign LUT_3[21099] = 32'b00000000000000011011101000100000;
assign LUT_3[21100] = 32'b00000000000000010000000011010101;
assign LUT_3[21101] = 32'b00000000000000010110101110110010;
assign LUT_3[21102] = 32'b00000000000000010010001010111001;
assign LUT_3[21103] = 32'b00000000000000011000110110010110;
assign LUT_3[21104] = 32'b00000000000000010000101111011100;
assign LUT_3[21105] = 32'b00000000000000010111011010111001;
assign LUT_3[21106] = 32'b00000000000000010010110111000000;
assign LUT_3[21107] = 32'b00000000000000011001100010011101;
assign LUT_3[21108] = 32'b00000000000000001101111101010010;
assign LUT_3[21109] = 32'b00000000000000010100101000101111;
assign LUT_3[21110] = 32'b00000000000000010000000100110110;
assign LUT_3[21111] = 32'b00000000000000010110110000010011;
assign LUT_3[21112] = 32'b00000000000000010110001000100010;
assign LUT_3[21113] = 32'b00000000000000011100110011111111;
assign LUT_3[21114] = 32'b00000000000000011000010000000110;
assign LUT_3[21115] = 32'b00000000000000011110111011100011;
assign LUT_3[21116] = 32'b00000000000000010011010110011000;
assign LUT_3[21117] = 32'b00000000000000011010000001110101;
assign LUT_3[21118] = 32'b00000000000000010101011101111100;
assign LUT_3[21119] = 32'b00000000000000011100001001011001;
assign LUT_3[21120] = 32'b00000000000000001110100000001100;
assign LUT_3[21121] = 32'b00000000000000010101001011101001;
assign LUT_3[21122] = 32'b00000000000000010000100111110000;
assign LUT_3[21123] = 32'b00000000000000010111010011001101;
assign LUT_3[21124] = 32'b00000000000000001011101110000010;
assign LUT_3[21125] = 32'b00000000000000010010011001011111;
assign LUT_3[21126] = 32'b00000000000000001101110101100110;
assign LUT_3[21127] = 32'b00000000000000010100100001000011;
assign LUT_3[21128] = 32'b00000000000000010011111001010010;
assign LUT_3[21129] = 32'b00000000000000011010100100101111;
assign LUT_3[21130] = 32'b00000000000000010110000000110110;
assign LUT_3[21131] = 32'b00000000000000011100101100010011;
assign LUT_3[21132] = 32'b00000000000000010001000111001000;
assign LUT_3[21133] = 32'b00000000000000010111110010100101;
assign LUT_3[21134] = 32'b00000000000000010011001110101100;
assign LUT_3[21135] = 32'b00000000000000011001111010001001;
assign LUT_3[21136] = 32'b00000000000000010001110011001111;
assign LUT_3[21137] = 32'b00000000000000011000011110101100;
assign LUT_3[21138] = 32'b00000000000000010011111010110011;
assign LUT_3[21139] = 32'b00000000000000011010100110010000;
assign LUT_3[21140] = 32'b00000000000000001111000001000101;
assign LUT_3[21141] = 32'b00000000000000010101101100100010;
assign LUT_3[21142] = 32'b00000000000000010001001000101001;
assign LUT_3[21143] = 32'b00000000000000010111110100000110;
assign LUT_3[21144] = 32'b00000000000000010111001100010101;
assign LUT_3[21145] = 32'b00000000000000011101110111110010;
assign LUT_3[21146] = 32'b00000000000000011001010011111001;
assign LUT_3[21147] = 32'b00000000000000011111111111010110;
assign LUT_3[21148] = 32'b00000000000000010100011010001011;
assign LUT_3[21149] = 32'b00000000000000011011000101101000;
assign LUT_3[21150] = 32'b00000000000000010110100001101111;
assign LUT_3[21151] = 32'b00000000000000011101001101001100;
assign LUT_3[21152] = 32'b00000000000000001111101110101100;
assign LUT_3[21153] = 32'b00000000000000010110011010001001;
assign LUT_3[21154] = 32'b00000000000000010001110110010000;
assign LUT_3[21155] = 32'b00000000000000011000100001101101;
assign LUT_3[21156] = 32'b00000000000000001100111100100010;
assign LUT_3[21157] = 32'b00000000000000010011100111111111;
assign LUT_3[21158] = 32'b00000000000000001111000100000110;
assign LUT_3[21159] = 32'b00000000000000010101101111100011;
assign LUT_3[21160] = 32'b00000000000000010101000111110010;
assign LUT_3[21161] = 32'b00000000000000011011110011001111;
assign LUT_3[21162] = 32'b00000000000000010111001111010110;
assign LUT_3[21163] = 32'b00000000000000011101111010110011;
assign LUT_3[21164] = 32'b00000000000000010010010101101000;
assign LUT_3[21165] = 32'b00000000000000011001000001000101;
assign LUT_3[21166] = 32'b00000000000000010100011101001100;
assign LUT_3[21167] = 32'b00000000000000011011001000101001;
assign LUT_3[21168] = 32'b00000000000000010011000001101111;
assign LUT_3[21169] = 32'b00000000000000011001101101001100;
assign LUT_3[21170] = 32'b00000000000000010101001001010011;
assign LUT_3[21171] = 32'b00000000000000011011110100110000;
assign LUT_3[21172] = 32'b00000000000000010000001111100101;
assign LUT_3[21173] = 32'b00000000000000010110111011000010;
assign LUT_3[21174] = 32'b00000000000000010010010111001001;
assign LUT_3[21175] = 32'b00000000000000011001000010100110;
assign LUT_3[21176] = 32'b00000000000000011000011010110101;
assign LUT_3[21177] = 32'b00000000000000011111000110010010;
assign LUT_3[21178] = 32'b00000000000000011010100010011001;
assign LUT_3[21179] = 32'b00000000000000100001001101110110;
assign LUT_3[21180] = 32'b00000000000000010101101000101011;
assign LUT_3[21181] = 32'b00000000000000011100010100001000;
assign LUT_3[21182] = 32'b00000000000000010111110000001111;
assign LUT_3[21183] = 32'b00000000000000011110011011101100;
assign LUT_3[21184] = 32'b00000000000000001110011000110111;
assign LUT_3[21185] = 32'b00000000000000010101000100010100;
assign LUT_3[21186] = 32'b00000000000000010000100000011011;
assign LUT_3[21187] = 32'b00000000000000010111001011111000;
assign LUT_3[21188] = 32'b00000000000000001011100110101101;
assign LUT_3[21189] = 32'b00000000000000010010010010001010;
assign LUT_3[21190] = 32'b00000000000000001101101110010001;
assign LUT_3[21191] = 32'b00000000000000010100011001101110;
assign LUT_3[21192] = 32'b00000000000000010011110001111101;
assign LUT_3[21193] = 32'b00000000000000011010011101011010;
assign LUT_3[21194] = 32'b00000000000000010101111001100001;
assign LUT_3[21195] = 32'b00000000000000011100100100111110;
assign LUT_3[21196] = 32'b00000000000000010000111111110011;
assign LUT_3[21197] = 32'b00000000000000010111101011010000;
assign LUT_3[21198] = 32'b00000000000000010011000111010111;
assign LUT_3[21199] = 32'b00000000000000011001110010110100;
assign LUT_3[21200] = 32'b00000000000000010001101011111010;
assign LUT_3[21201] = 32'b00000000000000011000010111010111;
assign LUT_3[21202] = 32'b00000000000000010011110011011110;
assign LUT_3[21203] = 32'b00000000000000011010011110111011;
assign LUT_3[21204] = 32'b00000000000000001110111001110000;
assign LUT_3[21205] = 32'b00000000000000010101100101001101;
assign LUT_3[21206] = 32'b00000000000000010001000001010100;
assign LUT_3[21207] = 32'b00000000000000010111101100110001;
assign LUT_3[21208] = 32'b00000000000000010111000101000000;
assign LUT_3[21209] = 32'b00000000000000011101110000011101;
assign LUT_3[21210] = 32'b00000000000000011001001100100100;
assign LUT_3[21211] = 32'b00000000000000011111111000000001;
assign LUT_3[21212] = 32'b00000000000000010100010010110110;
assign LUT_3[21213] = 32'b00000000000000011010111110010011;
assign LUT_3[21214] = 32'b00000000000000010110011010011010;
assign LUT_3[21215] = 32'b00000000000000011101000101110111;
assign LUT_3[21216] = 32'b00000000000000001111100111010111;
assign LUT_3[21217] = 32'b00000000000000010110010010110100;
assign LUT_3[21218] = 32'b00000000000000010001101110111011;
assign LUT_3[21219] = 32'b00000000000000011000011010011000;
assign LUT_3[21220] = 32'b00000000000000001100110101001101;
assign LUT_3[21221] = 32'b00000000000000010011100000101010;
assign LUT_3[21222] = 32'b00000000000000001110111100110001;
assign LUT_3[21223] = 32'b00000000000000010101101000001110;
assign LUT_3[21224] = 32'b00000000000000010101000000011101;
assign LUT_3[21225] = 32'b00000000000000011011101011111010;
assign LUT_3[21226] = 32'b00000000000000010111001000000001;
assign LUT_3[21227] = 32'b00000000000000011101110011011110;
assign LUT_3[21228] = 32'b00000000000000010010001110010011;
assign LUT_3[21229] = 32'b00000000000000011000111001110000;
assign LUT_3[21230] = 32'b00000000000000010100010101110111;
assign LUT_3[21231] = 32'b00000000000000011011000001010100;
assign LUT_3[21232] = 32'b00000000000000010010111010011010;
assign LUT_3[21233] = 32'b00000000000000011001100101110111;
assign LUT_3[21234] = 32'b00000000000000010101000001111110;
assign LUT_3[21235] = 32'b00000000000000011011101101011011;
assign LUT_3[21236] = 32'b00000000000000010000001000010000;
assign LUT_3[21237] = 32'b00000000000000010110110011101101;
assign LUT_3[21238] = 32'b00000000000000010010001111110100;
assign LUT_3[21239] = 32'b00000000000000011000111011010001;
assign LUT_3[21240] = 32'b00000000000000011000010011100000;
assign LUT_3[21241] = 32'b00000000000000011110111110111101;
assign LUT_3[21242] = 32'b00000000000000011010011011000100;
assign LUT_3[21243] = 32'b00000000000000100001000110100001;
assign LUT_3[21244] = 32'b00000000000000010101100001010110;
assign LUT_3[21245] = 32'b00000000000000011100001100110011;
assign LUT_3[21246] = 32'b00000000000000010111101000111010;
assign LUT_3[21247] = 32'b00000000000000011110010100010111;
assign LUT_3[21248] = 32'b00000000000000001000100100101111;
assign LUT_3[21249] = 32'b00000000000000001111010000001100;
assign LUT_3[21250] = 32'b00000000000000001010101100010011;
assign LUT_3[21251] = 32'b00000000000000010001010111110000;
assign LUT_3[21252] = 32'b00000000000000000101110010100101;
assign LUT_3[21253] = 32'b00000000000000001100011110000010;
assign LUT_3[21254] = 32'b00000000000000000111111010001001;
assign LUT_3[21255] = 32'b00000000000000001110100101100110;
assign LUT_3[21256] = 32'b00000000000000001101111101110101;
assign LUT_3[21257] = 32'b00000000000000010100101001010010;
assign LUT_3[21258] = 32'b00000000000000010000000101011001;
assign LUT_3[21259] = 32'b00000000000000010110110000110110;
assign LUT_3[21260] = 32'b00000000000000001011001011101011;
assign LUT_3[21261] = 32'b00000000000000010001110111001000;
assign LUT_3[21262] = 32'b00000000000000001101010011001111;
assign LUT_3[21263] = 32'b00000000000000010011111110101100;
assign LUT_3[21264] = 32'b00000000000000001011110111110010;
assign LUT_3[21265] = 32'b00000000000000010010100011001111;
assign LUT_3[21266] = 32'b00000000000000001101111111010110;
assign LUT_3[21267] = 32'b00000000000000010100101010110011;
assign LUT_3[21268] = 32'b00000000000000001001000101101000;
assign LUT_3[21269] = 32'b00000000000000001111110001000101;
assign LUT_3[21270] = 32'b00000000000000001011001101001100;
assign LUT_3[21271] = 32'b00000000000000010001111000101001;
assign LUT_3[21272] = 32'b00000000000000010001010000111000;
assign LUT_3[21273] = 32'b00000000000000010111111100010101;
assign LUT_3[21274] = 32'b00000000000000010011011000011100;
assign LUT_3[21275] = 32'b00000000000000011010000011111001;
assign LUT_3[21276] = 32'b00000000000000001110011110101110;
assign LUT_3[21277] = 32'b00000000000000010101001010001011;
assign LUT_3[21278] = 32'b00000000000000010000100110010010;
assign LUT_3[21279] = 32'b00000000000000010111010001101111;
assign LUT_3[21280] = 32'b00000000000000001001110011001111;
assign LUT_3[21281] = 32'b00000000000000010000011110101100;
assign LUT_3[21282] = 32'b00000000000000001011111010110011;
assign LUT_3[21283] = 32'b00000000000000010010100110010000;
assign LUT_3[21284] = 32'b00000000000000000111000001000101;
assign LUT_3[21285] = 32'b00000000000000001101101100100010;
assign LUT_3[21286] = 32'b00000000000000001001001000101001;
assign LUT_3[21287] = 32'b00000000000000001111110100000110;
assign LUT_3[21288] = 32'b00000000000000001111001100010101;
assign LUT_3[21289] = 32'b00000000000000010101110111110010;
assign LUT_3[21290] = 32'b00000000000000010001010011111001;
assign LUT_3[21291] = 32'b00000000000000010111111111010110;
assign LUT_3[21292] = 32'b00000000000000001100011010001011;
assign LUT_3[21293] = 32'b00000000000000010011000101101000;
assign LUT_3[21294] = 32'b00000000000000001110100001101111;
assign LUT_3[21295] = 32'b00000000000000010101001101001100;
assign LUT_3[21296] = 32'b00000000000000001101000110010010;
assign LUT_3[21297] = 32'b00000000000000010011110001101111;
assign LUT_3[21298] = 32'b00000000000000001111001101110110;
assign LUT_3[21299] = 32'b00000000000000010101111001010011;
assign LUT_3[21300] = 32'b00000000000000001010010100001000;
assign LUT_3[21301] = 32'b00000000000000010000111111100101;
assign LUT_3[21302] = 32'b00000000000000001100011011101100;
assign LUT_3[21303] = 32'b00000000000000010011000111001001;
assign LUT_3[21304] = 32'b00000000000000010010011111011000;
assign LUT_3[21305] = 32'b00000000000000011001001010110101;
assign LUT_3[21306] = 32'b00000000000000010100100110111100;
assign LUT_3[21307] = 32'b00000000000000011011010010011001;
assign LUT_3[21308] = 32'b00000000000000001111101101001110;
assign LUT_3[21309] = 32'b00000000000000010110011000101011;
assign LUT_3[21310] = 32'b00000000000000010001110100110010;
assign LUT_3[21311] = 32'b00000000000000011000100000001111;
assign LUT_3[21312] = 32'b00000000000000001000011101011010;
assign LUT_3[21313] = 32'b00000000000000001111001000110111;
assign LUT_3[21314] = 32'b00000000000000001010100100111110;
assign LUT_3[21315] = 32'b00000000000000010001010000011011;
assign LUT_3[21316] = 32'b00000000000000000101101011010000;
assign LUT_3[21317] = 32'b00000000000000001100010110101101;
assign LUT_3[21318] = 32'b00000000000000000111110010110100;
assign LUT_3[21319] = 32'b00000000000000001110011110010001;
assign LUT_3[21320] = 32'b00000000000000001101110110100000;
assign LUT_3[21321] = 32'b00000000000000010100100001111101;
assign LUT_3[21322] = 32'b00000000000000001111111110000100;
assign LUT_3[21323] = 32'b00000000000000010110101001100001;
assign LUT_3[21324] = 32'b00000000000000001011000100010110;
assign LUT_3[21325] = 32'b00000000000000010001101111110011;
assign LUT_3[21326] = 32'b00000000000000001101001011111010;
assign LUT_3[21327] = 32'b00000000000000010011110111010111;
assign LUT_3[21328] = 32'b00000000000000001011110000011101;
assign LUT_3[21329] = 32'b00000000000000010010011011111010;
assign LUT_3[21330] = 32'b00000000000000001101111000000001;
assign LUT_3[21331] = 32'b00000000000000010100100011011110;
assign LUT_3[21332] = 32'b00000000000000001000111110010011;
assign LUT_3[21333] = 32'b00000000000000001111101001110000;
assign LUT_3[21334] = 32'b00000000000000001011000101110111;
assign LUT_3[21335] = 32'b00000000000000010001110001010100;
assign LUT_3[21336] = 32'b00000000000000010001001001100011;
assign LUT_3[21337] = 32'b00000000000000010111110101000000;
assign LUT_3[21338] = 32'b00000000000000010011010001000111;
assign LUT_3[21339] = 32'b00000000000000011001111100100100;
assign LUT_3[21340] = 32'b00000000000000001110010111011001;
assign LUT_3[21341] = 32'b00000000000000010101000010110110;
assign LUT_3[21342] = 32'b00000000000000010000011110111101;
assign LUT_3[21343] = 32'b00000000000000010111001010011010;
assign LUT_3[21344] = 32'b00000000000000001001101011111010;
assign LUT_3[21345] = 32'b00000000000000010000010111010111;
assign LUT_3[21346] = 32'b00000000000000001011110011011110;
assign LUT_3[21347] = 32'b00000000000000010010011110111011;
assign LUT_3[21348] = 32'b00000000000000000110111001110000;
assign LUT_3[21349] = 32'b00000000000000001101100101001101;
assign LUT_3[21350] = 32'b00000000000000001001000001010100;
assign LUT_3[21351] = 32'b00000000000000001111101100110001;
assign LUT_3[21352] = 32'b00000000000000001111000101000000;
assign LUT_3[21353] = 32'b00000000000000010101110000011101;
assign LUT_3[21354] = 32'b00000000000000010001001100100100;
assign LUT_3[21355] = 32'b00000000000000010111111000000001;
assign LUT_3[21356] = 32'b00000000000000001100010010110110;
assign LUT_3[21357] = 32'b00000000000000010010111110010011;
assign LUT_3[21358] = 32'b00000000000000001110011010011010;
assign LUT_3[21359] = 32'b00000000000000010101000101110111;
assign LUT_3[21360] = 32'b00000000000000001100111110111101;
assign LUT_3[21361] = 32'b00000000000000010011101010011010;
assign LUT_3[21362] = 32'b00000000000000001111000110100001;
assign LUT_3[21363] = 32'b00000000000000010101110001111110;
assign LUT_3[21364] = 32'b00000000000000001010001100110011;
assign LUT_3[21365] = 32'b00000000000000010000111000010000;
assign LUT_3[21366] = 32'b00000000000000001100010100010111;
assign LUT_3[21367] = 32'b00000000000000010010111111110100;
assign LUT_3[21368] = 32'b00000000000000010010011000000011;
assign LUT_3[21369] = 32'b00000000000000011001000011100000;
assign LUT_3[21370] = 32'b00000000000000010100011111100111;
assign LUT_3[21371] = 32'b00000000000000011011001011000100;
assign LUT_3[21372] = 32'b00000000000000001111100101111001;
assign LUT_3[21373] = 32'b00000000000000010110010001010110;
assign LUT_3[21374] = 32'b00000000000000010001101101011101;
assign LUT_3[21375] = 32'b00000000000000011000011000111010;
assign LUT_3[21376] = 32'b00000000000000001010101111101101;
assign LUT_3[21377] = 32'b00000000000000010001011011001010;
assign LUT_3[21378] = 32'b00000000000000001100110111010001;
assign LUT_3[21379] = 32'b00000000000000010011100010101110;
assign LUT_3[21380] = 32'b00000000000000000111111101100011;
assign LUT_3[21381] = 32'b00000000000000001110101001000000;
assign LUT_3[21382] = 32'b00000000000000001010000101000111;
assign LUT_3[21383] = 32'b00000000000000010000110000100100;
assign LUT_3[21384] = 32'b00000000000000010000001000110011;
assign LUT_3[21385] = 32'b00000000000000010110110100010000;
assign LUT_3[21386] = 32'b00000000000000010010010000010111;
assign LUT_3[21387] = 32'b00000000000000011000111011110100;
assign LUT_3[21388] = 32'b00000000000000001101010110101001;
assign LUT_3[21389] = 32'b00000000000000010100000010000110;
assign LUT_3[21390] = 32'b00000000000000001111011110001101;
assign LUT_3[21391] = 32'b00000000000000010110001001101010;
assign LUT_3[21392] = 32'b00000000000000001110000010110000;
assign LUT_3[21393] = 32'b00000000000000010100101110001101;
assign LUT_3[21394] = 32'b00000000000000010000001010010100;
assign LUT_3[21395] = 32'b00000000000000010110110101110001;
assign LUT_3[21396] = 32'b00000000000000001011010000100110;
assign LUT_3[21397] = 32'b00000000000000010001111100000011;
assign LUT_3[21398] = 32'b00000000000000001101011000001010;
assign LUT_3[21399] = 32'b00000000000000010100000011100111;
assign LUT_3[21400] = 32'b00000000000000010011011011110110;
assign LUT_3[21401] = 32'b00000000000000011010000111010011;
assign LUT_3[21402] = 32'b00000000000000010101100011011010;
assign LUT_3[21403] = 32'b00000000000000011100001110110111;
assign LUT_3[21404] = 32'b00000000000000010000101001101100;
assign LUT_3[21405] = 32'b00000000000000010111010101001001;
assign LUT_3[21406] = 32'b00000000000000010010110001010000;
assign LUT_3[21407] = 32'b00000000000000011001011100101101;
assign LUT_3[21408] = 32'b00000000000000001011111110001101;
assign LUT_3[21409] = 32'b00000000000000010010101001101010;
assign LUT_3[21410] = 32'b00000000000000001110000101110001;
assign LUT_3[21411] = 32'b00000000000000010100110001001110;
assign LUT_3[21412] = 32'b00000000000000001001001100000011;
assign LUT_3[21413] = 32'b00000000000000001111110111100000;
assign LUT_3[21414] = 32'b00000000000000001011010011100111;
assign LUT_3[21415] = 32'b00000000000000010001111111000100;
assign LUT_3[21416] = 32'b00000000000000010001010111010011;
assign LUT_3[21417] = 32'b00000000000000011000000010110000;
assign LUT_3[21418] = 32'b00000000000000010011011110110111;
assign LUT_3[21419] = 32'b00000000000000011010001010010100;
assign LUT_3[21420] = 32'b00000000000000001110100101001001;
assign LUT_3[21421] = 32'b00000000000000010101010000100110;
assign LUT_3[21422] = 32'b00000000000000010000101100101101;
assign LUT_3[21423] = 32'b00000000000000010111011000001010;
assign LUT_3[21424] = 32'b00000000000000001111010001010000;
assign LUT_3[21425] = 32'b00000000000000010101111100101101;
assign LUT_3[21426] = 32'b00000000000000010001011000110100;
assign LUT_3[21427] = 32'b00000000000000011000000100010001;
assign LUT_3[21428] = 32'b00000000000000001100011111000110;
assign LUT_3[21429] = 32'b00000000000000010011001010100011;
assign LUT_3[21430] = 32'b00000000000000001110100110101010;
assign LUT_3[21431] = 32'b00000000000000010101010010000111;
assign LUT_3[21432] = 32'b00000000000000010100101010010110;
assign LUT_3[21433] = 32'b00000000000000011011010101110011;
assign LUT_3[21434] = 32'b00000000000000010110110001111010;
assign LUT_3[21435] = 32'b00000000000000011101011101010111;
assign LUT_3[21436] = 32'b00000000000000010001111000001100;
assign LUT_3[21437] = 32'b00000000000000011000100011101001;
assign LUT_3[21438] = 32'b00000000000000010011111111110000;
assign LUT_3[21439] = 32'b00000000000000011010101011001101;
assign LUT_3[21440] = 32'b00000000000000001010101000011000;
assign LUT_3[21441] = 32'b00000000000000010001010011110101;
assign LUT_3[21442] = 32'b00000000000000001100101111111100;
assign LUT_3[21443] = 32'b00000000000000010011011011011001;
assign LUT_3[21444] = 32'b00000000000000000111110110001110;
assign LUT_3[21445] = 32'b00000000000000001110100001101011;
assign LUT_3[21446] = 32'b00000000000000001001111101110010;
assign LUT_3[21447] = 32'b00000000000000010000101001001111;
assign LUT_3[21448] = 32'b00000000000000010000000001011110;
assign LUT_3[21449] = 32'b00000000000000010110101100111011;
assign LUT_3[21450] = 32'b00000000000000010010001001000010;
assign LUT_3[21451] = 32'b00000000000000011000110100011111;
assign LUT_3[21452] = 32'b00000000000000001101001111010100;
assign LUT_3[21453] = 32'b00000000000000010011111010110001;
assign LUT_3[21454] = 32'b00000000000000001111010110111000;
assign LUT_3[21455] = 32'b00000000000000010110000010010101;
assign LUT_3[21456] = 32'b00000000000000001101111011011011;
assign LUT_3[21457] = 32'b00000000000000010100100110111000;
assign LUT_3[21458] = 32'b00000000000000010000000010111111;
assign LUT_3[21459] = 32'b00000000000000010110101110011100;
assign LUT_3[21460] = 32'b00000000000000001011001001010001;
assign LUT_3[21461] = 32'b00000000000000010001110100101110;
assign LUT_3[21462] = 32'b00000000000000001101010000110101;
assign LUT_3[21463] = 32'b00000000000000010011111100010010;
assign LUT_3[21464] = 32'b00000000000000010011010100100001;
assign LUT_3[21465] = 32'b00000000000000011001111111111110;
assign LUT_3[21466] = 32'b00000000000000010101011100000101;
assign LUT_3[21467] = 32'b00000000000000011100000111100010;
assign LUT_3[21468] = 32'b00000000000000010000100010010111;
assign LUT_3[21469] = 32'b00000000000000010111001101110100;
assign LUT_3[21470] = 32'b00000000000000010010101001111011;
assign LUT_3[21471] = 32'b00000000000000011001010101011000;
assign LUT_3[21472] = 32'b00000000000000001011110110111000;
assign LUT_3[21473] = 32'b00000000000000010010100010010101;
assign LUT_3[21474] = 32'b00000000000000001101111110011100;
assign LUT_3[21475] = 32'b00000000000000010100101001111001;
assign LUT_3[21476] = 32'b00000000000000001001000100101110;
assign LUT_3[21477] = 32'b00000000000000001111110000001011;
assign LUT_3[21478] = 32'b00000000000000001011001100010010;
assign LUT_3[21479] = 32'b00000000000000010001110111101111;
assign LUT_3[21480] = 32'b00000000000000010001001111111110;
assign LUT_3[21481] = 32'b00000000000000010111111011011011;
assign LUT_3[21482] = 32'b00000000000000010011010111100010;
assign LUT_3[21483] = 32'b00000000000000011010000010111111;
assign LUT_3[21484] = 32'b00000000000000001110011101110100;
assign LUT_3[21485] = 32'b00000000000000010101001001010001;
assign LUT_3[21486] = 32'b00000000000000010000100101011000;
assign LUT_3[21487] = 32'b00000000000000010111010000110101;
assign LUT_3[21488] = 32'b00000000000000001111001001111011;
assign LUT_3[21489] = 32'b00000000000000010101110101011000;
assign LUT_3[21490] = 32'b00000000000000010001010001011111;
assign LUT_3[21491] = 32'b00000000000000010111111100111100;
assign LUT_3[21492] = 32'b00000000000000001100010111110001;
assign LUT_3[21493] = 32'b00000000000000010011000011001110;
assign LUT_3[21494] = 32'b00000000000000001110011111010101;
assign LUT_3[21495] = 32'b00000000000000010101001010110010;
assign LUT_3[21496] = 32'b00000000000000010100100011000001;
assign LUT_3[21497] = 32'b00000000000000011011001110011110;
assign LUT_3[21498] = 32'b00000000000000010110101010100101;
assign LUT_3[21499] = 32'b00000000000000011101010110000010;
assign LUT_3[21500] = 32'b00000000000000010001110000110111;
assign LUT_3[21501] = 32'b00000000000000011000011100010100;
assign LUT_3[21502] = 32'b00000000000000010011111000011011;
assign LUT_3[21503] = 32'b00000000000000011010100011111000;
assign LUT_3[21504] = 32'b00000000000000001111100100111111;
assign LUT_3[21505] = 32'b00000000000000010110010000011100;
assign LUT_3[21506] = 32'b00000000000000010001101100100011;
assign LUT_3[21507] = 32'b00000000000000011000011000000000;
assign LUT_3[21508] = 32'b00000000000000001100110010110101;
assign LUT_3[21509] = 32'b00000000000000010011011110010010;
assign LUT_3[21510] = 32'b00000000000000001110111010011001;
assign LUT_3[21511] = 32'b00000000000000010101100101110110;
assign LUT_3[21512] = 32'b00000000000000010100111110000101;
assign LUT_3[21513] = 32'b00000000000000011011101001100010;
assign LUT_3[21514] = 32'b00000000000000010111000101101001;
assign LUT_3[21515] = 32'b00000000000000011101110001000110;
assign LUT_3[21516] = 32'b00000000000000010010001011111011;
assign LUT_3[21517] = 32'b00000000000000011000110111011000;
assign LUT_3[21518] = 32'b00000000000000010100010011011111;
assign LUT_3[21519] = 32'b00000000000000011010111110111100;
assign LUT_3[21520] = 32'b00000000000000010010111000000010;
assign LUT_3[21521] = 32'b00000000000000011001100011011111;
assign LUT_3[21522] = 32'b00000000000000010100111111100110;
assign LUT_3[21523] = 32'b00000000000000011011101011000011;
assign LUT_3[21524] = 32'b00000000000000010000000101111000;
assign LUT_3[21525] = 32'b00000000000000010110110001010101;
assign LUT_3[21526] = 32'b00000000000000010010001101011100;
assign LUT_3[21527] = 32'b00000000000000011000111000111001;
assign LUT_3[21528] = 32'b00000000000000011000010001001000;
assign LUT_3[21529] = 32'b00000000000000011110111100100101;
assign LUT_3[21530] = 32'b00000000000000011010011000101100;
assign LUT_3[21531] = 32'b00000000000000100001000100001001;
assign LUT_3[21532] = 32'b00000000000000010101011110111110;
assign LUT_3[21533] = 32'b00000000000000011100001010011011;
assign LUT_3[21534] = 32'b00000000000000010111100110100010;
assign LUT_3[21535] = 32'b00000000000000011110010001111111;
assign LUT_3[21536] = 32'b00000000000000010000110011011111;
assign LUT_3[21537] = 32'b00000000000000010111011110111100;
assign LUT_3[21538] = 32'b00000000000000010010111011000011;
assign LUT_3[21539] = 32'b00000000000000011001100110100000;
assign LUT_3[21540] = 32'b00000000000000001110000001010101;
assign LUT_3[21541] = 32'b00000000000000010100101100110010;
assign LUT_3[21542] = 32'b00000000000000010000001000111001;
assign LUT_3[21543] = 32'b00000000000000010110110100010110;
assign LUT_3[21544] = 32'b00000000000000010110001100100101;
assign LUT_3[21545] = 32'b00000000000000011100111000000010;
assign LUT_3[21546] = 32'b00000000000000011000010100001001;
assign LUT_3[21547] = 32'b00000000000000011110111111100110;
assign LUT_3[21548] = 32'b00000000000000010011011010011011;
assign LUT_3[21549] = 32'b00000000000000011010000101111000;
assign LUT_3[21550] = 32'b00000000000000010101100001111111;
assign LUT_3[21551] = 32'b00000000000000011100001101011100;
assign LUT_3[21552] = 32'b00000000000000010100000110100010;
assign LUT_3[21553] = 32'b00000000000000011010110001111111;
assign LUT_3[21554] = 32'b00000000000000010110001110000110;
assign LUT_3[21555] = 32'b00000000000000011100111001100011;
assign LUT_3[21556] = 32'b00000000000000010001010100011000;
assign LUT_3[21557] = 32'b00000000000000010111111111110101;
assign LUT_3[21558] = 32'b00000000000000010011011011111100;
assign LUT_3[21559] = 32'b00000000000000011010000111011001;
assign LUT_3[21560] = 32'b00000000000000011001011111101000;
assign LUT_3[21561] = 32'b00000000000000100000001011000101;
assign LUT_3[21562] = 32'b00000000000000011011100111001100;
assign LUT_3[21563] = 32'b00000000000000100010010010101001;
assign LUT_3[21564] = 32'b00000000000000010110101101011110;
assign LUT_3[21565] = 32'b00000000000000011101011000111011;
assign LUT_3[21566] = 32'b00000000000000011000110101000010;
assign LUT_3[21567] = 32'b00000000000000011111100000011111;
assign LUT_3[21568] = 32'b00000000000000001111011101101010;
assign LUT_3[21569] = 32'b00000000000000010110001001000111;
assign LUT_3[21570] = 32'b00000000000000010001100101001110;
assign LUT_3[21571] = 32'b00000000000000011000010000101011;
assign LUT_3[21572] = 32'b00000000000000001100101011100000;
assign LUT_3[21573] = 32'b00000000000000010011010110111101;
assign LUT_3[21574] = 32'b00000000000000001110110011000100;
assign LUT_3[21575] = 32'b00000000000000010101011110100001;
assign LUT_3[21576] = 32'b00000000000000010100110110110000;
assign LUT_3[21577] = 32'b00000000000000011011100010001101;
assign LUT_3[21578] = 32'b00000000000000010110111110010100;
assign LUT_3[21579] = 32'b00000000000000011101101001110001;
assign LUT_3[21580] = 32'b00000000000000010010000100100110;
assign LUT_3[21581] = 32'b00000000000000011000110000000011;
assign LUT_3[21582] = 32'b00000000000000010100001100001010;
assign LUT_3[21583] = 32'b00000000000000011010110111100111;
assign LUT_3[21584] = 32'b00000000000000010010110000101101;
assign LUT_3[21585] = 32'b00000000000000011001011100001010;
assign LUT_3[21586] = 32'b00000000000000010100111000010001;
assign LUT_3[21587] = 32'b00000000000000011011100011101110;
assign LUT_3[21588] = 32'b00000000000000001111111110100011;
assign LUT_3[21589] = 32'b00000000000000010110101010000000;
assign LUT_3[21590] = 32'b00000000000000010010000110000111;
assign LUT_3[21591] = 32'b00000000000000011000110001100100;
assign LUT_3[21592] = 32'b00000000000000011000001001110011;
assign LUT_3[21593] = 32'b00000000000000011110110101010000;
assign LUT_3[21594] = 32'b00000000000000011010010001010111;
assign LUT_3[21595] = 32'b00000000000000100000111100110100;
assign LUT_3[21596] = 32'b00000000000000010101010111101001;
assign LUT_3[21597] = 32'b00000000000000011100000011000110;
assign LUT_3[21598] = 32'b00000000000000010111011111001101;
assign LUT_3[21599] = 32'b00000000000000011110001010101010;
assign LUT_3[21600] = 32'b00000000000000010000101100001010;
assign LUT_3[21601] = 32'b00000000000000010111010111100111;
assign LUT_3[21602] = 32'b00000000000000010010110011101110;
assign LUT_3[21603] = 32'b00000000000000011001011111001011;
assign LUT_3[21604] = 32'b00000000000000001101111010000000;
assign LUT_3[21605] = 32'b00000000000000010100100101011101;
assign LUT_3[21606] = 32'b00000000000000010000000001100100;
assign LUT_3[21607] = 32'b00000000000000010110101101000001;
assign LUT_3[21608] = 32'b00000000000000010110000101010000;
assign LUT_3[21609] = 32'b00000000000000011100110000101101;
assign LUT_3[21610] = 32'b00000000000000011000001100110100;
assign LUT_3[21611] = 32'b00000000000000011110111000010001;
assign LUT_3[21612] = 32'b00000000000000010011010011000110;
assign LUT_3[21613] = 32'b00000000000000011001111110100011;
assign LUT_3[21614] = 32'b00000000000000010101011010101010;
assign LUT_3[21615] = 32'b00000000000000011100000110000111;
assign LUT_3[21616] = 32'b00000000000000010011111111001101;
assign LUT_3[21617] = 32'b00000000000000011010101010101010;
assign LUT_3[21618] = 32'b00000000000000010110000110110001;
assign LUT_3[21619] = 32'b00000000000000011100110010001110;
assign LUT_3[21620] = 32'b00000000000000010001001101000011;
assign LUT_3[21621] = 32'b00000000000000010111111000100000;
assign LUT_3[21622] = 32'b00000000000000010011010100100111;
assign LUT_3[21623] = 32'b00000000000000011010000000000100;
assign LUT_3[21624] = 32'b00000000000000011001011000010011;
assign LUT_3[21625] = 32'b00000000000000100000000011110000;
assign LUT_3[21626] = 32'b00000000000000011011011111110111;
assign LUT_3[21627] = 32'b00000000000000100010001011010100;
assign LUT_3[21628] = 32'b00000000000000010110100110001001;
assign LUT_3[21629] = 32'b00000000000000011101010001100110;
assign LUT_3[21630] = 32'b00000000000000011000101101101101;
assign LUT_3[21631] = 32'b00000000000000011111011001001010;
assign LUT_3[21632] = 32'b00000000000000010001101111111101;
assign LUT_3[21633] = 32'b00000000000000011000011011011010;
assign LUT_3[21634] = 32'b00000000000000010011110111100001;
assign LUT_3[21635] = 32'b00000000000000011010100010111110;
assign LUT_3[21636] = 32'b00000000000000001110111101110011;
assign LUT_3[21637] = 32'b00000000000000010101101001010000;
assign LUT_3[21638] = 32'b00000000000000010001000101010111;
assign LUT_3[21639] = 32'b00000000000000010111110000110100;
assign LUT_3[21640] = 32'b00000000000000010111001001000011;
assign LUT_3[21641] = 32'b00000000000000011101110100100000;
assign LUT_3[21642] = 32'b00000000000000011001010000100111;
assign LUT_3[21643] = 32'b00000000000000011111111100000100;
assign LUT_3[21644] = 32'b00000000000000010100010110111001;
assign LUT_3[21645] = 32'b00000000000000011011000010010110;
assign LUT_3[21646] = 32'b00000000000000010110011110011101;
assign LUT_3[21647] = 32'b00000000000000011101001001111010;
assign LUT_3[21648] = 32'b00000000000000010101000011000000;
assign LUT_3[21649] = 32'b00000000000000011011101110011101;
assign LUT_3[21650] = 32'b00000000000000010111001010100100;
assign LUT_3[21651] = 32'b00000000000000011101110110000001;
assign LUT_3[21652] = 32'b00000000000000010010010000110110;
assign LUT_3[21653] = 32'b00000000000000011000111100010011;
assign LUT_3[21654] = 32'b00000000000000010100011000011010;
assign LUT_3[21655] = 32'b00000000000000011011000011110111;
assign LUT_3[21656] = 32'b00000000000000011010011100000110;
assign LUT_3[21657] = 32'b00000000000000100001000111100011;
assign LUT_3[21658] = 32'b00000000000000011100100011101010;
assign LUT_3[21659] = 32'b00000000000000100011001111000111;
assign LUT_3[21660] = 32'b00000000000000010111101001111100;
assign LUT_3[21661] = 32'b00000000000000011110010101011001;
assign LUT_3[21662] = 32'b00000000000000011001110001100000;
assign LUT_3[21663] = 32'b00000000000000100000011100111101;
assign LUT_3[21664] = 32'b00000000000000010010111110011101;
assign LUT_3[21665] = 32'b00000000000000011001101001111010;
assign LUT_3[21666] = 32'b00000000000000010101000110000001;
assign LUT_3[21667] = 32'b00000000000000011011110001011110;
assign LUT_3[21668] = 32'b00000000000000010000001100010011;
assign LUT_3[21669] = 32'b00000000000000010110110111110000;
assign LUT_3[21670] = 32'b00000000000000010010010011110111;
assign LUT_3[21671] = 32'b00000000000000011000111111010100;
assign LUT_3[21672] = 32'b00000000000000011000010111100011;
assign LUT_3[21673] = 32'b00000000000000011111000011000000;
assign LUT_3[21674] = 32'b00000000000000011010011111000111;
assign LUT_3[21675] = 32'b00000000000000100001001010100100;
assign LUT_3[21676] = 32'b00000000000000010101100101011001;
assign LUT_3[21677] = 32'b00000000000000011100010000110110;
assign LUT_3[21678] = 32'b00000000000000010111101100111101;
assign LUT_3[21679] = 32'b00000000000000011110011000011010;
assign LUT_3[21680] = 32'b00000000000000010110010001100000;
assign LUT_3[21681] = 32'b00000000000000011100111100111101;
assign LUT_3[21682] = 32'b00000000000000011000011001000100;
assign LUT_3[21683] = 32'b00000000000000011111000100100001;
assign LUT_3[21684] = 32'b00000000000000010011011111010110;
assign LUT_3[21685] = 32'b00000000000000011010001010110011;
assign LUT_3[21686] = 32'b00000000000000010101100110111010;
assign LUT_3[21687] = 32'b00000000000000011100010010010111;
assign LUT_3[21688] = 32'b00000000000000011011101010100110;
assign LUT_3[21689] = 32'b00000000000000100010010110000011;
assign LUT_3[21690] = 32'b00000000000000011101110010001010;
assign LUT_3[21691] = 32'b00000000000000100100011101100111;
assign LUT_3[21692] = 32'b00000000000000011000111000011100;
assign LUT_3[21693] = 32'b00000000000000011111100011111001;
assign LUT_3[21694] = 32'b00000000000000011011000000000000;
assign LUT_3[21695] = 32'b00000000000000100001101011011101;
assign LUT_3[21696] = 32'b00000000000000010001101000101000;
assign LUT_3[21697] = 32'b00000000000000011000010100000101;
assign LUT_3[21698] = 32'b00000000000000010011110000001100;
assign LUT_3[21699] = 32'b00000000000000011010011011101001;
assign LUT_3[21700] = 32'b00000000000000001110110110011110;
assign LUT_3[21701] = 32'b00000000000000010101100001111011;
assign LUT_3[21702] = 32'b00000000000000010000111110000010;
assign LUT_3[21703] = 32'b00000000000000010111101001011111;
assign LUT_3[21704] = 32'b00000000000000010111000001101110;
assign LUT_3[21705] = 32'b00000000000000011101101101001011;
assign LUT_3[21706] = 32'b00000000000000011001001001010010;
assign LUT_3[21707] = 32'b00000000000000011111110100101111;
assign LUT_3[21708] = 32'b00000000000000010100001111100100;
assign LUT_3[21709] = 32'b00000000000000011010111011000001;
assign LUT_3[21710] = 32'b00000000000000010110010111001000;
assign LUT_3[21711] = 32'b00000000000000011101000010100101;
assign LUT_3[21712] = 32'b00000000000000010100111011101011;
assign LUT_3[21713] = 32'b00000000000000011011100111001000;
assign LUT_3[21714] = 32'b00000000000000010111000011001111;
assign LUT_3[21715] = 32'b00000000000000011101101110101100;
assign LUT_3[21716] = 32'b00000000000000010010001001100001;
assign LUT_3[21717] = 32'b00000000000000011000110100111110;
assign LUT_3[21718] = 32'b00000000000000010100010001000101;
assign LUT_3[21719] = 32'b00000000000000011010111100100010;
assign LUT_3[21720] = 32'b00000000000000011010010100110001;
assign LUT_3[21721] = 32'b00000000000000100001000000001110;
assign LUT_3[21722] = 32'b00000000000000011100011100010101;
assign LUT_3[21723] = 32'b00000000000000100011000111110010;
assign LUT_3[21724] = 32'b00000000000000010111100010100111;
assign LUT_3[21725] = 32'b00000000000000011110001110000100;
assign LUT_3[21726] = 32'b00000000000000011001101010001011;
assign LUT_3[21727] = 32'b00000000000000100000010101101000;
assign LUT_3[21728] = 32'b00000000000000010010110111001000;
assign LUT_3[21729] = 32'b00000000000000011001100010100101;
assign LUT_3[21730] = 32'b00000000000000010100111110101100;
assign LUT_3[21731] = 32'b00000000000000011011101010001001;
assign LUT_3[21732] = 32'b00000000000000010000000100111110;
assign LUT_3[21733] = 32'b00000000000000010110110000011011;
assign LUT_3[21734] = 32'b00000000000000010010001100100010;
assign LUT_3[21735] = 32'b00000000000000011000110111111111;
assign LUT_3[21736] = 32'b00000000000000011000010000001110;
assign LUT_3[21737] = 32'b00000000000000011110111011101011;
assign LUT_3[21738] = 32'b00000000000000011010010111110010;
assign LUT_3[21739] = 32'b00000000000000100001000011001111;
assign LUT_3[21740] = 32'b00000000000000010101011110000100;
assign LUT_3[21741] = 32'b00000000000000011100001001100001;
assign LUT_3[21742] = 32'b00000000000000010111100101101000;
assign LUT_3[21743] = 32'b00000000000000011110010001000101;
assign LUT_3[21744] = 32'b00000000000000010110001010001011;
assign LUT_3[21745] = 32'b00000000000000011100110101101000;
assign LUT_3[21746] = 32'b00000000000000011000010001101111;
assign LUT_3[21747] = 32'b00000000000000011110111101001100;
assign LUT_3[21748] = 32'b00000000000000010011011000000001;
assign LUT_3[21749] = 32'b00000000000000011010000011011110;
assign LUT_3[21750] = 32'b00000000000000010101011111100101;
assign LUT_3[21751] = 32'b00000000000000011100001011000010;
assign LUT_3[21752] = 32'b00000000000000011011100011010001;
assign LUT_3[21753] = 32'b00000000000000100010001110101110;
assign LUT_3[21754] = 32'b00000000000000011101101010110101;
assign LUT_3[21755] = 32'b00000000000000100100010110010010;
assign LUT_3[21756] = 32'b00000000000000011000110001000111;
assign LUT_3[21757] = 32'b00000000000000011111011100100100;
assign LUT_3[21758] = 32'b00000000000000011010111000101011;
assign LUT_3[21759] = 32'b00000000000000100001100100001000;
assign LUT_3[21760] = 32'b00000000000000001011110100100000;
assign LUT_3[21761] = 32'b00000000000000010010011111111101;
assign LUT_3[21762] = 32'b00000000000000001101111100000100;
assign LUT_3[21763] = 32'b00000000000000010100100111100001;
assign LUT_3[21764] = 32'b00000000000000001001000010010110;
assign LUT_3[21765] = 32'b00000000000000001111101101110011;
assign LUT_3[21766] = 32'b00000000000000001011001001111010;
assign LUT_3[21767] = 32'b00000000000000010001110101010111;
assign LUT_3[21768] = 32'b00000000000000010001001101100110;
assign LUT_3[21769] = 32'b00000000000000010111111001000011;
assign LUT_3[21770] = 32'b00000000000000010011010101001010;
assign LUT_3[21771] = 32'b00000000000000011010000000100111;
assign LUT_3[21772] = 32'b00000000000000001110011011011100;
assign LUT_3[21773] = 32'b00000000000000010101000110111001;
assign LUT_3[21774] = 32'b00000000000000010000100011000000;
assign LUT_3[21775] = 32'b00000000000000010111001110011101;
assign LUT_3[21776] = 32'b00000000000000001111000111100011;
assign LUT_3[21777] = 32'b00000000000000010101110011000000;
assign LUT_3[21778] = 32'b00000000000000010001001111000111;
assign LUT_3[21779] = 32'b00000000000000010111111010100100;
assign LUT_3[21780] = 32'b00000000000000001100010101011001;
assign LUT_3[21781] = 32'b00000000000000010011000000110110;
assign LUT_3[21782] = 32'b00000000000000001110011100111101;
assign LUT_3[21783] = 32'b00000000000000010101001000011010;
assign LUT_3[21784] = 32'b00000000000000010100100000101001;
assign LUT_3[21785] = 32'b00000000000000011011001100000110;
assign LUT_3[21786] = 32'b00000000000000010110101000001101;
assign LUT_3[21787] = 32'b00000000000000011101010011101010;
assign LUT_3[21788] = 32'b00000000000000010001101110011111;
assign LUT_3[21789] = 32'b00000000000000011000011001111100;
assign LUT_3[21790] = 32'b00000000000000010011110110000011;
assign LUT_3[21791] = 32'b00000000000000011010100001100000;
assign LUT_3[21792] = 32'b00000000000000001101000011000000;
assign LUT_3[21793] = 32'b00000000000000010011101110011101;
assign LUT_3[21794] = 32'b00000000000000001111001010100100;
assign LUT_3[21795] = 32'b00000000000000010101110110000001;
assign LUT_3[21796] = 32'b00000000000000001010010000110110;
assign LUT_3[21797] = 32'b00000000000000010000111100010011;
assign LUT_3[21798] = 32'b00000000000000001100011000011010;
assign LUT_3[21799] = 32'b00000000000000010011000011110111;
assign LUT_3[21800] = 32'b00000000000000010010011100000110;
assign LUT_3[21801] = 32'b00000000000000011001000111100011;
assign LUT_3[21802] = 32'b00000000000000010100100011101010;
assign LUT_3[21803] = 32'b00000000000000011011001111000111;
assign LUT_3[21804] = 32'b00000000000000001111101001111100;
assign LUT_3[21805] = 32'b00000000000000010110010101011001;
assign LUT_3[21806] = 32'b00000000000000010001110001100000;
assign LUT_3[21807] = 32'b00000000000000011000011100111101;
assign LUT_3[21808] = 32'b00000000000000010000010110000011;
assign LUT_3[21809] = 32'b00000000000000010111000001100000;
assign LUT_3[21810] = 32'b00000000000000010010011101100111;
assign LUT_3[21811] = 32'b00000000000000011001001001000100;
assign LUT_3[21812] = 32'b00000000000000001101100011111001;
assign LUT_3[21813] = 32'b00000000000000010100001111010110;
assign LUT_3[21814] = 32'b00000000000000001111101011011101;
assign LUT_3[21815] = 32'b00000000000000010110010110111010;
assign LUT_3[21816] = 32'b00000000000000010101101111001001;
assign LUT_3[21817] = 32'b00000000000000011100011010100110;
assign LUT_3[21818] = 32'b00000000000000010111110110101101;
assign LUT_3[21819] = 32'b00000000000000011110100010001010;
assign LUT_3[21820] = 32'b00000000000000010010111100111111;
assign LUT_3[21821] = 32'b00000000000000011001101000011100;
assign LUT_3[21822] = 32'b00000000000000010101000100100011;
assign LUT_3[21823] = 32'b00000000000000011011110000000000;
assign LUT_3[21824] = 32'b00000000000000001011101101001011;
assign LUT_3[21825] = 32'b00000000000000010010011000101000;
assign LUT_3[21826] = 32'b00000000000000001101110100101111;
assign LUT_3[21827] = 32'b00000000000000010100100000001100;
assign LUT_3[21828] = 32'b00000000000000001000111011000001;
assign LUT_3[21829] = 32'b00000000000000001111100110011110;
assign LUT_3[21830] = 32'b00000000000000001011000010100101;
assign LUT_3[21831] = 32'b00000000000000010001101110000010;
assign LUT_3[21832] = 32'b00000000000000010001000110010001;
assign LUT_3[21833] = 32'b00000000000000010111110001101110;
assign LUT_3[21834] = 32'b00000000000000010011001101110101;
assign LUT_3[21835] = 32'b00000000000000011001111001010010;
assign LUT_3[21836] = 32'b00000000000000001110010100000111;
assign LUT_3[21837] = 32'b00000000000000010100111111100100;
assign LUT_3[21838] = 32'b00000000000000010000011011101011;
assign LUT_3[21839] = 32'b00000000000000010111000111001000;
assign LUT_3[21840] = 32'b00000000000000001111000000001110;
assign LUT_3[21841] = 32'b00000000000000010101101011101011;
assign LUT_3[21842] = 32'b00000000000000010001000111110010;
assign LUT_3[21843] = 32'b00000000000000010111110011001111;
assign LUT_3[21844] = 32'b00000000000000001100001110000100;
assign LUT_3[21845] = 32'b00000000000000010010111001100001;
assign LUT_3[21846] = 32'b00000000000000001110010101101000;
assign LUT_3[21847] = 32'b00000000000000010101000001000101;
assign LUT_3[21848] = 32'b00000000000000010100011001010100;
assign LUT_3[21849] = 32'b00000000000000011011000100110001;
assign LUT_3[21850] = 32'b00000000000000010110100000111000;
assign LUT_3[21851] = 32'b00000000000000011101001100010101;
assign LUT_3[21852] = 32'b00000000000000010001100111001010;
assign LUT_3[21853] = 32'b00000000000000011000010010100111;
assign LUT_3[21854] = 32'b00000000000000010011101110101110;
assign LUT_3[21855] = 32'b00000000000000011010011010001011;
assign LUT_3[21856] = 32'b00000000000000001100111011101011;
assign LUT_3[21857] = 32'b00000000000000010011100111001000;
assign LUT_3[21858] = 32'b00000000000000001111000011001111;
assign LUT_3[21859] = 32'b00000000000000010101101110101100;
assign LUT_3[21860] = 32'b00000000000000001010001001100001;
assign LUT_3[21861] = 32'b00000000000000010000110100111110;
assign LUT_3[21862] = 32'b00000000000000001100010001000101;
assign LUT_3[21863] = 32'b00000000000000010010111100100010;
assign LUT_3[21864] = 32'b00000000000000010010010100110001;
assign LUT_3[21865] = 32'b00000000000000011001000000001110;
assign LUT_3[21866] = 32'b00000000000000010100011100010101;
assign LUT_3[21867] = 32'b00000000000000011011000111110010;
assign LUT_3[21868] = 32'b00000000000000001111100010100111;
assign LUT_3[21869] = 32'b00000000000000010110001110000100;
assign LUT_3[21870] = 32'b00000000000000010001101010001011;
assign LUT_3[21871] = 32'b00000000000000011000010101101000;
assign LUT_3[21872] = 32'b00000000000000010000001110101110;
assign LUT_3[21873] = 32'b00000000000000010110111010001011;
assign LUT_3[21874] = 32'b00000000000000010010010110010010;
assign LUT_3[21875] = 32'b00000000000000011001000001101111;
assign LUT_3[21876] = 32'b00000000000000001101011100100100;
assign LUT_3[21877] = 32'b00000000000000010100001000000001;
assign LUT_3[21878] = 32'b00000000000000001111100100001000;
assign LUT_3[21879] = 32'b00000000000000010110001111100101;
assign LUT_3[21880] = 32'b00000000000000010101100111110100;
assign LUT_3[21881] = 32'b00000000000000011100010011010001;
assign LUT_3[21882] = 32'b00000000000000010111101111011000;
assign LUT_3[21883] = 32'b00000000000000011110011010110101;
assign LUT_3[21884] = 32'b00000000000000010010110101101010;
assign LUT_3[21885] = 32'b00000000000000011001100001000111;
assign LUT_3[21886] = 32'b00000000000000010100111101001110;
assign LUT_3[21887] = 32'b00000000000000011011101000101011;
assign LUT_3[21888] = 32'b00000000000000001101111111011110;
assign LUT_3[21889] = 32'b00000000000000010100101010111011;
assign LUT_3[21890] = 32'b00000000000000010000000111000010;
assign LUT_3[21891] = 32'b00000000000000010110110010011111;
assign LUT_3[21892] = 32'b00000000000000001011001101010100;
assign LUT_3[21893] = 32'b00000000000000010001111000110001;
assign LUT_3[21894] = 32'b00000000000000001101010100111000;
assign LUT_3[21895] = 32'b00000000000000010100000000010101;
assign LUT_3[21896] = 32'b00000000000000010011011000100100;
assign LUT_3[21897] = 32'b00000000000000011010000100000001;
assign LUT_3[21898] = 32'b00000000000000010101100000001000;
assign LUT_3[21899] = 32'b00000000000000011100001011100101;
assign LUT_3[21900] = 32'b00000000000000010000100110011010;
assign LUT_3[21901] = 32'b00000000000000010111010001110111;
assign LUT_3[21902] = 32'b00000000000000010010101101111110;
assign LUT_3[21903] = 32'b00000000000000011001011001011011;
assign LUT_3[21904] = 32'b00000000000000010001010010100001;
assign LUT_3[21905] = 32'b00000000000000010111111101111110;
assign LUT_3[21906] = 32'b00000000000000010011011010000101;
assign LUT_3[21907] = 32'b00000000000000011010000101100010;
assign LUT_3[21908] = 32'b00000000000000001110100000010111;
assign LUT_3[21909] = 32'b00000000000000010101001011110100;
assign LUT_3[21910] = 32'b00000000000000010000100111111011;
assign LUT_3[21911] = 32'b00000000000000010111010011011000;
assign LUT_3[21912] = 32'b00000000000000010110101011100111;
assign LUT_3[21913] = 32'b00000000000000011101010111000100;
assign LUT_3[21914] = 32'b00000000000000011000110011001011;
assign LUT_3[21915] = 32'b00000000000000011111011110101000;
assign LUT_3[21916] = 32'b00000000000000010011111001011101;
assign LUT_3[21917] = 32'b00000000000000011010100100111010;
assign LUT_3[21918] = 32'b00000000000000010110000001000001;
assign LUT_3[21919] = 32'b00000000000000011100101100011110;
assign LUT_3[21920] = 32'b00000000000000001111001101111110;
assign LUT_3[21921] = 32'b00000000000000010101111001011011;
assign LUT_3[21922] = 32'b00000000000000010001010101100010;
assign LUT_3[21923] = 32'b00000000000000011000000000111111;
assign LUT_3[21924] = 32'b00000000000000001100011011110100;
assign LUT_3[21925] = 32'b00000000000000010011000111010001;
assign LUT_3[21926] = 32'b00000000000000001110100011011000;
assign LUT_3[21927] = 32'b00000000000000010101001110110101;
assign LUT_3[21928] = 32'b00000000000000010100100111000100;
assign LUT_3[21929] = 32'b00000000000000011011010010100001;
assign LUT_3[21930] = 32'b00000000000000010110101110101000;
assign LUT_3[21931] = 32'b00000000000000011101011010000101;
assign LUT_3[21932] = 32'b00000000000000010001110100111010;
assign LUT_3[21933] = 32'b00000000000000011000100000010111;
assign LUT_3[21934] = 32'b00000000000000010011111100011110;
assign LUT_3[21935] = 32'b00000000000000011010100111111011;
assign LUT_3[21936] = 32'b00000000000000010010100001000001;
assign LUT_3[21937] = 32'b00000000000000011001001100011110;
assign LUT_3[21938] = 32'b00000000000000010100101000100101;
assign LUT_3[21939] = 32'b00000000000000011011010100000010;
assign LUT_3[21940] = 32'b00000000000000001111101110110111;
assign LUT_3[21941] = 32'b00000000000000010110011010010100;
assign LUT_3[21942] = 32'b00000000000000010001110110011011;
assign LUT_3[21943] = 32'b00000000000000011000100001111000;
assign LUT_3[21944] = 32'b00000000000000010111111010000111;
assign LUT_3[21945] = 32'b00000000000000011110100101100100;
assign LUT_3[21946] = 32'b00000000000000011010000001101011;
assign LUT_3[21947] = 32'b00000000000000100000101101001000;
assign LUT_3[21948] = 32'b00000000000000010101000111111101;
assign LUT_3[21949] = 32'b00000000000000011011110011011010;
assign LUT_3[21950] = 32'b00000000000000010111001111100001;
assign LUT_3[21951] = 32'b00000000000000011101111010111110;
assign LUT_3[21952] = 32'b00000000000000001101111000001001;
assign LUT_3[21953] = 32'b00000000000000010100100011100110;
assign LUT_3[21954] = 32'b00000000000000001111111111101101;
assign LUT_3[21955] = 32'b00000000000000010110101011001010;
assign LUT_3[21956] = 32'b00000000000000001011000101111111;
assign LUT_3[21957] = 32'b00000000000000010001110001011100;
assign LUT_3[21958] = 32'b00000000000000001101001101100011;
assign LUT_3[21959] = 32'b00000000000000010011111001000000;
assign LUT_3[21960] = 32'b00000000000000010011010001001111;
assign LUT_3[21961] = 32'b00000000000000011001111100101100;
assign LUT_3[21962] = 32'b00000000000000010101011000110011;
assign LUT_3[21963] = 32'b00000000000000011100000100010000;
assign LUT_3[21964] = 32'b00000000000000010000011111000101;
assign LUT_3[21965] = 32'b00000000000000010111001010100010;
assign LUT_3[21966] = 32'b00000000000000010010100110101001;
assign LUT_3[21967] = 32'b00000000000000011001010010000110;
assign LUT_3[21968] = 32'b00000000000000010001001011001100;
assign LUT_3[21969] = 32'b00000000000000010111110110101001;
assign LUT_3[21970] = 32'b00000000000000010011010010110000;
assign LUT_3[21971] = 32'b00000000000000011001111110001101;
assign LUT_3[21972] = 32'b00000000000000001110011001000010;
assign LUT_3[21973] = 32'b00000000000000010101000100011111;
assign LUT_3[21974] = 32'b00000000000000010000100000100110;
assign LUT_3[21975] = 32'b00000000000000010111001100000011;
assign LUT_3[21976] = 32'b00000000000000010110100100010010;
assign LUT_3[21977] = 32'b00000000000000011101001111101111;
assign LUT_3[21978] = 32'b00000000000000011000101011110110;
assign LUT_3[21979] = 32'b00000000000000011111010111010011;
assign LUT_3[21980] = 32'b00000000000000010011110010001000;
assign LUT_3[21981] = 32'b00000000000000011010011101100101;
assign LUT_3[21982] = 32'b00000000000000010101111001101100;
assign LUT_3[21983] = 32'b00000000000000011100100101001001;
assign LUT_3[21984] = 32'b00000000000000001111000110101001;
assign LUT_3[21985] = 32'b00000000000000010101110010000110;
assign LUT_3[21986] = 32'b00000000000000010001001110001101;
assign LUT_3[21987] = 32'b00000000000000010111111001101010;
assign LUT_3[21988] = 32'b00000000000000001100010100011111;
assign LUT_3[21989] = 32'b00000000000000010010111111111100;
assign LUT_3[21990] = 32'b00000000000000001110011100000011;
assign LUT_3[21991] = 32'b00000000000000010101000111100000;
assign LUT_3[21992] = 32'b00000000000000010100011111101111;
assign LUT_3[21993] = 32'b00000000000000011011001011001100;
assign LUT_3[21994] = 32'b00000000000000010110100111010011;
assign LUT_3[21995] = 32'b00000000000000011101010010110000;
assign LUT_3[21996] = 32'b00000000000000010001101101100101;
assign LUT_3[21997] = 32'b00000000000000011000011001000010;
assign LUT_3[21998] = 32'b00000000000000010011110101001001;
assign LUT_3[21999] = 32'b00000000000000011010100000100110;
assign LUT_3[22000] = 32'b00000000000000010010011001101100;
assign LUT_3[22001] = 32'b00000000000000011001000101001001;
assign LUT_3[22002] = 32'b00000000000000010100100001010000;
assign LUT_3[22003] = 32'b00000000000000011011001100101101;
assign LUT_3[22004] = 32'b00000000000000001111100111100010;
assign LUT_3[22005] = 32'b00000000000000010110010010111111;
assign LUT_3[22006] = 32'b00000000000000010001101111000110;
assign LUT_3[22007] = 32'b00000000000000011000011010100011;
assign LUT_3[22008] = 32'b00000000000000010111110010110010;
assign LUT_3[22009] = 32'b00000000000000011110011110001111;
assign LUT_3[22010] = 32'b00000000000000011001111010010110;
assign LUT_3[22011] = 32'b00000000000000100000100101110011;
assign LUT_3[22012] = 32'b00000000000000010101000000101000;
assign LUT_3[22013] = 32'b00000000000000011011101100000101;
assign LUT_3[22014] = 32'b00000000000000010111001000001100;
assign LUT_3[22015] = 32'b00000000000000011101110011101001;
assign LUT_3[22016] = 32'b00000000000000010010111010001011;
assign LUT_3[22017] = 32'b00000000000000011001100101101000;
assign LUT_3[22018] = 32'b00000000000000010101000001101111;
assign LUT_3[22019] = 32'b00000000000000011011101101001100;
assign LUT_3[22020] = 32'b00000000000000010000001000000001;
assign LUT_3[22021] = 32'b00000000000000010110110011011110;
assign LUT_3[22022] = 32'b00000000000000010010001111100101;
assign LUT_3[22023] = 32'b00000000000000011000111011000010;
assign LUT_3[22024] = 32'b00000000000000011000010011010001;
assign LUT_3[22025] = 32'b00000000000000011110111110101110;
assign LUT_3[22026] = 32'b00000000000000011010011010110101;
assign LUT_3[22027] = 32'b00000000000000100001000110010010;
assign LUT_3[22028] = 32'b00000000000000010101100001000111;
assign LUT_3[22029] = 32'b00000000000000011100001100100100;
assign LUT_3[22030] = 32'b00000000000000010111101000101011;
assign LUT_3[22031] = 32'b00000000000000011110010100001000;
assign LUT_3[22032] = 32'b00000000000000010110001101001110;
assign LUT_3[22033] = 32'b00000000000000011100111000101011;
assign LUT_3[22034] = 32'b00000000000000011000010100110010;
assign LUT_3[22035] = 32'b00000000000000011111000000001111;
assign LUT_3[22036] = 32'b00000000000000010011011011000100;
assign LUT_3[22037] = 32'b00000000000000011010000110100001;
assign LUT_3[22038] = 32'b00000000000000010101100010101000;
assign LUT_3[22039] = 32'b00000000000000011100001110000101;
assign LUT_3[22040] = 32'b00000000000000011011100110010100;
assign LUT_3[22041] = 32'b00000000000000100010010001110001;
assign LUT_3[22042] = 32'b00000000000000011101101101111000;
assign LUT_3[22043] = 32'b00000000000000100100011001010101;
assign LUT_3[22044] = 32'b00000000000000011000110100001010;
assign LUT_3[22045] = 32'b00000000000000011111011111100111;
assign LUT_3[22046] = 32'b00000000000000011010111011101110;
assign LUT_3[22047] = 32'b00000000000000100001100111001011;
assign LUT_3[22048] = 32'b00000000000000010100001000101011;
assign LUT_3[22049] = 32'b00000000000000011010110100001000;
assign LUT_3[22050] = 32'b00000000000000010110010000001111;
assign LUT_3[22051] = 32'b00000000000000011100111011101100;
assign LUT_3[22052] = 32'b00000000000000010001010110100001;
assign LUT_3[22053] = 32'b00000000000000011000000001111110;
assign LUT_3[22054] = 32'b00000000000000010011011110000101;
assign LUT_3[22055] = 32'b00000000000000011010001001100010;
assign LUT_3[22056] = 32'b00000000000000011001100001110001;
assign LUT_3[22057] = 32'b00000000000000100000001101001110;
assign LUT_3[22058] = 32'b00000000000000011011101001010101;
assign LUT_3[22059] = 32'b00000000000000100010010100110010;
assign LUT_3[22060] = 32'b00000000000000010110101111100111;
assign LUT_3[22061] = 32'b00000000000000011101011011000100;
assign LUT_3[22062] = 32'b00000000000000011000110111001011;
assign LUT_3[22063] = 32'b00000000000000011111100010101000;
assign LUT_3[22064] = 32'b00000000000000010111011011101110;
assign LUT_3[22065] = 32'b00000000000000011110000111001011;
assign LUT_3[22066] = 32'b00000000000000011001100011010010;
assign LUT_3[22067] = 32'b00000000000000100000001110101111;
assign LUT_3[22068] = 32'b00000000000000010100101001100100;
assign LUT_3[22069] = 32'b00000000000000011011010101000001;
assign LUT_3[22070] = 32'b00000000000000010110110001001000;
assign LUT_3[22071] = 32'b00000000000000011101011100100101;
assign LUT_3[22072] = 32'b00000000000000011100110100110100;
assign LUT_3[22073] = 32'b00000000000000100011100000010001;
assign LUT_3[22074] = 32'b00000000000000011110111100011000;
assign LUT_3[22075] = 32'b00000000000000100101100111110101;
assign LUT_3[22076] = 32'b00000000000000011010000010101010;
assign LUT_3[22077] = 32'b00000000000000100000101110000111;
assign LUT_3[22078] = 32'b00000000000000011100001010001110;
assign LUT_3[22079] = 32'b00000000000000100010110101101011;
assign LUT_3[22080] = 32'b00000000000000010010110010110110;
assign LUT_3[22081] = 32'b00000000000000011001011110010011;
assign LUT_3[22082] = 32'b00000000000000010100111010011010;
assign LUT_3[22083] = 32'b00000000000000011011100101110111;
assign LUT_3[22084] = 32'b00000000000000010000000000101100;
assign LUT_3[22085] = 32'b00000000000000010110101100001001;
assign LUT_3[22086] = 32'b00000000000000010010001000010000;
assign LUT_3[22087] = 32'b00000000000000011000110011101101;
assign LUT_3[22088] = 32'b00000000000000011000001011111100;
assign LUT_3[22089] = 32'b00000000000000011110110111011001;
assign LUT_3[22090] = 32'b00000000000000011010010011100000;
assign LUT_3[22091] = 32'b00000000000000100000111110111101;
assign LUT_3[22092] = 32'b00000000000000010101011001110010;
assign LUT_3[22093] = 32'b00000000000000011100000101001111;
assign LUT_3[22094] = 32'b00000000000000010111100001010110;
assign LUT_3[22095] = 32'b00000000000000011110001100110011;
assign LUT_3[22096] = 32'b00000000000000010110000101111001;
assign LUT_3[22097] = 32'b00000000000000011100110001010110;
assign LUT_3[22098] = 32'b00000000000000011000001101011101;
assign LUT_3[22099] = 32'b00000000000000011110111000111010;
assign LUT_3[22100] = 32'b00000000000000010011010011101111;
assign LUT_3[22101] = 32'b00000000000000011001111111001100;
assign LUT_3[22102] = 32'b00000000000000010101011011010011;
assign LUT_3[22103] = 32'b00000000000000011100000110110000;
assign LUT_3[22104] = 32'b00000000000000011011011110111111;
assign LUT_3[22105] = 32'b00000000000000100010001010011100;
assign LUT_3[22106] = 32'b00000000000000011101100110100011;
assign LUT_3[22107] = 32'b00000000000000100100010010000000;
assign LUT_3[22108] = 32'b00000000000000011000101100110101;
assign LUT_3[22109] = 32'b00000000000000011111011000010010;
assign LUT_3[22110] = 32'b00000000000000011010110100011001;
assign LUT_3[22111] = 32'b00000000000000100001011111110110;
assign LUT_3[22112] = 32'b00000000000000010100000001010110;
assign LUT_3[22113] = 32'b00000000000000011010101100110011;
assign LUT_3[22114] = 32'b00000000000000010110001000111010;
assign LUT_3[22115] = 32'b00000000000000011100110100010111;
assign LUT_3[22116] = 32'b00000000000000010001001111001100;
assign LUT_3[22117] = 32'b00000000000000010111111010101001;
assign LUT_3[22118] = 32'b00000000000000010011010110110000;
assign LUT_3[22119] = 32'b00000000000000011010000010001101;
assign LUT_3[22120] = 32'b00000000000000011001011010011100;
assign LUT_3[22121] = 32'b00000000000000100000000101111001;
assign LUT_3[22122] = 32'b00000000000000011011100010000000;
assign LUT_3[22123] = 32'b00000000000000100010001101011101;
assign LUT_3[22124] = 32'b00000000000000010110101000010010;
assign LUT_3[22125] = 32'b00000000000000011101010011101111;
assign LUT_3[22126] = 32'b00000000000000011000101111110110;
assign LUT_3[22127] = 32'b00000000000000011111011011010011;
assign LUT_3[22128] = 32'b00000000000000010111010100011001;
assign LUT_3[22129] = 32'b00000000000000011101111111110110;
assign LUT_3[22130] = 32'b00000000000000011001011011111101;
assign LUT_3[22131] = 32'b00000000000000100000000111011010;
assign LUT_3[22132] = 32'b00000000000000010100100010001111;
assign LUT_3[22133] = 32'b00000000000000011011001101101100;
assign LUT_3[22134] = 32'b00000000000000010110101001110011;
assign LUT_3[22135] = 32'b00000000000000011101010101010000;
assign LUT_3[22136] = 32'b00000000000000011100101101011111;
assign LUT_3[22137] = 32'b00000000000000100011011000111100;
assign LUT_3[22138] = 32'b00000000000000011110110101000011;
assign LUT_3[22139] = 32'b00000000000000100101100000100000;
assign LUT_3[22140] = 32'b00000000000000011001111011010101;
assign LUT_3[22141] = 32'b00000000000000100000100110110010;
assign LUT_3[22142] = 32'b00000000000000011100000010111001;
assign LUT_3[22143] = 32'b00000000000000100010101110010110;
assign LUT_3[22144] = 32'b00000000000000010101000101001001;
assign LUT_3[22145] = 32'b00000000000000011011110000100110;
assign LUT_3[22146] = 32'b00000000000000010111001100101101;
assign LUT_3[22147] = 32'b00000000000000011101111000001010;
assign LUT_3[22148] = 32'b00000000000000010010010010111111;
assign LUT_3[22149] = 32'b00000000000000011000111110011100;
assign LUT_3[22150] = 32'b00000000000000010100011010100011;
assign LUT_3[22151] = 32'b00000000000000011011000110000000;
assign LUT_3[22152] = 32'b00000000000000011010011110001111;
assign LUT_3[22153] = 32'b00000000000000100001001001101100;
assign LUT_3[22154] = 32'b00000000000000011100100101110011;
assign LUT_3[22155] = 32'b00000000000000100011010001010000;
assign LUT_3[22156] = 32'b00000000000000010111101100000101;
assign LUT_3[22157] = 32'b00000000000000011110010111100010;
assign LUT_3[22158] = 32'b00000000000000011001110011101001;
assign LUT_3[22159] = 32'b00000000000000100000011111000110;
assign LUT_3[22160] = 32'b00000000000000011000011000001100;
assign LUT_3[22161] = 32'b00000000000000011111000011101001;
assign LUT_3[22162] = 32'b00000000000000011010011111110000;
assign LUT_3[22163] = 32'b00000000000000100001001011001101;
assign LUT_3[22164] = 32'b00000000000000010101100110000010;
assign LUT_3[22165] = 32'b00000000000000011100010001011111;
assign LUT_3[22166] = 32'b00000000000000010111101101100110;
assign LUT_3[22167] = 32'b00000000000000011110011001000011;
assign LUT_3[22168] = 32'b00000000000000011101110001010010;
assign LUT_3[22169] = 32'b00000000000000100100011100101111;
assign LUT_3[22170] = 32'b00000000000000011111111000110110;
assign LUT_3[22171] = 32'b00000000000000100110100100010011;
assign LUT_3[22172] = 32'b00000000000000011010111111001000;
assign LUT_3[22173] = 32'b00000000000000100001101010100101;
assign LUT_3[22174] = 32'b00000000000000011101000110101100;
assign LUT_3[22175] = 32'b00000000000000100011110010001001;
assign LUT_3[22176] = 32'b00000000000000010110010011101001;
assign LUT_3[22177] = 32'b00000000000000011100111111000110;
assign LUT_3[22178] = 32'b00000000000000011000011011001101;
assign LUT_3[22179] = 32'b00000000000000011111000110101010;
assign LUT_3[22180] = 32'b00000000000000010011100001011111;
assign LUT_3[22181] = 32'b00000000000000011010001100111100;
assign LUT_3[22182] = 32'b00000000000000010101101001000011;
assign LUT_3[22183] = 32'b00000000000000011100010100100000;
assign LUT_3[22184] = 32'b00000000000000011011101100101111;
assign LUT_3[22185] = 32'b00000000000000100010011000001100;
assign LUT_3[22186] = 32'b00000000000000011101110100010011;
assign LUT_3[22187] = 32'b00000000000000100100011111110000;
assign LUT_3[22188] = 32'b00000000000000011000111010100101;
assign LUT_3[22189] = 32'b00000000000000011111100110000010;
assign LUT_3[22190] = 32'b00000000000000011011000010001001;
assign LUT_3[22191] = 32'b00000000000000100001101101100110;
assign LUT_3[22192] = 32'b00000000000000011001100110101100;
assign LUT_3[22193] = 32'b00000000000000100000010010001001;
assign LUT_3[22194] = 32'b00000000000000011011101110010000;
assign LUT_3[22195] = 32'b00000000000000100010011001101101;
assign LUT_3[22196] = 32'b00000000000000010110110100100010;
assign LUT_3[22197] = 32'b00000000000000011101011111111111;
assign LUT_3[22198] = 32'b00000000000000011000111100000110;
assign LUT_3[22199] = 32'b00000000000000011111100111100011;
assign LUT_3[22200] = 32'b00000000000000011110111111110010;
assign LUT_3[22201] = 32'b00000000000000100101101011001111;
assign LUT_3[22202] = 32'b00000000000000100001000111010110;
assign LUT_3[22203] = 32'b00000000000000100111110010110011;
assign LUT_3[22204] = 32'b00000000000000011100001101101000;
assign LUT_3[22205] = 32'b00000000000000100010111001000101;
assign LUT_3[22206] = 32'b00000000000000011110010101001100;
assign LUT_3[22207] = 32'b00000000000000100101000000101001;
assign LUT_3[22208] = 32'b00000000000000010100111101110100;
assign LUT_3[22209] = 32'b00000000000000011011101001010001;
assign LUT_3[22210] = 32'b00000000000000010111000101011000;
assign LUT_3[22211] = 32'b00000000000000011101110000110101;
assign LUT_3[22212] = 32'b00000000000000010010001011101010;
assign LUT_3[22213] = 32'b00000000000000011000110111000111;
assign LUT_3[22214] = 32'b00000000000000010100010011001110;
assign LUT_3[22215] = 32'b00000000000000011010111110101011;
assign LUT_3[22216] = 32'b00000000000000011010010110111010;
assign LUT_3[22217] = 32'b00000000000000100001000010010111;
assign LUT_3[22218] = 32'b00000000000000011100011110011110;
assign LUT_3[22219] = 32'b00000000000000100011001001111011;
assign LUT_3[22220] = 32'b00000000000000010111100100110000;
assign LUT_3[22221] = 32'b00000000000000011110010000001101;
assign LUT_3[22222] = 32'b00000000000000011001101100010100;
assign LUT_3[22223] = 32'b00000000000000100000010111110001;
assign LUT_3[22224] = 32'b00000000000000011000010000110111;
assign LUT_3[22225] = 32'b00000000000000011110111100010100;
assign LUT_3[22226] = 32'b00000000000000011010011000011011;
assign LUT_3[22227] = 32'b00000000000000100001000011111000;
assign LUT_3[22228] = 32'b00000000000000010101011110101101;
assign LUT_3[22229] = 32'b00000000000000011100001010001010;
assign LUT_3[22230] = 32'b00000000000000010111100110010001;
assign LUT_3[22231] = 32'b00000000000000011110010001101110;
assign LUT_3[22232] = 32'b00000000000000011101101001111101;
assign LUT_3[22233] = 32'b00000000000000100100010101011010;
assign LUT_3[22234] = 32'b00000000000000011111110001100001;
assign LUT_3[22235] = 32'b00000000000000100110011100111110;
assign LUT_3[22236] = 32'b00000000000000011010110111110011;
assign LUT_3[22237] = 32'b00000000000000100001100011010000;
assign LUT_3[22238] = 32'b00000000000000011100111111010111;
assign LUT_3[22239] = 32'b00000000000000100011101010110100;
assign LUT_3[22240] = 32'b00000000000000010110001100010100;
assign LUT_3[22241] = 32'b00000000000000011100110111110001;
assign LUT_3[22242] = 32'b00000000000000011000010011111000;
assign LUT_3[22243] = 32'b00000000000000011110111111010101;
assign LUT_3[22244] = 32'b00000000000000010011011010001010;
assign LUT_3[22245] = 32'b00000000000000011010000101100111;
assign LUT_3[22246] = 32'b00000000000000010101100001101110;
assign LUT_3[22247] = 32'b00000000000000011100001101001011;
assign LUT_3[22248] = 32'b00000000000000011011100101011010;
assign LUT_3[22249] = 32'b00000000000000100010010000110111;
assign LUT_3[22250] = 32'b00000000000000011101101100111110;
assign LUT_3[22251] = 32'b00000000000000100100011000011011;
assign LUT_3[22252] = 32'b00000000000000011000110011010000;
assign LUT_3[22253] = 32'b00000000000000011111011110101101;
assign LUT_3[22254] = 32'b00000000000000011010111010110100;
assign LUT_3[22255] = 32'b00000000000000100001100110010001;
assign LUT_3[22256] = 32'b00000000000000011001011111010111;
assign LUT_3[22257] = 32'b00000000000000100000001010110100;
assign LUT_3[22258] = 32'b00000000000000011011100110111011;
assign LUT_3[22259] = 32'b00000000000000100010010010011000;
assign LUT_3[22260] = 32'b00000000000000010110101101001101;
assign LUT_3[22261] = 32'b00000000000000011101011000101010;
assign LUT_3[22262] = 32'b00000000000000011000110100110001;
assign LUT_3[22263] = 32'b00000000000000011111100000001110;
assign LUT_3[22264] = 32'b00000000000000011110111000011101;
assign LUT_3[22265] = 32'b00000000000000100101100011111010;
assign LUT_3[22266] = 32'b00000000000000100001000000000001;
assign LUT_3[22267] = 32'b00000000000000100111101011011110;
assign LUT_3[22268] = 32'b00000000000000011100000110010011;
assign LUT_3[22269] = 32'b00000000000000100010110001110000;
assign LUT_3[22270] = 32'b00000000000000011110001101110111;
assign LUT_3[22271] = 32'b00000000000000100100111001010100;
assign LUT_3[22272] = 32'b00000000000000001111001001101100;
assign LUT_3[22273] = 32'b00000000000000010101110101001001;
assign LUT_3[22274] = 32'b00000000000000010001010001010000;
assign LUT_3[22275] = 32'b00000000000000010111111100101101;
assign LUT_3[22276] = 32'b00000000000000001100010111100010;
assign LUT_3[22277] = 32'b00000000000000010011000010111111;
assign LUT_3[22278] = 32'b00000000000000001110011111000110;
assign LUT_3[22279] = 32'b00000000000000010101001010100011;
assign LUT_3[22280] = 32'b00000000000000010100100010110010;
assign LUT_3[22281] = 32'b00000000000000011011001110001111;
assign LUT_3[22282] = 32'b00000000000000010110101010010110;
assign LUT_3[22283] = 32'b00000000000000011101010101110011;
assign LUT_3[22284] = 32'b00000000000000010001110000101000;
assign LUT_3[22285] = 32'b00000000000000011000011100000101;
assign LUT_3[22286] = 32'b00000000000000010011111000001100;
assign LUT_3[22287] = 32'b00000000000000011010100011101001;
assign LUT_3[22288] = 32'b00000000000000010010011100101111;
assign LUT_3[22289] = 32'b00000000000000011001001000001100;
assign LUT_3[22290] = 32'b00000000000000010100100100010011;
assign LUT_3[22291] = 32'b00000000000000011011001111110000;
assign LUT_3[22292] = 32'b00000000000000001111101010100101;
assign LUT_3[22293] = 32'b00000000000000010110010110000010;
assign LUT_3[22294] = 32'b00000000000000010001110010001001;
assign LUT_3[22295] = 32'b00000000000000011000011101100110;
assign LUT_3[22296] = 32'b00000000000000010111110101110101;
assign LUT_3[22297] = 32'b00000000000000011110100001010010;
assign LUT_3[22298] = 32'b00000000000000011001111101011001;
assign LUT_3[22299] = 32'b00000000000000100000101000110110;
assign LUT_3[22300] = 32'b00000000000000010101000011101011;
assign LUT_3[22301] = 32'b00000000000000011011101111001000;
assign LUT_3[22302] = 32'b00000000000000010111001011001111;
assign LUT_3[22303] = 32'b00000000000000011101110110101100;
assign LUT_3[22304] = 32'b00000000000000010000011000001100;
assign LUT_3[22305] = 32'b00000000000000010111000011101001;
assign LUT_3[22306] = 32'b00000000000000010010011111110000;
assign LUT_3[22307] = 32'b00000000000000011001001011001101;
assign LUT_3[22308] = 32'b00000000000000001101100110000010;
assign LUT_3[22309] = 32'b00000000000000010100010001011111;
assign LUT_3[22310] = 32'b00000000000000001111101101100110;
assign LUT_3[22311] = 32'b00000000000000010110011001000011;
assign LUT_3[22312] = 32'b00000000000000010101110001010010;
assign LUT_3[22313] = 32'b00000000000000011100011100101111;
assign LUT_3[22314] = 32'b00000000000000010111111000110110;
assign LUT_3[22315] = 32'b00000000000000011110100100010011;
assign LUT_3[22316] = 32'b00000000000000010010111111001000;
assign LUT_3[22317] = 32'b00000000000000011001101010100101;
assign LUT_3[22318] = 32'b00000000000000010101000110101100;
assign LUT_3[22319] = 32'b00000000000000011011110010001001;
assign LUT_3[22320] = 32'b00000000000000010011101011001111;
assign LUT_3[22321] = 32'b00000000000000011010010110101100;
assign LUT_3[22322] = 32'b00000000000000010101110010110011;
assign LUT_3[22323] = 32'b00000000000000011100011110010000;
assign LUT_3[22324] = 32'b00000000000000010000111001000101;
assign LUT_3[22325] = 32'b00000000000000010111100100100010;
assign LUT_3[22326] = 32'b00000000000000010011000000101001;
assign LUT_3[22327] = 32'b00000000000000011001101100000110;
assign LUT_3[22328] = 32'b00000000000000011001000100010101;
assign LUT_3[22329] = 32'b00000000000000011111101111110010;
assign LUT_3[22330] = 32'b00000000000000011011001011111001;
assign LUT_3[22331] = 32'b00000000000000100001110111010110;
assign LUT_3[22332] = 32'b00000000000000010110010010001011;
assign LUT_3[22333] = 32'b00000000000000011100111101101000;
assign LUT_3[22334] = 32'b00000000000000011000011001101111;
assign LUT_3[22335] = 32'b00000000000000011111000101001100;
assign LUT_3[22336] = 32'b00000000000000001111000010010111;
assign LUT_3[22337] = 32'b00000000000000010101101101110100;
assign LUT_3[22338] = 32'b00000000000000010001001001111011;
assign LUT_3[22339] = 32'b00000000000000010111110101011000;
assign LUT_3[22340] = 32'b00000000000000001100010000001101;
assign LUT_3[22341] = 32'b00000000000000010010111011101010;
assign LUT_3[22342] = 32'b00000000000000001110010111110001;
assign LUT_3[22343] = 32'b00000000000000010101000011001110;
assign LUT_3[22344] = 32'b00000000000000010100011011011101;
assign LUT_3[22345] = 32'b00000000000000011011000110111010;
assign LUT_3[22346] = 32'b00000000000000010110100011000001;
assign LUT_3[22347] = 32'b00000000000000011101001110011110;
assign LUT_3[22348] = 32'b00000000000000010001101001010011;
assign LUT_3[22349] = 32'b00000000000000011000010100110000;
assign LUT_3[22350] = 32'b00000000000000010011110000110111;
assign LUT_3[22351] = 32'b00000000000000011010011100010100;
assign LUT_3[22352] = 32'b00000000000000010010010101011010;
assign LUT_3[22353] = 32'b00000000000000011001000000110111;
assign LUT_3[22354] = 32'b00000000000000010100011100111110;
assign LUT_3[22355] = 32'b00000000000000011011001000011011;
assign LUT_3[22356] = 32'b00000000000000001111100011010000;
assign LUT_3[22357] = 32'b00000000000000010110001110101101;
assign LUT_3[22358] = 32'b00000000000000010001101010110100;
assign LUT_3[22359] = 32'b00000000000000011000010110010001;
assign LUT_3[22360] = 32'b00000000000000010111101110100000;
assign LUT_3[22361] = 32'b00000000000000011110011001111101;
assign LUT_3[22362] = 32'b00000000000000011001110110000100;
assign LUT_3[22363] = 32'b00000000000000100000100001100001;
assign LUT_3[22364] = 32'b00000000000000010100111100010110;
assign LUT_3[22365] = 32'b00000000000000011011100111110011;
assign LUT_3[22366] = 32'b00000000000000010111000011111010;
assign LUT_3[22367] = 32'b00000000000000011101101111010111;
assign LUT_3[22368] = 32'b00000000000000010000010000110111;
assign LUT_3[22369] = 32'b00000000000000010110111100010100;
assign LUT_3[22370] = 32'b00000000000000010010011000011011;
assign LUT_3[22371] = 32'b00000000000000011001000011111000;
assign LUT_3[22372] = 32'b00000000000000001101011110101101;
assign LUT_3[22373] = 32'b00000000000000010100001010001010;
assign LUT_3[22374] = 32'b00000000000000001111100110010001;
assign LUT_3[22375] = 32'b00000000000000010110010001101110;
assign LUT_3[22376] = 32'b00000000000000010101101001111101;
assign LUT_3[22377] = 32'b00000000000000011100010101011010;
assign LUT_3[22378] = 32'b00000000000000010111110001100001;
assign LUT_3[22379] = 32'b00000000000000011110011100111110;
assign LUT_3[22380] = 32'b00000000000000010010110111110011;
assign LUT_3[22381] = 32'b00000000000000011001100011010000;
assign LUT_3[22382] = 32'b00000000000000010100111111010111;
assign LUT_3[22383] = 32'b00000000000000011011101010110100;
assign LUT_3[22384] = 32'b00000000000000010011100011111010;
assign LUT_3[22385] = 32'b00000000000000011010001111010111;
assign LUT_3[22386] = 32'b00000000000000010101101011011110;
assign LUT_3[22387] = 32'b00000000000000011100010110111011;
assign LUT_3[22388] = 32'b00000000000000010000110001110000;
assign LUT_3[22389] = 32'b00000000000000010111011101001101;
assign LUT_3[22390] = 32'b00000000000000010010111001010100;
assign LUT_3[22391] = 32'b00000000000000011001100100110001;
assign LUT_3[22392] = 32'b00000000000000011000111101000000;
assign LUT_3[22393] = 32'b00000000000000011111101000011101;
assign LUT_3[22394] = 32'b00000000000000011011000100100100;
assign LUT_3[22395] = 32'b00000000000000100001110000000001;
assign LUT_3[22396] = 32'b00000000000000010110001010110110;
assign LUT_3[22397] = 32'b00000000000000011100110110010011;
assign LUT_3[22398] = 32'b00000000000000011000010010011010;
assign LUT_3[22399] = 32'b00000000000000011110111101110111;
assign LUT_3[22400] = 32'b00000000000000010001010100101010;
assign LUT_3[22401] = 32'b00000000000000011000000000000111;
assign LUT_3[22402] = 32'b00000000000000010011011100001110;
assign LUT_3[22403] = 32'b00000000000000011010000111101011;
assign LUT_3[22404] = 32'b00000000000000001110100010100000;
assign LUT_3[22405] = 32'b00000000000000010101001101111101;
assign LUT_3[22406] = 32'b00000000000000010000101010000100;
assign LUT_3[22407] = 32'b00000000000000010111010101100001;
assign LUT_3[22408] = 32'b00000000000000010110101101110000;
assign LUT_3[22409] = 32'b00000000000000011101011001001101;
assign LUT_3[22410] = 32'b00000000000000011000110101010100;
assign LUT_3[22411] = 32'b00000000000000011111100000110001;
assign LUT_3[22412] = 32'b00000000000000010011111011100110;
assign LUT_3[22413] = 32'b00000000000000011010100111000011;
assign LUT_3[22414] = 32'b00000000000000010110000011001010;
assign LUT_3[22415] = 32'b00000000000000011100101110100111;
assign LUT_3[22416] = 32'b00000000000000010100100111101101;
assign LUT_3[22417] = 32'b00000000000000011011010011001010;
assign LUT_3[22418] = 32'b00000000000000010110101111010001;
assign LUT_3[22419] = 32'b00000000000000011101011010101110;
assign LUT_3[22420] = 32'b00000000000000010001110101100011;
assign LUT_3[22421] = 32'b00000000000000011000100001000000;
assign LUT_3[22422] = 32'b00000000000000010011111101000111;
assign LUT_3[22423] = 32'b00000000000000011010101000100100;
assign LUT_3[22424] = 32'b00000000000000011010000000110011;
assign LUT_3[22425] = 32'b00000000000000100000101100010000;
assign LUT_3[22426] = 32'b00000000000000011100001000010111;
assign LUT_3[22427] = 32'b00000000000000100010110011110100;
assign LUT_3[22428] = 32'b00000000000000010111001110101001;
assign LUT_3[22429] = 32'b00000000000000011101111010000110;
assign LUT_3[22430] = 32'b00000000000000011001010110001101;
assign LUT_3[22431] = 32'b00000000000000100000000001101010;
assign LUT_3[22432] = 32'b00000000000000010010100011001010;
assign LUT_3[22433] = 32'b00000000000000011001001110100111;
assign LUT_3[22434] = 32'b00000000000000010100101010101110;
assign LUT_3[22435] = 32'b00000000000000011011010110001011;
assign LUT_3[22436] = 32'b00000000000000001111110001000000;
assign LUT_3[22437] = 32'b00000000000000010110011100011101;
assign LUT_3[22438] = 32'b00000000000000010001111000100100;
assign LUT_3[22439] = 32'b00000000000000011000100100000001;
assign LUT_3[22440] = 32'b00000000000000010111111100010000;
assign LUT_3[22441] = 32'b00000000000000011110100111101101;
assign LUT_3[22442] = 32'b00000000000000011010000011110100;
assign LUT_3[22443] = 32'b00000000000000100000101111010001;
assign LUT_3[22444] = 32'b00000000000000010101001010000110;
assign LUT_3[22445] = 32'b00000000000000011011110101100011;
assign LUT_3[22446] = 32'b00000000000000010111010001101010;
assign LUT_3[22447] = 32'b00000000000000011101111101000111;
assign LUT_3[22448] = 32'b00000000000000010101110110001101;
assign LUT_3[22449] = 32'b00000000000000011100100001101010;
assign LUT_3[22450] = 32'b00000000000000010111111101110001;
assign LUT_3[22451] = 32'b00000000000000011110101001001110;
assign LUT_3[22452] = 32'b00000000000000010011000100000011;
assign LUT_3[22453] = 32'b00000000000000011001101111100000;
assign LUT_3[22454] = 32'b00000000000000010101001011100111;
assign LUT_3[22455] = 32'b00000000000000011011110111000100;
assign LUT_3[22456] = 32'b00000000000000011011001111010011;
assign LUT_3[22457] = 32'b00000000000000100001111010110000;
assign LUT_3[22458] = 32'b00000000000000011101010110110111;
assign LUT_3[22459] = 32'b00000000000000100100000010010100;
assign LUT_3[22460] = 32'b00000000000000011000011101001001;
assign LUT_3[22461] = 32'b00000000000000011111001000100110;
assign LUT_3[22462] = 32'b00000000000000011010100100101101;
assign LUT_3[22463] = 32'b00000000000000100001010000001010;
assign LUT_3[22464] = 32'b00000000000000010001001101010101;
assign LUT_3[22465] = 32'b00000000000000010111111000110010;
assign LUT_3[22466] = 32'b00000000000000010011010100111001;
assign LUT_3[22467] = 32'b00000000000000011010000000010110;
assign LUT_3[22468] = 32'b00000000000000001110011011001011;
assign LUT_3[22469] = 32'b00000000000000010101000110101000;
assign LUT_3[22470] = 32'b00000000000000010000100010101111;
assign LUT_3[22471] = 32'b00000000000000010111001110001100;
assign LUT_3[22472] = 32'b00000000000000010110100110011011;
assign LUT_3[22473] = 32'b00000000000000011101010001111000;
assign LUT_3[22474] = 32'b00000000000000011000101101111111;
assign LUT_3[22475] = 32'b00000000000000011111011001011100;
assign LUT_3[22476] = 32'b00000000000000010011110100010001;
assign LUT_3[22477] = 32'b00000000000000011010011111101110;
assign LUT_3[22478] = 32'b00000000000000010101111011110101;
assign LUT_3[22479] = 32'b00000000000000011100100111010010;
assign LUT_3[22480] = 32'b00000000000000010100100000011000;
assign LUT_3[22481] = 32'b00000000000000011011001011110101;
assign LUT_3[22482] = 32'b00000000000000010110100111111100;
assign LUT_3[22483] = 32'b00000000000000011101010011011001;
assign LUT_3[22484] = 32'b00000000000000010001101110001110;
assign LUT_3[22485] = 32'b00000000000000011000011001101011;
assign LUT_3[22486] = 32'b00000000000000010011110101110010;
assign LUT_3[22487] = 32'b00000000000000011010100001001111;
assign LUT_3[22488] = 32'b00000000000000011001111001011110;
assign LUT_3[22489] = 32'b00000000000000100000100100111011;
assign LUT_3[22490] = 32'b00000000000000011100000001000010;
assign LUT_3[22491] = 32'b00000000000000100010101100011111;
assign LUT_3[22492] = 32'b00000000000000010111000111010100;
assign LUT_3[22493] = 32'b00000000000000011101110010110001;
assign LUT_3[22494] = 32'b00000000000000011001001110111000;
assign LUT_3[22495] = 32'b00000000000000011111111010010101;
assign LUT_3[22496] = 32'b00000000000000010010011011110101;
assign LUT_3[22497] = 32'b00000000000000011001000111010010;
assign LUT_3[22498] = 32'b00000000000000010100100011011001;
assign LUT_3[22499] = 32'b00000000000000011011001110110110;
assign LUT_3[22500] = 32'b00000000000000001111101001101011;
assign LUT_3[22501] = 32'b00000000000000010110010101001000;
assign LUT_3[22502] = 32'b00000000000000010001110001001111;
assign LUT_3[22503] = 32'b00000000000000011000011100101100;
assign LUT_3[22504] = 32'b00000000000000010111110100111011;
assign LUT_3[22505] = 32'b00000000000000011110100000011000;
assign LUT_3[22506] = 32'b00000000000000011001111100011111;
assign LUT_3[22507] = 32'b00000000000000100000100111111100;
assign LUT_3[22508] = 32'b00000000000000010101000010110001;
assign LUT_3[22509] = 32'b00000000000000011011101110001110;
assign LUT_3[22510] = 32'b00000000000000010111001010010101;
assign LUT_3[22511] = 32'b00000000000000011101110101110010;
assign LUT_3[22512] = 32'b00000000000000010101101110111000;
assign LUT_3[22513] = 32'b00000000000000011100011010010101;
assign LUT_3[22514] = 32'b00000000000000010111110110011100;
assign LUT_3[22515] = 32'b00000000000000011110100001111001;
assign LUT_3[22516] = 32'b00000000000000010010111100101110;
assign LUT_3[22517] = 32'b00000000000000011001101000001011;
assign LUT_3[22518] = 32'b00000000000000010101000100010010;
assign LUT_3[22519] = 32'b00000000000000011011101111101111;
assign LUT_3[22520] = 32'b00000000000000011011000111111110;
assign LUT_3[22521] = 32'b00000000000000100001110011011011;
assign LUT_3[22522] = 32'b00000000000000011101001111100010;
assign LUT_3[22523] = 32'b00000000000000100011111010111111;
assign LUT_3[22524] = 32'b00000000000000011000010101110100;
assign LUT_3[22525] = 32'b00000000000000011111000001010001;
assign LUT_3[22526] = 32'b00000000000000011010011101011000;
assign LUT_3[22527] = 32'b00000000000000100001001000110101;
assign LUT_3[22528] = 32'b00000000000000001010110110010000;
assign LUT_3[22529] = 32'b00000000000000010001100001101101;
assign LUT_3[22530] = 32'b00000000000000001100111101110100;
assign LUT_3[22531] = 32'b00000000000000010011101001010001;
assign LUT_3[22532] = 32'b00000000000000001000000100000110;
assign LUT_3[22533] = 32'b00000000000000001110101111100011;
assign LUT_3[22534] = 32'b00000000000000001010001011101010;
assign LUT_3[22535] = 32'b00000000000000010000110111000111;
assign LUT_3[22536] = 32'b00000000000000010000001111010110;
assign LUT_3[22537] = 32'b00000000000000010110111010110011;
assign LUT_3[22538] = 32'b00000000000000010010010110111010;
assign LUT_3[22539] = 32'b00000000000000011001000010010111;
assign LUT_3[22540] = 32'b00000000000000001101011101001100;
assign LUT_3[22541] = 32'b00000000000000010100001000101001;
assign LUT_3[22542] = 32'b00000000000000001111100100110000;
assign LUT_3[22543] = 32'b00000000000000010110010000001101;
assign LUT_3[22544] = 32'b00000000000000001110001001010011;
assign LUT_3[22545] = 32'b00000000000000010100110100110000;
assign LUT_3[22546] = 32'b00000000000000010000010000110111;
assign LUT_3[22547] = 32'b00000000000000010110111100010100;
assign LUT_3[22548] = 32'b00000000000000001011010111001001;
assign LUT_3[22549] = 32'b00000000000000010010000010100110;
assign LUT_3[22550] = 32'b00000000000000001101011110101101;
assign LUT_3[22551] = 32'b00000000000000010100001010001010;
assign LUT_3[22552] = 32'b00000000000000010011100010011001;
assign LUT_3[22553] = 32'b00000000000000011010001101110110;
assign LUT_3[22554] = 32'b00000000000000010101101001111101;
assign LUT_3[22555] = 32'b00000000000000011100010101011010;
assign LUT_3[22556] = 32'b00000000000000010000110000001111;
assign LUT_3[22557] = 32'b00000000000000010111011011101100;
assign LUT_3[22558] = 32'b00000000000000010010110111110011;
assign LUT_3[22559] = 32'b00000000000000011001100011010000;
assign LUT_3[22560] = 32'b00000000000000001100000100110000;
assign LUT_3[22561] = 32'b00000000000000010010110000001101;
assign LUT_3[22562] = 32'b00000000000000001110001100010100;
assign LUT_3[22563] = 32'b00000000000000010100110111110001;
assign LUT_3[22564] = 32'b00000000000000001001010010100110;
assign LUT_3[22565] = 32'b00000000000000001111111110000011;
assign LUT_3[22566] = 32'b00000000000000001011011010001010;
assign LUT_3[22567] = 32'b00000000000000010010000101100111;
assign LUT_3[22568] = 32'b00000000000000010001011101110110;
assign LUT_3[22569] = 32'b00000000000000011000001001010011;
assign LUT_3[22570] = 32'b00000000000000010011100101011010;
assign LUT_3[22571] = 32'b00000000000000011010010000110111;
assign LUT_3[22572] = 32'b00000000000000001110101011101100;
assign LUT_3[22573] = 32'b00000000000000010101010111001001;
assign LUT_3[22574] = 32'b00000000000000010000110011010000;
assign LUT_3[22575] = 32'b00000000000000010111011110101101;
assign LUT_3[22576] = 32'b00000000000000001111010111110011;
assign LUT_3[22577] = 32'b00000000000000010110000011010000;
assign LUT_3[22578] = 32'b00000000000000010001011111010111;
assign LUT_3[22579] = 32'b00000000000000011000001010110100;
assign LUT_3[22580] = 32'b00000000000000001100100101101001;
assign LUT_3[22581] = 32'b00000000000000010011010001000110;
assign LUT_3[22582] = 32'b00000000000000001110101101001101;
assign LUT_3[22583] = 32'b00000000000000010101011000101010;
assign LUT_3[22584] = 32'b00000000000000010100110000111001;
assign LUT_3[22585] = 32'b00000000000000011011011100010110;
assign LUT_3[22586] = 32'b00000000000000010110111000011101;
assign LUT_3[22587] = 32'b00000000000000011101100011111010;
assign LUT_3[22588] = 32'b00000000000000010001111110101111;
assign LUT_3[22589] = 32'b00000000000000011000101010001100;
assign LUT_3[22590] = 32'b00000000000000010100000110010011;
assign LUT_3[22591] = 32'b00000000000000011010110001110000;
assign LUT_3[22592] = 32'b00000000000000001010101110111011;
assign LUT_3[22593] = 32'b00000000000000010001011010011000;
assign LUT_3[22594] = 32'b00000000000000001100110110011111;
assign LUT_3[22595] = 32'b00000000000000010011100001111100;
assign LUT_3[22596] = 32'b00000000000000000111111100110001;
assign LUT_3[22597] = 32'b00000000000000001110101000001110;
assign LUT_3[22598] = 32'b00000000000000001010000100010101;
assign LUT_3[22599] = 32'b00000000000000010000101111110010;
assign LUT_3[22600] = 32'b00000000000000010000001000000001;
assign LUT_3[22601] = 32'b00000000000000010110110011011110;
assign LUT_3[22602] = 32'b00000000000000010010001111100101;
assign LUT_3[22603] = 32'b00000000000000011000111011000010;
assign LUT_3[22604] = 32'b00000000000000001101010101110111;
assign LUT_3[22605] = 32'b00000000000000010100000001010100;
assign LUT_3[22606] = 32'b00000000000000001111011101011011;
assign LUT_3[22607] = 32'b00000000000000010110001000111000;
assign LUT_3[22608] = 32'b00000000000000001110000001111110;
assign LUT_3[22609] = 32'b00000000000000010100101101011011;
assign LUT_3[22610] = 32'b00000000000000010000001001100010;
assign LUT_3[22611] = 32'b00000000000000010110110100111111;
assign LUT_3[22612] = 32'b00000000000000001011001111110100;
assign LUT_3[22613] = 32'b00000000000000010001111011010001;
assign LUT_3[22614] = 32'b00000000000000001101010111011000;
assign LUT_3[22615] = 32'b00000000000000010100000010110101;
assign LUT_3[22616] = 32'b00000000000000010011011011000100;
assign LUT_3[22617] = 32'b00000000000000011010000110100001;
assign LUT_3[22618] = 32'b00000000000000010101100010101000;
assign LUT_3[22619] = 32'b00000000000000011100001110000101;
assign LUT_3[22620] = 32'b00000000000000010000101000111010;
assign LUT_3[22621] = 32'b00000000000000010111010100010111;
assign LUT_3[22622] = 32'b00000000000000010010110000011110;
assign LUT_3[22623] = 32'b00000000000000011001011011111011;
assign LUT_3[22624] = 32'b00000000000000001011111101011011;
assign LUT_3[22625] = 32'b00000000000000010010101000111000;
assign LUT_3[22626] = 32'b00000000000000001110000100111111;
assign LUT_3[22627] = 32'b00000000000000010100110000011100;
assign LUT_3[22628] = 32'b00000000000000001001001011010001;
assign LUT_3[22629] = 32'b00000000000000001111110110101110;
assign LUT_3[22630] = 32'b00000000000000001011010010110101;
assign LUT_3[22631] = 32'b00000000000000010001111110010010;
assign LUT_3[22632] = 32'b00000000000000010001010110100001;
assign LUT_3[22633] = 32'b00000000000000011000000001111110;
assign LUT_3[22634] = 32'b00000000000000010011011110000101;
assign LUT_3[22635] = 32'b00000000000000011010001001100010;
assign LUT_3[22636] = 32'b00000000000000001110100100010111;
assign LUT_3[22637] = 32'b00000000000000010101001111110100;
assign LUT_3[22638] = 32'b00000000000000010000101011111011;
assign LUT_3[22639] = 32'b00000000000000010111010111011000;
assign LUT_3[22640] = 32'b00000000000000001111010000011110;
assign LUT_3[22641] = 32'b00000000000000010101111011111011;
assign LUT_3[22642] = 32'b00000000000000010001011000000010;
assign LUT_3[22643] = 32'b00000000000000011000000011011111;
assign LUT_3[22644] = 32'b00000000000000001100011110010100;
assign LUT_3[22645] = 32'b00000000000000010011001001110001;
assign LUT_3[22646] = 32'b00000000000000001110100101111000;
assign LUT_3[22647] = 32'b00000000000000010101010001010101;
assign LUT_3[22648] = 32'b00000000000000010100101001100100;
assign LUT_3[22649] = 32'b00000000000000011011010101000001;
assign LUT_3[22650] = 32'b00000000000000010110110001001000;
assign LUT_3[22651] = 32'b00000000000000011101011100100101;
assign LUT_3[22652] = 32'b00000000000000010001110111011010;
assign LUT_3[22653] = 32'b00000000000000011000100010110111;
assign LUT_3[22654] = 32'b00000000000000010011111110111110;
assign LUT_3[22655] = 32'b00000000000000011010101010011011;
assign LUT_3[22656] = 32'b00000000000000001101000001001110;
assign LUT_3[22657] = 32'b00000000000000010011101100101011;
assign LUT_3[22658] = 32'b00000000000000001111001000110010;
assign LUT_3[22659] = 32'b00000000000000010101110100001111;
assign LUT_3[22660] = 32'b00000000000000001010001111000100;
assign LUT_3[22661] = 32'b00000000000000010000111010100001;
assign LUT_3[22662] = 32'b00000000000000001100010110101000;
assign LUT_3[22663] = 32'b00000000000000010011000010000101;
assign LUT_3[22664] = 32'b00000000000000010010011010010100;
assign LUT_3[22665] = 32'b00000000000000011001000101110001;
assign LUT_3[22666] = 32'b00000000000000010100100001111000;
assign LUT_3[22667] = 32'b00000000000000011011001101010101;
assign LUT_3[22668] = 32'b00000000000000001111101000001010;
assign LUT_3[22669] = 32'b00000000000000010110010011100111;
assign LUT_3[22670] = 32'b00000000000000010001101111101110;
assign LUT_3[22671] = 32'b00000000000000011000011011001011;
assign LUT_3[22672] = 32'b00000000000000010000010100010001;
assign LUT_3[22673] = 32'b00000000000000010110111111101110;
assign LUT_3[22674] = 32'b00000000000000010010011011110101;
assign LUT_3[22675] = 32'b00000000000000011001000111010010;
assign LUT_3[22676] = 32'b00000000000000001101100010000111;
assign LUT_3[22677] = 32'b00000000000000010100001101100100;
assign LUT_3[22678] = 32'b00000000000000001111101001101011;
assign LUT_3[22679] = 32'b00000000000000010110010101001000;
assign LUT_3[22680] = 32'b00000000000000010101101101010111;
assign LUT_3[22681] = 32'b00000000000000011100011000110100;
assign LUT_3[22682] = 32'b00000000000000010111110100111011;
assign LUT_3[22683] = 32'b00000000000000011110100000011000;
assign LUT_3[22684] = 32'b00000000000000010010111011001101;
assign LUT_3[22685] = 32'b00000000000000011001100110101010;
assign LUT_3[22686] = 32'b00000000000000010101000010110001;
assign LUT_3[22687] = 32'b00000000000000011011101110001110;
assign LUT_3[22688] = 32'b00000000000000001110001111101110;
assign LUT_3[22689] = 32'b00000000000000010100111011001011;
assign LUT_3[22690] = 32'b00000000000000010000010111010010;
assign LUT_3[22691] = 32'b00000000000000010111000010101111;
assign LUT_3[22692] = 32'b00000000000000001011011101100100;
assign LUT_3[22693] = 32'b00000000000000010010001001000001;
assign LUT_3[22694] = 32'b00000000000000001101100101001000;
assign LUT_3[22695] = 32'b00000000000000010100010000100101;
assign LUT_3[22696] = 32'b00000000000000010011101000110100;
assign LUT_3[22697] = 32'b00000000000000011010010100010001;
assign LUT_3[22698] = 32'b00000000000000010101110000011000;
assign LUT_3[22699] = 32'b00000000000000011100011011110101;
assign LUT_3[22700] = 32'b00000000000000010000110110101010;
assign LUT_3[22701] = 32'b00000000000000010111100010000111;
assign LUT_3[22702] = 32'b00000000000000010010111110001110;
assign LUT_3[22703] = 32'b00000000000000011001101001101011;
assign LUT_3[22704] = 32'b00000000000000010001100010110001;
assign LUT_3[22705] = 32'b00000000000000011000001110001110;
assign LUT_3[22706] = 32'b00000000000000010011101010010101;
assign LUT_3[22707] = 32'b00000000000000011010010101110010;
assign LUT_3[22708] = 32'b00000000000000001110110000100111;
assign LUT_3[22709] = 32'b00000000000000010101011100000100;
assign LUT_3[22710] = 32'b00000000000000010000111000001011;
assign LUT_3[22711] = 32'b00000000000000010111100011101000;
assign LUT_3[22712] = 32'b00000000000000010110111011110111;
assign LUT_3[22713] = 32'b00000000000000011101100111010100;
assign LUT_3[22714] = 32'b00000000000000011001000011011011;
assign LUT_3[22715] = 32'b00000000000000011111101110111000;
assign LUT_3[22716] = 32'b00000000000000010100001001101101;
assign LUT_3[22717] = 32'b00000000000000011010110101001010;
assign LUT_3[22718] = 32'b00000000000000010110010001010001;
assign LUT_3[22719] = 32'b00000000000000011100111100101110;
assign LUT_3[22720] = 32'b00000000000000001100111001111001;
assign LUT_3[22721] = 32'b00000000000000010011100101010110;
assign LUT_3[22722] = 32'b00000000000000001111000001011101;
assign LUT_3[22723] = 32'b00000000000000010101101100111010;
assign LUT_3[22724] = 32'b00000000000000001010000111101111;
assign LUT_3[22725] = 32'b00000000000000010000110011001100;
assign LUT_3[22726] = 32'b00000000000000001100001111010011;
assign LUT_3[22727] = 32'b00000000000000010010111010110000;
assign LUT_3[22728] = 32'b00000000000000010010010010111111;
assign LUT_3[22729] = 32'b00000000000000011000111110011100;
assign LUT_3[22730] = 32'b00000000000000010100011010100011;
assign LUT_3[22731] = 32'b00000000000000011011000110000000;
assign LUT_3[22732] = 32'b00000000000000001111100000110101;
assign LUT_3[22733] = 32'b00000000000000010110001100010010;
assign LUT_3[22734] = 32'b00000000000000010001101000011001;
assign LUT_3[22735] = 32'b00000000000000011000010011110110;
assign LUT_3[22736] = 32'b00000000000000010000001100111100;
assign LUT_3[22737] = 32'b00000000000000010110111000011001;
assign LUT_3[22738] = 32'b00000000000000010010010100100000;
assign LUT_3[22739] = 32'b00000000000000011000111111111101;
assign LUT_3[22740] = 32'b00000000000000001101011010110010;
assign LUT_3[22741] = 32'b00000000000000010100000110001111;
assign LUT_3[22742] = 32'b00000000000000001111100010010110;
assign LUT_3[22743] = 32'b00000000000000010110001101110011;
assign LUT_3[22744] = 32'b00000000000000010101100110000010;
assign LUT_3[22745] = 32'b00000000000000011100010001011111;
assign LUT_3[22746] = 32'b00000000000000010111101101100110;
assign LUT_3[22747] = 32'b00000000000000011110011001000011;
assign LUT_3[22748] = 32'b00000000000000010010110011111000;
assign LUT_3[22749] = 32'b00000000000000011001011111010101;
assign LUT_3[22750] = 32'b00000000000000010100111011011100;
assign LUT_3[22751] = 32'b00000000000000011011100110111001;
assign LUT_3[22752] = 32'b00000000000000001110001000011001;
assign LUT_3[22753] = 32'b00000000000000010100110011110110;
assign LUT_3[22754] = 32'b00000000000000010000001111111101;
assign LUT_3[22755] = 32'b00000000000000010110111011011010;
assign LUT_3[22756] = 32'b00000000000000001011010110001111;
assign LUT_3[22757] = 32'b00000000000000010010000001101100;
assign LUT_3[22758] = 32'b00000000000000001101011101110011;
assign LUT_3[22759] = 32'b00000000000000010100001001010000;
assign LUT_3[22760] = 32'b00000000000000010011100001011111;
assign LUT_3[22761] = 32'b00000000000000011010001100111100;
assign LUT_3[22762] = 32'b00000000000000010101101001000011;
assign LUT_3[22763] = 32'b00000000000000011100010100100000;
assign LUT_3[22764] = 32'b00000000000000010000101111010101;
assign LUT_3[22765] = 32'b00000000000000010111011010110010;
assign LUT_3[22766] = 32'b00000000000000010010110110111001;
assign LUT_3[22767] = 32'b00000000000000011001100010010110;
assign LUT_3[22768] = 32'b00000000000000010001011011011100;
assign LUT_3[22769] = 32'b00000000000000011000000110111001;
assign LUT_3[22770] = 32'b00000000000000010011100011000000;
assign LUT_3[22771] = 32'b00000000000000011010001110011101;
assign LUT_3[22772] = 32'b00000000000000001110101001010010;
assign LUT_3[22773] = 32'b00000000000000010101010100101111;
assign LUT_3[22774] = 32'b00000000000000010000110000110110;
assign LUT_3[22775] = 32'b00000000000000010111011100010011;
assign LUT_3[22776] = 32'b00000000000000010110110100100010;
assign LUT_3[22777] = 32'b00000000000000011101011111111111;
assign LUT_3[22778] = 32'b00000000000000011000111100000110;
assign LUT_3[22779] = 32'b00000000000000011111100111100011;
assign LUT_3[22780] = 32'b00000000000000010100000010011000;
assign LUT_3[22781] = 32'b00000000000000011010101101110101;
assign LUT_3[22782] = 32'b00000000000000010110001001111100;
assign LUT_3[22783] = 32'b00000000000000011100110101011001;
assign LUT_3[22784] = 32'b00000000000000000111000101110001;
assign LUT_3[22785] = 32'b00000000000000001101110001001110;
assign LUT_3[22786] = 32'b00000000000000001001001101010101;
assign LUT_3[22787] = 32'b00000000000000001111111000110010;
assign LUT_3[22788] = 32'b00000000000000000100010011100111;
assign LUT_3[22789] = 32'b00000000000000001010111111000100;
assign LUT_3[22790] = 32'b00000000000000000110011011001011;
assign LUT_3[22791] = 32'b00000000000000001101000110101000;
assign LUT_3[22792] = 32'b00000000000000001100011110110111;
assign LUT_3[22793] = 32'b00000000000000010011001010010100;
assign LUT_3[22794] = 32'b00000000000000001110100110011011;
assign LUT_3[22795] = 32'b00000000000000010101010001111000;
assign LUT_3[22796] = 32'b00000000000000001001101100101101;
assign LUT_3[22797] = 32'b00000000000000010000011000001010;
assign LUT_3[22798] = 32'b00000000000000001011110100010001;
assign LUT_3[22799] = 32'b00000000000000010010011111101110;
assign LUT_3[22800] = 32'b00000000000000001010011000110100;
assign LUT_3[22801] = 32'b00000000000000010001000100010001;
assign LUT_3[22802] = 32'b00000000000000001100100000011000;
assign LUT_3[22803] = 32'b00000000000000010011001011110101;
assign LUT_3[22804] = 32'b00000000000000000111100110101010;
assign LUT_3[22805] = 32'b00000000000000001110010010000111;
assign LUT_3[22806] = 32'b00000000000000001001101110001110;
assign LUT_3[22807] = 32'b00000000000000010000011001101011;
assign LUT_3[22808] = 32'b00000000000000001111110001111010;
assign LUT_3[22809] = 32'b00000000000000010110011101010111;
assign LUT_3[22810] = 32'b00000000000000010001111001011110;
assign LUT_3[22811] = 32'b00000000000000011000100100111011;
assign LUT_3[22812] = 32'b00000000000000001100111111110000;
assign LUT_3[22813] = 32'b00000000000000010011101011001101;
assign LUT_3[22814] = 32'b00000000000000001111000111010100;
assign LUT_3[22815] = 32'b00000000000000010101110010110001;
assign LUT_3[22816] = 32'b00000000000000001000010100010001;
assign LUT_3[22817] = 32'b00000000000000001110111111101110;
assign LUT_3[22818] = 32'b00000000000000001010011011110101;
assign LUT_3[22819] = 32'b00000000000000010001000111010010;
assign LUT_3[22820] = 32'b00000000000000000101100010000111;
assign LUT_3[22821] = 32'b00000000000000001100001101100100;
assign LUT_3[22822] = 32'b00000000000000000111101001101011;
assign LUT_3[22823] = 32'b00000000000000001110010101001000;
assign LUT_3[22824] = 32'b00000000000000001101101101010111;
assign LUT_3[22825] = 32'b00000000000000010100011000110100;
assign LUT_3[22826] = 32'b00000000000000001111110100111011;
assign LUT_3[22827] = 32'b00000000000000010110100000011000;
assign LUT_3[22828] = 32'b00000000000000001010111011001101;
assign LUT_3[22829] = 32'b00000000000000010001100110101010;
assign LUT_3[22830] = 32'b00000000000000001101000010110001;
assign LUT_3[22831] = 32'b00000000000000010011101110001110;
assign LUT_3[22832] = 32'b00000000000000001011100111010100;
assign LUT_3[22833] = 32'b00000000000000010010010010110001;
assign LUT_3[22834] = 32'b00000000000000001101101110111000;
assign LUT_3[22835] = 32'b00000000000000010100011010010101;
assign LUT_3[22836] = 32'b00000000000000001000110101001010;
assign LUT_3[22837] = 32'b00000000000000001111100000100111;
assign LUT_3[22838] = 32'b00000000000000001010111100101110;
assign LUT_3[22839] = 32'b00000000000000010001101000001011;
assign LUT_3[22840] = 32'b00000000000000010001000000011010;
assign LUT_3[22841] = 32'b00000000000000010111101011110111;
assign LUT_3[22842] = 32'b00000000000000010011000111111110;
assign LUT_3[22843] = 32'b00000000000000011001110011011011;
assign LUT_3[22844] = 32'b00000000000000001110001110010000;
assign LUT_3[22845] = 32'b00000000000000010100111001101101;
assign LUT_3[22846] = 32'b00000000000000010000010101110100;
assign LUT_3[22847] = 32'b00000000000000010111000001010001;
assign LUT_3[22848] = 32'b00000000000000000110111110011100;
assign LUT_3[22849] = 32'b00000000000000001101101001111001;
assign LUT_3[22850] = 32'b00000000000000001001000110000000;
assign LUT_3[22851] = 32'b00000000000000001111110001011101;
assign LUT_3[22852] = 32'b00000000000000000100001100010010;
assign LUT_3[22853] = 32'b00000000000000001010110111101111;
assign LUT_3[22854] = 32'b00000000000000000110010011110110;
assign LUT_3[22855] = 32'b00000000000000001100111111010011;
assign LUT_3[22856] = 32'b00000000000000001100010111100010;
assign LUT_3[22857] = 32'b00000000000000010011000010111111;
assign LUT_3[22858] = 32'b00000000000000001110011111000110;
assign LUT_3[22859] = 32'b00000000000000010101001010100011;
assign LUT_3[22860] = 32'b00000000000000001001100101011000;
assign LUT_3[22861] = 32'b00000000000000010000010000110101;
assign LUT_3[22862] = 32'b00000000000000001011101100111100;
assign LUT_3[22863] = 32'b00000000000000010010011000011001;
assign LUT_3[22864] = 32'b00000000000000001010010001011111;
assign LUT_3[22865] = 32'b00000000000000010000111100111100;
assign LUT_3[22866] = 32'b00000000000000001100011001000011;
assign LUT_3[22867] = 32'b00000000000000010011000100100000;
assign LUT_3[22868] = 32'b00000000000000000111011111010101;
assign LUT_3[22869] = 32'b00000000000000001110001010110010;
assign LUT_3[22870] = 32'b00000000000000001001100110111001;
assign LUT_3[22871] = 32'b00000000000000010000010010010110;
assign LUT_3[22872] = 32'b00000000000000001111101010100101;
assign LUT_3[22873] = 32'b00000000000000010110010110000010;
assign LUT_3[22874] = 32'b00000000000000010001110010001001;
assign LUT_3[22875] = 32'b00000000000000011000011101100110;
assign LUT_3[22876] = 32'b00000000000000001100111000011011;
assign LUT_3[22877] = 32'b00000000000000010011100011111000;
assign LUT_3[22878] = 32'b00000000000000001110111111111111;
assign LUT_3[22879] = 32'b00000000000000010101101011011100;
assign LUT_3[22880] = 32'b00000000000000001000001100111100;
assign LUT_3[22881] = 32'b00000000000000001110111000011001;
assign LUT_3[22882] = 32'b00000000000000001010010100100000;
assign LUT_3[22883] = 32'b00000000000000010000111111111101;
assign LUT_3[22884] = 32'b00000000000000000101011010110010;
assign LUT_3[22885] = 32'b00000000000000001100000110001111;
assign LUT_3[22886] = 32'b00000000000000000111100010010110;
assign LUT_3[22887] = 32'b00000000000000001110001101110011;
assign LUT_3[22888] = 32'b00000000000000001101100110000010;
assign LUT_3[22889] = 32'b00000000000000010100010001011111;
assign LUT_3[22890] = 32'b00000000000000001111101101100110;
assign LUT_3[22891] = 32'b00000000000000010110011001000011;
assign LUT_3[22892] = 32'b00000000000000001010110011111000;
assign LUT_3[22893] = 32'b00000000000000010001011111010101;
assign LUT_3[22894] = 32'b00000000000000001100111011011100;
assign LUT_3[22895] = 32'b00000000000000010011100110111001;
assign LUT_3[22896] = 32'b00000000000000001011011111111111;
assign LUT_3[22897] = 32'b00000000000000010010001011011100;
assign LUT_3[22898] = 32'b00000000000000001101100111100011;
assign LUT_3[22899] = 32'b00000000000000010100010011000000;
assign LUT_3[22900] = 32'b00000000000000001000101101110101;
assign LUT_3[22901] = 32'b00000000000000001111011001010010;
assign LUT_3[22902] = 32'b00000000000000001010110101011001;
assign LUT_3[22903] = 32'b00000000000000010001100000110110;
assign LUT_3[22904] = 32'b00000000000000010000111001000101;
assign LUT_3[22905] = 32'b00000000000000010111100100100010;
assign LUT_3[22906] = 32'b00000000000000010011000000101001;
assign LUT_3[22907] = 32'b00000000000000011001101100000110;
assign LUT_3[22908] = 32'b00000000000000001110000110111011;
assign LUT_3[22909] = 32'b00000000000000010100110010011000;
assign LUT_3[22910] = 32'b00000000000000010000001110011111;
assign LUT_3[22911] = 32'b00000000000000010110111001111100;
assign LUT_3[22912] = 32'b00000000000000001001010000101111;
assign LUT_3[22913] = 32'b00000000000000001111111100001100;
assign LUT_3[22914] = 32'b00000000000000001011011000010011;
assign LUT_3[22915] = 32'b00000000000000010010000011110000;
assign LUT_3[22916] = 32'b00000000000000000110011110100101;
assign LUT_3[22917] = 32'b00000000000000001101001010000010;
assign LUT_3[22918] = 32'b00000000000000001000100110001001;
assign LUT_3[22919] = 32'b00000000000000001111010001100110;
assign LUT_3[22920] = 32'b00000000000000001110101001110101;
assign LUT_3[22921] = 32'b00000000000000010101010101010010;
assign LUT_3[22922] = 32'b00000000000000010000110001011001;
assign LUT_3[22923] = 32'b00000000000000010111011100110110;
assign LUT_3[22924] = 32'b00000000000000001011110111101011;
assign LUT_3[22925] = 32'b00000000000000010010100011001000;
assign LUT_3[22926] = 32'b00000000000000001101111111001111;
assign LUT_3[22927] = 32'b00000000000000010100101010101100;
assign LUT_3[22928] = 32'b00000000000000001100100011110010;
assign LUT_3[22929] = 32'b00000000000000010011001111001111;
assign LUT_3[22930] = 32'b00000000000000001110101011010110;
assign LUT_3[22931] = 32'b00000000000000010101010110110011;
assign LUT_3[22932] = 32'b00000000000000001001110001101000;
assign LUT_3[22933] = 32'b00000000000000010000011101000101;
assign LUT_3[22934] = 32'b00000000000000001011111001001100;
assign LUT_3[22935] = 32'b00000000000000010010100100101001;
assign LUT_3[22936] = 32'b00000000000000010001111100111000;
assign LUT_3[22937] = 32'b00000000000000011000101000010101;
assign LUT_3[22938] = 32'b00000000000000010100000100011100;
assign LUT_3[22939] = 32'b00000000000000011010101111111001;
assign LUT_3[22940] = 32'b00000000000000001111001010101110;
assign LUT_3[22941] = 32'b00000000000000010101110110001011;
assign LUT_3[22942] = 32'b00000000000000010001010010010010;
assign LUT_3[22943] = 32'b00000000000000010111111101101111;
assign LUT_3[22944] = 32'b00000000000000001010011111001111;
assign LUT_3[22945] = 32'b00000000000000010001001010101100;
assign LUT_3[22946] = 32'b00000000000000001100100110110011;
assign LUT_3[22947] = 32'b00000000000000010011010010010000;
assign LUT_3[22948] = 32'b00000000000000000111101101000101;
assign LUT_3[22949] = 32'b00000000000000001110011000100010;
assign LUT_3[22950] = 32'b00000000000000001001110100101001;
assign LUT_3[22951] = 32'b00000000000000010000100000000110;
assign LUT_3[22952] = 32'b00000000000000001111111000010101;
assign LUT_3[22953] = 32'b00000000000000010110100011110010;
assign LUT_3[22954] = 32'b00000000000000010001111111111001;
assign LUT_3[22955] = 32'b00000000000000011000101011010110;
assign LUT_3[22956] = 32'b00000000000000001101000110001011;
assign LUT_3[22957] = 32'b00000000000000010011110001101000;
assign LUT_3[22958] = 32'b00000000000000001111001101101111;
assign LUT_3[22959] = 32'b00000000000000010101111001001100;
assign LUT_3[22960] = 32'b00000000000000001101110010010010;
assign LUT_3[22961] = 32'b00000000000000010100011101101111;
assign LUT_3[22962] = 32'b00000000000000001111111001110110;
assign LUT_3[22963] = 32'b00000000000000010110100101010011;
assign LUT_3[22964] = 32'b00000000000000001011000000001000;
assign LUT_3[22965] = 32'b00000000000000010001101011100101;
assign LUT_3[22966] = 32'b00000000000000001101000111101100;
assign LUT_3[22967] = 32'b00000000000000010011110011001001;
assign LUT_3[22968] = 32'b00000000000000010011001011011000;
assign LUT_3[22969] = 32'b00000000000000011001110110110101;
assign LUT_3[22970] = 32'b00000000000000010101010010111100;
assign LUT_3[22971] = 32'b00000000000000011011111110011001;
assign LUT_3[22972] = 32'b00000000000000010000011001001110;
assign LUT_3[22973] = 32'b00000000000000010111000100101011;
assign LUT_3[22974] = 32'b00000000000000010010100000110010;
assign LUT_3[22975] = 32'b00000000000000011001001100001111;
assign LUT_3[22976] = 32'b00000000000000001001001001011010;
assign LUT_3[22977] = 32'b00000000000000001111110100110111;
assign LUT_3[22978] = 32'b00000000000000001011010000111110;
assign LUT_3[22979] = 32'b00000000000000010001111100011011;
assign LUT_3[22980] = 32'b00000000000000000110010111010000;
assign LUT_3[22981] = 32'b00000000000000001101000010101101;
assign LUT_3[22982] = 32'b00000000000000001000011110110100;
assign LUT_3[22983] = 32'b00000000000000001111001010010001;
assign LUT_3[22984] = 32'b00000000000000001110100010100000;
assign LUT_3[22985] = 32'b00000000000000010101001101111101;
assign LUT_3[22986] = 32'b00000000000000010000101010000100;
assign LUT_3[22987] = 32'b00000000000000010111010101100001;
assign LUT_3[22988] = 32'b00000000000000001011110000010110;
assign LUT_3[22989] = 32'b00000000000000010010011011110011;
assign LUT_3[22990] = 32'b00000000000000001101110111111010;
assign LUT_3[22991] = 32'b00000000000000010100100011010111;
assign LUT_3[22992] = 32'b00000000000000001100011100011101;
assign LUT_3[22993] = 32'b00000000000000010011000111111010;
assign LUT_3[22994] = 32'b00000000000000001110100100000001;
assign LUT_3[22995] = 32'b00000000000000010101001111011110;
assign LUT_3[22996] = 32'b00000000000000001001101010010011;
assign LUT_3[22997] = 32'b00000000000000010000010101110000;
assign LUT_3[22998] = 32'b00000000000000001011110001110111;
assign LUT_3[22999] = 32'b00000000000000010010011101010100;
assign LUT_3[23000] = 32'b00000000000000010001110101100011;
assign LUT_3[23001] = 32'b00000000000000011000100001000000;
assign LUT_3[23002] = 32'b00000000000000010011111101000111;
assign LUT_3[23003] = 32'b00000000000000011010101000100100;
assign LUT_3[23004] = 32'b00000000000000001111000011011001;
assign LUT_3[23005] = 32'b00000000000000010101101110110110;
assign LUT_3[23006] = 32'b00000000000000010001001010111101;
assign LUT_3[23007] = 32'b00000000000000010111110110011010;
assign LUT_3[23008] = 32'b00000000000000001010010111111010;
assign LUT_3[23009] = 32'b00000000000000010001000011010111;
assign LUT_3[23010] = 32'b00000000000000001100011111011110;
assign LUT_3[23011] = 32'b00000000000000010011001010111011;
assign LUT_3[23012] = 32'b00000000000000000111100101110000;
assign LUT_3[23013] = 32'b00000000000000001110010001001101;
assign LUT_3[23014] = 32'b00000000000000001001101101010100;
assign LUT_3[23015] = 32'b00000000000000010000011000110001;
assign LUT_3[23016] = 32'b00000000000000001111110001000000;
assign LUT_3[23017] = 32'b00000000000000010110011100011101;
assign LUT_3[23018] = 32'b00000000000000010001111000100100;
assign LUT_3[23019] = 32'b00000000000000011000100100000001;
assign LUT_3[23020] = 32'b00000000000000001100111110110110;
assign LUT_3[23021] = 32'b00000000000000010011101010010011;
assign LUT_3[23022] = 32'b00000000000000001111000110011010;
assign LUT_3[23023] = 32'b00000000000000010101110001110111;
assign LUT_3[23024] = 32'b00000000000000001101101010111101;
assign LUT_3[23025] = 32'b00000000000000010100010110011010;
assign LUT_3[23026] = 32'b00000000000000001111110010100001;
assign LUT_3[23027] = 32'b00000000000000010110011101111110;
assign LUT_3[23028] = 32'b00000000000000001010111000110011;
assign LUT_3[23029] = 32'b00000000000000010001100100010000;
assign LUT_3[23030] = 32'b00000000000000001101000000010111;
assign LUT_3[23031] = 32'b00000000000000010011101011110100;
assign LUT_3[23032] = 32'b00000000000000010011000100000011;
assign LUT_3[23033] = 32'b00000000000000011001101111100000;
assign LUT_3[23034] = 32'b00000000000000010101001011100111;
assign LUT_3[23035] = 32'b00000000000000011011110111000100;
assign LUT_3[23036] = 32'b00000000000000010000010001111001;
assign LUT_3[23037] = 32'b00000000000000010110111101010110;
assign LUT_3[23038] = 32'b00000000000000010010011001011101;
assign LUT_3[23039] = 32'b00000000000000011001000100111010;
assign LUT_3[23040] = 32'b00000000000000001110001011011100;
assign LUT_3[23041] = 32'b00000000000000010100110110111001;
assign LUT_3[23042] = 32'b00000000000000010000010011000000;
assign LUT_3[23043] = 32'b00000000000000010110111110011101;
assign LUT_3[23044] = 32'b00000000000000001011011001010010;
assign LUT_3[23045] = 32'b00000000000000010010000100101111;
assign LUT_3[23046] = 32'b00000000000000001101100000110110;
assign LUT_3[23047] = 32'b00000000000000010100001100010011;
assign LUT_3[23048] = 32'b00000000000000010011100100100010;
assign LUT_3[23049] = 32'b00000000000000011010001111111111;
assign LUT_3[23050] = 32'b00000000000000010101101100000110;
assign LUT_3[23051] = 32'b00000000000000011100010111100011;
assign LUT_3[23052] = 32'b00000000000000010000110010011000;
assign LUT_3[23053] = 32'b00000000000000010111011101110101;
assign LUT_3[23054] = 32'b00000000000000010010111001111100;
assign LUT_3[23055] = 32'b00000000000000011001100101011001;
assign LUT_3[23056] = 32'b00000000000000010001011110011111;
assign LUT_3[23057] = 32'b00000000000000011000001001111100;
assign LUT_3[23058] = 32'b00000000000000010011100110000011;
assign LUT_3[23059] = 32'b00000000000000011010010001100000;
assign LUT_3[23060] = 32'b00000000000000001110101100010101;
assign LUT_3[23061] = 32'b00000000000000010101010111110010;
assign LUT_3[23062] = 32'b00000000000000010000110011111001;
assign LUT_3[23063] = 32'b00000000000000010111011111010110;
assign LUT_3[23064] = 32'b00000000000000010110110111100101;
assign LUT_3[23065] = 32'b00000000000000011101100011000010;
assign LUT_3[23066] = 32'b00000000000000011000111111001001;
assign LUT_3[23067] = 32'b00000000000000011111101010100110;
assign LUT_3[23068] = 32'b00000000000000010100000101011011;
assign LUT_3[23069] = 32'b00000000000000011010110000111000;
assign LUT_3[23070] = 32'b00000000000000010110001100111111;
assign LUT_3[23071] = 32'b00000000000000011100111000011100;
assign LUT_3[23072] = 32'b00000000000000001111011001111100;
assign LUT_3[23073] = 32'b00000000000000010110000101011001;
assign LUT_3[23074] = 32'b00000000000000010001100001100000;
assign LUT_3[23075] = 32'b00000000000000011000001100111101;
assign LUT_3[23076] = 32'b00000000000000001100100111110010;
assign LUT_3[23077] = 32'b00000000000000010011010011001111;
assign LUT_3[23078] = 32'b00000000000000001110101111010110;
assign LUT_3[23079] = 32'b00000000000000010101011010110011;
assign LUT_3[23080] = 32'b00000000000000010100110011000010;
assign LUT_3[23081] = 32'b00000000000000011011011110011111;
assign LUT_3[23082] = 32'b00000000000000010110111010100110;
assign LUT_3[23083] = 32'b00000000000000011101100110000011;
assign LUT_3[23084] = 32'b00000000000000010010000000111000;
assign LUT_3[23085] = 32'b00000000000000011000101100010101;
assign LUT_3[23086] = 32'b00000000000000010100001000011100;
assign LUT_3[23087] = 32'b00000000000000011010110011111001;
assign LUT_3[23088] = 32'b00000000000000010010101100111111;
assign LUT_3[23089] = 32'b00000000000000011001011000011100;
assign LUT_3[23090] = 32'b00000000000000010100110100100011;
assign LUT_3[23091] = 32'b00000000000000011011100000000000;
assign LUT_3[23092] = 32'b00000000000000001111111010110101;
assign LUT_3[23093] = 32'b00000000000000010110100110010010;
assign LUT_3[23094] = 32'b00000000000000010010000010011001;
assign LUT_3[23095] = 32'b00000000000000011000101101110110;
assign LUT_3[23096] = 32'b00000000000000011000000110000101;
assign LUT_3[23097] = 32'b00000000000000011110110001100010;
assign LUT_3[23098] = 32'b00000000000000011010001101101001;
assign LUT_3[23099] = 32'b00000000000000100000111001000110;
assign LUT_3[23100] = 32'b00000000000000010101010011111011;
assign LUT_3[23101] = 32'b00000000000000011011111111011000;
assign LUT_3[23102] = 32'b00000000000000010111011011011111;
assign LUT_3[23103] = 32'b00000000000000011110000110111100;
assign LUT_3[23104] = 32'b00000000000000001110000100000111;
assign LUT_3[23105] = 32'b00000000000000010100101111100100;
assign LUT_3[23106] = 32'b00000000000000010000001011101011;
assign LUT_3[23107] = 32'b00000000000000010110110111001000;
assign LUT_3[23108] = 32'b00000000000000001011010001111101;
assign LUT_3[23109] = 32'b00000000000000010001111101011010;
assign LUT_3[23110] = 32'b00000000000000001101011001100001;
assign LUT_3[23111] = 32'b00000000000000010100000100111110;
assign LUT_3[23112] = 32'b00000000000000010011011101001101;
assign LUT_3[23113] = 32'b00000000000000011010001000101010;
assign LUT_3[23114] = 32'b00000000000000010101100100110001;
assign LUT_3[23115] = 32'b00000000000000011100010000001110;
assign LUT_3[23116] = 32'b00000000000000010000101011000011;
assign LUT_3[23117] = 32'b00000000000000010111010110100000;
assign LUT_3[23118] = 32'b00000000000000010010110010100111;
assign LUT_3[23119] = 32'b00000000000000011001011110000100;
assign LUT_3[23120] = 32'b00000000000000010001010111001010;
assign LUT_3[23121] = 32'b00000000000000011000000010100111;
assign LUT_3[23122] = 32'b00000000000000010011011110101110;
assign LUT_3[23123] = 32'b00000000000000011010001010001011;
assign LUT_3[23124] = 32'b00000000000000001110100101000000;
assign LUT_3[23125] = 32'b00000000000000010101010000011101;
assign LUT_3[23126] = 32'b00000000000000010000101100100100;
assign LUT_3[23127] = 32'b00000000000000010111011000000001;
assign LUT_3[23128] = 32'b00000000000000010110110000010000;
assign LUT_3[23129] = 32'b00000000000000011101011011101101;
assign LUT_3[23130] = 32'b00000000000000011000110111110100;
assign LUT_3[23131] = 32'b00000000000000011111100011010001;
assign LUT_3[23132] = 32'b00000000000000010011111110000110;
assign LUT_3[23133] = 32'b00000000000000011010101001100011;
assign LUT_3[23134] = 32'b00000000000000010110000101101010;
assign LUT_3[23135] = 32'b00000000000000011100110001000111;
assign LUT_3[23136] = 32'b00000000000000001111010010100111;
assign LUT_3[23137] = 32'b00000000000000010101111110000100;
assign LUT_3[23138] = 32'b00000000000000010001011010001011;
assign LUT_3[23139] = 32'b00000000000000011000000101101000;
assign LUT_3[23140] = 32'b00000000000000001100100000011101;
assign LUT_3[23141] = 32'b00000000000000010011001011111010;
assign LUT_3[23142] = 32'b00000000000000001110101000000001;
assign LUT_3[23143] = 32'b00000000000000010101010011011110;
assign LUT_3[23144] = 32'b00000000000000010100101011101101;
assign LUT_3[23145] = 32'b00000000000000011011010111001010;
assign LUT_3[23146] = 32'b00000000000000010110110011010001;
assign LUT_3[23147] = 32'b00000000000000011101011110101110;
assign LUT_3[23148] = 32'b00000000000000010001111001100011;
assign LUT_3[23149] = 32'b00000000000000011000100101000000;
assign LUT_3[23150] = 32'b00000000000000010100000001000111;
assign LUT_3[23151] = 32'b00000000000000011010101100100100;
assign LUT_3[23152] = 32'b00000000000000010010100101101010;
assign LUT_3[23153] = 32'b00000000000000011001010001000111;
assign LUT_3[23154] = 32'b00000000000000010100101101001110;
assign LUT_3[23155] = 32'b00000000000000011011011000101011;
assign LUT_3[23156] = 32'b00000000000000001111110011100000;
assign LUT_3[23157] = 32'b00000000000000010110011110111101;
assign LUT_3[23158] = 32'b00000000000000010001111011000100;
assign LUT_3[23159] = 32'b00000000000000011000100110100001;
assign LUT_3[23160] = 32'b00000000000000010111111110110000;
assign LUT_3[23161] = 32'b00000000000000011110101010001101;
assign LUT_3[23162] = 32'b00000000000000011010000110010100;
assign LUT_3[23163] = 32'b00000000000000100000110001110001;
assign LUT_3[23164] = 32'b00000000000000010101001100100110;
assign LUT_3[23165] = 32'b00000000000000011011111000000011;
assign LUT_3[23166] = 32'b00000000000000010111010100001010;
assign LUT_3[23167] = 32'b00000000000000011101111111100111;
assign LUT_3[23168] = 32'b00000000000000010000010110011010;
assign LUT_3[23169] = 32'b00000000000000010111000001110111;
assign LUT_3[23170] = 32'b00000000000000010010011101111110;
assign LUT_3[23171] = 32'b00000000000000011001001001011011;
assign LUT_3[23172] = 32'b00000000000000001101100100010000;
assign LUT_3[23173] = 32'b00000000000000010100001111101101;
assign LUT_3[23174] = 32'b00000000000000001111101011110100;
assign LUT_3[23175] = 32'b00000000000000010110010111010001;
assign LUT_3[23176] = 32'b00000000000000010101101111100000;
assign LUT_3[23177] = 32'b00000000000000011100011010111101;
assign LUT_3[23178] = 32'b00000000000000010111110111000100;
assign LUT_3[23179] = 32'b00000000000000011110100010100001;
assign LUT_3[23180] = 32'b00000000000000010010111101010110;
assign LUT_3[23181] = 32'b00000000000000011001101000110011;
assign LUT_3[23182] = 32'b00000000000000010101000100111010;
assign LUT_3[23183] = 32'b00000000000000011011110000010111;
assign LUT_3[23184] = 32'b00000000000000010011101001011101;
assign LUT_3[23185] = 32'b00000000000000011010010100111010;
assign LUT_3[23186] = 32'b00000000000000010101110001000001;
assign LUT_3[23187] = 32'b00000000000000011100011100011110;
assign LUT_3[23188] = 32'b00000000000000010000110111010011;
assign LUT_3[23189] = 32'b00000000000000010111100010110000;
assign LUT_3[23190] = 32'b00000000000000010010111110110111;
assign LUT_3[23191] = 32'b00000000000000011001101010010100;
assign LUT_3[23192] = 32'b00000000000000011001000010100011;
assign LUT_3[23193] = 32'b00000000000000011111101110000000;
assign LUT_3[23194] = 32'b00000000000000011011001010000111;
assign LUT_3[23195] = 32'b00000000000000100001110101100100;
assign LUT_3[23196] = 32'b00000000000000010110010000011001;
assign LUT_3[23197] = 32'b00000000000000011100111011110110;
assign LUT_3[23198] = 32'b00000000000000011000010111111101;
assign LUT_3[23199] = 32'b00000000000000011111000011011010;
assign LUT_3[23200] = 32'b00000000000000010001100100111010;
assign LUT_3[23201] = 32'b00000000000000011000010000010111;
assign LUT_3[23202] = 32'b00000000000000010011101100011110;
assign LUT_3[23203] = 32'b00000000000000011010010111111011;
assign LUT_3[23204] = 32'b00000000000000001110110010110000;
assign LUT_3[23205] = 32'b00000000000000010101011110001101;
assign LUT_3[23206] = 32'b00000000000000010000111010010100;
assign LUT_3[23207] = 32'b00000000000000010111100101110001;
assign LUT_3[23208] = 32'b00000000000000010110111110000000;
assign LUT_3[23209] = 32'b00000000000000011101101001011101;
assign LUT_3[23210] = 32'b00000000000000011001000101100100;
assign LUT_3[23211] = 32'b00000000000000011111110001000001;
assign LUT_3[23212] = 32'b00000000000000010100001011110110;
assign LUT_3[23213] = 32'b00000000000000011010110111010011;
assign LUT_3[23214] = 32'b00000000000000010110010011011010;
assign LUT_3[23215] = 32'b00000000000000011100111110110111;
assign LUT_3[23216] = 32'b00000000000000010100110111111101;
assign LUT_3[23217] = 32'b00000000000000011011100011011010;
assign LUT_3[23218] = 32'b00000000000000010110111111100001;
assign LUT_3[23219] = 32'b00000000000000011101101010111110;
assign LUT_3[23220] = 32'b00000000000000010010000101110011;
assign LUT_3[23221] = 32'b00000000000000011000110001010000;
assign LUT_3[23222] = 32'b00000000000000010100001101010111;
assign LUT_3[23223] = 32'b00000000000000011010111000110100;
assign LUT_3[23224] = 32'b00000000000000011010010001000011;
assign LUT_3[23225] = 32'b00000000000000100000111100100000;
assign LUT_3[23226] = 32'b00000000000000011100011000100111;
assign LUT_3[23227] = 32'b00000000000000100011000100000100;
assign LUT_3[23228] = 32'b00000000000000010111011110111001;
assign LUT_3[23229] = 32'b00000000000000011110001010010110;
assign LUT_3[23230] = 32'b00000000000000011001100110011101;
assign LUT_3[23231] = 32'b00000000000000100000010001111010;
assign LUT_3[23232] = 32'b00000000000000010000001111000101;
assign LUT_3[23233] = 32'b00000000000000010110111010100010;
assign LUT_3[23234] = 32'b00000000000000010010010110101001;
assign LUT_3[23235] = 32'b00000000000000011001000010000110;
assign LUT_3[23236] = 32'b00000000000000001101011100111011;
assign LUT_3[23237] = 32'b00000000000000010100001000011000;
assign LUT_3[23238] = 32'b00000000000000001111100100011111;
assign LUT_3[23239] = 32'b00000000000000010110001111111100;
assign LUT_3[23240] = 32'b00000000000000010101101000001011;
assign LUT_3[23241] = 32'b00000000000000011100010011101000;
assign LUT_3[23242] = 32'b00000000000000010111101111101111;
assign LUT_3[23243] = 32'b00000000000000011110011011001100;
assign LUT_3[23244] = 32'b00000000000000010010110110000001;
assign LUT_3[23245] = 32'b00000000000000011001100001011110;
assign LUT_3[23246] = 32'b00000000000000010100111101100101;
assign LUT_3[23247] = 32'b00000000000000011011101001000010;
assign LUT_3[23248] = 32'b00000000000000010011100010001000;
assign LUT_3[23249] = 32'b00000000000000011010001101100101;
assign LUT_3[23250] = 32'b00000000000000010101101001101100;
assign LUT_3[23251] = 32'b00000000000000011100010101001001;
assign LUT_3[23252] = 32'b00000000000000010000101111111110;
assign LUT_3[23253] = 32'b00000000000000010111011011011011;
assign LUT_3[23254] = 32'b00000000000000010010110111100010;
assign LUT_3[23255] = 32'b00000000000000011001100010111111;
assign LUT_3[23256] = 32'b00000000000000011000111011001110;
assign LUT_3[23257] = 32'b00000000000000011111100110101011;
assign LUT_3[23258] = 32'b00000000000000011011000010110010;
assign LUT_3[23259] = 32'b00000000000000100001101110001111;
assign LUT_3[23260] = 32'b00000000000000010110001001000100;
assign LUT_3[23261] = 32'b00000000000000011100110100100001;
assign LUT_3[23262] = 32'b00000000000000011000010000101000;
assign LUT_3[23263] = 32'b00000000000000011110111100000101;
assign LUT_3[23264] = 32'b00000000000000010001011101100101;
assign LUT_3[23265] = 32'b00000000000000011000001001000010;
assign LUT_3[23266] = 32'b00000000000000010011100101001001;
assign LUT_3[23267] = 32'b00000000000000011010010000100110;
assign LUT_3[23268] = 32'b00000000000000001110101011011011;
assign LUT_3[23269] = 32'b00000000000000010101010110111000;
assign LUT_3[23270] = 32'b00000000000000010000110010111111;
assign LUT_3[23271] = 32'b00000000000000010111011110011100;
assign LUT_3[23272] = 32'b00000000000000010110110110101011;
assign LUT_3[23273] = 32'b00000000000000011101100010001000;
assign LUT_3[23274] = 32'b00000000000000011000111110001111;
assign LUT_3[23275] = 32'b00000000000000011111101001101100;
assign LUT_3[23276] = 32'b00000000000000010100000100100001;
assign LUT_3[23277] = 32'b00000000000000011010101111111110;
assign LUT_3[23278] = 32'b00000000000000010110001100000101;
assign LUT_3[23279] = 32'b00000000000000011100110111100010;
assign LUT_3[23280] = 32'b00000000000000010100110000101000;
assign LUT_3[23281] = 32'b00000000000000011011011100000101;
assign LUT_3[23282] = 32'b00000000000000010110111000001100;
assign LUT_3[23283] = 32'b00000000000000011101100011101001;
assign LUT_3[23284] = 32'b00000000000000010001111110011110;
assign LUT_3[23285] = 32'b00000000000000011000101001111011;
assign LUT_3[23286] = 32'b00000000000000010100000110000010;
assign LUT_3[23287] = 32'b00000000000000011010110001011111;
assign LUT_3[23288] = 32'b00000000000000011010001001101110;
assign LUT_3[23289] = 32'b00000000000000100000110101001011;
assign LUT_3[23290] = 32'b00000000000000011100010001010010;
assign LUT_3[23291] = 32'b00000000000000100010111100101111;
assign LUT_3[23292] = 32'b00000000000000010111010111100100;
assign LUT_3[23293] = 32'b00000000000000011110000011000001;
assign LUT_3[23294] = 32'b00000000000000011001011111001000;
assign LUT_3[23295] = 32'b00000000000000100000001010100101;
assign LUT_3[23296] = 32'b00000000000000001010011010111101;
assign LUT_3[23297] = 32'b00000000000000010001000110011010;
assign LUT_3[23298] = 32'b00000000000000001100100010100001;
assign LUT_3[23299] = 32'b00000000000000010011001101111110;
assign LUT_3[23300] = 32'b00000000000000000111101000110011;
assign LUT_3[23301] = 32'b00000000000000001110010100010000;
assign LUT_3[23302] = 32'b00000000000000001001110000010111;
assign LUT_3[23303] = 32'b00000000000000010000011011110100;
assign LUT_3[23304] = 32'b00000000000000001111110100000011;
assign LUT_3[23305] = 32'b00000000000000010110011111100000;
assign LUT_3[23306] = 32'b00000000000000010001111011100111;
assign LUT_3[23307] = 32'b00000000000000011000100111000100;
assign LUT_3[23308] = 32'b00000000000000001101000001111001;
assign LUT_3[23309] = 32'b00000000000000010011101101010110;
assign LUT_3[23310] = 32'b00000000000000001111001001011101;
assign LUT_3[23311] = 32'b00000000000000010101110100111010;
assign LUT_3[23312] = 32'b00000000000000001101101110000000;
assign LUT_3[23313] = 32'b00000000000000010100011001011101;
assign LUT_3[23314] = 32'b00000000000000001111110101100100;
assign LUT_3[23315] = 32'b00000000000000010110100001000001;
assign LUT_3[23316] = 32'b00000000000000001010111011110110;
assign LUT_3[23317] = 32'b00000000000000010001100111010011;
assign LUT_3[23318] = 32'b00000000000000001101000011011010;
assign LUT_3[23319] = 32'b00000000000000010011101110110111;
assign LUT_3[23320] = 32'b00000000000000010011000111000110;
assign LUT_3[23321] = 32'b00000000000000011001110010100011;
assign LUT_3[23322] = 32'b00000000000000010101001110101010;
assign LUT_3[23323] = 32'b00000000000000011011111010000111;
assign LUT_3[23324] = 32'b00000000000000010000010100111100;
assign LUT_3[23325] = 32'b00000000000000010111000000011001;
assign LUT_3[23326] = 32'b00000000000000010010011100100000;
assign LUT_3[23327] = 32'b00000000000000011001000111111101;
assign LUT_3[23328] = 32'b00000000000000001011101001011101;
assign LUT_3[23329] = 32'b00000000000000010010010100111010;
assign LUT_3[23330] = 32'b00000000000000001101110001000001;
assign LUT_3[23331] = 32'b00000000000000010100011100011110;
assign LUT_3[23332] = 32'b00000000000000001000110111010011;
assign LUT_3[23333] = 32'b00000000000000001111100010110000;
assign LUT_3[23334] = 32'b00000000000000001010111110110111;
assign LUT_3[23335] = 32'b00000000000000010001101010010100;
assign LUT_3[23336] = 32'b00000000000000010001000010100011;
assign LUT_3[23337] = 32'b00000000000000010111101110000000;
assign LUT_3[23338] = 32'b00000000000000010011001010000111;
assign LUT_3[23339] = 32'b00000000000000011001110101100100;
assign LUT_3[23340] = 32'b00000000000000001110010000011001;
assign LUT_3[23341] = 32'b00000000000000010100111011110110;
assign LUT_3[23342] = 32'b00000000000000010000010111111101;
assign LUT_3[23343] = 32'b00000000000000010111000011011010;
assign LUT_3[23344] = 32'b00000000000000001110111100100000;
assign LUT_3[23345] = 32'b00000000000000010101100111111101;
assign LUT_3[23346] = 32'b00000000000000010001000100000100;
assign LUT_3[23347] = 32'b00000000000000010111101111100001;
assign LUT_3[23348] = 32'b00000000000000001100001010010110;
assign LUT_3[23349] = 32'b00000000000000010010110101110011;
assign LUT_3[23350] = 32'b00000000000000001110010001111010;
assign LUT_3[23351] = 32'b00000000000000010100111101010111;
assign LUT_3[23352] = 32'b00000000000000010100010101100110;
assign LUT_3[23353] = 32'b00000000000000011011000001000011;
assign LUT_3[23354] = 32'b00000000000000010110011101001010;
assign LUT_3[23355] = 32'b00000000000000011101001000100111;
assign LUT_3[23356] = 32'b00000000000000010001100011011100;
assign LUT_3[23357] = 32'b00000000000000011000001110111001;
assign LUT_3[23358] = 32'b00000000000000010011101011000000;
assign LUT_3[23359] = 32'b00000000000000011010010110011101;
assign LUT_3[23360] = 32'b00000000000000001010010011101000;
assign LUT_3[23361] = 32'b00000000000000010000111111000101;
assign LUT_3[23362] = 32'b00000000000000001100011011001100;
assign LUT_3[23363] = 32'b00000000000000010011000110101001;
assign LUT_3[23364] = 32'b00000000000000000111100001011110;
assign LUT_3[23365] = 32'b00000000000000001110001100111011;
assign LUT_3[23366] = 32'b00000000000000001001101001000010;
assign LUT_3[23367] = 32'b00000000000000010000010100011111;
assign LUT_3[23368] = 32'b00000000000000001111101100101110;
assign LUT_3[23369] = 32'b00000000000000010110011000001011;
assign LUT_3[23370] = 32'b00000000000000010001110100010010;
assign LUT_3[23371] = 32'b00000000000000011000011111101111;
assign LUT_3[23372] = 32'b00000000000000001100111010100100;
assign LUT_3[23373] = 32'b00000000000000010011100110000001;
assign LUT_3[23374] = 32'b00000000000000001111000010001000;
assign LUT_3[23375] = 32'b00000000000000010101101101100101;
assign LUT_3[23376] = 32'b00000000000000001101100110101011;
assign LUT_3[23377] = 32'b00000000000000010100010010001000;
assign LUT_3[23378] = 32'b00000000000000001111101110001111;
assign LUT_3[23379] = 32'b00000000000000010110011001101100;
assign LUT_3[23380] = 32'b00000000000000001010110100100001;
assign LUT_3[23381] = 32'b00000000000000010001011111111110;
assign LUT_3[23382] = 32'b00000000000000001100111100000101;
assign LUT_3[23383] = 32'b00000000000000010011100111100010;
assign LUT_3[23384] = 32'b00000000000000010010111111110001;
assign LUT_3[23385] = 32'b00000000000000011001101011001110;
assign LUT_3[23386] = 32'b00000000000000010101000111010101;
assign LUT_3[23387] = 32'b00000000000000011011110010110010;
assign LUT_3[23388] = 32'b00000000000000010000001101100111;
assign LUT_3[23389] = 32'b00000000000000010110111001000100;
assign LUT_3[23390] = 32'b00000000000000010010010101001011;
assign LUT_3[23391] = 32'b00000000000000011001000000101000;
assign LUT_3[23392] = 32'b00000000000000001011100010001000;
assign LUT_3[23393] = 32'b00000000000000010010001101100101;
assign LUT_3[23394] = 32'b00000000000000001101101001101100;
assign LUT_3[23395] = 32'b00000000000000010100010101001001;
assign LUT_3[23396] = 32'b00000000000000001000101111111110;
assign LUT_3[23397] = 32'b00000000000000001111011011011011;
assign LUT_3[23398] = 32'b00000000000000001010110111100010;
assign LUT_3[23399] = 32'b00000000000000010001100010111111;
assign LUT_3[23400] = 32'b00000000000000010000111011001110;
assign LUT_3[23401] = 32'b00000000000000010111100110101011;
assign LUT_3[23402] = 32'b00000000000000010011000010110010;
assign LUT_3[23403] = 32'b00000000000000011001101110001111;
assign LUT_3[23404] = 32'b00000000000000001110001001000100;
assign LUT_3[23405] = 32'b00000000000000010100110100100001;
assign LUT_3[23406] = 32'b00000000000000010000010000101000;
assign LUT_3[23407] = 32'b00000000000000010110111100000101;
assign LUT_3[23408] = 32'b00000000000000001110110101001011;
assign LUT_3[23409] = 32'b00000000000000010101100000101000;
assign LUT_3[23410] = 32'b00000000000000010000111100101111;
assign LUT_3[23411] = 32'b00000000000000010111101000001100;
assign LUT_3[23412] = 32'b00000000000000001100000011000001;
assign LUT_3[23413] = 32'b00000000000000010010101110011110;
assign LUT_3[23414] = 32'b00000000000000001110001010100101;
assign LUT_3[23415] = 32'b00000000000000010100110110000010;
assign LUT_3[23416] = 32'b00000000000000010100001110010001;
assign LUT_3[23417] = 32'b00000000000000011010111001101110;
assign LUT_3[23418] = 32'b00000000000000010110010101110101;
assign LUT_3[23419] = 32'b00000000000000011101000001010010;
assign LUT_3[23420] = 32'b00000000000000010001011100000111;
assign LUT_3[23421] = 32'b00000000000000011000000111100100;
assign LUT_3[23422] = 32'b00000000000000010011100011101011;
assign LUT_3[23423] = 32'b00000000000000011010001111001000;
assign LUT_3[23424] = 32'b00000000000000001100100101111011;
assign LUT_3[23425] = 32'b00000000000000010011010001011000;
assign LUT_3[23426] = 32'b00000000000000001110101101011111;
assign LUT_3[23427] = 32'b00000000000000010101011000111100;
assign LUT_3[23428] = 32'b00000000000000001001110011110001;
assign LUT_3[23429] = 32'b00000000000000010000011111001110;
assign LUT_3[23430] = 32'b00000000000000001011111011010101;
assign LUT_3[23431] = 32'b00000000000000010010100110110010;
assign LUT_3[23432] = 32'b00000000000000010001111111000001;
assign LUT_3[23433] = 32'b00000000000000011000101010011110;
assign LUT_3[23434] = 32'b00000000000000010100000110100101;
assign LUT_3[23435] = 32'b00000000000000011010110010000010;
assign LUT_3[23436] = 32'b00000000000000001111001100110111;
assign LUT_3[23437] = 32'b00000000000000010101111000010100;
assign LUT_3[23438] = 32'b00000000000000010001010100011011;
assign LUT_3[23439] = 32'b00000000000000010111111111111000;
assign LUT_3[23440] = 32'b00000000000000001111111000111110;
assign LUT_3[23441] = 32'b00000000000000010110100100011011;
assign LUT_3[23442] = 32'b00000000000000010010000000100010;
assign LUT_3[23443] = 32'b00000000000000011000101011111111;
assign LUT_3[23444] = 32'b00000000000000001101000110110100;
assign LUT_3[23445] = 32'b00000000000000010011110010010001;
assign LUT_3[23446] = 32'b00000000000000001111001110011000;
assign LUT_3[23447] = 32'b00000000000000010101111001110101;
assign LUT_3[23448] = 32'b00000000000000010101010010000100;
assign LUT_3[23449] = 32'b00000000000000011011111101100001;
assign LUT_3[23450] = 32'b00000000000000010111011001101000;
assign LUT_3[23451] = 32'b00000000000000011110000101000101;
assign LUT_3[23452] = 32'b00000000000000010010011111111010;
assign LUT_3[23453] = 32'b00000000000000011001001011010111;
assign LUT_3[23454] = 32'b00000000000000010100100111011110;
assign LUT_3[23455] = 32'b00000000000000011011010010111011;
assign LUT_3[23456] = 32'b00000000000000001101110100011011;
assign LUT_3[23457] = 32'b00000000000000010100011111111000;
assign LUT_3[23458] = 32'b00000000000000001111111011111111;
assign LUT_3[23459] = 32'b00000000000000010110100111011100;
assign LUT_3[23460] = 32'b00000000000000001011000010010001;
assign LUT_3[23461] = 32'b00000000000000010001101101101110;
assign LUT_3[23462] = 32'b00000000000000001101001001110101;
assign LUT_3[23463] = 32'b00000000000000010011110101010010;
assign LUT_3[23464] = 32'b00000000000000010011001101100001;
assign LUT_3[23465] = 32'b00000000000000011001111000111110;
assign LUT_3[23466] = 32'b00000000000000010101010101000101;
assign LUT_3[23467] = 32'b00000000000000011100000000100010;
assign LUT_3[23468] = 32'b00000000000000010000011011010111;
assign LUT_3[23469] = 32'b00000000000000010111000110110100;
assign LUT_3[23470] = 32'b00000000000000010010100010111011;
assign LUT_3[23471] = 32'b00000000000000011001001110011000;
assign LUT_3[23472] = 32'b00000000000000010001000111011110;
assign LUT_3[23473] = 32'b00000000000000010111110010111011;
assign LUT_3[23474] = 32'b00000000000000010011001111000010;
assign LUT_3[23475] = 32'b00000000000000011001111010011111;
assign LUT_3[23476] = 32'b00000000000000001110010101010100;
assign LUT_3[23477] = 32'b00000000000000010101000000110001;
assign LUT_3[23478] = 32'b00000000000000010000011100111000;
assign LUT_3[23479] = 32'b00000000000000010111001000010101;
assign LUT_3[23480] = 32'b00000000000000010110100000100100;
assign LUT_3[23481] = 32'b00000000000000011101001100000001;
assign LUT_3[23482] = 32'b00000000000000011000101000001000;
assign LUT_3[23483] = 32'b00000000000000011111010011100101;
assign LUT_3[23484] = 32'b00000000000000010011101110011010;
assign LUT_3[23485] = 32'b00000000000000011010011001110111;
assign LUT_3[23486] = 32'b00000000000000010101110101111110;
assign LUT_3[23487] = 32'b00000000000000011100100001011011;
assign LUT_3[23488] = 32'b00000000000000001100011110100110;
assign LUT_3[23489] = 32'b00000000000000010011001010000011;
assign LUT_3[23490] = 32'b00000000000000001110100110001010;
assign LUT_3[23491] = 32'b00000000000000010101010001100111;
assign LUT_3[23492] = 32'b00000000000000001001101100011100;
assign LUT_3[23493] = 32'b00000000000000010000010111111001;
assign LUT_3[23494] = 32'b00000000000000001011110100000000;
assign LUT_3[23495] = 32'b00000000000000010010011111011101;
assign LUT_3[23496] = 32'b00000000000000010001110111101100;
assign LUT_3[23497] = 32'b00000000000000011000100011001001;
assign LUT_3[23498] = 32'b00000000000000010011111111010000;
assign LUT_3[23499] = 32'b00000000000000011010101010101101;
assign LUT_3[23500] = 32'b00000000000000001111000101100010;
assign LUT_3[23501] = 32'b00000000000000010101110000111111;
assign LUT_3[23502] = 32'b00000000000000010001001101000110;
assign LUT_3[23503] = 32'b00000000000000010111111000100011;
assign LUT_3[23504] = 32'b00000000000000001111110001101001;
assign LUT_3[23505] = 32'b00000000000000010110011101000110;
assign LUT_3[23506] = 32'b00000000000000010001111001001101;
assign LUT_3[23507] = 32'b00000000000000011000100100101010;
assign LUT_3[23508] = 32'b00000000000000001100111111011111;
assign LUT_3[23509] = 32'b00000000000000010011101010111100;
assign LUT_3[23510] = 32'b00000000000000001111000111000011;
assign LUT_3[23511] = 32'b00000000000000010101110010100000;
assign LUT_3[23512] = 32'b00000000000000010101001010101111;
assign LUT_3[23513] = 32'b00000000000000011011110110001100;
assign LUT_3[23514] = 32'b00000000000000010111010010010011;
assign LUT_3[23515] = 32'b00000000000000011101111101110000;
assign LUT_3[23516] = 32'b00000000000000010010011000100101;
assign LUT_3[23517] = 32'b00000000000000011001000100000010;
assign LUT_3[23518] = 32'b00000000000000010100100000001001;
assign LUT_3[23519] = 32'b00000000000000011011001011100110;
assign LUT_3[23520] = 32'b00000000000000001101101101000110;
assign LUT_3[23521] = 32'b00000000000000010100011000100011;
assign LUT_3[23522] = 32'b00000000000000001111110100101010;
assign LUT_3[23523] = 32'b00000000000000010110100000000111;
assign LUT_3[23524] = 32'b00000000000000001010111010111100;
assign LUT_3[23525] = 32'b00000000000000010001100110011001;
assign LUT_3[23526] = 32'b00000000000000001101000010100000;
assign LUT_3[23527] = 32'b00000000000000010011101101111101;
assign LUT_3[23528] = 32'b00000000000000010011000110001100;
assign LUT_3[23529] = 32'b00000000000000011001110001101001;
assign LUT_3[23530] = 32'b00000000000000010101001101110000;
assign LUT_3[23531] = 32'b00000000000000011011111001001101;
assign LUT_3[23532] = 32'b00000000000000010000010100000010;
assign LUT_3[23533] = 32'b00000000000000010110111111011111;
assign LUT_3[23534] = 32'b00000000000000010010011011100110;
assign LUT_3[23535] = 32'b00000000000000011001000111000011;
assign LUT_3[23536] = 32'b00000000000000010001000000001001;
assign LUT_3[23537] = 32'b00000000000000010111101011100110;
assign LUT_3[23538] = 32'b00000000000000010011000111101101;
assign LUT_3[23539] = 32'b00000000000000011001110011001010;
assign LUT_3[23540] = 32'b00000000000000001110001101111111;
assign LUT_3[23541] = 32'b00000000000000010100111001011100;
assign LUT_3[23542] = 32'b00000000000000010000010101100011;
assign LUT_3[23543] = 32'b00000000000000010111000001000000;
assign LUT_3[23544] = 32'b00000000000000010110011001001111;
assign LUT_3[23545] = 32'b00000000000000011101000100101100;
assign LUT_3[23546] = 32'b00000000000000011000100000110011;
assign LUT_3[23547] = 32'b00000000000000011111001100010000;
assign LUT_3[23548] = 32'b00000000000000010011100111000101;
assign LUT_3[23549] = 32'b00000000000000011010010010100010;
assign LUT_3[23550] = 32'b00000000000000010101101110101001;
assign LUT_3[23551] = 32'b00000000000000011100011010000110;
assign LUT_3[23552] = 32'b00000000000000010001011011001101;
assign LUT_3[23553] = 32'b00000000000000011000000110101010;
assign LUT_3[23554] = 32'b00000000000000010011100010110001;
assign LUT_3[23555] = 32'b00000000000000011010001110001110;
assign LUT_3[23556] = 32'b00000000000000001110101001000011;
assign LUT_3[23557] = 32'b00000000000000010101010100100000;
assign LUT_3[23558] = 32'b00000000000000010000110000100111;
assign LUT_3[23559] = 32'b00000000000000010111011100000100;
assign LUT_3[23560] = 32'b00000000000000010110110100010011;
assign LUT_3[23561] = 32'b00000000000000011101011111110000;
assign LUT_3[23562] = 32'b00000000000000011000111011110111;
assign LUT_3[23563] = 32'b00000000000000011111100111010100;
assign LUT_3[23564] = 32'b00000000000000010100000010001001;
assign LUT_3[23565] = 32'b00000000000000011010101101100110;
assign LUT_3[23566] = 32'b00000000000000010110001001101101;
assign LUT_3[23567] = 32'b00000000000000011100110101001010;
assign LUT_3[23568] = 32'b00000000000000010100101110010000;
assign LUT_3[23569] = 32'b00000000000000011011011001101101;
assign LUT_3[23570] = 32'b00000000000000010110110101110100;
assign LUT_3[23571] = 32'b00000000000000011101100001010001;
assign LUT_3[23572] = 32'b00000000000000010001111100000110;
assign LUT_3[23573] = 32'b00000000000000011000100111100011;
assign LUT_3[23574] = 32'b00000000000000010100000011101010;
assign LUT_3[23575] = 32'b00000000000000011010101111000111;
assign LUT_3[23576] = 32'b00000000000000011010000111010110;
assign LUT_3[23577] = 32'b00000000000000100000110010110011;
assign LUT_3[23578] = 32'b00000000000000011100001110111010;
assign LUT_3[23579] = 32'b00000000000000100010111010010111;
assign LUT_3[23580] = 32'b00000000000000010111010101001100;
assign LUT_3[23581] = 32'b00000000000000011110000000101001;
assign LUT_3[23582] = 32'b00000000000000011001011100110000;
assign LUT_3[23583] = 32'b00000000000000100000001000001101;
assign LUT_3[23584] = 32'b00000000000000010010101001101101;
assign LUT_3[23585] = 32'b00000000000000011001010101001010;
assign LUT_3[23586] = 32'b00000000000000010100110001010001;
assign LUT_3[23587] = 32'b00000000000000011011011100101110;
assign LUT_3[23588] = 32'b00000000000000001111110111100011;
assign LUT_3[23589] = 32'b00000000000000010110100011000000;
assign LUT_3[23590] = 32'b00000000000000010001111111000111;
assign LUT_3[23591] = 32'b00000000000000011000101010100100;
assign LUT_3[23592] = 32'b00000000000000011000000010110011;
assign LUT_3[23593] = 32'b00000000000000011110101110010000;
assign LUT_3[23594] = 32'b00000000000000011010001010010111;
assign LUT_3[23595] = 32'b00000000000000100000110101110100;
assign LUT_3[23596] = 32'b00000000000000010101010000101001;
assign LUT_3[23597] = 32'b00000000000000011011111100000110;
assign LUT_3[23598] = 32'b00000000000000010111011000001101;
assign LUT_3[23599] = 32'b00000000000000011110000011101010;
assign LUT_3[23600] = 32'b00000000000000010101111100110000;
assign LUT_3[23601] = 32'b00000000000000011100101000001101;
assign LUT_3[23602] = 32'b00000000000000011000000100010100;
assign LUT_3[23603] = 32'b00000000000000011110101111110001;
assign LUT_3[23604] = 32'b00000000000000010011001010100110;
assign LUT_3[23605] = 32'b00000000000000011001110110000011;
assign LUT_3[23606] = 32'b00000000000000010101010010001010;
assign LUT_3[23607] = 32'b00000000000000011011111101100111;
assign LUT_3[23608] = 32'b00000000000000011011010101110110;
assign LUT_3[23609] = 32'b00000000000000100010000001010011;
assign LUT_3[23610] = 32'b00000000000000011101011101011010;
assign LUT_3[23611] = 32'b00000000000000100100001000110111;
assign LUT_3[23612] = 32'b00000000000000011000100011101100;
assign LUT_3[23613] = 32'b00000000000000011111001111001001;
assign LUT_3[23614] = 32'b00000000000000011010101011010000;
assign LUT_3[23615] = 32'b00000000000000100001010110101101;
assign LUT_3[23616] = 32'b00000000000000010001010011111000;
assign LUT_3[23617] = 32'b00000000000000010111111111010101;
assign LUT_3[23618] = 32'b00000000000000010011011011011100;
assign LUT_3[23619] = 32'b00000000000000011010000110111001;
assign LUT_3[23620] = 32'b00000000000000001110100001101110;
assign LUT_3[23621] = 32'b00000000000000010101001101001011;
assign LUT_3[23622] = 32'b00000000000000010000101001010010;
assign LUT_3[23623] = 32'b00000000000000010111010100101111;
assign LUT_3[23624] = 32'b00000000000000010110101100111110;
assign LUT_3[23625] = 32'b00000000000000011101011000011011;
assign LUT_3[23626] = 32'b00000000000000011000110100100010;
assign LUT_3[23627] = 32'b00000000000000011111011111111111;
assign LUT_3[23628] = 32'b00000000000000010011111010110100;
assign LUT_3[23629] = 32'b00000000000000011010100110010001;
assign LUT_3[23630] = 32'b00000000000000010110000010011000;
assign LUT_3[23631] = 32'b00000000000000011100101101110101;
assign LUT_3[23632] = 32'b00000000000000010100100110111011;
assign LUT_3[23633] = 32'b00000000000000011011010010011000;
assign LUT_3[23634] = 32'b00000000000000010110101110011111;
assign LUT_3[23635] = 32'b00000000000000011101011001111100;
assign LUT_3[23636] = 32'b00000000000000010001110100110001;
assign LUT_3[23637] = 32'b00000000000000011000100000001110;
assign LUT_3[23638] = 32'b00000000000000010011111100010101;
assign LUT_3[23639] = 32'b00000000000000011010100111110010;
assign LUT_3[23640] = 32'b00000000000000011010000000000001;
assign LUT_3[23641] = 32'b00000000000000100000101011011110;
assign LUT_3[23642] = 32'b00000000000000011100000111100101;
assign LUT_3[23643] = 32'b00000000000000100010110011000010;
assign LUT_3[23644] = 32'b00000000000000010111001101110111;
assign LUT_3[23645] = 32'b00000000000000011101111001010100;
assign LUT_3[23646] = 32'b00000000000000011001010101011011;
assign LUT_3[23647] = 32'b00000000000000100000000000111000;
assign LUT_3[23648] = 32'b00000000000000010010100010011000;
assign LUT_3[23649] = 32'b00000000000000011001001101110101;
assign LUT_3[23650] = 32'b00000000000000010100101001111100;
assign LUT_3[23651] = 32'b00000000000000011011010101011001;
assign LUT_3[23652] = 32'b00000000000000001111110000001110;
assign LUT_3[23653] = 32'b00000000000000010110011011101011;
assign LUT_3[23654] = 32'b00000000000000010001110111110010;
assign LUT_3[23655] = 32'b00000000000000011000100011001111;
assign LUT_3[23656] = 32'b00000000000000010111111011011110;
assign LUT_3[23657] = 32'b00000000000000011110100110111011;
assign LUT_3[23658] = 32'b00000000000000011010000011000010;
assign LUT_3[23659] = 32'b00000000000000100000101110011111;
assign LUT_3[23660] = 32'b00000000000000010101001001010100;
assign LUT_3[23661] = 32'b00000000000000011011110100110001;
assign LUT_3[23662] = 32'b00000000000000010111010000111000;
assign LUT_3[23663] = 32'b00000000000000011101111100010101;
assign LUT_3[23664] = 32'b00000000000000010101110101011011;
assign LUT_3[23665] = 32'b00000000000000011100100000111000;
assign LUT_3[23666] = 32'b00000000000000010111111100111111;
assign LUT_3[23667] = 32'b00000000000000011110101000011100;
assign LUT_3[23668] = 32'b00000000000000010011000011010001;
assign LUT_3[23669] = 32'b00000000000000011001101110101110;
assign LUT_3[23670] = 32'b00000000000000010101001010110101;
assign LUT_3[23671] = 32'b00000000000000011011110110010010;
assign LUT_3[23672] = 32'b00000000000000011011001110100001;
assign LUT_3[23673] = 32'b00000000000000100001111001111110;
assign LUT_3[23674] = 32'b00000000000000011101010110000101;
assign LUT_3[23675] = 32'b00000000000000100100000001100010;
assign LUT_3[23676] = 32'b00000000000000011000011100010111;
assign LUT_3[23677] = 32'b00000000000000011111000111110100;
assign LUT_3[23678] = 32'b00000000000000011010100011111011;
assign LUT_3[23679] = 32'b00000000000000100001001111011000;
assign LUT_3[23680] = 32'b00000000000000010011100110001011;
assign LUT_3[23681] = 32'b00000000000000011010010001101000;
assign LUT_3[23682] = 32'b00000000000000010101101101101111;
assign LUT_3[23683] = 32'b00000000000000011100011001001100;
assign LUT_3[23684] = 32'b00000000000000010000110100000001;
assign LUT_3[23685] = 32'b00000000000000010111011111011110;
assign LUT_3[23686] = 32'b00000000000000010010111011100101;
assign LUT_3[23687] = 32'b00000000000000011001100111000010;
assign LUT_3[23688] = 32'b00000000000000011000111111010001;
assign LUT_3[23689] = 32'b00000000000000011111101010101110;
assign LUT_3[23690] = 32'b00000000000000011011000110110101;
assign LUT_3[23691] = 32'b00000000000000100001110010010010;
assign LUT_3[23692] = 32'b00000000000000010110001101000111;
assign LUT_3[23693] = 32'b00000000000000011100111000100100;
assign LUT_3[23694] = 32'b00000000000000011000010100101011;
assign LUT_3[23695] = 32'b00000000000000011111000000001000;
assign LUT_3[23696] = 32'b00000000000000010110111001001110;
assign LUT_3[23697] = 32'b00000000000000011101100100101011;
assign LUT_3[23698] = 32'b00000000000000011001000000110010;
assign LUT_3[23699] = 32'b00000000000000011111101100001111;
assign LUT_3[23700] = 32'b00000000000000010100000111000100;
assign LUT_3[23701] = 32'b00000000000000011010110010100001;
assign LUT_3[23702] = 32'b00000000000000010110001110101000;
assign LUT_3[23703] = 32'b00000000000000011100111010000101;
assign LUT_3[23704] = 32'b00000000000000011100010010010100;
assign LUT_3[23705] = 32'b00000000000000100010111101110001;
assign LUT_3[23706] = 32'b00000000000000011110011001111000;
assign LUT_3[23707] = 32'b00000000000000100101000101010101;
assign LUT_3[23708] = 32'b00000000000000011001100000001010;
assign LUT_3[23709] = 32'b00000000000000100000001011100111;
assign LUT_3[23710] = 32'b00000000000000011011100111101110;
assign LUT_3[23711] = 32'b00000000000000100010010011001011;
assign LUT_3[23712] = 32'b00000000000000010100110100101011;
assign LUT_3[23713] = 32'b00000000000000011011100000001000;
assign LUT_3[23714] = 32'b00000000000000010110111100001111;
assign LUT_3[23715] = 32'b00000000000000011101100111101100;
assign LUT_3[23716] = 32'b00000000000000010010000010100001;
assign LUT_3[23717] = 32'b00000000000000011000101101111110;
assign LUT_3[23718] = 32'b00000000000000010100001010000101;
assign LUT_3[23719] = 32'b00000000000000011010110101100010;
assign LUT_3[23720] = 32'b00000000000000011010001101110001;
assign LUT_3[23721] = 32'b00000000000000100000111001001110;
assign LUT_3[23722] = 32'b00000000000000011100010101010101;
assign LUT_3[23723] = 32'b00000000000000100011000000110010;
assign LUT_3[23724] = 32'b00000000000000010111011011100111;
assign LUT_3[23725] = 32'b00000000000000011110000111000100;
assign LUT_3[23726] = 32'b00000000000000011001100011001011;
assign LUT_3[23727] = 32'b00000000000000100000001110101000;
assign LUT_3[23728] = 32'b00000000000000011000000111101110;
assign LUT_3[23729] = 32'b00000000000000011110110011001011;
assign LUT_3[23730] = 32'b00000000000000011010001111010010;
assign LUT_3[23731] = 32'b00000000000000100000111010101111;
assign LUT_3[23732] = 32'b00000000000000010101010101100100;
assign LUT_3[23733] = 32'b00000000000000011100000001000001;
assign LUT_3[23734] = 32'b00000000000000010111011101001000;
assign LUT_3[23735] = 32'b00000000000000011110001000100101;
assign LUT_3[23736] = 32'b00000000000000011101100000110100;
assign LUT_3[23737] = 32'b00000000000000100100001100010001;
assign LUT_3[23738] = 32'b00000000000000011111101000011000;
assign LUT_3[23739] = 32'b00000000000000100110010011110101;
assign LUT_3[23740] = 32'b00000000000000011010101110101010;
assign LUT_3[23741] = 32'b00000000000000100001011010000111;
assign LUT_3[23742] = 32'b00000000000000011100110110001110;
assign LUT_3[23743] = 32'b00000000000000100011100001101011;
assign LUT_3[23744] = 32'b00000000000000010011011110110110;
assign LUT_3[23745] = 32'b00000000000000011010001010010011;
assign LUT_3[23746] = 32'b00000000000000010101100110011010;
assign LUT_3[23747] = 32'b00000000000000011100010001110111;
assign LUT_3[23748] = 32'b00000000000000010000101100101100;
assign LUT_3[23749] = 32'b00000000000000010111011000001001;
assign LUT_3[23750] = 32'b00000000000000010010110100010000;
assign LUT_3[23751] = 32'b00000000000000011001011111101101;
assign LUT_3[23752] = 32'b00000000000000011000110111111100;
assign LUT_3[23753] = 32'b00000000000000011111100011011001;
assign LUT_3[23754] = 32'b00000000000000011010111111100000;
assign LUT_3[23755] = 32'b00000000000000100001101010111101;
assign LUT_3[23756] = 32'b00000000000000010110000101110010;
assign LUT_3[23757] = 32'b00000000000000011100110001001111;
assign LUT_3[23758] = 32'b00000000000000011000001101010110;
assign LUT_3[23759] = 32'b00000000000000011110111000110011;
assign LUT_3[23760] = 32'b00000000000000010110110001111001;
assign LUT_3[23761] = 32'b00000000000000011101011101010110;
assign LUT_3[23762] = 32'b00000000000000011000111001011101;
assign LUT_3[23763] = 32'b00000000000000011111100100111010;
assign LUT_3[23764] = 32'b00000000000000010011111111101111;
assign LUT_3[23765] = 32'b00000000000000011010101011001100;
assign LUT_3[23766] = 32'b00000000000000010110000111010011;
assign LUT_3[23767] = 32'b00000000000000011100110010110000;
assign LUT_3[23768] = 32'b00000000000000011100001010111111;
assign LUT_3[23769] = 32'b00000000000000100010110110011100;
assign LUT_3[23770] = 32'b00000000000000011110010010100011;
assign LUT_3[23771] = 32'b00000000000000100100111110000000;
assign LUT_3[23772] = 32'b00000000000000011001011000110101;
assign LUT_3[23773] = 32'b00000000000000100000000100010010;
assign LUT_3[23774] = 32'b00000000000000011011100000011001;
assign LUT_3[23775] = 32'b00000000000000100010001011110110;
assign LUT_3[23776] = 32'b00000000000000010100101101010110;
assign LUT_3[23777] = 32'b00000000000000011011011000110011;
assign LUT_3[23778] = 32'b00000000000000010110110100111010;
assign LUT_3[23779] = 32'b00000000000000011101100000010111;
assign LUT_3[23780] = 32'b00000000000000010001111011001100;
assign LUT_3[23781] = 32'b00000000000000011000100110101001;
assign LUT_3[23782] = 32'b00000000000000010100000010110000;
assign LUT_3[23783] = 32'b00000000000000011010101110001101;
assign LUT_3[23784] = 32'b00000000000000011010000110011100;
assign LUT_3[23785] = 32'b00000000000000100000110001111001;
assign LUT_3[23786] = 32'b00000000000000011100001110000000;
assign LUT_3[23787] = 32'b00000000000000100010111001011101;
assign LUT_3[23788] = 32'b00000000000000010111010100010010;
assign LUT_3[23789] = 32'b00000000000000011101111111101111;
assign LUT_3[23790] = 32'b00000000000000011001011011110110;
assign LUT_3[23791] = 32'b00000000000000100000000111010011;
assign LUT_3[23792] = 32'b00000000000000011000000000011001;
assign LUT_3[23793] = 32'b00000000000000011110101011110110;
assign LUT_3[23794] = 32'b00000000000000011010000111111101;
assign LUT_3[23795] = 32'b00000000000000100000110011011010;
assign LUT_3[23796] = 32'b00000000000000010101001110001111;
assign LUT_3[23797] = 32'b00000000000000011011111001101100;
assign LUT_3[23798] = 32'b00000000000000010111010101110011;
assign LUT_3[23799] = 32'b00000000000000011110000001010000;
assign LUT_3[23800] = 32'b00000000000000011101011001011111;
assign LUT_3[23801] = 32'b00000000000000100100000100111100;
assign LUT_3[23802] = 32'b00000000000000011111100001000011;
assign LUT_3[23803] = 32'b00000000000000100110001100100000;
assign LUT_3[23804] = 32'b00000000000000011010100111010101;
assign LUT_3[23805] = 32'b00000000000000100001010010110010;
assign LUT_3[23806] = 32'b00000000000000011100101110111001;
assign LUT_3[23807] = 32'b00000000000000100011011010010110;
assign LUT_3[23808] = 32'b00000000000000001101101010101110;
assign LUT_3[23809] = 32'b00000000000000010100010110001011;
assign LUT_3[23810] = 32'b00000000000000001111110010010010;
assign LUT_3[23811] = 32'b00000000000000010110011101101111;
assign LUT_3[23812] = 32'b00000000000000001010111000100100;
assign LUT_3[23813] = 32'b00000000000000010001100100000001;
assign LUT_3[23814] = 32'b00000000000000001101000000001000;
assign LUT_3[23815] = 32'b00000000000000010011101011100101;
assign LUT_3[23816] = 32'b00000000000000010011000011110100;
assign LUT_3[23817] = 32'b00000000000000011001101111010001;
assign LUT_3[23818] = 32'b00000000000000010101001011011000;
assign LUT_3[23819] = 32'b00000000000000011011110110110101;
assign LUT_3[23820] = 32'b00000000000000010000010001101010;
assign LUT_3[23821] = 32'b00000000000000010110111101000111;
assign LUT_3[23822] = 32'b00000000000000010010011001001110;
assign LUT_3[23823] = 32'b00000000000000011001000100101011;
assign LUT_3[23824] = 32'b00000000000000010000111101110001;
assign LUT_3[23825] = 32'b00000000000000010111101001001110;
assign LUT_3[23826] = 32'b00000000000000010011000101010101;
assign LUT_3[23827] = 32'b00000000000000011001110000110010;
assign LUT_3[23828] = 32'b00000000000000001110001011100111;
assign LUT_3[23829] = 32'b00000000000000010100110111000100;
assign LUT_3[23830] = 32'b00000000000000010000010011001011;
assign LUT_3[23831] = 32'b00000000000000010110111110101000;
assign LUT_3[23832] = 32'b00000000000000010110010110110111;
assign LUT_3[23833] = 32'b00000000000000011101000010010100;
assign LUT_3[23834] = 32'b00000000000000011000011110011011;
assign LUT_3[23835] = 32'b00000000000000011111001001111000;
assign LUT_3[23836] = 32'b00000000000000010011100100101101;
assign LUT_3[23837] = 32'b00000000000000011010010000001010;
assign LUT_3[23838] = 32'b00000000000000010101101100010001;
assign LUT_3[23839] = 32'b00000000000000011100010111101110;
assign LUT_3[23840] = 32'b00000000000000001110111001001110;
assign LUT_3[23841] = 32'b00000000000000010101100100101011;
assign LUT_3[23842] = 32'b00000000000000010001000000110010;
assign LUT_3[23843] = 32'b00000000000000010111101100001111;
assign LUT_3[23844] = 32'b00000000000000001100000111000100;
assign LUT_3[23845] = 32'b00000000000000010010110010100001;
assign LUT_3[23846] = 32'b00000000000000001110001110101000;
assign LUT_3[23847] = 32'b00000000000000010100111010000101;
assign LUT_3[23848] = 32'b00000000000000010100010010010100;
assign LUT_3[23849] = 32'b00000000000000011010111101110001;
assign LUT_3[23850] = 32'b00000000000000010110011001111000;
assign LUT_3[23851] = 32'b00000000000000011101000101010101;
assign LUT_3[23852] = 32'b00000000000000010001100000001010;
assign LUT_3[23853] = 32'b00000000000000011000001011100111;
assign LUT_3[23854] = 32'b00000000000000010011100111101110;
assign LUT_3[23855] = 32'b00000000000000011010010011001011;
assign LUT_3[23856] = 32'b00000000000000010010001100010001;
assign LUT_3[23857] = 32'b00000000000000011000110111101110;
assign LUT_3[23858] = 32'b00000000000000010100010011110101;
assign LUT_3[23859] = 32'b00000000000000011010111111010010;
assign LUT_3[23860] = 32'b00000000000000001111011010000111;
assign LUT_3[23861] = 32'b00000000000000010110000101100100;
assign LUT_3[23862] = 32'b00000000000000010001100001101011;
assign LUT_3[23863] = 32'b00000000000000011000001101001000;
assign LUT_3[23864] = 32'b00000000000000010111100101010111;
assign LUT_3[23865] = 32'b00000000000000011110010000110100;
assign LUT_3[23866] = 32'b00000000000000011001101100111011;
assign LUT_3[23867] = 32'b00000000000000100000011000011000;
assign LUT_3[23868] = 32'b00000000000000010100110011001101;
assign LUT_3[23869] = 32'b00000000000000011011011110101010;
assign LUT_3[23870] = 32'b00000000000000010110111010110001;
assign LUT_3[23871] = 32'b00000000000000011101100110001110;
assign LUT_3[23872] = 32'b00000000000000001101100011011001;
assign LUT_3[23873] = 32'b00000000000000010100001110110110;
assign LUT_3[23874] = 32'b00000000000000001111101010111101;
assign LUT_3[23875] = 32'b00000000000000010110010110011010;
assign LUT_3[23876] = 32'b00000000000000001010110001001111;
assign LUT_3[23877] = 32'b00000000000000010001011100101100;
assign LUT_3[23878] = 32'b00000000000000001100111000110011;
assign LUT_3[23879] = 32'b00000000000000010011100100010000;
assign LUT_3[23880] = 32'b00000000000000010010111100011111;
assign LUT_3[23881] = 32'b00000000000000011001100111111100;
assign LUT_3[23882] = 32'b00000000000000010101000100000011;
assign LUT_3[23883] = 32'b00000000000000011011101111100000;
assign LUT_3[23884] = 32'b00000000000000010000001010010101;
assign LUT_3[23885] = 32'b00000000000000010110110101110010;
assign LUT_3[23886] = 32'b00000000000000010010010001111001;
assign LUT_3[23887] = 32'b00000000000000011000111101010110;
assign LUT_3[23888] = 32'b00000000000000010000110110011100;
assign LUT_3[23889] = 32'b00000000000000010111100001111001;
assign LUT_3[23890] = 32'b00000000000000010010111110000000;
assign LUT_3[23891] = 32'b00000000000000011001101001011101;
assign LUT_3[23892] = 32'b00000000000000001110000100010010;
assign LUT_3[23893] = 32'b00000000000000010100101111101111;
assign LUT_3[23894] = 32'b00000000000000010000001011110110;
assign LUT_3[23895] = 32'b00000000000000010110110111010011;
assign LUT_3[23896] = 32'b00000000000000010110001111100010;
assign LUT_3[23897] = 32'b00000000000000011100111010111111;
assign LUT_3[23898] = 32'b00000000000000011000010111000110;
assign LUT_3[23899] = 32'b00000000000000011111000010100011;
assign LUT_3[23900] = 32'b00000000000000010011011101011000;
assign LUT_3[23901] = 32'b00000000000000011010001000110101;
assign LUT_3[23902] = 32'b00000000000000010101100100111100;
assign LUT_3[23903] = 32'b00000000000000011100010000011001;
assign LUT_3[23904] = 32'b00000000000000001110110001111001;
assign LUT_3[23905] = 32'b00000000000000010101011101010110;
assign LUT_3[23906] = 32'b00000000000000010000111001011101;
assign LUT_3[23907] = 32'b00000000000000010111100100111010;
assign LUT_3[23908] = 32'b00000000000000001011111111101111;
assign LUT_3[23909] = 32'b00000000000000010010101011001100;
assign LUT_3[23910] = 32'b00000000000000001110000111010011;
assign LUT_3[23911] = 32'b00000000000000010100110010110000;
assign LUT_3[23912] = 32'b00000000000000010100001010111111;
assign LUT_3[23913] = 32'b00000000000000011010110110011100;
assign LUT_3[23914] = 32'b00000000000000010110010010100011;
assign LUT_3[23915] = 32'b00000000000000011100111110000000;
assign LUT_3[23916] = 32'b00000000000000010001011000110101;
assign LUT_3[23917] = 32'b00000000000000011000000100010010;
assign LUT_3[23918] = 32'b00000000000000010011100000011001;
assign LUT_3[23919] = 32'b00000000000000011010001011110110;
assign LUT_3[23920] = 32'b00000000000000010010000100111100;
assign LUT_3[23921] = 32'b00000000000000011000110000011001;
assign LUT_3[23922] = 32'b00000000000000010100001100100000;
assign LUT_3[23923] = 32'b00000000000000011010110111111101;
assign LUT_3[23924] = 32'b00000000000000001111010010110010;
assign LUT_3[23925] = 32'b00000000000000010101111110001111;
assign LUT_3[23926] = 32'b00000000000000010001011010010110;
assign LUT_3[23927] = 32'b00000000000000011000000101110011;
assign LUT_3[23928] = 32'b00000000000000010111011110000010;
assign LUT_3[23929] = 32'b00000000000000011110001001011111;
assign LUT_3[23930] = 32'b00000000000000011001100101100110;
assign LUT_3[23931] = 32'b00000000000000100000010001000011;
assign LUT_3[23932] = 32'b00000000000000010100101011111000;
assign LUT_3[23933] = 32'b00000000000000011011010111010101;
assign LUT_3[23934] = 32'b00000000000000010110110011011100;
assign LUT_3[23935] = 32'b00000000000000011101011110111001;
assign LUT_3[23936] = 32'b00000000000000001111110101101100;
assign LUT_3[23937] = 32'b00000000000000010110100001001001;
assign LUT_3[23938] = 32'b00000000000000010001111101010000;
assign LUT_3[23939] = 32'b00000000000000011000101000101101;
assign LUT_3[23940] = 32'b00000000000000001101000011100010;
assign LUT_3[23941] = 32'b00000000000000010011101110111111;
assign LUT_3[23942] = 32'b00000000000000001111001011000110;
assign LUT_3[23943] = 32'b00000000000000010101110110100011;
assign LUT_3[23944] = 32'b00000000000000010101001110110010;
assign LUT_3[23945] = 32'b00000000000000011011111010001111;
assign LUT_3[23946] = 32'b00000000000000010111010110010110;
assign LUT_3[23947] = 32'b00000000000000011110000001110011;
assign LUT_3[23948] = 32'b00000000000000010010011100101000;
assign LUT_3[23949] = 32'b00000000000000011001001000000101;
assign LUT_3[23950] = 32'b00000000000000010100100100001100;
assign LUT_3[23951] = 32'b00000000000000011011001111101001;
assign LUT_3[23952] = 32'b00000000000000010011001000101111;
assign LUT_3[23953] = 32'b00000000000000011001110100001100;
assign LUT_3[23954] = 32'b00000000000000010101010000010011;
assign LUT_3[23955] = 32'b00000000000000011011111011110000;
assign LUT_3[23956] = 32'b00000000000000010000010110100101;
assign LUT_3[23957] = 32'b00000000000000010111000010000010;
assign LUT_3[23958] = 32'b00000000000000010010011110001001;
assign LUT_3[23959] = 32'b00000000000000011001001001100110;
assign LUT_3[23960] = 32'b00000000000000011000100001110101;
assign LUT_3[23961] = 32'b00000000000000011111001101010010;
assign LUT_3[23962] = 32'b00000000000000011010101001011001;
assign LUT_3[23963] = 32'b00000000000000100001010100110110;
assign LUT_3[23964] = 32'b00000000000000010101101111101011;
assign LUT_3[23965] = 32'b00000000000000011100011011001000;
assign LUT_3[23966] = 32'b00000000000000010111110111001111;
assign LUT_3[23967] = 32'b00000000000000011110100010101100;
assign LUT_3[23968] = 32'b00000000000000010001000100001100;
assign LUT_3[23969] = 32'b00000000000000010111101111101001;
assign LUT_3[23970] = 32'b00000000000000010011001011110000;
assign LUT_3[23971] = 32'b00000000000000011001110111001101;
assign LUT_3[23972] = 32'b00000000000000001110010010000010;
assign LUT_3[23973] = 32'b00000000000000010100111101011111;
assign LUT_3[23974] = 32'b00000000000000010000011001100110;
assign LUT_3[23975] = 32'b00000000000000010111000101000011;
assign LUT_3[23976] = 32'b00000000000000010110011101010010;
assign LUT_3[23977] = 32'b00000000000000011101001000101111;
assign LUT_3[23978] = 32'b00000000000000011000100100110110;
assign LUT_3[23979] = 32'b00000000000000011111010000010011;
assign LUT_3[23980] = 32'b00000000000000010011101011001000;
assign LUT_3[23981] = 32'b00000000000000011010010110100101;
assign LUT_3[23982] = 32'b00000000000000010101110010101100;
assign LUT_3[23983] = 32'b00000000000000011100011110001001;
assign LUT_3[23984] = 32'b00000000000000010100010111001111;
assign LUT_3[23985] = 32'b00000000000000011011000010101100;
assign LUT_3[23986] = 32'b00000000000000010110011110110011;
assign LUT_3[23987] = 32'b00000000000000011101001010010000;
assign LUT_3[23988] = 32'b00000000000000010001100101000101;
assign LUT_3[23989] = 32'b00000000000000011000010000100010;
assign LUT_3[23990] = 32'b00000000000000010011101100101001;
assign LUT_3[23991] = 32'b00000000000000011010011000000110;
assign LUT_3[23992] = 32'b00000000000000011001110000010101;
assign LUT_3[23993] = 32'b00000000000000100000011011110010;
assign LUT_3[23994] = 32'b00000000000000011011110111111001;
assign LUT_3[23995] = 32'b00000000000000100010100011010110;
assign LUT_3[23996] = 32'b00000000000000010110111110001011;
assign LUT_3[23997] = 32'b00000000000000011101101001101000;
assign LUT_3[23998] = 32'b00000000000000011001000101101111;
assign LUT_3[23999] = 32'b00000000000000011111110001001100;
assign LUT_3[24000] = 32'b00000000000000001111101110010111;
assign LUT_3[24001] = 32'b00000000000000010110011001110100;
assign LUT_3[24002] = 32'b00000000000000010001110101111011;
assign LUT_3[24003] = 32'b00000000000000011000100001011000;
assign LUT_3[24004] = 32'b00000000000000001100111100001101;
assign LUT_3[24005] = 32'b00000000000000010011100111101010;
assign LUT_3[24006] = 32'b00000000000000001111000011110001;
assign LUT_3[24007] = 32'b00000000000000010101101111001110;
assign LUT_3[24008] = 32'b00000000000000010101000111011101;
assign LUT_3[24009] = 32'b00000000000000011011110010111010;
assign LUT_3[24010] = 32'b00000000000000010111001111000001;
assign LUT_3[24011] = 32'b00000000000000011101111010011110;
assign LUT_3[24012] = 32'b00000000000000010010010101010011;
assign LUT_3[24013] = 32'b00000000000000011001000000110000;
assign LUT_3[24014] = 32'b00000000000000010100011100110111;
assign LUT_3[24015] = 32'b00000000000000011011001000010100;
assign LUT_3[24016] = 32'b00000000000000010011000001011010;
assign LUT_3[24017] = 32'b00000000000000011001101100110111;
assign LUT_3[24018] = 32'b00000000000000010101001000111110;
assign LUT_3[24019] = 32'b00000000000000011011110100011011;
assign LUT_3[24020] = 32'b00000000000000010000001111010000;
assign LUT_3[24021] = 32'b00000000000000010110111010101101;
assign LUT_3[24022] = 32'b00000000000000010010010110110100;
assign LUT_3[24023] = 32'b00000000000000011001000010010001;
assign LUT_3[24024] = 32'b00000000000000011000011010100000;
assign LUT_3[24025] = 32'b00000000000000011111000101111101;
assign LUT_3[24026] = 32'b00000000000000011010100010000100;
assign LUT_3[24027] = 32'b00000000000000100001001101100001;
assign LUT_3[24028] = 32'b00000000000000010101101000010110;
assign LUT_3[24029] = 32'b00000000000000011100010011110011;
assign LUT_3[24030] = 32'b00000000000000010111101111111010;
assign LUT_3[24031] = 32'b00000000000000011110011011010111;
assign LUT_3[24032] = 32'b00000000000000010000111100110111;
assign LUT_3[24033] = 32'b00000000000000010111101000010100;
assign LUT_3[24034] = 32'b00000000000000010011000100011011;
assign LUT_3[24035] = 32'b00000000000000011001101111111000;
assign LUT_3[24036] = 32'b00000000000000001110001010101101;
assign LUT_3[24037] = 32'b00000000000000010100110110001010;
assign LUT_3[24038] = 32'b00000000000000010000010010010001;
assign LUT_3[24039] = 32'b00000000000000010110111101101110;
assign LUT_3[24040] = 32'b00000000000000010110010101111101;
assign LUT_3[24041] = 32'b00000000000000011101000001011010;
assign LUT_3[24042] = 32'b00000000000000011000011101100001;
assign LUT_3[24043] = 32'b00000000000000011111001000111110;
assign LUT_3[24044] = 32'b00000000000000010011100011110011;
assign LUT_3[24045] = 32'b00000000000000011010001111010000;
assign LUT_3[24046] = 32'b00000000000000010101101011010111;
assign LUT_3[24047] = 32'b00000000000000011100010110110100;
assign LUT_3[24048] = 32'b00000000000000010100001111111010;
assign LUT_3[24049] = 32'b00000000000000011010111011010111;
assign LUT_3[24050] = 32'b00000000000000010110010111011110;
assign LUT_3[24051] = 32'b00000000000000011101000010111011;
assign LUT_3[24052] = 32'b00000000000000010001011101110000;
assign LUT_3[24053] = 32'b00000000000000011000001001001101;
assign LUT_3[24054] = 32'b00000000000000010011100101010100;
assign LUT_3[24055] = 32'b00000000000000011010010000110001;
assign LUT_3[24056] = 32'b00000000000000011001101001000000;
assign LUT_3[24057] = 32'b00000000000000100000010100011101;
assign LUT_3[24058] = 32'b00000000000000011011110000100100;
assign LUT_3[24059] = 32'b00000000000000100010011100000001;
assign LUT_3[24060] = 32'b00000000000000010110110110110110;
assign LUT_3[24061] = 32'b00000000000000011101100010010011;
assign LUT_3[24062] = 32'b00000000000000011000111110011010;
assign LUT_3[24063] = 32'b00000000000000011111101001110111;
assign LUT_3[24064] = 32'b00000000000000010100110000011001;
assign LUT_3[24065] = 32'b00000000000000011011011011110110;
assign LUT_3[24066] = 32'b00000000000000010110110111111101;
assign LUT_3[24067] = 32'b00000000000000011101100011011010;
assign LUT_3[24068] = 32'b00000000000000010001111110001111;
assign LUT_3[24069] = 32'b00000000000000011000101001101100;
assign LUT_3[24070] = 32'b00000000000000010100000101110011;
assign LUT_3[24071] = 32'b00000000000000011010110001010000;
assign LUT_3[24072] = 32'b00000000000000011010001001011111;
assign LUT_3[24073] = 32'b00000000000000100000110100111100;
assign LUT_3[24074] = 32'b00000000000000011100010001000011;
assign LUT_3[24075] = 32'b00000000000000100010111100100000;
assign LUT_3[24076] = 32'b00000000000000010111010111010101;
assign LUT_3[24077] = 32'b00000000000000011110000010110010;
assign LUT_3[24078] = 32'b00000000000000011001011110111001;
assign LUT_3[24079] = 32'b00000000000000100000001010010110;
assign LUT_3[24080] = 32'b00000000000000011000000011011100;
assign LUT_3[24081] = 32'b00000000000000011110101110111001;
assign LUT_3[24082] = 32'b00000000000000011010001011000000;
assign LUT_3[24083] = 32'b00000000000000100000110110011101;
assign LUT_3[24084] = 32'b00000000000000010101010001010010;
assign LUT_3[24085] = 32'b00000000000000011011111100101111;
assign LUT_3[24086] = 32'b00000000000000010111011000110110;
assign LUT_3[24087] = 32'b00000000000000011110000100010011;
assign LUT_3[24088] = 32'b00000000000000011101011100100010;
assign LUT_3[24089] = 32'b00000000000000100100000111111111;
assign LUT_3[24090] = 32'b00000000000000011111100100000110;
assign LUT_3[24091] = 32'b00000000000000100110001111100011;
assign LUT_3[24092] = 32'b00000000000000011010101010011000;
assign LUT_3[24093] = 32'b00000000000000100001010101110101;
assign LUT_3[24094] = 32'b00000000000000011100110001111100;
assign LUT_3[24095] = 32'b00000000000000100011011101011001;
assign LUT_3[24096] = 32'b00000000000000010101111110111001;
assign LUT_3[24097] = 32'b00000000000000011100101010010110;
assign LUT_3[24098] = 32'b00000000000000011000000110011101;
assign LUT_3[24099] = 32'b00000000000000011110110001111010;
assign LUT_3[24100] = 32'b00000000000000010011001100101111;
assign LUT_3[24101] = 32'b00000000000000011001111000001100;
assign LUT_3[24102] = 32'b00000000000000010101010100010011;
assign LUT_3[24103] = 32'b00000000000000011011111111110000;
assign LUT_3[24104] = 32'b00000000000000011011010111111111;
assign LUT_3[24105] = 32'b00000000000000100010000011011100;
assign LUT_3[24106] = 32'b00000000000000011101011111100011;
assign LUT_3[24107] = 32'b00000000000000100100001011000000;
assign LUT_3[24108] = 32'b00000000000000011000100101110101;
assign LUT_3[24109] = 32'b00000000000000011111010001010010;
assign LUT_3[24110] = 32'b00000000000000011010101101011001;
assign LUT_3[24111] = 32'b00000000000000100001011000110110;
assign LUT_3[24112] = 32'b00000000000000011001010001111100;
assign LUT_3[24113] = 32'b00000000000000011111111101011001;
assign LUT_3[24114] = 32'b00000000000000011011011001100000;
assign LUT_3[24115] = 32'b00000000000000100010000100111101;
assign LUT_3[24116] = 32'b00000000000000010110011111110010;
assign LUT_3[24117] = 32'b00000000000000011101001011001111;
assign LUT_3[24118] = 32'b00000000000000011000100111010110;
assign LUT_3[24119] = 32'b00000000000000011111010010110011;
assign LUT_3[24120] = 32'b00000000000000011110101011000010;
assign LUT_3[24121] = 32'b00000000000000100101010110011111;
assign LUT_3[24122] = 32'b00000000000000100000110010100110;
assign LUT_3[24123] = 32'b00000000000000100111011110000011;
assign LUT_3[24124] = 32'b00000000000000011011111000111000;
assign LUT_3[24125] = 32'b00000000000000100010100100010101;
assign LUT_3[24126] = 32'b00000000000000011110000000011100;
assign LUT_3[24127] = 32'b00000000000000100100101011111001;
assign LUT_3[24128] = 32'b00000000000000010100101001000100;
assign LUT_3[24129] = 32'b00000000000000011011010100100001;
assign LUT_3[24130] = 32'b00000000000000010110110000101000;
assign LUT_3[24131] = 32'b00000000000000011101011100000101;
assign LUT_3[24132] = 32'b00000000000000010001110110111010;
assign LUT_3[24133] = 32'b00000000000000011000100010010111;
assign LUT_3[24134] = 32'b00000000000000010011111110011110;
assign LUT_3[24135] = 32'b00000000000000011010101001111011;
assign LUT_3[24136] = 32'b00000000000000011010000010001010;
assign LUT_3[24137] = 32'b00000000000000100000101101100111;
assign LUT_3[24138] = 32'b00000000000000011100001001101110;
assign LUT_3[24139] = 32'b00000000000000100010110101001011;
assign LUT_3[24140] = 32'b00000000000000010111010000000000;
assign LUT_3[24141] = 32'b00000000000000011101111011011101;
assign LUT_3[24142] = 32'b00000000000000011001010111100100;
assign LUT_3[24143] = 32'b00000000000000100000000011000001;
assign LUT_3[24144] = 32'b00000000000000010111111100000111;
assign LUT_3[24145] = 32'b00000000000000011110100111100100;
assign LUT_3[24146] = 32'b00000000000000011010000011101011;
assign LUT_3[24147] = 32'b00000000000000100000101111001000;
assign LUT_3[24148] = 32'b00000000000000010101001001111101;
assign LUT_3[24149] = 32'b00000000000000011011110101011010;
assign LUT_3[24150] = 32'b00000000000000010111010001100001;
assign LUT_3[24151] = 32'b00000000000000011101111100111110;
assign LUT_3[24152] = 32'b00000000000000011101010101001101;
assign LUT_3[24153] = 32'b00000000000000100100000000101010;
assign LUT_3[24154] = 32'b00000000000000011111011100110001;
assign LUT_3[24155] = 32'b00000000000000100110001000001110;
assign LUT_3[24156] = 32'b00000000000000011010100011000011;
assign LUT_3[24157] = 32'b00000000000000100001001110100000;
assign LUT_3[24158] = 32'b00000000000000011100101010100111;
assign LUT_3[24159] = 32'b00000000000000100011010110000100;
assign LUT_3[24160] = 32'b00000000000000010101110111100100;
assign LUT_3[24161] = 32'b00000000000000011100100011000001;
assign LUT_3[24162] = 32'b00000000000000010111111111001000;
assign LUT_3[24163] = 32'b00000000000000011110101010100101;
assign LUT_3[24164] = 32'b00000000000000010011000101011010;
assign LUT_3[24165] = 32'b00000000000000011001110000110111;
assign LUT_3[24166] = 32'b00000000000000010101001100111110;
assign LUT_3[24167] = 32'b00000000000000011011111000011011;
assign LUT_3[24168] = 32'b00000000000000011011010000101010;
assign LUT_3[24169] = 32'b00000000000000100001111100000111;
assign LUT_3[24170] = 32'b00000000000000011101011000001110;
assign LUT_3[24171] = 32'b00000000000000100100000011101011;
assign LUT_3[24172] = 32'b00000000000000011000011110100000;
assign LUT_3[24173] = 32'b00000000000000011111001001111101;
assign LUT_3[24174] = 32'b00000000000000011010100110000100;
assign LUT_3[24175] = 32'b00000000000000100001010001100001;
assign LUT_3[24176] = 32'b00000000000000011001001010100111;
assign LUT_3[24177] = 32'b00000000000000011111110110000100;
assign LUT_3[24178] = 32'b00000000000000011011010010001011;
assign LUT_3[24179] = 32'b00000000000000100001111101101000;
assign LUT_3[24180] = 32'b00000000000000010110011000011101;
assign LUT_3[24181] = 32'b00000000000000011101000011111010;
assign LUT_3[24182] = 32'b00000000000000011000100000000001;
assign LUT_3[24183] = 32'b00000000000000011111001011011110;
assign LUT_3[24184] = 32'b00000000000000011110100011101101;
assign LUT_3[24185] = 32'b00000000000000100101001111001010;
assign LUT_3[24186] = 32'b00000000000000100000101011010001;
assign LUT_3[24187] = 32'b00000000000000100111010110101110;
assign LUT_3[24188] = 32'b00000000000000011011110001100011;
assign LUT_3[24189] = 32'b00000000000000100010011101000000;
assign LUT_3[24190] = 32'b00000000000000011101111001000111;
assign LUT_3[24191] = 32'b00000000000000100100100100100100;
assign LUT_3[24192] = 32'b00000000000000010110111011010111;
assign LUT_3[24193] = 32'b00000000000000011101100110110100;
assign LUT_3[24194] = 32'b00000000000000011001000010111011;
assign LUT_3[24195] = 32'b00000000000000011111101110011000;
assign LUT_3[24196] = 32'b00000000000000010100001001001101;
assign LUT_3[24197] = 32'b00000000000000011010110100101010;
assign LUT_3[24198] = 32'b00000000000000010110010000110001;
assign LUT_3[24199] = 32'b00000000000000011100111100001110;
assign LUT_3[24200] = 32'b00000000000000011100010100011101;
assign LUT_3[24201] = 32'b00000000000000100010111111111010;
assign LUT_3[24202] = 32'b00000000000000011110011100000001;
assign LUT_3[24203] = 32'b00000000000000100101000111011110;
assign LUT_3[24204] = 32'b00000000000000011001100010010011;
assign LUT_3[24205] = 32'b00000000000000100000001101110000;
assign LUT_3[24206] = 32'b00000000000000011011101001110111;
assign LUT_3[24207] = 32'b00000000000000100010010101010100;
assign LUT_3[24208] = 32'b00000000000000011010001110011010;
assign LUT_3[24209] = 32'b00000000000000100000111001110111;
assign LUT_3[24210] = 32'b00000000000000011100010101111110;
assign LUT_3[24211] = 32'b00000000000000100011000001011011;
assign LUT_3[24212] = 32'b00000000000000010111011100010000;
assign LUT_3[24213] = 32'b00000000000000011110000111101101;
assign LUT_3[24214] = 32'b00000000000000011001100011110100;
assign LUT_3[24215] = 32'b00000000000000100000001111010001;
assign LUT_3[24216] = 32'b00000000000000011111100111100000;
assign LUT_3[24217] = 32'b00000000000000100110010010111101;
assign LUT_3[24218] = 32'b00000000000000100001101111000100;
assign LUT_3[24219] = 32'b00000000000000101000011010100001;
assign LUT_3[24220] = 32'b00000000000000011100110101010110;
assign LUT_3[24221] = 32'b00000000000000100011100000110011;
assign LUT_3[24222] = 32'b00000000000000011110111100111010;
assign LUT_3[24223] = 32'b00000000000000100101101000010111;
assign LUT_3[24224] = 32'b00000000000000011000001001110111;
assign LUT_3[24225] = 32'b00000000000000011110110101010100;
assign LUT_3[24226] = 32'b00000000000000011010010001011011;
assign LUT_3[24227] = 32'b00000000000000100000111100111000;
assign LUT_3[24228] = 32'b00000000000000010101010111101101;
assign LUT_3[24229] = 32'b00000000000000011100000011001010;
assign LUT_3[24230] = 32'b00000000000000010111011111010001;
assign LUT_3[24231] = 32'b00000000000000011110001010101110;
assign LUT_3[24232] = 32'b00000000000000011101100010111101;
assign LUT_3[24233] = 32'b00000000000000100100001110011010;
assign LUT_3[24234] = 32'b00000000000000011111101010100001;
assign LUT_3[24235] = 32'b00000000000000100110010101111110;
assign LUT_3[24236] = 32'b00000000000000011010110000110011;
assign LUT_3[24237] = 32'b00000000000000100001011100010000;
assign LUT_3[24238] = 32'b00000000000000011100111000010111;
assign LUT_3[24239] = 32'b00000000000000100011100011110100;
assign LUT_3[24240] = 32'b00000000000000011011011100111010;
assign LUT_3[24241] = 32'b00000000000000100010001000010111;
assign LUT_3[24242] = 32'b00000000000000011101100100011110;
assign LUT_3[24243] = 32'b00000000000000100100001111111011;
assign LUT_3[24244] = 32'b00000000000000011000101010110000;
assign LUT_3[24245] = 32'b00000000000000011111010110001101;
assign LUT_3[24246] = 32'b00000000000000011010110010010100;
assign LUT_3[24247] = 32'b00000000000000100001011101110001;
assign LUT_3[24248] = 32'b00000000000000100000110110000000;
assign LUT_3[24249] = 32'b00000000000000100111100001011101;
assign LUT_3[24250] = 32'b00000000000000100010111101100100;
assign LUT_3[24251] = 32'b00000000000000101001101001000001;
assign LUT_3[24252] = 32'b00000000000000011110000011110110;
assign LUT_3[24253] = 32'b00000000000000100100101111010011;
assign LUT_3[24254] = 32'b00000000000000100000001011011010;
assign LUT_3[24255] = 32'b00000000000000100110110110110111;
assign LUT_3[24256] = 32'b00000000000000010110110100000010;
assign LUT_3[24257] = 32'b00000000000000011101011111011111;
assign LUT_3[24258] = 32'b00000000000000011000111011100110;
assign LUT_3[24259] = 32'b00000000000000011111100111000011;
assign LUT_3[24260] = 32'b00000000000000010100000001111000;
assign LUT_3[24261] = 32'b00000000000000011010101101010101;
assign LUT_3[24262] = 32'b00000000000000010110001001011100;
assign LUT_3[24263] = 32'b00000000000000011100110100111001;
assign LUT_3[24264] = 32'b00000000000000011100001101001000;
assign LUT_3[24265] = 32'b00000000000000100010111000100101;
assign LUT_3[24266] = 32'b00000000000000011110010100101100;
assign LUT_3[24267] = 32'b00000000000000100101000000001001;
assign LUT_3[24268] = 32'b00000000000000011001011010111110;
assign LUT_3[24269] = 32'b00000000000000100000000110011011;
assign LUT_3[24270] = 32'b00000000000000011011100010100010;
assign LUT_3[24271] = 32'b00000000000000100010001101111111;
assign LUT_3[24272] = 32'b00000000000000011010000111000101;
assign LUT_3[24273] = 32'b00000000000000100000110010100010;
assign LUT_3[24274] = 32'b00000000000000011100001110101001;
assign LUT_3[24275] = 32'b00000000000000100010111010000110;
assign LUT_3[24276] = 32'b00000000000000010111010100111011;
assign LUT_3[24277] = 32'b00000000000000011110000000011000;
assign LUT_3[24278] = 32'b00000000000000011001011100011111;
assign LUT_3[24279] = 32'b00000000000000100000000111111100;
assign LUT_3[24280] = 32'b00000000000000011111100000001011;
assign LUT_3[24281] = 32'b00000000000000100110001011101000;
assign LUT_3[24282] = 32'b00000000000000100001100111101111;
assign LUT_3[24283] = 32'b00000000000000101000010011001100;
assign LUT_3[24284] = 32'b00000000000000011100101110000001;
assign LUT_3[24285] = 32'b00000000000000100011011001011110;
assign LUT_3[24286] = 32'b00000000000000011110110101100101;
assign LUT_3[24287] = 32'b00000000000000100101100001000010;
assign LUT_3[24288] = 32'b00000000000000011000000010100010;
assign LUT_3[24289] = 32'b00000000000000011110101101111111;
assign LUT_3[24290] = 32'b00000000000000011010001010000110;
assign LUT_3[24291] = 32'b00000000000000100000110101100011;
assign LUT_3[24292] = 32'b00000000000000010101010000011000;
assign LUT_3[24293] = 32'b00000000000000011011111011110101;
assign LUT_3[24294] = 32'b00000000000000010111010111111100;
assign LUT_3[24295] = 32'b00000000000000011110000011011001;
assign LUT_3[24296] = 32'b00000000000000011101011011101000;
assign LUT_3[24297] = 32'b00000000000000100100000111000101;
assign LUT_3[24298] = 32'b00000000000000011111100011001100;
assign LUT_3[24299] = 32'b00000000000000100110001110101001;
assign LUT_3[24300] = 32'b00000000000000011010101001011110;
assign LUT_3[24301] = 32'b00000000000000100001010100111011;
assign LUT_3[24302] = 32'b00000000000000011100110001000010;
assign LUT_3[24303] = 32'b00000000000000100011011100011111;
assign LUT_3[24304] = 32'b00000000000000011011010101100101;
assign LUT_3[24305] = 32'b00000000000000100010000001000010;
assign LUT_3[24306] = 32'b00000000000000011101011101001001;
assign LUT_3[24307] = 32'b00000000000000100100001000100110;
assign LUT_3[24308] = 32'b00000000000000011000100011011011;
assign LUT_3[24309] = 32'b00000000000000011111001110111000;
assign LUT_3[24310] = 32'b00000000000000011010101010111111;
assign LUT_3[24311] = 32'b00000000000000100001010110011100;
assign LUT_3[24312] = 32'b00000000000000100000101110101011;
assign LUT_3[24313] = 32'b00000000000000100111011010001000;
assign LUT_3[24314] = 32'b00000000000000100010110110001111;
assign LUT_3[24315] = 32'b00000000000000101001100001101100;
assign LUT_3[24316] = 32'b00000000000000011101111100100001;
assign LUT_3[24317] = 32'b00000000000000100100100111111110;
assign LUT_3[24318] = 32'b00000000000000100000000100000101;
assign LUT_3[24319] = 32'b00000000000000100110101111100010;
assign LUT_3[24320] = 32'b00000000000000010000111111111010;
assign LUT_3[24321] = 32'b00000000000000010111101011010111;
assign LUT_3[24322] = 32'b00000000000000010011000111011110;
assign LUT_3[24323] = 32'b00000000000000011001110010111011;
assign LUT_3[24324] = 32'b00000000000000001110001101110000;
assign LUT_3[24325] = 32'b00000000000000010100111001001101;
assign LUT_3[24326] = 32'b00000000000000010000010101010100;
assign LUT_3[24327] = 32'b00000000000000010111000000110001;
assign LUT_3[24328] = 32'b00000000000000010110011001000000;
assign LUT_3[24329] = 32'b00000000000000011101000100011101;
assign LUT_3[24330] = 32'b00000000000000011000100000100100;
assign LUT_3[24331] = 32'b00000000000000011111001100000001;
assign LUT_3[24332] = 32'b00000000000000010011100110110110;
assign LUT_3[24333] = 32'b00000000000000011010010010010011;
assign LUT_3[24334] = 32'b00000000000000010101101110011010;
assign LUT_3[24335] = 32'b00000000000000011100011001110111;
assign LUT_3[24336] = 32'b00000000000000010100010010111101;
assign LUT_3[24337] = 32'b00000000000000011010111110011010;
assign LUT_3[24338] = 32'b00000000000000010110011010100001;
assign LUT_3[24339] = 32'b00000000000000011101000101111110;
assign LUT_3[24340] = 32'b00000000000000010001100000110011;
assign LUT_3[24341] = 32'b00000000000000011000001100010000;
assign LUT_3[24342] = 32'b00000000000000010011101000010111;
assign LUT_3[24343] = 32'b00000000000000011010010011110100;
assign LUT_3[24344] = 32'b00000000000000011001101100000011;
assign LUT_3[24345] = 32'b00000000000000100000010111100000;
assign LUT_3[24346] = 32'b00000000000000011011110011100111;
assign LUT_3[24347] = 32'b00000000000000100010011111000100;
assign LUT_3[24348] = 32'b00000000000000010110111001111001;
assign LUT_3[24349] = 32'b00000000000000011101100101010110;
assign LUT_3[24350] = 32'b00000000000000011001000001011101;
assign LUT_3[24351] = 32'b00000000000000011111101100111010;
assign LUT_3[24352] = 32'b00000000000000010010001110011010;
assign LUT_3[24353] = 32'b00000000000000011000111001110111;
assign LUT_3[24354] = 32'b00000000000000010100010101111110;
assign LUT_3[24355] = 32'b00000000000000011011000001011011;
assign LUT_3[24356] = 32'b00000000000000001111011100010000;
assign LUT_3[24357] = 32'b00000000000000010110000111101101;
assign LUT_3[24358] = 32'b00000000000000010001100011110100;
assign LUT_3[24359] = 32'b00000000000000011000001111010001;
assign LUT_3[24360] = 32'b00000000000000010111100111100000;
assign LUT_3[24361] = 32'b00000000000000011110010010111101;
assign LUT_3[24362] = 32'b00000000000000011001101111000100;
assign LUT_3[24363] = 32'b00000000000000100000011010100001;
assign LUT_3[24364] = 32'b00000000000000010100110101010110;
assign LUT_3[24365] = 32'b00000000000000011011100000110011;
assign LUT_3[24366] = 32'b00000000000000010110111100111010;
assign LUT_3[24367] = 32'b00000000000000011101101000010111;
assign LUT_3[24368] = 32'b00000000000000010101100001011101;
assign LUT_3[24369] = 32'b00000000000000011100001100111010;
assign LUT_3[24370] = 32'b00000000000000010111101001000001;
assign LUT_3[24371] = 32'b00000000000000011110010100011110;
assign LUT_3[24372] = 32'b00000000000000010010101111010011;
assign LUT_3[24373] = 32'b00000000000000011001011010110000;
assign LUT_3[24374] = 32'b00000000000000010100110110110111;
assign LUT_3[24375] = 32'b00000000000000011011100010010100;
assign LUT_3[24376] = 32'b00000000000000011010111010100011;
assign LUT_3[24377] = 32'b00000000000000100001100110000000;
assign LUT_3[24378] = 32'b00000000000000011101000010000111;
assign LUT_3[24379] = 32'b00000000000000100011101101100100;
assign LUT_3[24380] = 32'b00000000000000011000001000011001;
assign LUT_3[24381] = 32'b00000000000000011110110011110110;
assign LUT_3[24382] = 32'b00000000000000011010001111111101;
assign LUT_3[24383] = 32'b00000000000000100000111011011010;
assign LUT_3[24384] = 32'b00000000000000010000111000100101;
assign LUT_3[24385] = 32'b00000000000000010111100100000010;
assign LUT_3[24386] = 32'b00000000000000010011000000001001;
assign LUT_3[24387] = 32'b00000000000000011001101011100110;
assign LUT_3[24388] = 32'b00000000000000001110000110011011;
assign LUT_3[24389] = 32'b00000000000000010100110001111000;
assign LUT_3[24390] = 32'b00000000000000010000001101111111;
assign LUT_3[24391] = 32'b00000000000000010110111001011100;
assign LUT_3[24392] = 32'b00000000000000010110010001101011;
assign LUT_3[24393] = 32'b00000000000000011100111101001000;
assign LUT_3[24394] = 32'b00000000000000011000011001001111;
assign LUT_3[24395] = 32'b00000000000000011111000100101100;
assign LUT_3[24396] = 32'b00000000000000010011011111100001;
assign LUT_3[24397] = 32'b00000000000000011010001010111110;
assign LUT_3[24398] = 32'b00000000000000010101100111000101;
assign LUT_3[24399] = 32'b00000000000000011100010010100010;
assign LUT_3[24400] = 32'b00000000000000010100001011101000;
assign LUT_3[24401] = 32'b00000000000000011010110111000101;
assign LUT_3[24402] = 32'b00000000000000010110010011001100;
assign LUT_3[24403] = 32'b00000000000000011100111110101001;
assign LUT_3[24404] = 32'b00000000000000010001011001011110;
assign LUT_3[24405] = 32'b00000000000000011000000100111011;
assign LUT_3[24406] = 32'b00000000000000010011100001000010;
assign LUT_3[24407] = 32'b00000000000000011010001100011111;
assign LUT_3[24408] = 32'b00000000000000011001100100101110;
assign LUT_3[24409] = 32'b00000000000000100000010000001011;
assign LUT_3[24410] = 32'b00000000000000011011101100010010;
assign LUT_3[24411] = 32'b00000000000000100010010111101111;
assign LUT_3[24412] = 32'b00000000000000010110110010100100;
assign LUT_3[24413] = 32'b00000000000000011101011110000001;
assign LUT_3[24414] = 32'b00000000000000011000111010001000;
assign LUT_3[24415] = 32'b00000000000000011111100101100101;
assign LUT_3[24416] = 32'b00000000000000010010000111000101;
assign LUT_3[24417] = 32'b00000000000000011000110010100010;
assign LUT_3[24418] = 32'b00000000000000010100001110101001;
assign LUT_3[24419] = 32'b00000000000000011010111010000110;
assign LUT_3[24420] = 32'b00000000000000001111010100111011;
assign LUT_3[24421] = 32'b00000000000000010110000000011000;
assign LUT_3[24422] = 32'b00000000000000010001011100011111;
assign LUT_3[24423] = 32'b00000000000000011000000111111100;
assign LUT_3[24424] = 32'b00000000000000010111100000001011;
assign LUT_3[24425] = 32'b00000000000000011110001011101000;
assign LUT_3[24426] = 32'b00000000000000011001100111101111;
assign LUT_3[24427] = 32'b00000000000000100000010011001100;
assign LUT_3[24428] = 32'b00000000000000010100101110000001;
assign LUT_3[24429] = 32'b00000000000000011011011001011110;
assign LUT_3[24430] = 32'b00000000000000010110110101100101;
assign LUT_3[24431] = 32'b00000000000000011101100001000010;
assign LUT_3[24432] = 32'b00000000000000010101011010001000;
assign LUT_3[24433] = 32'b00000000000000011100000101100101;
assign LUT_3[24434] = 32'b00000000000000010111100001101100;
assign LUT_3[24435] = 32'b00000000000000011110001101001001;
assign LUT_3[24436] = 32'b00000000000000010010100111111110;
assign LUT_3[24437] = 32'b00000000000000011001010011011011;
assign LUT_3[24438] = 32'b00000000000000010100101111100010;
assign LUT_3[24439] = 32'b00000000000000011011011010111111;
assign LUT_3[24440] = 32'b00000000000000011010110011001110;
assign LUT_3[24441] = 32'b00000000000000100001011110101011;
assign LUT_3[24442] = 32'b00000000000000011100111010110010;
assign LUT_3[24443] = 32'b00000000000000100011100110001111;
assign LUT_3[24444] = 32'b00000000000000011000000001000100;
assign LUT_3[24445] = 32'b00000000000000011110101100100001;
assign LUT_3[24446] = 32'b00000000000000011010001000101000;
assign LUT_3[24447] = 32'b00000000000000100000110100000101;
assign LUT_3[24448] = 32'b00000000000000010011001010111000;
assign LUT_3[24449] = 32'b00000000000000011001110110010101;
assign LUT_3[24450] = 32'b00000000000000010101010010011100;
assign LUT_3[24451] = 32'b00000000000000011011111101111001;
assign LUT_3[24452] = 32'b00000000000000010000011000101110;
assign LUT_3[24453] = 32'b00000000000000010111000100001011;
assign LUT_3[24454] = 32'b00000000000000010010100000010010;
assign LUT_3[24455] = 32'b00000000000000011001001011101111;
assign LUT_3[24456] = 32'b00000000000000011000100011111110;
assign LUT_3[24457] = 32'b00000000000000011111001111011011;
assign LUT_3[24458] = 32'b00000000000000011010101011100010;
assign LUT_3[24459] = 32'b00000000000000100001010110111111;
assign LUT_3[24460] = 32'b00000000000000010101110001110100;
assign LUT_3[24461] = 32'b00000000000000011100011101010001;
assign LUT_3[24462] = 32'b00000000000000010111111001011000;
assign LUT_3[24463] = 32'b00000000000000011110100100110101;
assign LUT_3[24464] = 32'b00000000000000010110011101111011;
assign LUT_3[24465] = 32'b00000000000000011101001001011000;
assign LUT_3[24466] = 32'b00000000000000011000100101011111;
assign LUT_3[24467] = 32'b00000000000000011111010000111100;
assign LUT_3[24468] = 32'b00000000000000010011101011110001;
assign LUT_3[24469] = 32'b00000000000000011010010111001110;
assign LUT_3[24470] = 32'b00000000000000010101110011010101;
assign LUT_3[24471] = 32'b00000000000000011100011110110010;
assign LUT_3[24472] = 32'b00000000000000011011110111000001;
assign LUT_3[24473] = 32'b00000000000000100010100010011110;
assign LUT_3[24474] = 32'b00000000000000011101111110100101;
assign LUT_3[24475] = 32'b00000000000000100100101010000010;
assign LUT_3[24476] = 32'b00000000000000011001000100110111;
assign LUT_3[24477] = 32'b00000000000000011111110000010100;
assign LUT_3[24478] = 32'b00000000000000011011001100011011;
assign LUT_3[24479] = 32'b00000000000000100001110111111000;
assign LUT_3[24480] = 32'b00000000000000010100011001011000;
assign LUT_3[24481] = 32'b00000000000000011011000100110101;
assign LUT_3[24482] = 32'b00000000000000010110100000111100;
assign LUT_3[24483] = 32'b00000000000000011101001100011001;
assign LUT_3[24484] = 32'b00000000000000010001100111001110;
assign LUT_3[24485] = 32'b00000000000000011000010010101011;
assign LUT_3[24486] = 32'b00000000000000010011101110110010;
assign LUT_3[24487] = 32'b00000000000000011010011010001111;
assign LUT_3[24488] = 32'b00000000000000011001110010011110;
assign LUT_3[24489] = 32'b00000000000000100000011101111011;
assign LUT_3[24490] = 32'b00000000000000011011111010000010;
assign LUT_3[24491] = 32'b00000000000000100010100101011111;
assign LUT_3[24492] = 32'b00000000000000010111000000010100;
assign LUT_3[24493] = 32'b00000000000000011101101011110001;
assign LUT_3[24494] = 32'b00000000000000011001000111111000;
assign LUT_3[24495] = 32'b00000000000000011111110011010101;
assign LUT_3[24496] = 32'b00000000000000010111101100011011;
assign LUT_3[24497] = 32'b00000000000000011110010111111000;
assign LUT_3[24498] = 32'b00000000000000011001110011111111;
assign LUT_3[24499] = 32'b00000000000000100000011111011100;
assign LUT_3[24500] = 32'b00000000000000010100111010010001;
assign LUT_3[24501] = 32'b00000000000000011011100101101110;
assign LUT_3[24502] = 32'b00000000000000010111000001110101;
assign LUT_3[24503] = 32'b00000000000000011101101101010010;
assign LUT_3[24504] = 32'b00000000000000011101000101100001;
assign LUT_3[24505] = 32'b00000000000000100011110000111110;
assign LUT_3[24506] = 32'b00000000000000011111001101000101;
assign LUT_3[24507] = 32'b00000000000000100101111000100010;
assign LUT_3[24508] = 32'b00000000000000011010010011010111;
assign LUT_3[24509] = 32'b00000000000000100000111110110100;
assign LUT_3[24510] = 32'b00000000000000011100011010111011;
assign LUT_3[24511] = 32'b00000000000000100011000110011000;
assign LUT_3[24512] = 32'b00000000000000010011000011100011;
assign LUT_3[24513] = 32'b00000000000000011001101111000000;
assign LUT_3[24514] = 32'b00000000000000010101001011000111;
assign LUT_3[24515] = 32'b00000000000000011011110110100100;
assign LUT_3[24516] = 32'b00000000000000010000010001011001;
assign LUT_3[24517] = 32'b00000000000000010110111100110110;
assign LUT_3[24518] = 32'b00000000000000010010011000111101;
assign LUT_3[24519] = 32'b00000000000000011001000100011010;
assign LUT_3[24520] = 32'b00000000000000011000011100101001;
assign LUT_3[24521] = 32'b00000000000000011111001000000110;
assign LUT_3[24522] = 32'b00000000000000011010100100001101;
assign LUT_3[24523] = 32'b00000000000000100001001111101010;
assign LUT_3[24524] = 32'b00000000000000010101101010011111;
assign LUT_3[24525] = 32'b00000000000000011100010101111100;
assign LUT_3[24526] = 32'b00000000000000010111110010000011;
assign LUT_3[24527] = 32'b00000000000000011110011101100000;
assign LUT_3[24528] = 32'b00000000000000010110010110100110;
assign LUT_3[24529] = 32'b00000000000000011101000010000011;
assign LUT_3[24530] = 32'b00000000000000011000011110001010;
assign LUT_3[24531] = 32'b00000000000000011111001001100111;
assign LUT_3[24532] = 32'b00000000000000010011100100011100;
assign LUT_3[24533] = 32'b00000000000000011010001111111001;
assign LUT_3[24534] = 32'b00000000000000010101101100000000;
assign LUT_3[24535] = 32'b00000000000000011100010111011101;
assign LUT_3[24536] = 32'b00000000000000011011101111101100;
assign LUT_3[24537] = 32'b00000000000000100010011011001001;
assign LUT_3[24538] = 32'b00000000000000011101110111010000;
assign LUT_3[24539] = 32'b00000000000000100100100010101101;
assign LUT_3[24540] = 32'b00000000000000011000111101100010;
assign LUT_3[24541] = 32'b00000000000000011111101000111111;
assign LUT_3[24542] = 32'b00000000000000011011000101000110;
assign LUT_3[24543] = 32'b00000000000000100001110000100011;
assign LUT_3[24544] = 32'b00000000000000010100010010000011;
assign LUT_3[24545] = 32'b00000000000000011010111101100000;
assign LUT_3[24546] = 32'b00000000000000010110011001100111;
assign LUT_3[24547] = 32'b00000000000000011101000101000100;
assign LUT_3[24548] = 32'b00000000000000010001011111111001;
assign LUT_3[24549] = 32'b00000000000000011000001011010110;
assign LUT_3[24550] = 32'b00000000000000010011100111011101;
assign LUT_3[24551] = 32'b00000000000000011010010010111010;
assign LUT_3[24552] = 32'b00000000000000011001101011001001;
assign LUT_3[24553] = 32'b00000000000000100000010110100110;
assign LUT_3[24554] = 32'b00000000000000011011110010101101;
assign LUT_3[24555] = 32'b00000000000000100010011110001010;
assign LUT_3[24556] = 32'b00000000000000010110111000111111;
assign LUT_3[24557] = 32'b00000000000000011101100100011100;
assign LUT_3[24558] = 32'b00000000000000011001000000100011;
assign LUT_3[24559] = 32'b00000000000000011111101100000000;
assign LUT_3[24560] = 32'b00000000000000010111100101000110;
assign LUT_3[24561] = 32'b00000000000000011110010000100011;
assign LUT_3[24562] = 32'b00000000000000011001101100101010;
assign LUT_3[24563] = 32'b00000000000000100000011000000111;
assign LUT_3[24564] = 32'b00000000000000010100110010111100;
assign LUT_3[24565] = 32'b00000000000000011011011110011001;
assign LUT_3[24566] = 32'b00000000000000010110111010100000;
assign LUT_3[24567] = 32'b00000000000000011101100101111101;
assign LUT_3[24568] = 32'b00000000000000011100111110001100;
assign LUT_3[24569] = 32'b00000000000000100011101001101001;
assign LUT_3[24570] = 32'b00000000000000011111000101110000;
assign LUT_3[24571] = 32'b00000000000000100101110001001101;
assign LUT_3[24572] = 32'b00000000000000011010001100000010;
assign LUT_3[24573] = 32'b00000000000000100000110111011111;
assign LUT_3[24574] = 32'b00000000000000011100010011100110;
assign LUT_3[24575] = 32'b00000000000000100010111111000011;
assign LUT_3[24576] = 32'b00000000000000001011000100000010;
assign LUT_3[24577] = 32'b00000000000000010001101111011111;
assign LUT_3[24578] = 32'b00000000000000001101001011100110;
assign LUT_3[24579] = 32'b00000000000000010011110111000011;
assign LUT_3[24580] = 32'b00000000000000001000010001111000;
assign LUT_3[24581] = 32'b00000000000000001110111101010101;
assign LUT_3[24582] = 32'b00000000000000001010011001011100;
assign LUT_3[24583] = 32'b00000000000000010001000100111001;
assign LUT_3[24584] = 32'b00000000000000010000011101001000;
assign LUT_3[24585] = 32'b00000000000000010111001000100101;
assign LUT_3[24586] = 32'b00000000000000010010100100101100;
assign LUT_3[24587] = 32'b00000000000000011001010000001001;
assign LUT_3[24588] = 32'b00000000000000001101101010111110;
assign LUT_3[24589] = 32'b00000000000000010100010110011011;
assign LUT_3[24590] = 32'b00000000000000001111110010100010;
assign LUT_3[24591] = 32'b00000000000000010110011101111111;
assign LUT_3[24592] = 32'b00000000000000001110010111000101;
assign LUT_3[24593] = 32'b00000000000000010101000010100010;
assign LUT_3[24594] = 32'b00000000000000010000011110101001;
assign LUT_3[24595] = 32'b00000000000000010111001010000110;
assign LUT_3[24596] = 32'b00000000000000001011100100111011;
assign LUT_3[24597] = 32'b00000000000000010010010000011000;
assign LUT_3[24598] = 32'b00000000000000001101101100011111;
assign LUT_3[24599] = 32'b00000000000000010100010111111100;
assign LUT_3[24600] = 32'b00000000000000010011110000001011;
assign LUT_3[24601] = 32'b00000000000000011010011011101000;
assign LUT_3[24602] = 32'b00000000000000010101110111101111;
assign LUT_3[24603] = 32'b00000000000000011100100011001100;
assign LUT_3[24604] = 32'b00000000000000010000111110000001;
assign LUT_3[24605] = 32'b00000000000000010111101001011110;
assign LUT_3[24606] = 32'b00000000000000010011000101100101;
assign LUT_3[24607] = 32'b00000000000000011001110001000010;
assign LUT_3[24608] = 32'b00000000000000001100010010100010;
assign LUT_3[24609] = 32'b00000000000000010010111101111111;
assign LUT_3[24610] = 32'b00000000000000001110011010000110;
assign LUT_3[24611] = 32'b00000000000000010101000101100011;
assign LUT_3[24612] = 32'b00000000000000001001100000011000;
assign LUT_3[24613] = 32'b00000000000000010000001011110101;
assign LUT_3[24614] = 32'b00000000000000001011100111111100;
assign LUT_3[24615] = 32'b00000000000000010010010011011001;
assign LUT_3[24616] = 32'b00000000000000010001101011101000;
assign LUT_3[24617] = 32'b00000000000000011000010111000101;
assign LUT_3[24618] = 32'b00000000000000010011110011001100;
assign LUT_3[24619] = 32'b00000000000000011010011110101001;
assign LUT_3[24620] = 32'b00000000000000001110111001011110;
assign LUT_3[24621] = 32'b00000000000000010101100100111011;
assign LUT_3[24622] = 32'b00000000000000010001000001000010;
assign LUT_3[24623] = 32'b00000000000000010111101100011111;
assign LUT_3[24624] = 32'b00000000000000001111100101100101;
assign LUT_3[24625] = 32'b00000000000000010110010001000010;
assign LUT_3[24626] = 32'b00000000000000010001101101001001;
assign LUT_3[24627] = 32'b00000000000000011000011000100110;
assign LUT_3[24628] = 32'b00000000000000001100110011011011;
assign LUT_3[24629] = 32'b00000000000000010011011110111000;
assign LUT_3[24630] = 32'b00000000000000001110111010111111;
assign LUT_3[24631] = 32'b00000000000000010101100110011100;
assign LUT_3[24632] = 32'b00000000000000010100111110101011;
assign LUT_3[24633] = 32'b00000000000000011011101010001000;
assign LUT_3[24634] = 32'b00000000000000010111000110001111;
assign LUT_3[24635] = 32'b00000000000000011101110001101100;
assign LUT_3[24636] = 32'b00000000000000010010001100100001;
assign LUT_3[24637] = 32'b00000000000000011000110111111110;
assign LUT_3[24638] = 32'b00000000000000010100010100000101;
assign LUT_3[24639] = 32'b00000000000000011010111111100010;
assign LUT_3[24640] = 32'b00000000000000001010111100101101;
assign LUT_3[24641] = 32'b00000000000000010001101000001010;
assign LUT_3[24642] = 32'b00000000000000001101000100010001;
assign LUT_3[24643] = 32'b00000000000000010011101111101110;
assign LUT_3[24644] = 32'b00000000000000001000001010100011;
assign LUT_3[24645] = 32'b00000000000000001110110110000000;
assign LUT_3[24646] = 32'b00000000000000001010010010000111;
assign LUT_3[24647] = 32'b00000000000000010000111101100100;
assign LUT_3[24648] = 32'b00000000000000010000010101110011;
assign LUT_3[24649] = 32'b00000000000000010111000001010000;
assign LUT_3[24650] = 32'b00000000000000010010011101010111;
assign LUT_3[24651] = 32'b00000000000000011001001000110100;
assign LUT_3[24652] = 32'b00000000000000001101100011101001;
assign LUT_3[24653] = 32'b00000000000000010100001111000110;
assign LUT_3[24654] = 32'b00000000000000001111101011001101;
assign LUT_3[24655] = 32'b00000000000000010110010110101010;
assign LUT_3[24656] = 32'b00000000000000001110001111110000;
assign LUT_3[24657] = 32'b00000000000000010100111011001101;
assign LUT_3[24658] = 32'b00000000000000010000010111010100;
assign LUT_3[24659] = 32'b00000000000000010111000010110001;
assign LUT_3[24660] = 32'b00000000000000001011011101100110;
assign LUT_3[24661] = 32'b00000000000000010010001001000011;
assign LUT_3[24662] = 32'b00000000000000001101100101001010;
assign LUT_3[24663] = 32'b00000000000000010100010000100111;
assign LUT_3[24664] = 32'b00000000000000010011101000110110;
assign LUT_3[24665] = 32'b00000000000000011010010100010011;
assign LUT_3[24666] = 32'b00000000000000010101110000011010;
assign LUT_3[24667] = 32'b00000000000000011100011011110111;
assign LUT_3[24668] = 32'b00000000000000010000110110101100;
assign LUT_3[24669] = 32'b00000000000000010111100010001001;
assign LUT_3[24670] = 32'b00000000000000010010111110010000;
assign LUT_3[24671] = 32'b00000000000000011001101001101101;
assign LUT_3[24672] = 32'b00000000000000001100001011001101;
assign LUT_3[24673] = 32'b00000000000000010010110110101010;
assign LUT_3[24674] = 32'b00000000000000001110010010110001;
assign LUT_3[24675] = 32'b00000000000000010100111110001110;
assign LUT_3[24676] = 32'b00000000000000001001011001000011;
assign LUT_3[24677] = 32'b00000000000000010000000100100000;
assign LUT_3[24678] = 32'b00000000000000001011100000100111;
assign LUT_3[24679] = 32'b00000000000000010010001100000100;
assign LUT_3[24680] = 32'b00000000000000010001100100010011;
assign LUT_3[24681] = 32'b00000000000000011000001111110000;
assign LUT_3[24682] = 32'b00000000000000010011101011110111;
assign LUT_3[24683] = 32'b00000000000000011010010111010100;
assign LUT_3[24684] = 32'b00000000000000001110110010001001;
assign LUT_3[24685] = 32'b00000000000000010101011101100110;
assign LUT_3[24686] = 32'b00000000000000010000111001101101;
assign LUT_3[24687] = 32'b00000000000000010111100101001010;
assign LUT_3[24688] = 32'b00000000000000001111011110010000;
assign LUT_3[24689] = 32'b00000000000000010110001001101101;
assign LUT_3[24690] = 32'b00000000000000010001100101110100;
assign LUT_3[24691] = 32'b00000000000000011000010001010001;
assign LUT_3[24692] = 32'b00000000000000001100101100000110;
assign LUT_3[24693] = 32'b00000000000000010011010111100011;
assign LUT_3[24694] = 32'b00000000000000001110110011101010;
assign LUT_3[24695] = 32'b00000000000000010101011111000111;
assign LUT_3[24696] = 32'b00000000000000010100110111010110;
assign LUT_3[24697] = 32'b00000000000000011011100010110011;
assign LUT_3[24698] = 32'b00000000000000010110111110111010;
assign LUT_3[24699] = 32'b00000000000000011101101010010111;
assign LUT_3[24700] = 32'b00000000000000010010000101001100;
assign LUT_3[24701] = 32'b00000000000000011000110000101001;
assign LUT_3[24702] = 32'b00000000000000010100001100110000;
assign LUT_3[24703] = 32'b00000000000000011010111000001101;
assign LUT_3[24704] = 32'b00000000000000001101001111000000;
assign LUT_3[24705] = 32'b00000000000000010011111010011101;
assign LUT_3[24706] = 32'b00000000000000001111010110100100;
assign LUT_3[24707] = 32'b00000000000000010110000010000001;
assign LUT_3[24708] = 32'b00000000000000001010011100110110;
assign LUT_3[24709] = 32'b00000000000000010001001000010011;
assign LUT_3[24710] = 32'b00000000000000001100100100011010;
assign LUT_3[24711] = 32'b00000000000000010011001111110111;
assign LUT_3[24712] = 32'b00000000000000010010101000000110;
assign LUT_3[24713] = 32'b00000000000000011001010011100011;
assign LUT_3[24714] = 32'b00000000000000010100101111101010;
assign LUT_3[24715] = 32'b00000000000000011011011011000111;
assign LUT_3[24716] = 32'b00000000000000001111110101111100;
assign LUT_3[24717] = 32'b00000000000000010110100001011001;
assign LUT_3[24718] = 32'b00000000000000010001111101100000;
assign LUT_3[24719] = 32'b00000000000000011000101000111101;
assign LUT_3[24720] = 32'b00000000000000010000100010000011;
assign LUT_3[24721] = 32'b00000000000000010111001101100000;
assign LUT_3[24722] = 32'b00000000000000010010101001100111;
assign LUT_3[24723] = 32'b00000000000000011001010101000100;
assign LUT_3[24724] = 32'b00000000000000001101101111111001;
assign LUT_3[24725] = 32'b00000000000000010100011011010110;
assign LUT_3[24726] = 32'b00000000000000001111110111011101;
assign LUT_3[24727] = 32'b00000000000000010110100010111010;
assign LUT_3[24728] = 32'b00000000000000010101111011001001;
assign LUT_3[24729] = 32'b00000000000000011100100110100110;
assign LUT_3[24730] = 32'b00000000000000011000000010101101;
assign LUT_3[24731] = 32'b00000000000000011110101110001010;
assign LUT_3[24732] = 32'b00000000000000010011001000111111;
assign LUT_3[24733] = 32'b00000000000000011001110100011100;
assign LUT_3[24734] = 32'b00000000000000010101010000100011;
assign LUT_3[24735] = 32'b00000000000000011011111100000000;
assign LUT_3[24736] = 32'b00000000000000001110011101100000;
assign LUT_3[24737] = 32'b00000000000000010101001000111101;
assign LUT_3[24738] = 32'b00000000000000010000100101000100;
assign LUT_3[24739] = 32'b00000000000000010111010000100001;
assign LUT_3[24740] = 32'b00000000000000001011101011010110;
assign LUT_3[24741] = 32'b00000000000000010010010110110011;
assign LUT_3[24742] = 32'b00000000000000001101110010111010;
assign LUT_3[24743] = 32'b00000000000000010100011110010111;
assign LUT_3[24744] = 32'b00000000000000010011110110100110;
assign LUT_3[24745] = 32'b00000000000000011010100010000011;
assign LUT_3[24746] = 32'b00000000000000010101111110001010;
assign LUT_3[24747] = 32'b00000000000000011100101001100111;
assign LUT_3[24748] = 32'b00000000000000010001000100011100;
assign LUT_3[24749] = 32'b00000000000000010111101111111001;
assign LUT_3[24750] = 32'b00000000000000010011001100000000;
assign LUT_3[24751] = 32'b00000000000000011001110111011101;
assign LUT_3[24752] = 32'b00000000000000010001110000100011;
assign LUT_3[24753] = 32'b00000000000000011000011100000000;
assign LUT_3[24754] = 32'b00000000000000010011111000000111;
assign LUT_3[24755] = 32'b00000000000000011010100011100100;
assign LUT_3[24756] = 32'b00000000000000001110111110011001;
assign LUT_3[24757] = 32'b00000000000000010101101001110110;
assign LUT_3[24758] = 32'b00000000000000010001000101111101;
assign LUT_3[24759] = 32'b00000000000000010111110001011010;
assign LUT_3[24760] = 32'b00000000000000010111001001101001;
assign LUT_3[24761] = 32'b00000000000000011101110101000110;
assign LUT_3[24762] = 32'b00000000000000011001010001001101;
assign LUT_3[24763] = 32'b00000000000000011111111100101010;
assign LUT_3[24764] = 32'b00000000000000010100010111011111;
assign LUT_3[24765] = 32'b00000000000000011011000010111100;
assign LUT_3[24766] = 32'b00000000000000010110011111000011;
assign LUT_3[24767] = 32'b00000000000000011101001010100000;
assign LUT_3[24768] = 32'b00000000000000001101000111101011;
assign LUT_3[24769] = 32'b00000000000000010011110011001000;
assign LUT_3[24770] = 32'b00000000000000001111001111001111;
assign LUT_3[24771] = 32'b00000000000000010101111010101100;
assign LUT_3[24772] = 32'b00000000000000001010010101100001;
assign LUT_3[24773] = 32'b00000000000000010001000000111110;
assign LUT_3[24774] = 32'b00000000000000001100011101000101;
assign LUT_3[24775] = 32'b00000000000000010011001000100010;
assign LUT_3[24776] = 32'b00000000000000010010100000110001;
assign LUT_3[24777] = 32'b00000000000000011001001100001110;
assign LUT_3[24778] = 32'b00000000000000010100101000010101;
assign LUT_3[24779] = 32'b00000000000000011011010011110010;
assign LUT_3[24780] = 32'b00000000000000001111101110100111;
assign LUT_3[24781] = 32'b00000000000000010110011010000100;
assign LUT_3[24782] = 32'b00000000000000010001110110001011;
assign LUT_3[24783] = 32'b00000000000000011000100001101000;
assign LUT_3[24784] = 32'b00000000000000010000011010101110;
assign LUT_3[24785] = 32'b00000000000000010111000110001011;
assign LUT_3[24786] = 32'b00000000000000010010100010010010;
assign LUT_3[24787] = 32'b00000000000000011001001101101111;
assign LUT_3[24788] = 32'b00000000000000001101101000100100;
assign LUT_3[24789] = 32'b00000000000000010100010100000001;
assign LUT_3[24790] = 32'b00000000000000001111110000001000;
assign LUT_3[24791] = 32'b00000000000000010110011011100101;
assign LUT_3[24792] = 32'b00000000000000010101110011110100;
assign LUT_3[24793] = 32'b00000000000000011100011111010001;
assign LUT_3[24794] = 32'b00000000000000010111111011011000;
assign LUT_3[24795] = 32'b00000000000000011110100110110101;
assign LUT_3[24796] = 32'b00000000000000010011000001101010;
assign LUT_3[24797] = 32'b00000000000000011001101101000111;
assign LUT_3[24798] = 32'b00000000000000010101001001001110;
assign LUT_3[24799] = 32'b00000000000000011011110100101011;
assign LUT_3[24800] = 32'b00000000000000001110010110001011;
assign LUT_3[24801] = 32'b00000000000000010101000001101000;
assign LUT_3[24802] = 32'b00000000000000010000011101101111;
assign LUT_3[24803] = 32'b00000000000000010111001001001100;
assign LUT_3[24804] = 32'b00000000000000001011100100000001;
assign LUT_3[24805] = 32'b00000000000000010010001111011110;
assign LUT_3[24806] = 32'b00000000000000001101101011100101;
assign LUT_3[24807] = 32'b00000000000000010100010111000010;
assign LUT_3[24808] = 32'b00000000000000010011101111010001;
assign LUT_3[24809] = 32'b00000000000000011010011010101110;
assign LUT_3[24810] = 32'b00000000000000010101110110110101;
assign LUT_3[24811] = 32'b00000000000000011100100010010010;
assign LUT_3[24812] = 32'b00000000000000010000111101000111;
assign LUT_3[24813] = 32'b00000000000000010111101000100100;
assign LUT_3[24814] = 32'b00000000000000010011000100101011;
assign LUT_3[24815] = 32'b00000000000000011001110000001000;
assign LUT_3[24816] = 32'b00000000000000010001101001001110;
assign LUT_3[24817] = 32'b00000000000000011000010100101011;
assign LUT_3[24818] = 32'b00000000000000010011110000110010;
assign LUT_3[24819] = 32'b00000000000000011010011100001111;
assign LUT_3[24820] = 32'b00000000000000001110110111000100;
assign LUT_3[24821] = 32'b00000000000000010101100010100001;
assign LUT_3[24822] = 32'b00000000000000010000111110101000;
assign LUT_3[24823] = 32'b00000000000000010111101010000101;
assign LUT_3[24824] = 32'b00000000000000010111000010010100;
assign LUT_3[24825] = 32'b00000000000000011101101101110001;
assign LUT_3[24826] = 32'b00000000000000011001001001111000;
assign LUT_3[24827] = 32'b00000000000000011111110101010101;
assign LUT_3[24828] = 32'b00000000000000010100010000001010;
assign LUT_3[24829] = 32'b00000000000000011010111011100111;
assign LUT_3[24830] = 32'b00000000000000010110010111101110;
assign LUT_3[24831] = 32'b00000000000000011101000011001011;
assign LUT_3[24832] = 32'b00000000000000000111010011100011;
assign LUT_3[24833] = 32'b00000000000000001101111111000000;
assign LUT_3[24834] = 32'b00000000000000001001011011000111;
assign LUT_3[24835] = 32'b00000000000000010000000110100100;
assign LUT_3[24836] = 32'b00000000000000000100100001011001;
assign LUT_3[24837] = 32'b00000000000000001011001100110110;
assign LUT_3[24838] = 32'b00000000000000000110101000111101;
assign LUT_3[24839] = 32'b00000000000000001101010100011010;
assign LUT_3[24840] = 32'b00000000000000001100101100101001;
assign LUT_3[24841] = 32'b00000000000000010011011000000110;
assign LUT_3[24842] = 32'b00000000000000001110110100001101;
assign LUT_3[24843] = 32'b00000000000000010101011111101010;
assign LUT_3[24844] = 32'b00000000000000001001111010011111;
assign LUT_3[24845] = 32'b00000000000000010000100101111100;
assign LUT_3[24846] = 32'b00000000000000001100000010000011;
assign LUT_3[24847] = 32'b00000000000000010010101101100000;
assign LUT_3[24848] = 32'b00000000000000001010100110100110;
assign LUT_3[24849] = 32'b00000000000000010001010010000011;
assign LUT_3[24850] = 32'b00000000000000001100101110001010;
assign LUT_3[24851] = 32'b00000000000000010011011001100111;
assign LUT_3[24852] = 32'b00000000000000000111110100011100;
assign LUT_3[24853] = 32'b00000000000000001110011111111001;
assign LUT_3[24854] = 32'b00000000000000001001111100000000;
assign LUT_3[24855] = 32'b00000000000000010000100111011101;
assign LUT_3[24856] = 32'b00000000000000001111111111101100;
assign LUT_3[24857] = 32'b00000000000000010110101011001001;
assign LUT_3[24858] = 32'b00000000000000010010000111010000;
assign LUT_3[24859] = 32'b00000000000000011000110010101101;
assign LUT_3[24860] = 32'b00000000000000001101001101100010;
assign LUT_3[24861] = 32'b00000000000000010011111000111111;
assign LUT_3[24862] = 32'b00000000000000001111010101000110;
assign LUT_3[24863] = 32'b00000000000000010110000000100011;
assign LUT_3[24864] = 32'b00000000000000001000100010000011;
assign LUT_3[24865] = 32'b00000000000000001111001101100000;
assign LUT_3[24866] = 32'b00000000000000001010101001100111;
assign LUT_3[24867] = 32'b00000000000000010001010101000100;
assign LUT_3[24868] = 32'b00000000000000000101101111111001;
assign LUT_3[24869] = 32'b00000000000000001100011011010110;
assign LUT_3[24870] = 32'b00000000000000000111110111011101;
assign LUT_3[24871] = 32'b00000000000000001110100010111010;
assign LUT_3[24872] = 32'b00000000000000001101111011001001;
assign LUT_3[24873] = 32'b00000000000000010100100110100110;
assign LUT_3[24874] = 32'b00000000000000010000000010101101;
assign LUT_3[24875] = 32'b00000000000000010110101110001010;
assign LUT_3[24876] = 32'b00000000000000001011001000111111;
assign LUT_3[24877] = 32'b00000000000000010001110100011100;
assign LUT_3[24878] = 32'b00000000000000001101010000100011;
assign LUT_3[24879] = 32'b00000000000000010011111100000000;
assign LUT_3[24880] = 32'b00000000000000001011110101000110;
assign LUT_3[24881] = 32'b00000000000000010010100000100011;
assign LUT_3[24882] = 32'b00000000000000001101111100101010;
assign LUT_3[24883] = 32'b00000000000000010100101000000111;
assign LUT_3[24884] = 32'b00000000000000001001000010111100;
assign LUT_3[24885] = 32'b00000000000000001111101110011001;
assign LUT_3[24886] = 32'b00000000000000001011001010100000;
assign LUT_3[24887] = 32'b00000000000000010001110101111101;
assign LUT_3[24888] = 32'b00000000000000010001001110001100;
assign LUT_3[24889] = 32'b00000000000000010111111001101001;
assign LUT_3[24890] = 32'b00000000000000010011010101110000;
assign LUT_3[24891] = 32'b00000000000000011010000001001101;
assign LUT_3[24892] = 32'b00000000000000001110011100000010;
assign LUT_3[24893] = 32'b00000000000000010101000111011111;
assign LUT_3[24894] = 32'b00000000000000010000100011100110;
assign LUT_3[24895] = 32'b00000000000000010111001111000011;
assign LUT_3[24896] = 32'b00000000000000000111001100001110;
assign LUT_3[24897] = 32'b00000000000000001101110111101011;
assign LUT_3[24898] = 32'b00000000000000001001010011110010;
assign LUT_3[24899] = 32'b00000000000000001111111111001111;
assign LUT_3[24900] = 32'b00000000000000000100011010000100;
assign LUT_3[24901] = 32'b00000000000000001011000101100001;
assign LUT_3[24902] = 32'b00000000000000000110100001101000;
assign LUT_3[24903] = 32'b00000000000000001101001101000101;
assign LUT_3[24904] = 32'b00000000000000001100100101010100;
assign LUT_3[24905] = 32'b00000000000000010011010000110001;
assign LUT_3[24906] = 32'b00000000000000001110101100111000;
assign LUT_3[24907] = 32'b00000000000000010101011000010101;
assign LUT_3[24908] = 32'b00000000000000001001110011001010;
assign LUT_3[24909] = 32'b00000000000000010000011110100111;
assign LUT_3[24910] = 32'b00000000000000001011111010101110;
assign LUT_3[24911] = 32'b00000000000000010010100110001011;
assign LUT_3[24912] = 32'b00000000000000001010011111010001;
assign LUT_3[24913] = 32'b00000000000000010001001010101110;
assign LUT_3[24914] = 32'b00000000000000001100100110110101;
assign LUT_3[24915] = 32'b00000000000000010011010010010010;
assign LUT_3[24916] = 32'b00000000000000000111101101000111;
assign LUT_3[24917] = 32'b00000000000000001110011000100100;
assign LUT_3[24918] = 32'b00000000000000001001110100101011;
assign LUT_3[24919] = 32'b00000000000000010000100000001000;
assign LUT_3[24920] = 32'b00000000000000001111111000010111;
assign LUT_3[24921] = 32'b00000000000000010110100011110100;
assign LUT_3[24922] = 32'b00000000000000010001111111111011;
assign LUT_3[24923] = 32'b00000000000000011000101011011000;
assign LUT_3[24924] = 32'b00000000000000001101000110001101;
assign LUT_3[24925] = 32'b00000000000000010011110001101010;
assign LUT_3[24926] = 32'b00000000000000001111001101110001;
assign LUT_3[24927] = 32'b00000000000000010101111001001110;
assign LUT_3[24928] = 32'b00000000000000001000011010101110;
assign LUT_3[24929] = 32'b00000000000000001111000110001011;
assign LUT_3[24930] = 32'b00000000000000001010100010010010;
assign LUT_3[24931] = 32'b00000000000000010001001101101111;
assign LUT_3[24932] = 32'b00000000000000000101101000100100;
assign LUT_3[24933] = 32'b00000000000000001100010100000001;
assign LUT_3[24934] = 32'b00000000000000000111110000001000;
assign LUT_3[24935] = 32'b00000000000000001110011011100101;
assign LUT_3[24936] = 32'b00000000000000001101110011110100;
assign LUT_3[24937] = 32'b00000000000000010100011111010001;
assign LUT_3[24938] = 32'b00000000000000001111111011011000;
assign LUT_3[24939] = 32'b00000000000000010110100110110101;
assign LUT_3[24940] = 32'b00000000000000001011000001101010;
assign LUT_3[24941] = 32'b00000000000000010001101101000111;
assign LUT_3[24942] = 32'b00000000000000001101001001001110;
assign LUT_3[24943] = 32'b00000000000000010011110100101011;
assign LUT_3[24944] = 32'b00000000000000001011101101110001;
assign LUT_3[24945] = 32'b00000000000000010010011001001110;
assign LUT_3[24946] = 32'b00000000000000001101110101010101;
assign LUT_3[24947] = 32'b00000000000000010100100000110010;
assign LUT_3[24948] = 32'b00000000000000001000111011100111;
assign LUT_3[24949] = 32'b00000000000000001111100111000100;
assign LUT_3[24950] = 32'b00000000000000001011000011001011;
assign LUT_3[24951] = 32'b00000000000000010001101110101000;
assign LUT_3[24952] = 32'b00000000000000010001000110110111;
assign LUT_3[24953] = 32'b00000000000000010111110010010100;
assign LUT_3[24954] = 32'b00000000000000010011001110011011;
assign LUT_3[24955] = 32'b00000000000000011001111001111000;
assign LUT_3[24956] = 32'b00000000000000001110010100101101;
assign LUT_3[24957] = 32'b00000000000000010101000000001010;
assign LUT_3[24958] = 32'b00000000000000010000011100010001;
assign LUT_3[24959] = 32'b00000000000000010111000111101110;
assign LUT_3[24960] = 32'b00000000000000001001011110100001;
assign LUT_3[24961] = 32'b00000000000000010000001001111110;
assign LUT_3[24962] = 32'b00000000000000001011100110000101;
assign LUT_3[24963] = 32'b00000000000000010010010001100010;
assign LUT_3[24964] = 32'b00000000000000000110101100010111;
assign LUT_3[24965] = 32'b00000000000000001101010111110100;
assign LUT_3[24966] = 32'b00000000000000001000110011111011;
assign LUT_3[24967] = 32'b00000000000000001111011111011000;
assign LUT_3[24968] = 32'b00000000000000001110110111100111;
assign LUT_3[24969] = 32'b00000000000000010101100011000100;
assign LUT_3[24970] = 32'b00000000000000010000111111001011;
assign LUT_3[24971] = 32'b00000000000000010111101010101000;
assign LUT_3[24972] = 32'b00000000000000001100000101011101;
assign LUT_3[24973] = 32'b00000000000000010010110000111010;
assign LUT_3[24974] = 32'b00000000000000001110001101000001;
assign LUT_3[24975] = 32'b00000000000000010100111000011110;
assign LUT_3[24976] = 32'b00000000000000001100110001100100;
assign LUT_3[24977] = 32'b00000000000000010011011101000001;
assign LUT_3[24978] = 32'b00000000000000001110111001001000;
assign LUT_3[24979] = 32'b00000000000000010101100100100101;
assign LUT_3[24980] = 32'b00000000000000001001111111011010;
assign LUT_3[24981] = 32'b00000000000000010000101010110111;
assign LUT_3[24982] = 32'b00000000000000001100000110111110;
assign LUT_3[24983] = 32'b00000000000000010010110010011011;
assign LUT_3[24984] = 32'b00000000000000010010001010101010;
assign LUT_3[24985] = 32'b00000000000000011000110110000111;
assign LUT_3[24986] = 32'b00000000000000010100010010001110;
assign LUT_3[24987] = 32'b00000000000000011010111101101011;
assign LUT_3[24988] = 32'b00000000000000001111011000100000;
assign LUT_3[24989] = 32'b00000000000000010110000011111101;
assign LUT_3[24990] = 32'b00000000000000010001100000000100;
assign LUT_3[24991] = 32'b00000000000000011000001011100001;
assign LUT_3[24992] = 32'b00000000000000001010101101000001;
assign LUT_3[24993] = 32'b00000000000000010001011000011110;
assign LUT_3[24994] = 32'b00000000000000001100110100100101;
assign LUT_3[24995] = 32'b00000000000000010011100000000010;
assign LUT_3[24996] = 32'b00000000000000000111111010110111;
assign LUT_3[24997] = 32'b00000000000000001110100110010100;
assign LUT_3[24998] = 32'b00000000000000001010000010011011;
assign LUT_3[24999] = 32'b00000000000000010000101101111000;
assign LUT_3[25000] = 32'b00000000000000010000000110000111;
assign LUT_3[25001] = 32'b00000000000000010110110001100100;
assign LUT_3[25002] = 32'b00000000000000010010001101101011;
assign LUT_3[25003] = 32'b00000000000000011000111001001000;
assign LUT_3[25004] = 32'b00000000000000001101010011111101;
assign LUT_3[25005] = 32'b00000000000000010011111111011010;
assign LUT_3[25006] = 32'b00000000000000001111011011100001;
assign LUT_3[25007] = 32'b00000000000000010110000110111110;
assign LUT_3[25008] = 32'b00000000000000001110000000000100;
assign LUT_3[25009] = 32'b00000000000000010100101011100001;
assign LUT_3[25010] = 32'b00000000000000010000000111101000;
assign LUT_3[25011] = 32'b00000000000000010110110011000101;
assign LUT_3[25012] = 32'b00000000000000001011001101111010;
assign LUT_3[25013] = 32'b00000000000000010001111001010111;
assign LUT_3[25014] = 32'b00000000000000001101010101011110;
assign LUT_3[25015] = 32'b00000000000000010100000000111011;
assign LUT_3[25016] = 32'b00000000000000010011011001001010;
assign LUT_3[25017] = 32'b00000000000000011010000100100111;
assign LUT_3[25018] = 32'b00000000000000010101100000101110;
assign LUT_3[25019] = 32'b00000000000000011100001100001011;
assign LUT_3[25020] = 32'b00000000000000010000100111000000;
assign LUT_3[25021] = 32'b00000000000000010111010010011101;
assign LUT_3[25022] = 32'b00000000000000010010101110100100;
assign LUT_3[25023] = 32'b00000000000000011001011010000001;
assign LUT_3[25024] = 32'b00000000000000001001010111001100;
assign LUT_3[25025] = 32'b00000000000000010000000010101001;
assign LUT_3[25026] = 32'b00000000000000001011011110110000;
assign LUT_3[25027] = 32'b00000000000000010010001010001101;
assign LUT_3[25028] = 32'b00000000000000000110100101000010;
assign LUT_3[25029] = 32'b00000000000000001101010000011111;
assign LUT_3[25030] = 32'b00000000000000001000101100100110;
assign LUT_3[25031] = 32'b00000000000000001111011000000011;
assign LUT_3[25032] = 32'b00000000000000001110110000010010;
assign LUT_3[25033] = 32'b00000000000000010101011011101111;
assign LUT_3[25034] = 32'b00000000000000010000110111110110;
assign LUT_3[25035] = 32'b00000000000000010111100011010011;
assign LUT_3[25036] = 32'b00000000000000001011111110001000;
assign LUT_3[25037] = 32'b00000000000000010010101001100101;
assign LUT_3[25038] = 32'b00000000000000001110000101101100;
assign LUT_3[25039] = 32'b00000000000000010100110001001001;
assign LUT_3[25040] = 32'b00000000000000001100101010001111;
assign LUT_3[25041] = 32'b00000000000000010011010101101100;
assign LUT_3[25042] = 32'b00000000000000001110110001110011;
assign LUT_3[25043] = 32'b00000000000000010101011101010000;
assign LUT_3[25044] = 32'b00000000000000001001111000000101;
assign LUT_3[25045] = 32'b00000000000000010000100011100010;
assign LUT_3[25046] = 32'b00000000000000001011111111101001;
assign LUT_3[25047] = 32'b00000000000000010010101011000110;
assign LUT_3[25048] = 32'b00000000000000010010000011010101;
assign LUT_3[25049] = 32'b00000000000000011000101110110010;
assign LUT_3[25050] = 32'b00000000000000010100001010111001;
assign LUT_3[25051] = 32'b00000000000000011010110110010110;
assign LUT_3[25052] = 32'b00000000000000001111010001001011;
assign LUT_3[25053] = 32'b00000000000000010101111100101000;
assign LUT_3[25054] = 32'b00000000000000010001011000101111;
assign LUT_3[25055] = 32'b00000000000000011000000100001100;
assign LUT_3[25056] = 32'b00000000000000001010100101101100;
assign LUT_3[25057] = 32'b00000000000000010001010001001001;
assign LUT_3[25058] = 32'b00000000000000001100101101010000;
assign LUT_3[25059] = 32'b00000000000000010011011000101101;
assign LUT_3[25060] = 32'b00000000000000000111110011100010;
assign LUT_3[25061] = 32'b00000000000000001110011110111111;
assign LUT_3[25062] = 32'b00000000000000001001111011000110;
assign LUT_3[25063] = 32'b00000000000000010000100110100011;
assign LUT_3[25064] = 32'b00000000000000001111111110110010;
assign LUT_3[25065] = 32'b00000000000000010110101010001111;
assign LUT_3[25066] = 32'b00000000000000010010000110010110;
assign LUT_3[25067] = 32'b00000000000000011000110001110011;
assign LUT_3[25068] = 32'b00000000000000001101001100101000;
assign LUT_3[25069] = 32'b00000000000000010011111000000101;
assign LUT_3[25070] = 32'b00000000000000001111010100001100;
assign LUT_3[25071] = 32'b00000000000000010101111111101001;
assign LUT_3[25072] = 32'b00000000000000001101111000101111;
assign LUT_3[25073] = 32'b00000000000000010100100100001100;
assign LUT_3[25074] = 32'b00000000000000010000000000010011;
assign LUT_3[25075] = 32'b00000000000000010110101011110000;
assign LUT_3[25076] = 32'b00000000000000001011000110100101;
assign LUT_3[25077] = 32'b00000000000000010001110010000010;
assign LUT_3[25078] = 32'b00000000000000001101001110001001;
assign LUT_3[25079] = 32'b00000000000000010011111001100110;
assign LUT_3[25080] = 32'b00000000000000010011010001110101;
assign LUT_3[25081] = 32'b00000000000000011001111101010010;
assign LUT_3[25082] = 32'b00000000000000010101011001011001;
assign LUT_3[25083] = 32'b00000000000000011100000100110110;
assign LUT_3[25084] = 32'b00000000000000010000011111101011;
assign LUT_3[25085] = 32'b00000000000000010111001011001000;
assign LUT_3[25086] = 32'b00000000000000010010100111001111;
assign LUT_3[25087] = 32'b00000000000000011001010010101100;
assign LUT_3[25088] = 32'b00000000000000001110011001001110;
assign LUT_3[25089] = 32'b00000000000000010101000100101011;
assign LUT_3[25090] = 32'b00000000000000010000100000110010;
assign LUT_3[25091] = 32'b00000000000000010111001100001111;
assign LUT_3[25092] = 32'b00000000000000001011100111000100;
assign LUT_3[25093] = 32'b00000000000000010010010010100001;
assign LUT_3[25094] = 32'b00000000000000001101101110101000;
assign LUT_3[25095] = 32'b00000000000000010100011010000101;
assign LUT_3[25096] = 32'b00000000000000010011110010010100;
assign LUT_3[25097] = 32'b00000000000000011010011101110001;
assign LUT_3[25098] = 32'b00000000000000010101111001111000;
assign LUT_3[25099] = 32'b00000000000000011100100101010101;
assign LUT_3[25100] = 32'b00000000000000010001000000001010;
assign LUT_3[25101] = 32'b00000000000000010111101011100111;
assign LUT_3[25102] = 32'b00000000000000010011000111101110;
assign LUT_3[25103] = 32'b00000000000000011001110011001011;
assign LUT_3[25104] = 32'b00000000000000010001101100010001;
assign LUT_3[25105] = 32'b00000000000000011000010111101110;
assign LUT_3[25106] = 32'b00000000000000010011110011110101;
assign LUT_3[25107] = 32'b00000000000000011010011111010010;
assign LUT_3[25108] = 32'b00000000000000001110111010000111;
assign LUT_3[25109] = 32'b00000000000000010101100101100100;
assign LUT_3[25110] = 32'b00000000000000010001000001101011;
assign LUT_3[25111] = 32'b00000000000000010111101101001000;
assign LUT_3[25112] = 32'b00000000000000010111000101010111;
assign LUT_3[25113] = 32'b00000000000000011101110000110100;
assign LUT_3[25114] = 32'b00000000000000011001001100111011;
assign LUT_3[25115] = 32'b00000000000000011111111000011000;
assign LUT_3[25116] = 32'b00000000000000010100010011001101;
assign LUT_3[25117] = 32'b00000000000000011010111110101010;
assign LUT_3[25118] = 32'b00000000000000010110011010110001;
assign LUT_3[25119] = 32'b00000000000000011101000110001110;
assign LUT_3[25120] = 32'b00000000000000001111100111101110;
assign LUT_3[25121] = 32'b00000000000000010110010011001011;
assign LUT_3[25122] = 32'b00000000000000010001101111010010;
assign LUT_3[25123] = 32'b00000000000000011000011010101111;
assign LUT_3[25124] = 32'b00000000000000001100110101100100;
assign LUT_3[25125] = 32'b00000000000000010011100001000001;
assign LUT_3[25126] = 32'b00000000000000001110111101001000;
assign LUT_3[25127] = 32'b00000000000000010101101000100101;
assign LUT_3[25128] = 32'b00000000000000010101000000110100;
assign LUT_3[25129] = 32'b00000000000000011011101100010001;
assign LUT_3[25130] = 32'b00000000000000010111001000011000;
assign LUT_3[25131] = 32'b00000000000000011101110011110101;
assign LUT_3[25132] = 32'b00000000000000010010001110101010;
assign LUT_3[25133] = 32'b00000000000000011000111010000111;
assign LUT_3[25134] = 32'b00000000000000010100010110001110;
assign LUT_3[25135] = 32'b00000000000000011011000001101011;
assign LUT_3[25136] = 32'b00000000000000010010111010110001;
assign LUT_3[25137] = 32'b00000000000000011001100110001110;
assign LUT_3[25138] = 32'b00000000000000010101000010010101;
assign LUT_3[25139] = 32'b00000000000000011011101101110010;
assign LUT_3[25140] = 32'b00000000000000010000001000100111;
assign LUT_3[25141] = 32'b00000000000000010110110100000100;
assign LUT_3[25142] = 32'b00000000000000010010010000001011;
assign LUT_3[25143] = 32'b00000000000000011000111011101000;
assign LUT_3[25144] = 32'b00000000000000011000010011110111;
assign LUT_3[25145] = 32'b00000000000000011110111111010100;
assign LUT_3[25146] = 32'b00000000000000011010011011011011;
assign LUT_3[25147] = 32'b00000000000000100001000110111000;
assign LUT_3[25148] = 32'b00000000000000010101100001101101;
assign LUT_3[25149] = 32'b00000000000000011100001101001010;
assign LUT_3[25150] = 32'b00000000000000010111101001010001;
assign LUT_3[25151] = 32'b00000000000000011110010100101110;
assign LUT_3[25152] = 32'b00000000000000001110010001111001;
assign LUT_3[25153] = 32'b00000000000000010100111101010110;
assign LUT_3[25154] = 32'b00000000000000010000011001011101;
assign LUT_3[25155] = 32'b00000000000000010111000100111010;
assign LUT_3[25156] = 32'b00000000000000001011011111101111;
assign LUT_3[25157] = 32'b00000000000000010010001011001100;
assign LUT_3[25158] = 32'b00000000000000001101100111010011;
assign LUT_3[25159] = 32'b00000000000000010100010010110000;
assign LUT_3[25160] = 32'b00000000000000010011101010111111;
assign LUT_3[25161] = 32'b00000000000000011010010110011100;
assign LUT_3[25162] = 32'b00000000000000010101110010100011;
assign LUT_3[25163] = 32'b00000000000000011100011110000000;
assign LUT_3[25164] = 32'b00000000000000010000111000110101;
assign LUT_3[25165] = 32'b00000000000000010111100100010010;
assign LUT_3[25166] = 32'b00000000000000010011000000011001;
assign LUT_3[25167] = 32'b00000000000000011001101011110110;
assign LUT_3[25168] = 32'b00000000000000010001100100111100;
assign LUT_3[25169] = 32'b00000000000000011000010000011001;
assign LUT_3[25170] = 32'b00000000000000010011101100100000;
assign LUT_3[25171] = 32'b00000000000000011010010111111101;
assign LUT_3[25172] = 32'b00000000000000001110110010110010;
assign LUT_3[25173] = 32'b00000000000000010101011110001111;
assign LUT_3[25174] = 32'b00000000000000010000111010010110;
assign LUT_3[25175] = 32'b00000000000000010111100101110011;
assign LUT_3[25176] = 32'b00000000000000010110111110000010;
assign LUT_3[25177] = 32'b00000000000000011101101001011111;
assign LUT_3[25178] = 32'b00000000000000011001000101100110;
assign LUT_3[25179] = 32'b00000000000000011111110001000011;
assign LUT_3[25180] = 32'b00000000000000010100001011111000;
assign LUT_3[25181] = 32'b00000000000000011010110111010101;
assign LUT_3[25182] = 32'b00000000000000010110010011011100;
assign LUT_3[25183] = 32'b00000000000000011100111110111001;
assign LUT_3[25184] = 32'b00000000000000001111100000011001;
assign LUT_3[25185] = 32'b00000000000000010110001011110110;
assign LUT_3[25186] = 32'b00000000000000010001100111111101;
assign LUT_3[25187] = 32'b00000000000000011000010011011010;
assign LUT_3[25188] = 32'b00000000000000001100101110001111;
assign LUT_3[25189] = 32'b00000000000000010011011001101100;
assign LUT_3[25190] = 32'b00000000000000001110110101110011;
assign LUT_3[25191] = 32'b00000000000000010101100001010000;
assign LUT_3[25192] = 32'b00000000000000010100111001011111;
assign LUT_3[25193] = 32'b00000000000000011011100100111100;
assign LUT_3[25194] = 32'b00000000000000010111000001000011;
assign LUT_3[25195] = 32'b00000000000000011101101100100000;
assign LUT_3[25196] = 32'b00000000000000010010000111010101;
assign LUT_3[25197] = 32'b00000000000000011000110010110010;
assign LUT_3[25198] = 32'b00000000000000010100001110111001;
assign LUT_3[25199] = 32'b00000000000000011010111010010110;
assign LUT_3[25200] = 32'b00000000000000010010110011011100;
assign LUT_3[25201] = 32'b00000000000000011001011110111001;
assign LUT_3[25202] = 32'b00000000000000010100111011000000;
assign LUT_3[25203] = 32'b00000000000000011011100110011101;
assign LUT_3[25204] = 32'b00000000000000010000000001010010;
assign LUT_3[25205] = 32'b00000000000000010110101100101111;
assign LUT_3[25206] = 32'b00000000000000010010001000110110;
assign LUT_3[25207] = 32'b00000000000000011000110100010011;
assign LUT_3[25208] = 32'b00000000000000011000001100100010;
assign LUT_3[25209] = 32'b00000000000000011110110111111111;
assign LUT_3[25210] = 32'b00000000000000011010010100000110;
assign LUT_3[25211] = 32'b00000000000000100000111111100011;
assign LUT_3[25212] = 32'b00000000000000010101011010011000;
assign LUT_3[25213] = 32'b00000000000000011100000101110101;
assign LUT_3[25214] = 32'b00000000000000010111100001111100;
assign LUT_3[25215] = 32'b00000000000000011110001101011001;
assign LUT_3[25216] = 32'b00000000000000010000100100001100;
assign LUT_3[25217] = 32'b00000000000000010111001111101001;
assign LUT_3[25218] = 32'b00000000000000010010101011110000;
assign LUT_3[25219] = 32'b00000000000000011001010111001101;
assign LUT_3[25220] = 32'b00000000000000001101110010000010;
assign LUT_3[25221] = 32'b00000000000000010100011101011111;
assign LUT_3[25222] = 32'b00000000000000001111111001100110;
assign LUT_3[25223] = 32'b00000000000000010110100101000011;
assign LUT_3[25224] = 32'b00000000000000010101111101010010;
assign LUT_3[25225] = 32'b00000000000000011100101000101111;
assign LUT_3[25226] = 32'b00000000000000011000000100110110;
assign LUT_3[25227] = 32'b00000000000000011110110000010011;
assign LUT_3[25228] = 32'b00000000000000010011001011001000;
assign LUT_3[25229] = 32'b00000000000000011001110110100101;
assign LUT_3[25230] = 32'b00000000000000010101010010101100;
assign LUT_3[25231] = 32'b00000000000000011011111110001001;
assign LUT_3[25232] = 32'b00000000000000010011110111001111;
assign LUT_3[25233] = 32'b00000000000000011010100010101100;
assign LUT_3[25234] = 32'b00000000000000010101111110110011;
assign LUT_3[25235] = 32'b00000000000000011100101010010000;
assign LUT_3[25236] = 32'b00000000000000010001000101000101;
assign LUT_3[25237] = 32'b00000000000000010111110000100010;
assign LUT_3[25238] = 32'b00000000000000010011001100101001;
assign LUT_3[25239] = 32'b00000000000000011001111000000110;
assign LUT_3[25240] = 32'b00000000000000011001010000010101;
assign LUT_3[25241] = 32'b00000000000000011111111011110010;
assign LUT_3[25242] = 32'b00000000000000011011010111111001;
assign LUT_3[25243] = 32'b00000000000000100010000011010110;
assign LUT_3[25244] = 32'b00000000000000010110011110001011;
assign LUT_3[25245] = 32'b00000000000000011101001001101000;
assign LUT_3[25246] = 32'b00000000000000011000100101101111;
assign LUT_3[25247] = 32'b00000000000000011111010001001100;
assign LUT_3[25248] = 32'b00000000000000010001110010101100;
assign LUT_3[25249] = 32'b00000000000000011000011110001001;
assign LUT_3[25250] = 32'b00000000000000010011111010010000;
assign LUT_3[25251] = 32'b00000000000000011010100101101101;
assign LUT_3[25252] = 32'b00000000000000001111000000100010;
assign LUT_3[25253] = 32'b00000000000000010101101011111111;
assign LUT_3[25254] = 32'b00000000000000010001001000000110;
assign LUT_3[25255] = 32'b00000000000000010111110011100011;
assign LUT_3[25256] = 32'b00000000000000010111001011110010;
assign LUT_3[25257] = 32'b00000000000000011101110111001111;
assign LUT_3[25258] = 32'b00000000000000011001010011010110;
assign LUT_3[25259] = 32'b00000000000000011111111110110011;
assign LUT_3[25260] = 32'b00000000000000010100011001101000;
assign LUT_3[25261] = 32'b00000000000000011011000101000101;
assign LUT_3[25262] = 32'b00000000000000010110100001001100;
assign LUT_3[25263] = 32'b00000000000000011101001100101001;
assign LUT_3[25264] = 32'b00000000000000010101000101101111;
assign LUT_3[25265] = 32'b00000000000000011011110001001100;
assign LUT_3[25266] = 32'b00000000000000010111001101010011;
assign LUT_3[25267] = 32'b00000000000000011101111000110000;
assign LUT_3[25268] = 32'b00000000000000010010010011100101;
assign LUT_3[25269] = 32'b00000000000000011000111111000010;
assign LUT_3[25270] = 32'b00000000000000010100011011001001;
assign LUT_3[25271] = 32'b00000000000000011011000110100110;
assign LUT_3[25272] = 32'b00000000000000011010011110110101;
assign LUT_3[25273] = 32'b00000000000000100001001010010010;
assign LUT_3[25274] = 32'b00000000000000011100100110011001;
assign LUT_3[25275] = 32'b00000000000000100011010001110110;
assign LUT_3[25276] = 32'b00000000000000010111101100101011;
assign LUT_3[25277] = 32'b00000000000000011110011000001000;
assign LUT_3[25278] = 32'b00000000000000011001110100001111;
assign LUT_3[25279] = 32'b00000000000000100000011111101100;
assign LUT_3[25280] = 32'b00000000000000010000011100110111;
assign LUT_3[25281] = 32'b00000000000000010111001000010100;
assign LUT_3[25282] = 32'b00000000000000010010100100011011;
assign LUT_3[25283] = 32'b00000000000000011001001111111000;
assign LUT_3[25284] = 32'b00000000000000001101101010101101;
assign LUT_3[25285] = 32'b00000000000000010100010110001010;
assign LUT_3[25286] = 32'b00000000000000001111110010010001;
assign LUT_3[25287] = 32'b00000000000000010110011101101110;
assign LUT_3[25288] = 32'b00000000000000010101110101111101;
assign LUT_3[25289] = 32'b00000000000000011100100001011010;
assign LUT_3[25290] = 32'b00000000000000010111111101100001;
assign LUT_3[25291] = 32'b00000000000000011110101000111110;
assign LUT_3[25292] = 32'b00000000000000010011000011110011;
assign LUT_3[25293] = 32'b00000000000000011001101111010000;
assign LUT_3[25294] = 32'b00000000000000010101001011010111;
assign LUT_3[25295] = 32'b00000000000000011011110110110100;
assign LUT_3[25296] = 32'b00000000000000010011101111111010;
assign LUT_3[25297] = 32'b00000000000000011010011011010111;
assign LUT_3[25298] = 32'b00000000000000010101110111011110;
assign LUT_3[25299] = 32'b00000000000000011100100010111011;
assign LUT_3[25300] = 32'b00000000000000010000111101110000;
assign LUT_3[25301] = 32'b00000000000000010111101001001101;
assign LUT_3[25302] = 32'b00000000000000010011000101010100;
assign LUT_3[25303] = 32'b00000000000000011001110000110001;
assign LUT_3[25304] = 32'b00000000000000011001001001000000;
assign LUT_3[25305] = 32'b00000000000000011111110100011101;
assign LUT_3[25306] = 32'b00000000000000011011010000100100;
assign LUT_3[25307] = 32'b00000000000000100001111100000001;
assign LUT_3[25308] = 32'b00000000000000010110010110110110;
assign LUT_3[25309] = 32'b00000000000000011101000010010011;
assign LUT_3[25310] = 32'b00000000000000011000011110011010;
assign LUT_3[25311] = 32'b00000000000000011111001001110111;
assign LUT_3[25312] = 32'b00000000000000010001101011010111;
assign LUT_3[25313] = 32'b00000000000000011000010110110100;
assign LUT_3[25314] = 32'b00000000000000010011110010111011;
assign LUT_3[25315] = 32'b00000000000000011010011110011000;
assign LUT_3[25316] = 32'b00000000000000001110111001001101;
assign LUT_3[25317] = 32'b00000000000000010101100100101010;
assign LUT_3[25318] = 32'b00000000000000010001000000110001;
assign LUT_3[25319] = 32'b00000000000000010111101100001110;
assign LUT_3[25320] = 32'b00000000000000010111000100011101;
assign LUT_3[25321] = 32'b00000000000000011101101111111010;
assign LUT_3[25322] = 32'b00000000000000011001001100000001;
assign LUT_3[25323] = 32'b00000000000000011111110111011110;
assign LUT_3[25324] = 32'b00000000000000010100010010010011;
assign LUT_3[25325] = 32'b00000000000000011010111101110000;
assign LUT_3[25326] = 32'b00000000000000010110011001110111;
assign LUT_3[25327] = 32'b00000000000000011101000101010100;
assign LUT_3[25328] = 32'b00000000000000010100111110011010;
assign LUT_3[25329] = 32'b00000000000000011011101001110111;
assign LUT_3[25330] = 32'b00000000000000010111000101111110;
assign LUT_3[25331] = 32'b00000000000000011101110001011011;
assign LUT_3[25332] = 32'b00000000000000010010001100010000;
assign LUT_3[25333] = 32'b00000000000000011000110111101101;
assign LUT_3[25334] = 32'b00000000000000010100010011110100;
assign LUT_3[25335] = 32'b00000000000000011010111111010001;
assign LUT_3[25336] = 32'b00000000000000011010010111100000;
assign LUT_3[25337] = 32'b00000000000000100001000010111101;
assign LUT_3[25338] = 32'b00000000000000011100011111000100;
assign LUT_3[25339] = 32'b00000000000000100011001010100001;
assign LUT_3[25340] = 32'b00000000000000010111100101010110;
assign LUT_3[25341] = 32'b00000000000000011110010000110011;
assign LUT_3[25342] = 32'b00000000000000011001101100111010;
assign LUT_3[25343] = 32'b00000000000000100000011000010111;
assign LUT_3[25344] = 32'b00000000000000001010101000101111;
assign LUT_3[25345] = 32'b00000000000000010001010100001100;
assign LUT_3[25346] = 32'b00000000000000001100110000010011;
assign LUT_3[25347] = 32'b00000000000000010011011011110000;
assign LUT_3[25348] = 32'b00000000000000000111110110100101;
assign LUT_3[25349] = 32'b00000000000000001110100010000010;
assign LUT_3[25350] = 32'b00000000000000001001111110001001;
assign LUT_3[25351] = 32'b00000000000000010000101001100110;
assign LUT_3[25352] = 32'b00000000000000010000000001110101;
assign LUT_3[25353] = 32'b00000000000000010110101101010010;
assign LUT_3[25354] = 32'b00000000000000010010001001011001;
assign LUT_3[25355] = 32'b00000000000000011000110100110110;
assign LUT_3[25356] = 32'b00000000000000001101001111101011;
assign LUT_3[25357] = 32'b00000000000000010011111011001000;
assign LUT_3[25358] = 32'b00000000000000001111010111001111;
assign LUT_3[25359] = 32'b00000000000000010110000010101100;
assign LUT_3[25360] = 32'b00000000000000001101111011110010;
assign LUT_3[25361] = 32'b00000000000000010100100111001111;
assign LUT_3[25362] = 32'b00000000000000010000000011010110;
assign LUT_3[25363] = 32'b00000000000000010110101110110011;
assign LUT_3[25364] = 32'b00000000000000001011001001101000;
assign LUT_3[25365] = 32'b00000000000000010001110101000101;
assign LUT_3[25366] = 32'b00000000000000001101010001001100;
assign LUT_3[25367] = 32'b00000000000000010011111100101001;
assign LUT_3[25368] = 32'b00000000000000010011010100111000;
assign LUT_3[25369] = 32'b00000000000000011010000000010101;
assign LUT_3[25370] = 32'b00000000000000010101011100011100;
assign LUT_3[25371] = 32'b00000000000000011100000111111001;
assign LUT_3[25372] = 32'b00000000000000010000100010101110;
assign LUT_3[25373] = 32'b00000000000000010111001110001011;
assign LUT_3[25374] = 32'b00000000000000010010101010010010;
assign LUT_3[25375] = 32'b00000000000000011001010101101111;
assign LUT_3[25376] = 32'b00000000000000001011110111001111;
assign LUT_3[25377] = 32'b00000000000000010010100010101100;
assign LUT_3[25378] = 32'b00000000000000001101111110110011;
assign LUT_3[25379] = 32'b00000000000000010100101010010000;
assign LUT_3[25380] = 32'b00000000000000001001000101000101;
assign LUT_3[25381] = 32'b00000000000000001111110000100010;
assign LUT_3[25382] = 32'b00000000000000001011001100101001;
assign LUT_3[25383] = 32'b00000000000000010001111000000110;
assign LUT_3[25384] = 32'b00000000000000010001010000010101;
assign LUT_3[25385] = 32'b00000000000000010111111011110010;
assign LUT_3[25386] = 32'b00000000000000010011010111111001;
assign LUT_3[25387] = 32'b00000000000000011010000011010110;
assign LUT_3[25388] = 32'b00000000000000001110011110001011;
assign LUT_3[25389] = 32'b00000000000000010101001001101000;
assign LUT_3[25390] = 32'b00000000000000010000100101101111;
assign LUT_3[25391] = 32'b00000000000000010111010001001100;
assign LUT_3[25392] = 32'b00000000000000001111001010010010;
assign LUT_3[25393] = 32'b00000000000000010101110101101111;
assign LUT_3[25394] = 32'b00000000000000010001010001110110;
assign LUT_3[25395] = 32'b00000000000000010111111101010011;
assign LUT_3[25396] = 32'b00000000000000001100011000001000;
assign LUT_3[25397] = 32'b00000000000000010011000011100101;
assign LUT_3[25398] = 32'b00000000000000001110011111101100;
assign LUT_3[25399] = 32'b00000000000000010101001011001001;
assign LUT_3[25400] = 32'b00000000000000010100100011011000;
assign LUT_3[25401] = 32'b00000000000000011011001110110101;
assign LUT_3[25402] = 32'b00000000000000010110101010111100;
assign LUT_3[25403] = 32'b00000000000000011101010110011001;
assign LUT_3[25404] = 32'b00000000000000010001110001001110;
assign LUT_3[25405] = 32'b00000000000000011000011100101011;
assign LUT_3[25406] = 32'b00000000000000010011111000110010;
assign LUT_3[25407] = 32'b00000000000000011010100100001111;
assign LUT_3[25408] = 32'b00000000000000001010100001011010;
assign LUT_3[25409] = 32'b00000000000000010001001100110111;
assign LUT_3[25410] = 32'b00000000000000001100101000111110;
assign LUT_3[25411] = 32'b00000000000000010011010100011011;
assign LUT_3[25412] = 32'b00000000000000000111101111010000;
assign LUT_3[25413] = 32'b00000000000000001110011010101101;
assign LUT_3[25414] = 32'b00000000000000001001110110110100;
assign LUT_3[25415] = 32'b00000000000000010000100010010001;
assign LUT_3[25416] = 32'b00000000000000001111111010100000;
assign LUT_3[25417] = 32'b00000000000000010110100101111101;
assign LUT_3[25418] = 32'b00000000000000010010000010000100;
assign LUT_3[25419] = 32'b00000000000000011000101101100001;
assign LUT_3[25420] = 32'b00000000000000001101001000010110;
assign LUT_3[25421] = 32'b00000000000000010011110011110011;
assign LUT_3[25422] = 32'b00000000000000001111001111111010;
assign LUT_3[25423] = 32'b00000000000000010101111011010111;
assign LUT_3[25424] = 32'b00000000000000001101110100011101;
assign LUT_3[25425] = 32'b00000000000000010100011111111010;
assign LUT_3[25426] = 32'b00000000000000001111111100000001;
assign LUT_3[25427] = 32'b00000000000000010110100111011110;
assign LUT_3[25428] = 32'b00000000000000001011000010010011;
assign LUT_3[25429] = 32'b00000000000000010001101101110000;
assign LUT_3[25430] = 32'b00000000000000001101001001110111;
assign LUT_3[25431] = 32'b00000000000000010011110101010100;
assign LUT_3[25432] = 32'b00000000000000010011001101100011;
assign LUT_3[25433] = 32'b00000000000000011001111001000000;
assign LUT_3[25434] = 32'b00000000000000010101010101000111;
assign LUT_3[25435] = 32'b00000000000000011100000000100100;
assign LUT_3[25436] = 32'b00000000000000010000011011011001;
assign LUT_3[25437] = 32'b00000000000000010111000110110110;
assign LUT_3[25438] = 32'b00000000000000010010100010111101;
assign LUT_3[25439] = 32'b00000000000000011001001110011010;
assign LUT_3[25440] = 32'b00000000000000001011101111111010;
assign LUT_3[25441] = 32'b00000000000000010010011011010111;
assign LUT_3[25442] = 32'b00000000000000001101110111011110;
assign LUT_3[25443] = 32'b00000000000000010100100010111011;
assign LUT_3[25444] = 32'b00000000000000001000111101110000;
assign LUT_3[25445] = 32'b00000000000000001111101001001101;
assign LUT_3[25446] = 32'b00000000000000001011000101010100;
assign LUT_3[25447] = 32'b00000000000000010001110000110001;
assign LUT_3[25448] = 32'b00000000000000010001001001000000;
assign LUT_3[25449] = 32'b00000000000000010111110100011101;
assign LUT_3[25450] = 32'b00000000000000010011010000100100;
assign LUT_3[25451] = 32'b00000000000000011001111100000001;
assign LUT_3[25452] = 32'b00000000000000001110010110110110;
assign LUT_3[25453] = 32'b00000000000000010101000010010011;
assign LUT_3[25454] = 32'b00000000000000010000011110011010;
assign LUT_3[25455] = 32'b00000000000000010111001001110111;
assign LUT_3[25456] = 32'b00000000000000001111000010111101;
assign LUT_3[25457] = 32'b00000000000000010101101110011010;
assign LUT_3[25458] = 32'b00000000000000010001001010100001;
assign LUT_3[25459] = 32'b00000000000000010111110101111110;
assign LUT_3[25460] = 32'b00000000000000001100010000110011;
assign LUT_3[25461] = 32'b00000000000000010010111100010000;
assign LUT_3[25462] = 32'b00000000000000001110011000010111;
assign LUT_3[25463] = 32'b00000000000000010101000011110100;
assign LUT_3[25464] = 32'b00000000000000010100011100000011;
assign LUT_3[25465] = 32'b00000000000000011011000111100000;
assign LUT_3[25466] = 32'b00000000000000010110100011100111;
assign LUT_3[25467] = 32'b00000000000000011101001111000100;
assign LUT_3[25468] = 32'b00000000000000010001101001111001;
assign LUT_3[25469] = 32'b00000000000000011000010101010110;
assign LUT_3[25470] = 32'b00000000000000010011110001011101;
assign LUT_3[25471] = 32'b00000000000000011010011100111010;
assign LUT_3[25472] = 32'b00000000000000001100110011101101;
assign LUT_3[25473] = 32'b00000000000000010011011111001010;
assign LUT_3[25474] = 32'b00000000000000001110111011010001;
assign LUT_3[25475] = 32'b00000000000000010101100110101110;
assign LUT_3[25476] = 32'b00000000000000001010000001100011;
assign LUT_3[25477] = 32'b00000000000000010000101101000000;
assign LUT_3[25478] = 32'b00000000000000001100001001000111;
assign LUT_3[25479] = 32'b00000000000000010010110100100100;
assign LUT_3[25480] = 32'b00000000000000010010001100110011;
assign LUT_3[25481] = 32'b00000000000000011000111000010000;
assign LUT_3[25482] = 32'b00000000000000010100010100010111;
assign LUT_3[25483] = 32'b00000000000000011010111111110100;
assign LUT_3[25484] = 32'b00000000000000001111011010101001;
assign LUT_3[25485] = 32'b00000000000000010110000110000110;
assign LUT_3[25486] = 32'b00000000000000010001100010001101;
assign LUT_3[25487] = 32'b00000000000000011000001101101010;
assign LUT_3[25488] = 32'b00000000000000010000000110110000;
assign LUT_3[25489] = 32'b00000000000000010110110010001101;
assign LUT_3[25490] = 32'b00000000000000010010001110010100;
assign LUT_3[25491] = 32'b00000000000000011000111001110001;
assign LUT_3[25492] = 32'b00000000000000001101010100100110;
assign LUT_3[25493] = 32'b00000000000000010100000000000011;
assign LUT_3[25494] = 32'b00000000000000001111011100001010;
assign LUT_3[25495] = 32'b00000000000000010110000111100111;
assign LUT_3[25496] = 32'b00000000000000010101011111110110;
assign LUT_3[25497] = 32'b00000000000000011100001011010011;
assign LUT_3[25498] = 32'b00000000000000010111100111011010;
assign LUT_3[25499] = 32'b00000000000000011110010010110111;
assign LUT_3[25500] = 32'b00000000000000010010101101101100;
assign LUT_3[25501] = 32'b00000000000000011001011001001001;
assign LUT_3[25502] = 32'b00000000000000010100110101010000;
assign LUT_3[25503] = 32'b00000000000000011011100000101101;
assign LUT_3[25504] = 32'b00000000000000001110000010001101;
assign LUT_3[25505] = 32'b00000000000000010100101101101010;
assign LUT_3[25506] = 32'b00000000000000010000001001110001;
assign LUT_3[25507] = 32'b00000000000000010110110101001110;
assign LUT_3[25508] = 32'b00000000000000001011010000000011;
assign LUT_3[25509] = 32'b00000000000000010001111011100000;
assign LUT_3[25510] = 32'b00000000000000001101010111100111;
assign LUT_3[25511] = 32'b00000000000000010100000011000100;
assign LUT_3[25512] = 32'b00000000000000010011011011010011;
assign LUT_3[25513] = 32'b00000000000000011010000110110000;
assign LUT_3[25514] = 32'b00000000000000010101100010110111;
assign LUT_3[25515] = 32'b00000000000000011100001110010100;
assign LUT_3[25516] = 32'b00000000000000010000101001001001;
assign LUT_3[25517] = 32'b00000000000000010111010100100110;
assign LUT_3[25518] = 32'b00000000000000010010110000101101;
assign LUT_3[25519] = 32'b00000000000000011001011100001010;
assign LUT_3[25520] = 32'b00000000000000010001010101010000;
assign LUT_3[25521] = 32'b00000000000000011000000000101101;
assign LUT_3[25522] = 32'b00000000000000010011011100110100;
assign LUT_3[25523] = 32'b00000000000000011010001000010001;
assign LUT_3[25524] = 32'b00000000000000001110100011000110;
assign LUT_3[25525] = 32'b00000000000000010101001110100011;
assign LUT_3[25526] = 32'b00000000000000010000101010101010;
assign LUT_3[25527] = 32'b00000000000000010111010110000111;
assign LUT_3[25528] = 32'b00000000000000010110101110010110;
assign LUT_3[25529] = 32'b00000000000000011101011001110011;
assign LUT_3[25530] = 32'b00000000000000011000110101111010;
assign LUT_3[25531] = 32'b00000000000000011111100001010111;
assign LUT_3[25532] = 32'b00000000000000010011111100001100;
assign LUT_3[25533] = 32'b00000000000000011010100111101001;
assign LUT_3[25534] = 32'b00000000000000010110000011110000;
assign LUT_3[25535] = 32'b00000000000000011100101111001101;
assign LUT_3[25536] = 32'b00000000000000001100101100011000;
assign LUT_3[25537] = 32'b00000000000000010011010111110101;
assign LUT_3[25538] = 32'b00000000000000001110110011111100;
assign LUT_3[25539] = 32'b00000000000000010101011111011001;
assign LUT_3[25540] = 32'b00000000000000001001111010001110;
assign LUT_3[25541] = 32'b00000000000000010000100101101011;
assign LUT_3[25542] = 32'b00000000000000001100000001110010;
assign LUT_3[25543] = 32'b00000000000000010010101101001111;
assign LUT_3[25544] = 32'b00000000000000010010000101011110;
assign LUT_3[25545] = 32'b00000000000000011000110000111011;
assign LUT_3[25546] = 32'b00000000000000010100001101000010;
assign LUT_3[25547] = 32'b00000000000000011010111000011111;
assign LUT_3[25548] = 32'b00000000000000001111010011010100;
assign LUT_3[25549] = 32'b00000000000000010101111110110001;
assign LUT_3[25550] = 32'b00000000000000010001011010111000;
assign LUT_3[25551] = 32'b00000000000000011000000110010101;
assign LUT_3[25552] = 32'b00000000000000001111111111011011;
assign LUT_3[25553] = 32'b00000000000000010110101010111000;
assign LUT_3[25554] = 32'b00000000000000010010000110111111;
assign LUT_3[25555] = 32'b00000000000000011000110010011100;
assign LUT_3[25556] = 32'b00000000000000001101001101010001;
assign LUT_3[25557] = 32'b00000000000000010011111000101110;
assign LUT_3[25558] = 32'b00000000000000001111010100110101;
assign LUT_3[25559] = 32'b00000000000000010110000000010010;
assign LUT_3[25560] = 32'b00000000000000010101011000100001;
assign LUT_3[25561] = 32'b00000000000000011100000011111110;
assign LUT_3[25562] = 32'b00000000000000010111100000000101;
assign LUT_3[25563] = 32'b00000000000000011110001011100010;
assign LUT_3[25564] = 32'b00000000000000010010100110010111;
assign LUT_3[25565] = 32'b00000000000000011001010001110100;
assign LUT_3[25566] = 32'b00000000000000010100101101111011;
assign LUT_3[25567] = 32'b00000000000000011011011001011000;
assign LUT_3[25568] = 32'b00000000000000001101111010111000;
assign LUT_3[25569] = 32'b00000000000000010100100110010101;
assign LUT_3[25570] = 32'b00000000000000010000000010011100;
assign LUT_3[25571] = 32'b00000000000000010110101101111001;
assign LUT_3[25572] = 32'b00000000000000001011001000101110;
assign LUT_3[25573] = 32'b00000000000000010001110100001011;
assign LUT_3[25574] = 32'b00000000000000001101010000010010;
assign LUT_3[25575] = 32'b00000000000000010011111011101111;
assign LUT_3[25576] = 32'b00000000000000010011010011111110;
assign LUT_3[25577] = 32'b00000000000000011001111111011011;
assign LUT_3[25578] = 32'b00000000000000010101011011100010;
assign LUT_3[25579] = 32'b00000000000000011100000110111111;
assign LUT_3[25580] = 32'b00000000000000010000100001110100;
assign LUT_3[25581] = 32'b00000000000000010111001101010001;
assign LUT_3[25582] = 32'b00000000000000010010101001011000;
assign LUT_3[25583] = 32'b00000000000000011001010100110101;
assign LUT_3[25584] = 32'b00000000000000010001001101111011;
assign LUT_3[25585] = 32'b00000000000000010111111001011000;
assign LUT_3[25586] = 32'b00000000000000010011010101011111;
assign LUT_3[25587] = 32'b00000000000000011010000000111100;
assign LUT_3[25588] = 32'b00000000000000001110011011110001;
assign LUT_3[25589] = 32'b00000000000000010101000111001110;
assign LUT_3[25590] = 32'b00000000000000010000100011010101;
assign LUT_3[25591] = 32'b00000000000000010111001110110010;
assign LUT_3[25592] = 32'b00000000000000010110100111000001;
assign LUT_3[25593] = 32'b00000000000000011101010010011110;
assign LUT_3[25594] = 32'b00000000000000011000101110100101;
assign LUT_3[25595] = 32'b00000000000000011111011010000010;
assign LUT_3[25596] = 32'b00000000000000010011110100110111;
assign LUT_3[25597] = 32'b00000000000000011010100000010100;
assign LUT_3[25598] = 32'b00000000000000010101111100011011;
assign LUT_3[25599] = 32'b00000000000000011100100111111000;
assign LUT_3[25600] = 32'b00000000000000010001101000111111;
assign LUT_3[25601] = 32'b00000000000000011000010100011100;
assign LUT_3[25602] = 32'b00000000000000010011110000100011;
assign LUT_3[25603] = 32'b00000000000000011010011100000000;
assign LUT_3[25604] = 32'b00000000000000001110110110110101;
assign LUT_3[25605] = 32'b00000000000000010101100010010010;
assign LUT_3[25606] = 32'b00000000000000010000111110011001;
assign LUT_3[25607] = 32'b00000000000000010111101001110110;
assign LUT_3[25608] = 32'b00000000000000010111000010000101;
assign LUT_3[25609] = 32'b00000000000000011101101101100010;
assign LUT_3[25610] = 32'b00000000000000011001001001101001;
assign LUT_3[25611] = 32'b00000000000000011111110101000110;
assign LUT_3[25612] = 32'b00000000000000010100001111111011;
assign LUT_3[25613] = 32'b00000000000000011010111011011000;
assign LUT_3[25614] = 32'b00000000000000010110010111011111;
assign LUT_3[25615] = 32'b00000000000000011101000010111100;
assign LUT_3[25616] = 32'b00000000000000010100111100000010;
assign LUT_3[25617] = 32'b00000000000000011011100111011111;
assign LUT_3[25618] = 32'b00000000000000010111000011100110;
assign LUT_3[25619] = 32'b00000000000000011101101111000011;
assign LUT_3[25620] = 32'b00000000000000010010001001111000;
assign LUT_3[25621] = 32'b00000000000000011000110101010101;
assign LUT_3[25622] = 32'b00000000000000010100010001011100;
assign LUT_3[25623] = 32'b00000000000000011010111100111001;
assign LUT_3[25624] = 32'b00000000000000011010010101001000;
assign LUT_3[25625] = 32'b00000000000000100001000000100101;
assign LUT_3[25626] = 32'b00000000000000011100011100101100;
assign LUT_3[25627] = 32'b00000000000000100011001000001001;
assign LUT_3[25628] = 32'b00000000000000010111100010111110;
assign LUT_3[25629] = 32'b00000000000000011110001110011011;
assign LUT_3[25630] = 32'b00000000000000011001101010100010;
assign LUT_3[25631] = 32'b00000000000000100000010101111111;
assign LUT_3[25632] = 32'b00000000000000010010110111011111;
assign LUT_3[25633] = 32'b00000000000000011001100010111100;
assign LUT_3[25634] = 32'b00000000000000010100111111000011;
assign LUT_3[25635] = 32'b00000000000000011011101010100000;
assign LUT_3[25636] = 32'b00000000000000010000000101010101;
assign LUT_3[25637] = 32'b00000000000000010110110000110010;
assign LUT_3[25638] = 32'b00000000000000010010001100111001;
assign LUT_3[25639] = 32'b00000000000000011000111000010110;
assign LUT_3[25640] = 32'b00000000000000011000010000100101;
assign LUT_3[25641] = 32'b00000000000000011110111100000010;
assign LUT_3[25642] = 32'b00000000000000011010011000001001;
assign LUT_3[25643] = 32'b00000000000000100001000011100110;
assign LUT_3[25644] = 32'b00000000000000010101011110011011;
assign LUT_3[25645] = 32'b00000000000000011100001001111000;
assign LUT_3[25646] = 32'b00000000000000010111100101111111;
assign LUT_3[25647] = 32'b00000000000000011110010001011100;
assign LUT_3[25648] = 32'b00000000000000010110001010100010;
assign LUT_3[25649] = 32'b00000000000000011100110101111111;
assign LUT_3[25650] = 32'b00000000000000011000010010000110;
assign LUT_3[25651] = 32'b00000000000000011110111101100011;
assign LUT_3[25652] = 32'b00000000000000010011011000011000;
assign LUT_3[25653] = 32'b00000000000000011010000011110101;
assign LUT_3[25654] = 32'b00000000000000010101011111111100;
assign LUT_3[25655] = 32'b00000000000000011100001011011001;
assign LUT_3[25656] = 32'b00000000000000011011100011101000;
assign LUT_3[25657] = 32'b00000000000000100010001111000101;
assign LUT_3[25658] = 32'b00000000000000011101101011001100;
assign LUT_3[25659] = 32'b00000000000000100100010110101001;
assign LUT_3[25660] = 32'b00000000000000011000110001011110;
assign LUT_3[25661] = 32'b00000000000000011111011100111011;
assign LUT_3[25662] = 32'b00000000000000011010111001000010;
assign LUT_3[25663] = 32'b00000000000000100001100100011111;
assign LUT_3[25664] = 32'b00000000000000010001100001101010;
assign LUT_3[25665] = 32'b00000000000000011000001101000111;
assign LUT_3[25666] = 32'b00000000000000010011101001001110;
assign LUT_3[25667] = 32'b00000000000000011010010100101011;
assign LUT_3[25668] = 32'b00000000000000001110101111100000;
assign LUT_3[25669] = 32'b00000000000000010101011010111101;
assign LUT_3[25670] = 32'b00000000000000010000110111000100;
assign LUT_3[25671] = 32'b00000000000000010111100010100001;
assign LUT_3[25672] = 32'b00000000000000010110111010110000;
assign LUT_3[25673] = 32'b00000000000000011101100110001101;
assign LUT_3[25674] = 32'b00000000000000011001000010010100;
assign LUT_3[25675] = 32'b00000000000000011111101101110001;
assign LUT_3[25676] = 32'b00000000000000010100001000100110;
assign LUT_3[25677] = 32'b00000000000000011010110100000011;
assign LUT_3[25678] = 32'b00000000000000010110010000001010;
assign LUT_3[25679] = 32'b00000000000000011100111011100111;
assign LUT_3[25680] = 32'b00000000000000010100110100101101;
assign LUT_3[25681] = 32'b00000000000000011011100000001010;
assign LUT_3[25682] = 32'b00000000000000010110111100010001;
assign LUT_3[25683] = 32'b00000000000000011101100111101110;
assign LUT_3[25684] = 32'b00000000000000010010000010100011;
assign LUT_3[25685] = 32'b00000000000000011000101110000000;
assign LUT_3[25686] = 32'b00000000000000010100001010000111;
assign LUT_3[25687] = 32'b00000000000000011010110101100100;
assign LUT_3[25688] = 32'b00000000000000011010001101110011;
assign LUT_3[25689] = 32'b00000000000000100000111001010000;
assign LUT_3[25690] = 32'b00000000000000011100010101010111;
assign LUT_3[25691] = 32'b00000000000000100011000000110100;
assign LUT_3[25692] = 32'b00000000000000010111011011101001;
assign LUT_3[25693] = 32'b00000000000000011110000111000110;
assign LUT_3[25694] = 32'b00000000000000011001100011001101;
assign LUT_3[25695] = 32'b00000000000000100000001110101010;
assign LUT_3[25696] = 32'b00000000000000010010110000001010;
assign LUT_3[25697] = 32'b00000000000000011001011011100111;
assign LUT_3[25698] = 32'b00000000000000010100110111101110;
assign LUT_3[25699] = 32'b00000000000000011011100011001011;
assign LUT_3[25700] = 32'b00000000000000001111111110000000;
assign LUT_3[25701] = 32'b00000000000000010110101001011101;
assign LUT_3[25702] = 32'b00000000000000010010000101100100;
assign LUT_3[25703] = 32'b00000000000000011000110001000001;
assign LUT_3[25704] = 32'b00000000000000011000001001010000;
assign LUT_3[25705] = 32'b00000000000000011110110100101101;
assign LUT_3[25706] = 32'b00000000000000011010010000110100;
assign LUT_3[25707] = 32'b00000000000000100000111100010001;
assign LUT_3[25708] = 32'b00000000000000010101010111000110;
assign LUT_3[25709] = 32'b00000000000000011100000010100011;
assign LUT_3[25710] = 32'b00000000000000010111011110101010;
assign LUT_3[25711] = 32'b00000000000000011110001010000111;
assign LUT_3[25712] = 32'b00000000000000010110000011001101;
assign LUT_3[25713] = 32'b00000000000000011100101110101010;
assign LUT_3[25714] = 32'b00000000000000011000001010110001;
assign LUT_3[25715] = 32'b00000000000000011110110110001110;
assign LUT_3[25716] = 32'b00000000000000010011010001000011;
assign LUT_3[25717] = 32'b00000000000000011001111100100000;
assign LUT_3[25718] = 32'b00000000000000010101011000100111;
assign LUT_3[25719] = 32'b00000000000000011100000100000100;
assign LUT_3[25720] = 32'b00000000000000011011011100010011;
assign LUT_3[25721] = 32'b00000000000000100010000111110000;
assign LUT_3[25722] = 32'b00000000000000011101100011110111;
assign LUT_3[25723] = 32'b00000000000000100100001111010100;
assign LUT_3[25724] = 32'b00000000000000011000101010001001;
assign LUT_3[25725] = 32'b00000000000000011111010101100110;
assign LUT_3[25726] = 32'b00000000000000011010110001101101;
assign LUT_3[25727] = 32'b00000000000000100001011101001010;
assign LUT_3[25728] = 32'b00000000000000010011110011111101;
assign LUT_3[25729] = 32'b00000000000000011010011111011010;
assign LUT_3[25730] = 32'b00000000000000010101111011100001;
assign LUT_3[25731] = 32'b00000000000000011100100110111110;
assign LUT_3[25732] = 32'b00000000000000010001000001110011;
assign LUT_3[25733] = 32'b00000000000000010111101101010000;
assign LUT_3[25734] = 32'b00000000000000010011001001010111;
assign LUT_3[25735] = 32'b00000000000000011001110100110100;
assign LUT_3[25736] = 32'b00000000000000011001001101000011;
assign LUT_3[25737] = 32'b00000000000000011111111000100000;
assign LUT_3[25738] = 32'b00000000000000011011010100100111;
assign LUT_3[25739] = 32'b00000000000000100010000000000100;
assign LUT_3[25740] = 32'b00000000000000010110011010111001;
assign LUT_3[25741] = 32'b00000000000000011101000110010110;
assign LUT_3[25742] = 32'b00000000000000011000100010011101;
assign LUT_3[25743] = 32'b00000000000000011111001101111010;
assign LUT_3[25744] = 32'b00000000000000010111000111000000;
assign LUT_3[25745] = 32'b00000000000000011101110010011101;
assign LUT_3[25746] = 32'b00000000000000011001001110100100;
assign LUT_3[25747] = 32'b00000000000000011111111010000001;
assign LUT_3[25748] = 32'b00000000000000010100010100110110;
assign LUT_3[25749] = 32'b00000000000000011011000000010011;
assign LUT_3[25750] = 32'b00000000000000010110011100011010;
assign LUT_3[25751] = 32'b00000000000000011101000111110111;
assign LUT_3[25752] = 32'b00000000000000011100100000000110;
assign LUT_3[25753] = 32'b00000000000000100011001011100011;
assign LUT_3[25754] = 32'b00000000000000011110100111101010;
assign LUT_3[25755] = 32'b00000000000000100101010011000111;
assign LUT_3[25756] = 32'b00000000000000011001101101111100;
assign LUT_3[25757] = 32'b00000000000000100000011001011001;
assign LUT_3[25758] = 32'b00000000000000011011110101100000;
assign LUT_3[25759] = 32'b00000000000000100010100000111101;
assign LUT_3[25760] = 32'b00000000000000010101000010011101;
assign LUT_3[25761] = 32'b00000000000000011011101101111010;
assign LUT_3[25762] = 32'b00000000000000010111001010000001;
assign LUT_3[25763] = 32'b00000000000000011101110101011110;
assign LUT_3[25764] = 32'b00000000000000010010010000010011;
assign LUT_3[25765] = 32'b00000000000000011000111011110000;
assign LUT_3[25766] = 32'b00000000000000010100010111110111;
assign LUT_3[25767] = 32'b00000000000000011011000011010100;
assign LUT_3[25768] = 32'b00000000000000011010011011100011;
assign LUT_3[25769] = 32'b00000000000000100001000111000000;
assign LUT_3[25770] = 32'b00000000000000011100100011000111;
assign LUT_3[25771] = 32'b00000000000000100011001110100100;
assign LUT_3[25772] = 32'b00000000000000010111101001011001;
assign LUT_3[25773] = 32'b00000000000000011110010100110110;
assign LUT_3[25774] = 32'b00000000000000011001110000111101;
assign LUT_3[25775] = 32'b00000000000000100000011100011010;
assign LUT_3[25776] = 32'b00000000000000011000010101100000;
assign LUT_3[25777] = 32'b00000000000000011111000000111101;
assign LUT_3[25778] = 32'b00000000000000011010011101000100;
assign LUT_3[25779] = 32'b00000000000000100001001000100001;
assign LUT_3[25780] = 32'b00000000000000010101100011010110;
assign LUT_3[25781] = 32'b00000000000000011100001110110011;
assign LUT_3[25782] = 32'b00000000000000010111101010111010;
assign LUT_3[25783] = 32'b00000000000000011110010110010111;
assign LUT_3[25784] = 32'b00000000000000011101101110100110;
assign LUT_3[25785] = 32'b00000000000000100100011010000011;
assign LUT_3[25786] = 32'b00000000000000011111110110001010;
assign LUT_3[25787] = 32'b00000000000000100110100001100111;
assign LUT_3[25788] = 32'b00000000000000011010111100011100;
assign LUT_3[25789] = 32'b00000000000000100001100111111001;
assign LUT_3[25790] = 32'b00000000000000011101000100000000;
assign LUT_3[25791] = 32'b00000000000000100011101111011101;
assign LUT_3[25792] = 32'b00000000000000010011101100101000;
assign LUT_3[25793] = 32'b00000000000000011010011000000101;
assign LUT_3[25794] = 32'b00000000000000010101110100001100;
assign LUT_3[25795] = 32'b00000000000000011100011111101001;
assign LUT_3[25796] = 32'b00000000000000010000111010011110;
assign LUT_3[25797] = 32'b00000000000000010111100101111011;
assign LUT_3[25798] = 32'b00000000000000010011000010000010;
assign LUT_3[25799] = 32'b00000000000000011001101101011111;
assign LUT_3[25800] = 32'b00000000000000011001000101101110;
assign LUT_3[25801] = 32'b00000000000000011111110001001011;
assign LUT_3[25802] = 32'b00000000000000011011001101010010;
assign LUT_3[25803] = 32'b00000000000000100001111000101111;
assign LUT_3[25804] = 32'b00000000000000010110010011100100;
assign LUT_3[25805] = 32'b00000000000000011100111111000001;
assign LUT_3[25806] = 32'b00000000000000011000011011001000;
assign LUT_3[25807] = 32'b00000000000000011111000110100101;
assign LUT_3[25808] = 32'b00000000000000010110111111101011;
assign LUT_3[25809] = 32'b00000000000000011101101011001000;
assign LUT_3[25810] = 32'b00000000000000011001000111001111;
assign LUT_3[25811] = 32'b00000000000000011111110010101100;
assign LUT_3[25812] = 32'b00000000000000010100001101100001;
assign LUT_3[25813] = 32'b00000000000000011010111000111110;
assign LUT_3[25814] = 32'b00000000000000010110010101000101;
assign LUT_3[25815] = 32'b00000000000000011101000000100010;
assign LUT_3[25816] = 32'b00000000000000011100011000110001;
assign LUT_3[25817] = 32'b00000000000000100011000100001110;
assign LUT_3[25818] = 32'b00000000000000011110100000010101;
assign LUT_3[25819] = 32'b00000000000000100101001011110010;
assign LUT_3[25820] = 32'b00000000000000011001100110100111;
assign LUT_3[25821] = 32'b00000000000000100000010010000100;
assign LUT_3[25822] = 32'b00000000000000011011101110001011;
assign LUT_3[25823] = 32'b00000000000000100010011001101000;
assign LUT_3[25824] = 32'b00000000000000010100111011001000;
assign LUT_3[25825] = 32'b00000000000000011011100110100101;
assign LUT_3[25826] = 32'b00000000000000010111000010101100;
assign LUT_3[25827] = 32'b00000000000000011101101110001001;
assign LUT_3[25828] = 32'b00000000000000010010001000111110;
assign LUT_3[25829] = 32'b00000000000000011000110100011011;
assign LUT_3[25830] = 32'b00000000000000010100010000100010;
assign LUT_3[25831] = 32'b00000000000000011010111011111111;
assign LUT_3[25832] = 32'b00000000000000011010010100001110;
assign LUT_3[25833] = 32'b00000000000000100000111111101011;
assign LUT_3[25834] = 32'b00000000000000011100011011110010;
assign LUT_3[25835] = 32'b00000000000000100011000111001111;
assign LUT_3[25836] = 32'b00000000000000010111100010000100;
assign LUT_3[25837] = 32'b00000000000000011110001101100001;
assign LUT_3[25838] = 32'b00000000000000011001101001101000;
assign LUT_3[25839] = 32'b00000000000000100000010101000101;
assign LUT_3[25840] = 32'b00000000000000011000001110001011;
assign LUT_3[25841] = 32'b00000000000000011110111001101000;
assign LUT_3[25842] = 32'b00000000000000011010010101101111;
assign LUT_3[25843] = 32'b00000000000000100001000001001100;
assign LUT_3[25844] = 32'b00000000000000010101011100000001;
assign LUT_3[25845] = 32'b00000000000000011100000111011110;
assign LUT_3[25846] = 32'b00000000000000010111100011100101;
assign LUT_3[25847] = 32'b00000000000000011110001111000010;
assign LUT_3[25848] = 32'b00000000000000011101100111010001;
assign LUT_3[25849] = 32'b00000000000000100100010010101110;
assign LUT_3[25850] = 32'b00000000000000011111101110110101;
assign LUT_3[25851] = 32'b00000000000000100110011010010010;
assign LUT_3[25852] = 32'b00000000000000011010110101000111;
assign LUT_3[25853] = 32'b00000000000000100001100000100100;
assign LUT_3[25854] = 32'b00000000000000011100111100101011;
assign LUT_3[25855] = 32'b00000000000000100011101000001000;
assign LUT_3[25856] = 32'b00000000000000001101111000100000;
assign LUT_3[25857] = 32'b00000000000000010100100011111101;
assign LUT_3[25858] = 32'b00000000000000010000000000000100;
assign LUT_3[25859] = 32'b00000000000000010110101011100001;
assign LUT_3[25860] = 32'b00000000000000001011000110010110;
assign LUT_3[25861] = 32'b00000000000000010001110001110011;
assign LUT_3[25862] = 32'b00000000000000001101001101111010;
assign LUT_3[25863] = 32'b00000000000000010011111001010111;
assign LUT_3[25864] = 32'b00000000000000010011010001100110;
assign LUT_3[25865] = 32'b00000000000000011001111101000011;
assign LUT_3[25866] = 32'b00000000000000010101011001001010;
assign LUT_3[25867] = 32'b00000000000000011100000100100111;
assign LUT_3[25868] = 32'b00000000000000010000011111011100;
assign LUT_3[25869] = 32'b00000000000000010111001010111001;
assign LUT_3[25870] = 32'b00000000000000010010100111000000;
assign LUT_3[25871] = 32'b00000000000000011001010010011101;
assign LUT_3[25872] = 32'b00000000000000010001001011100011;
assign LUT_3[25873] = 32'b00000000000000010111110111000000;
assign LUT_3[25874] = 32'b00000000000000010011010011000111;
assign LUT_3[25875] = 32'b00000000000000011001111110100100;
assign LUT_3[25876] = 32'b00000000000000001110011001011001;
assign LUT_3[25877] = 32'b00000000000000010101000100110110;
assign LUT_3[25878] = 32'b00000000000000010000100000111101;
assign LUT_3[25879] = 32'b00000000000000010111001100011010;
assign LUT_3[25880] = 32'b00000000000000010110100100101001;
assign LUT_3[25881] = 32'b00000000000000011101010000000110;
assign LUT_3[25882] = 32'b00000000000000011000101100001101;
assign LUT_3[25883] = 32'b00000000000000011111010111101010;
assign LUT_3[25884] = 32'b00000000000000010011110010011111;
assign LUT_3[25885] = 32'b00000000000000011010011101111100;
assign LUT_3[25886] = 32'b00000000000000010101111010000011;
assign LUT_3[25887] = 32'b00000000000000011100100101100000;
assign LUT_3[25888] = 32'b00000000000000001111000111000000;
assign LUT_3[25889] = 32'b00000000000000010101110010011101;
assign LUT_3[25890] = 32'b00000000000000010001001110100100;
assign LUT_3[25891] = 32'b00000000000000010111111010000001;
assign LUT_3[25892] = 32'b00000000000000001100010100110110;
assign LUT_3[25893] = 32'b00000000000000010011000000010011;
assign LUT_3[25894] = 32'b00000000000000001110011100011010;
assign LUT_3[25895] = 32'b00000000000000010101000111110111;
assign LUT_3[25896] = 32'b00000000000000010100100000000110;
assign LUT_3[25897] = 32'b00000000000000011011001011100011;
assign LUT_3[25898] = 32'b00000000000000010110100111101010;
assign LUT_3[25899] = 32'b00000000000000011101010011000111;
assign LUT_3[25900] = 32'b00000000000000010001101101111100;
assign LUT_3[25901] = 32'b00000000000000011000011001011001;
assign LUT_3[25902] = 32'b00000000000000010011110101100000;
assign LUT_3[25903] = 32'b00000000000000011010100000111101;
assign LUT_3[25904] = 32'b00000000000000010010011010000011;
assign LUT_3[25905] = 32'b00000000000000011001000101100000;
assign LUT_3[25906] = 32'b00000000000000010100100001100111;
assign LUT_3[25907] = 32'b00000000000000011011001101000100;
assign LUT_3[25908] = 32'b00000000000000001111100111111001;
assign LUT_3[25909] = 32'b00000000000000010110010011010110;
assign LUT_3[25910] = 32'b00000000000000010001101111011101;
assign LUT_3[25911] = 32'b00000000000000011000011010111010;
assign LUT_3[25912] = 32'b00000000000000010111110011001001;
assign LUT_3[25913] = 32'b00000000000000011110011110100110;
assign LUT_3[25914] = 32'b00000000000000011001111010101101;
assign LUT_3[25915] = 32'b00000000000000100000100110001010;
assign LUT_3[25916] = 32'b00000000000000010101000000111111;
assign LUT_3[25917] = 32'b00000000000000011011101100011100;
assign LUT_3[25918] = 32'b00000000000000010111001000100011;
assign LUT_3[25919] = 32'b00000000000000011101110100000000;
assign LUT_3[25920] = 32'b00000000000000001101110001001011;
assign LUT_3[25921] = 32'b00000000000000010100011100101000;
assign LUT_3[25922] = 32'b00000000000000001111111000101111;
assign LUT_3[25923] = 32'b00000000000000010110100100001100;
assign LUT_3[25924] = 32'b00000000000000001010111111000001;
assign LUT_3[25925] = 32'b00000000000000010001101010011110;
assign LUT_3[25926] = 32'b00000000000000001101000110100101;
assign LUT_3[25927] = 32'b00000000000000010011110010000010;
assign LUT_3[25928] = 32'b00000000000000010011001010010001;
assign LUT_3[25929] = 32'b00000000000000011001110101101110;
assign LUT_3[25930] = 32'b00000000000000010101010001110101;
assign LUT_3[25931] = 32'b00000000000000011011111101010010;
assign LUT_3[25932] = 32'b00000000000000010000011000000111;
assign LUT_3[25933] = 32'b00000000000000010111000011100100;
assign LUT_3[25934] = 32'b00000000000000010010011111101011;
assign LUT_3[25935] = 32'b00000000000000011001001011001000;
assign LUT_3[25936] = 32'b00000000000000010001000100001110;
assign LUT_3[25937] = 32'b00000000000000010111101111101011;
assign LUT_3[25938] = 32'b00000000000000010011001011110010;
assign LUT_3[25939] = 32'b00000000000000011001110111001111;
assign LUT_3[25940] = 32'b00000000000000001110010010000100;
assign LUT_3[25941] = 32'b00000000000000010100111101100001;
assign LUT_3[25942] = 32'b00000000000000010000011001101000;
assign LUT_3[25943] = 32'b00000000000000010111000101000101;
assign LUT_3[25944] = 32'b00000000000000010110011101010100;
assign LUT_3[25945] = 32'b00000000000000011101001000110001;
assign LUT_3[25946] = 32'b00000000000000011000100100111000;
assign LUT_3[25947] = 32'b00000000000000011111010000010101;
assign LUT_3[25948] = 32'b00000000000000010011101011001010;
assign LUT_3[25949] = 32'b00000000000000011010010110100111;
assign LUT_3[25950] = 32'b00000000000000010101110010101110;
assign LUT_3[25951] = 32'b00000000000000011100011110001011;
assign LUT_3[25952] = 32'b00000000000000001110111111101011;
assign LUT_3[25953] = 32'b00000000000000010101101011001000;
assign LUT_3[25954] = 32'b00000000000000010001000111001111;
assign LUT_3[25955] = 32'b00000000000000010111110010101100;
assign LUT_3[25956] = 32'b00000000000000001100001101100001;
assign LUT_3[25957] = 32'b00000000000000010010111000111110;
assign LUT_3[25958] = 32'b00000000000000001110010101000101;
assign LUT_3[25959] = 32'b00000000000000010101000000100010;
assign LUT_3[25960] = 32'b00000000000000010100011000110001;
assign LUT_3[25961] = 32'b00000000000000011011000100001110;
assign LUT_3[25962] = 32'b00000000000000010110100000010101;
assign LUT_3[25963] = 32'b00000000000000011101001011110010;
assign LUT_3[25964] = 32'b00000000000000010001100110100111;
assign LUT_3[25965] = 32'b00000000000000011000010010000100;
assign LUT_3[25966] = 32'b00000000000000010011101110001011;
assign LUT_3[25967] = 32'b00000000000000011010011001101000;
assign LUT_3[25968] = 32'b00000000000000010010010010101110;
assign LUT_3[25969] = 32'b00000000000000011000111110001011;
assign LUT_3[25970] = 32'b00000000000000010100011010010010;
assign LUT_3[25971] = 32'b00000000000000011011000101101111;
assign LUT_3[25972] = 32'b00000000000000001111100000100100;
assign LUT_3[25973] = 32'b00000000000000010110001100000001;
assign LUT_3[25974] = 32'b00000000000000010001101000001000;
assign LUT_3[25975] = 32'b00000000000000011000010011100101;
assign LUT_3[25976] = 32'b00000000000000010111101011110100;
assign LUT_3[25977] = 32'b00000000000000011110010111010001;
assign LUT_3[25978] = 32'b00000000000000011001110011011000;
assign LUT_3[25979] = 32'b00000000000000100000011110110101;
assign LUT_3[25980] = 32'b00000000000000010100111001101010;
assign LUT_3[25981] = 32'b00000000000000011011100101000111;
assign LUT_3[25982] = 32'b00000000000000010111000001001110;
assign LUT_3[25983] = 32'b00000000000000011101101100101011;
assign LUT_3[25984] = 32'b00000000000000010000000011011110;
assign LUT_3[25985] = 32'b00000000000000010110101110111011;
assign LUT_3[25986] = 32'b00000000000000010010001011000010;
assign LUT_3[25987] = 32'b00000000000000011000110110011111;
assign LUT_3[25988] = 32'b00000000000000001101010001010100;
assign LUT_3[25989] = 32'b00000000000000010011111100110001;
assign LUT_3[25990] = 32'b00000000000000001111011000111000;
assign LUT_3[25991] = 32'b00000000000000010110000100010101;
assign LUT_3[25992] = 32'b00000000000000010101011100100100;
assign LUT_3[25993] = 32'b00000000000000011100001000000001;
assign LUT_3[25994] = 32'b00000000000000010111100100001000;
assign LUT_3[25995] = 32'b00000000000000011110001111100101;
assign LUT_3[25996] = 32'b00000000000000010010101010011010;
assign LUT_3[25997] = 32'b00000000000000011001010101110111;
assign LUT_3[25998] = 32'b00000000000000010100110001111110;
assign LUT_3[25999] = 32'b00000000000000011011011101011011;
assign LUT_3[26000] = 32'b00000000000000010011010110100001;
assign LUT_3[26001] = 32'b00000000000000011010000001111110;
assign LUT_3[26002] = 32'b00000000000000010101011110000101;
assign LUT_3[26003] = 32'b00000000000000011100001001100010;
assign LUT_3[26004] = 32'b00000000000000010000100100010111;
assign LUT_3[26005] = 32'b00000000000000010111001111110100;
assign LUT_3[26006] = 32'b00000000000000010010101011111011;
assign LUT_3[26007] = 32'b00000000000000011001010111011000;
assign LUT_3[26008] = 32'b00000000000000011000101111100111;
assign LUT_3[26009] = 32'b00000000000000011111011011000100;
assign LUT_3[26010] = 32'b00000000000000011010110111001011;
assign LUT_3[26011] = 32'b00000000000000100001100010101000;
assign LUT_3[26012] = 32'b00000000000000010101111101011101;
assign LUT_3[26013] = 32'b00000000000000011100101000111010;
assign LUT_3[26014] = 32'b00000000000000011000000101000001;
assign LUT_3[26015] = 32'b00000000000000011110110000011110;
assign LUT_3[26016] = 32'b00000000000000010001010001111110;
assign LUT_3[26017] = 32'b00000000000000010111111101011011;
assign LUT_3[26018] = 32'b00000000000000010011011001100010;
assign LUT_3[26019] = 32'b00000000000000011010000100111111;
assign LUT_3[26020] = 32'b00000000000000001110011111110100;
assign LUT_3[26021] = 32'b00000000000000010101001011010001;
assign LUT_3[26022] = 32'b00000000000000010000100111011000;
assign LUT_3[26023] = 32'b00000000000000010111010010110101;
assign LUT_3[26024] = 32'b00000000000000010110101011000100;
assign LUT_3[26025] = 32'b00000000000000011101010110100001;
assign LUT_3[26026] = 32'b00000000000000011000110010101000;
assign LUT_3[26027] = 32'b00000000000000011111011110000101;
assign LUT_3[26028] = 32'b00000000000000010011111000111010;
assign LUT_3[26029] = 32'b00000000000000011010100100010111;
assign LUT_3[26030] = 32'b00000000000000010110000000011110;
assign LUT_3[26031] = 32'b00000000000000011100101011111011;
assign LUT_3[26032] = 32'b00000000000000010100100101000001;
assign LUT_3[26033] = 32'b00000000000000011011010000011110;
assign LUT_3[26034] = 32'b00000000000000010110101100100101;
assign LUT_3[26035] = 32'b00000000000000011101011000000010;
assign LUT_3[26036] = 32'b00000000000000010001110010110111;
assign LUT_3[26037] = 32'b00000000000000011000011110010100;
assign LUT_3[26038] = 32'b00000000000000010011111010011011;
assign LUT_3[26039] = 32'b00000000000000011010100101111000;
assign LUT_3[26040] = 32'b00000000000000011001111110000111;
assign LUT_3[26041] = 32'b00000000000000100000101001100100;
assign LUT_3[26042] = 32'b00000000000000011100000101101011;
assign LUT_3[26043] = 32'b00000000000000100010110001001000;
assign LUT_3[26044] = 32'b00000000000000010111001011111101;
assign LUT_3[26045] = 32'b00000000000000011101110111011010;
assign LUT_3[26046] = 32'b00000000000000011001010011100001;
assign LUT_3[26047] = 32'b00000000000000011111111110111110;
assign LUT_3[26048] = 32'b00000000000000001111111100001001;
assign LUT_3[26049] = 32'b00000000000000010110100111100110;
assign LUT_3[26050] = 32'b00000000000000010010000011101101;
assign LUT_3[26051] = 32'b00000000000000011000101111001010;
assign LUT_3[26052] = 32'b00000000000000001101001001111111;
assign LUT_3[26053] = 32'b00000000000000010011110101011100;
assign LUT_3[26054] = 32'b00000000000000001111010001100011;
assign LUT_3[26055] = 32'b00000000000000010101111101000000;
assign LUT_3[26056] = 32'b00000000000000010101010101001111;
assign LUT_3[26057] = 32'b00000000000000011100000000101100;
assign LUT_3[26058] = 32'b00000000000000010111011100110011;
assign LUT_3[26059] = 32'b00000000000000011110001000010000;
assign LUT_3[26060] = 32'b00000000000000010010100011000101;
assign LUT_3[26061] = 32'b00000000000000011001001110100010;
assign LUT_3[26062] = 32'b00000000000000010100101010101001;
assign LUT_3[26063] = 32'b00000000000000011011010110000110;
assign LUT_3[26064] = 32'b00000000000000010011001111001100;
assign LUT_3[26065] = 32'b00000000000000011001111010101001;
assign LUT_3[26066] = 32'b00000000000000010101010110110000;
assign LUT_3[26067] = 32'b00000000000000011100000010001101;
assign LUT_3[26068] = 32'b00000000000000010000011101000010;
assign LUT_3[26069] = 32'b00000000000000010111001000011111;
assign LUT_3[26070] = 32'b00000000000000010010100100100110;
assign LUT_3[26071] = 32'b00000000000000011001010000000011;
assign LUT_3[26072] = 32'b00000000000000011000101000010010;
assign LUT_3[26073] = 32'b00000000000000011111010011101111;
assign LUT_3[26074] = 32'b00000000000000011010101111110110;
assign LUT_3[26075] = 32'b00000000000000100001011011010011;
assign LUT_3[26076] = 32'b00000000000000010101110110001000;
assign LUT_3[26077] = 32'b00000000000000011100100001100101;
assign LUT_3[26078] = 32'b00000000000000010111111101101100;
assign LUT_3[26079] = 32'b00000000000000011110101001001001;
assign LUT_3[26080] = 32'b00000000000000010001001010101001;
assign LUT_3[26081] = 32'b00000000000000010111110110000110;
assign LUT_3[26082] = 32'b00000000000000010011010010001101;
assign LUT_3[26083] = 32'b00000000000000011001111101101010;
assign LUT_3[26084] = 32'b00000000000000001110011000011111;
assign LUT_3[26085] = 32'b00000000000000010101000011111100;
assign LUT_3[26086] = 32'b00000000000000010000100000000011;
assign LUT_3[26087] = 32'b00000000000000010111001011100000;
assign LUT_3[26088] = 32'b00000000000000010110100011101111;
assign LUT_3[26089] = 32'b00000000000000011101001111001100;
assign LUT_3[26090] = 32'b00000000000000011000101011010011;
assign LUT_3[26091] = 32'b00000000000000011111010110110000;
assign LUT_3[26092] = 32'b00000000000000010011110001100101;
assign LUT_3[26093] = 32'b00000000000000011010011101000010;
assign LUT_3[26094] = 32'b00000000000000010101111001001001;
assign LUT_3[26095] = 32'b00000000000000011100100100100110;
assign LUT_3[26096] = 32'b00000000000000010100011101101100;
assign LUT_3[26097] = 32'b00000000000000011011001001001001;
assign LUT_3[26098] = 32'b00000000000000010110100101010000;
assign LUT_3[26099] = 32'b00000000000000011101010000101101;
assign LUT_3[26100] = 32'b00000000000000010001101011100010;
assign LUT_3[26101] = 32'b00000000000000011000010110111111;
assign LUT_3[26102] = 32'b00000000000000010011110011000110;
assign LUT_3[26103] = 32'b00000000000000011010011110100011;
assign LUT_3[26104] = 32'b00000000000000011001110110110010;
assign LUT_3[26105] = 32'b00000000000000100000100010001111;
assign LUT_3[26106] = 32'b00000000000000011011111110010110;
assign LUT_3[26107] = 32'b00000000000000100010101001110011;
assign LUT_3[26108] = 32'b00000000000000010111000100101000;
assign LUT_3[26109] = 32'b00000000000000011101110000000101;
assign LUT_3[26110] = 32'b00000000000000011001001100001100;
assign LUT_3[26111] = 32'b00000000000000011111110111101001;
assign LUT_3[26112] = 32'b00000000000000010100111110001011;
assign LUT_3[26113] = 32'b00000000000000011011101001101000;
assign LUT_3[26114] = 32'b00000000000000010111000101101111;
assign LUT_3[26115] = 32'b00000000000000011101110001001100;
assign LUT_3[26116] = 32'b00000000000000010010001100000001;
assign LUT_3[26117] = 32'b00000000000000011000110111011110;
assign LUT_3[26118] = 32'b00000000000000010100010011100101;
assign LUT_3[26119] = 32'b00000000000000011010111111000010;
assign LUT_3[26120] = 32'b00000000000000011010010111010001;
assign LUT_3[26121] = 32'b00000000000000100001000010101110;
assign LUT_3[26122] = 32'b00000000000000011100011110110101;
assign LUT_3[26123] = 32'b00000000000000100011001010010010;
assign LUT_3[26124] = 32'b00000000000000010111100101000111;
assign LUT_3[26125] = 32'b00000000000000011110010000100100;
assign LUT_3[26126] = 32'b00000000000000011001101100101011;
assign LUT_3[26127] = 32'b00000000000000100000011000001000;
assign LUT_3[26128] = 32'b00000000000000011000010001001110;
assign LUT_3[26129] = 32'b00000000000000011110111100101011;
assign LUT_3[26130] = 32'b00000000000000011010011000110010;
assign LUT_3[26131] = 32'b00000000000000100001000100001111;
assign LUT_3[26132] = 32'b00000000000000010101011111000100;
assign LUT_3[26133] = 32'b00000000000000011100001010100001;
assign LUT_3[26134] = 32'b00000000000000010111100110101000;
assign LUT_3[26135] = 32'b00000000000000011110010010000101;
assign LUT_3[26136] = 32'b00000000000000011101101010010100;
assign LUT_3[26137] = 32'b00000000000000100100010101110001;
assign LUT_3[26138] = 32'b00000000000000011111110001111000;
assign LUT_3[26139] = 32'b00000000000000100110011101010101;
assign LUT_3[26140] = 32'b00000000000000011010111000001010;
assign LUT_3[26141] = 32'b00000000000000100001100011100111;
assign LUT_3[26142] = 32'b00000000000000011100111111101110;
assign LUT_3[26143] = 32'b00000000000000100011101011001011;
assign LUT_3[26144] = 32'b00000000000000010110001100101011;
assign LUT_3[26145] = 32'b00000000000000011100111000001000;
assign LUT_3[26146] = 32'b00000000000000011000010100001111;
assign LUT_3[26147] = 32'b00000000000000011110111111101100;
assign LUT_3[26148] = 32'b00000000000000010011011010100001;
assign LUT_3[26149] = 32'b00000000000000011010000101111110;
assign LUT_3[26150] = 32'b00000000000000010101100010000101;
assign LUT_3[26151] = 32'b00000000000000011100001101100010;
assign LUT_3[26152] = 32'b00000000000000011011100101110001;
assign LUT_3[26153] = 32'b00000000000000100010010001001110;
assign LUT_3[26154] = 32'b00000000000000011101101101010101;
assign LUT_3[26155] = 32'b00000000000000100100011000110010;
assign LUT_3[26156] = 32'b00000000000000011000110011100111;
assign LUT_3[26157] = 32'b00000000000000011111011111000100;
assign LUT_3[26158] = 32'b00000000000000011010111011001011;
assign LUT_3[26159] = 32'b00000000000000100001100110101000;
assign LUT_3[26160] = 32'b00000000000000011001011111101110;
assign LUT_3[26161] = 32'b00000000000000100000001011001011;
assign LUT_3[26162] = 32'b00000000000000011011100111010010;
assign LUT_3[26163] = 32'b00000000000000100010010010101111;
assign LUT_3[26164] = 32'b00000000000000010110101101100100;
assign LUT_3[26165] = 32'b00000000000000011101011001000001;
assign LUT_3[26166] = 32'b00000000000000011000110101001000;
assign LUT_3[26167] = 32'b00000000000000011111100000100101;
assign LUT_3[26168] = 32'b00000000000000011110111000110100;
assign LUT_3[26169] = 32'b00000000000000100101100100010001;
assign LUT_3[26170] = 32'b00000000000000100001000000011000;
assign LUT_3[26171] = 32'b00000000000000100111101011110101;
assign LUT_3[26172] = 32'b00000000000000011100000110101010;
assign LUT_3[26173] = 32'b00000000000000100010110010000111;
assign LUT_3[26174] = 32'b00000000000000011110001110001110;
assign LUT_3[26175] = 32'b00000000000000100100111001101011;
assign LUT_3[26176] = 32'b00000000000000010100110110110110;
assign LUT_3[26177] = 32'b00000000000000011011100010010011;
assign LUT_3[26178] = 32'b00000000000000010110111110011010;
assign LUT_3[26179] = 32'b00000000000000011101101001110111;
assign LUT_3[26180] = 32'b00000000000000010010000100101100;
assign LUT_3[26181] = 32'b00000000000000011000110000001001;
assign LUT_3[26182] = 32'b00000000000000010100001100010000;
assign LUT_3[26183] = 32'b00000000000000011010110111101101;
assign LUT_3[26184] = 32'b00000000000000011010001111111100;
assign LUT_3[26185] = 32'b00000000000000100000111011011001;
assign LUT_3[26186] = 32'b00000000000000011100010111100000;
assign LUT_3[26187] = 32'b00000000000000100011000010111101;
assign LUT_3[26188] = 32'b00000000000000010111011101110010;
assign LUT_3[26189] = 32'b00000000000000011110001001001111;
assign LUT_3[26190] = 32'b00000000000000011001100101010110;
assign LUT_3[26191] = 32'b00000000000000100000010000110011;
assign LUT_3[26192] = 32'b00000000000000011000001001111001;
assign LUT_3[26193] = 32'b00000000000000011110110101010110;
assign LUT_3[26194] = 32'b00000000000000011010010001011101;
assign LUT_3[26195] = 32'b00000000000000100000111100111010;
assign LUT_3[26196] = 32'b00000000000000010101010111101111;
assign LUT_3[26197] = 32'b00000000000000011100000011001100;
assign LUT_3[26198] = 32'b00000000000000010111011111010011;
assign LUT_3[26199] = 32'b00000000000000011110001010110000;
assign LUT_3[26200] = 32'b00000000000000011101100010111111;
assign LUT_3[26201] = 32'b00000000000000100100001110011100;
assign LUT_3[26202] = 32'b00000000000000011111101010100011;
assign LUT_3[26203] = 32'b00000000000000100110010110000000;
assign LUT_3[26204] = 32'b00000000000000011010110000110101;
assign LUT_3[26205] = 32'b00000000000000100001011100010010;
assign LUT_3[26206] = 32'b00000000000000011100111000011001;
assign LUT_3[26207] = 32'b00000000000000100011100011110110;
assign LUT_3[26208] = 32'b00000000000000010110000101010110;
assign LUT_3[26209] = 32'b00000000000000011100110000110011;
assign LUT_3[26210] = 32'b00000000000000011000001100111010;
assign LUT_3[26211] = 32'b00000000000000011110111000010111;
assign LUT_3[26212] = 32'b00000000000000010011010011001100;
assign LUT_3[26213] = 32'b00000000000000011001111110101001;
assign LUT_3[26214] = 32'b00000000000000010101011010110000;
assign LUT_3[26215] = 32'b00000000000000011100000110001101;
assign LUT_3[26216] = 32'b00000000000000011011011110011100;
assign LUT_3[26217] = 32'b00000000000000100010001001111001;
assign LUT_3[26218] = 32'b00000000000000011101100110000000;
assign LUT_3[26219] = 32'b00000000000000100100010001011101;
assign LUT_3[26220] = 32'b00000000000000011000101100010010;
assign LUT_3[26221] = 32'b00000000000000011111010111101111;
assign LUT_3[26222] = 32'b00000000000000011010110011110110;
assign LUT_3[26223] = 32'b00000000000000100001011111010011;
assign LUT_3[26224] = 32'b00000000000000011001011000011001;
assign LUT_3[26225] = 32'b00000000000000100000000011110110;
assign LUT_3[26226] = 32'b00000000000000011011011111111101;
assign LUT_3[26227] = 32'b00000000000000100010001011011010;
assign LUT_3[26228] = 32'b00000000000000010110100110001111;
assign LUT_3[26229] = 32'b00000000000000011101010001101100;
assign LUT_3[26230] = 32'b00000000000000011000101101110011;
assign LUT_3[26231] = 32'b00000000000000011111011001010000;
assign LUT_3[26232] = 32'b00000000000000011110110001011111;
assign LUT_3[26233] = 32'b00000000000000100101011100111100;
assign LUT_3[26234] = 32'b00000000000000100000111001000011;
assign LUT_3[26235] = 32'b00000000000000100111100100100000;
assign LUT_3[26236] = 32'b00000000000000011011111111010101;
assign LUT_3[26237] = 32'b00000000000000100010101010110010;
assign LUT_3[26238] = 32'b00000000000000011110000110111001;
assign LUT_3[26239] = 32'b00000000000000100100110010010110;
assign LUT_3[26240] = 32'b00000000000000010111001001001001;
assign LUT_3[26241] = 32'b00000000000000011101110100100110;
assign LUT_3[26242] = 32'b00000000000000011001010000101101;
assign LUT_3[26243] = 32'b00000000000000011111111100001010;
assign LUT_3[26244] = 32'b00000000000000010100010110111111;
assign LUT_3[26245] = 32'b00000000000000011011000010011100;
assign LUT_3[26246] = 32'b00000000000000010110011110100011;
assign LUT_3[26247] = 32'b00000000000000011101001010000000;
assign LUT_3[26248] = 32'b00000000000000011100100010001111;
assign LUT_3[26249] = 32'b00000000000000100011001101101100;
assign LUT_3[26250] = 32'b00000000000000011110101001110011;
assign LUT_3[26251] = 32'b00000000000000100101010101010000;
assign LUT_3[26252] = 32'b00000000000000011001110000000101;
assign LUT_3[26253] = 32'b00000000000000100000011011100010;
assign LUT_3[26254] = 32'b00000000000000011011110111101001;
assign LUT_3[26255] = 32'b00000000000000100010100011000110;
assign LUT_3[26256] = 32'b00000000000000011010011100001100;
assign LUT_3[26257] = 32'b00000000000000100001000111101001;
assign LUT_3[26258] = 32'b00000000000000011100100011110000;
assign LUT_3[26259] = 32'b00000000000000100011001111001101;
assign LUT_3[26260] = 32'b00000000000000010111101010000010;
assign LUT_3[26261] = 32'b00000000000000011110010101011111;
assign LUT_3[26262] = 32'b00000000000000011001110001100110;
assign LUT_3[26263] = 32'b00000000000000100000011101000011;
assign LUT_3[26264] = 32'b00000000000000011111110101010010;
assign LUT_3[26265] = 32'b00000000000000100110100000101111;
assign LUT_3[26266] = 32'b00000000000000100001111100110110;
assign LUT_3[26267] = 32'b00000000000000101000101000010011;
assign LUT_3[26268] = 32'b00000000000000011101000011001000;
assign LUT_3[26269] = 32'b00000000000000100011101110100101;
assign LUT_3[26270] = 32'b00000000000000011111001010101100;
assign LUT_3[26271] = 32'b00000000000000100101110110001001;
assign LUT_3[26272] = 32'b00000000000000011000010111101001;
assign LUT_3[26273] = 32'b00000000000000011111000011000110;
assign LUT_3[26274] = 32'b00000000000000011010011111001101;
assign LUT_3[26275] = 32'b00000000000000100001001010101010;
assign LUT_3[26276] = 32'b00000000000000010101100101011111;
assign LUT_3[26277] = 32'b00000000000000011100010000111100;
assign LUT_3[26278] = 32'b00000000000000010111101101000011;
assign LUT_3[26279] = 32'b00000000000000011110011000100000;
assign LUT_3[26280] = 32'b00000000000000011101110000101111;
assign LUT_3[26281] = 32'b00000000000000100100011100001100;
assign LUT_3[26282] = 32'b00000000000000011111111000010011;
assign LUT_3[26283] = 32'b00000000000000100110100011110000;
assign LUT_3[26284] = 32'b00000000000000011010111110100101;
assign LUT_3[26285] = 32'b00000000000000100001101010000010;
assign LUT_3[26286] = 32'b00000000000000011101000110001001;
assign LUT_3[26287] = 32'b00000000000000100011110001100110;
assign LUT_3[26288] = 32'b00000000000000011011101010101100;
assign LUT_3[26289] = 32'b00000000000000100010010110001001;
assign LUT_3[26290] = 32'b00000000000000011101110010010000;
assign LUT_3[26291] = 32'b00000000000000100100011101101101;
assign LUT_3[26292] = 32'b00000000000000011000111000100010;
assign LUT_3[26293] = 32'b00000000000000011111100011111111;
assign LUT_3[26294] = 32'b00000000000000011011000000000110;
assign LUT_3[26295] = 32'b00000000000000100001101011100011;
assign LUT_3[26296] = 32'b00000000000000100001000011110010;
assign LUT_3[26297] = 32'b00000000000000100111101111001111;
assign LUT_3[26298] = 32'b00000000000000100011001011010110;
assign LUT_3[26299] = 32'b00000000000000101001110110110011;
assign LUT_3[26300] = 32'b00000000000000011110010001101000;
assign LUT_3[26301] = 32'b00000000000000100100111101000101;
assign LUT_3[26302] = 32'b00000000000000100000011001001100;
assign LUT_3[26303] = 32'b00000000000000100111000100101001;
assign LUT_3[26304] = 32'b00000000000000010111000001110100;
assign LUT_3[26305] = 32'b00000000000000011101101101010001;
assign LUT_3[26306] = 32'b00000000000000011001001001011000;
assign LUT_3[26307] = 32'b00000000000000011111110100110101;
assign LUT_3[26308] = 32'b00000000000000010100001111101010;
assign LUT_3[26309] = 32'b00000000000000011010111011000111;
assign LUT_3[26310] = 32'b00000000000000010110010111001110;
assign LUT_3[26311] = 32'b00000000000000011101000010101011;
assign LUT_3[26312] = 32'b00000000000000011100011010111010;
assign LUT_3[26313] = 32'b00000000000000100011000110010111;
assign LUT_3[26314] = 32'b00000000000000011110100010011110;
assign LUT_3[26315] = 32'b00000000000000100101001101111011;
assign LUT_3[26316] = 32'b00000000000000011001101000110000;
assign LUT_3[26317] = 32'b00000000000000100000010100001101;
assign LUT_3[26318] = 32'b00000000000000011011110000010100;
assign LUT_3[26319] = 32'b00000000000000100010011011110001;
assign LUT_3[26320] = 32'b00000000000000011010010100110111;
assign LUT_3[26321] = 32'b00000000000000100001000000010100;
assign LUT_3[26322] = 32'b00000000000000011100011100011011;
assign LUT_3[26323] = 32'b00000000000000100011000111111000;
assign LUT_3[26324] = 32'b00000000000000010111100010101101;
assign LUT_3[26325] = 32'b00000000000000011110001110001010;
assign LUT_3[26326] = 32'b00000000000000011001101010010001;
assign LUT_3[26327] = 32'b00000000000000100000010101101110;
assign LUT_3[26328] = 32'b00000000000000011111101101111101;
assign LUT_3[26329] = 32'b00000000000000100110011001011010;
assign LUT_3[26330] = 32'b00000000000000100001110101100001;
assign LUT_3[26331] = 32'b00000000000000101000100000111110;
assign LUT_3[26332] = 32'b00000000000000011100111011110011;
assign LUT_3[26333] = 32'b00000000000000100011100111010000;
assign LUT_3[26334] = 32'b00000000000000011111000011010111;
assign LUT_3[26335] = 32'b00000000000000100101101110110100;
assign LUT_3[26336] = 32'b00000000000000011000010000010100;
assign LUT_3[26337] = 32'b00000000000000011110111011110001;
assign LUT_3[26338] = 32'b00000000000000011010010111111000;
assign LUT_3[26339] = 32'b00000000000000100001000011010101;
assign LUT_3[26340] = 32'b00000000000000010101011110001010;
assign LUT_3[26341] = 32'b00000000000000011100001001100111;
assign LUT_3[26342] = 32'b00000000000000010111100101101110;
assign LUT_3[26343] = 32'b00000000000000011110010001001011;
assign LUT_3[26344] = 32'b00000000000000011101101001011010;
assign LUT_3[26345] = 32'b00000000000000100100010100110111;
assign LUT_3[26346] = 32'b00000000000000011111110000111110;
assign LUT_3[26347] = 32'b00000000000000100110011100011011;
assign LUT_3[26348] = 32'b00000000000000011010110111010000;
assign LUT_3[26349] = 32'b00000000000000100001100010101101;
assign LUT_3[26350] = 32'b00000000000000011100111110110100;
assign LUT_3[26351] = 32'b00000000000000100011101010010001;
assign LUT_3[26352] = 32'b00000000000000011011100011010111;
assign LUT_3[26353] = 32'b00000000000000100010001110110100;
assign LUT_3[26354] = 32'b00000000000000011101101010111011;
assign LUT_3[26355] = 32'b00000000000000100100010110011000;
assign LUT_3[26356] = 32'b00000000000000011000110001001101;
assign LUT_3[26357] = 32'b00000000000000011111011100101010;
assign LUT_3[26358] = 32'b00000000000000011010111000110001;
assign LUT_3[26359] = 32'b00000000000000100001100100001110;
assign LUT_3[26360] = 32'b00000000000000100000111100011101;
assign LUT_3[26361] = 32'b00000000000000100111100111111010;
assign LUT_3[26362] = 32'b00000000000000100011000100000001;
assign LUT_3[26363] = 32'b00000000000000101001101111011110;
assign LUT_3[26364] = 32'b00000000000000011110001010010011;
assign LUT_3[26365] = 32'b00000000000000100100110101110000;
assign LUT_3[26366] = 32'b00000000000000100000010001110111;
assign LUT_3[26367] = 32'b00000000000000100110111101010100;
assign LUT_3[26368] = 32'b00000000000000010001001101101100;
assign LUT_3[26369] = 32'b00000000000000010111111001001001;
assign LUT_3[26370] = 32'b00000000000000010011010101010000;
assign LUT_3[26371] = 32'b00000000000000011010000000101101;
assign LUT_3[26372] = 32'b00000000000000001110011011100010;
assign LUT_3[26373] = 32'b00000000000000010101000110111111;
assign LUT_3[26374] = 32'b00000000000000010000100011000110;
assign LUT_3[26375] = 32'b00000000000000010111001110100011;
assign LUT_3[26376] = 32'b00000000000000010110100110110010;
assign LUT_3[26377] = 32'b00000000000000011101010010001111;
assign LUT_3[26378] = 32'b00000000000000011000101110010110;
assign LUT_3[26379] = 32'b00000000000000011111011001110011;
assign LUT_3[26380] = 32'b00000000000000010011110100101000;
assign LUT_3[26381] = 32'b00000000000000011010100000000101;
assign LUT_3[26382] = 32'b00000000000000010101111100001100;
assign LUT_3[26383] = 32'b00000000000000011100100111101001;
assign LUT_3[26384] = 32'b00000000000000010100100000101111;
assign LUT_3[26385] = 32'b00000000000000011011001100001100;
assign LUT_3[26386] = 32'b00000000000000010110101000010011;
assign LUT_3[26387] = 32'b00000000000000011101010011110000;
assign LUT_3[26388] = 32'b00000000000000010001101110100101;
assign LUT_3[26389] = 32'b00000000000000011000011010000010;
assign LUT_3[26390] = 32'b00000000000000010011110110001001;
assign LUT_3[26391] = 32'b00000000000000011010100001100110;
assign LUT_3[26392] = 32'b00000000000000011001111001110101;
assign LUT_3[26393] = 32'b00000000000000100000100101010010;
assign LUT_3[26394] = 32'b00000000000000011100000001011001;
assign LUT_3[26395] = 32'b00000000000000100010101100110110;
assign LUT_3[26396] = 32'b00000000000000010111000111101011;
assign LUT_3[26397] = 32'b00000000000000011101110011001000;
assign LUT_3[26398] = 32'b00000000000000011001001111001111;
assign LUT_3[26399] = 32'b00000000000000011111111010101100;
assign LUT_3[26400] = 32'b00000000000000010010011100001100;
assign LUT_3[26401] = 32'b00000000000000011001000111101001;
assign LUT_3[26402] = 32'b00000000000000010100100011110000;
assign LUT_3[26403] = 32'b00000000000000011011001111001101;
assign LUT_3[26404] = 32'b00000000000000001111101010000010;
assign LUT_3[26405] = 32'b00000000000000010110010101011111;
assign LUT_3[26406] = 32'b00000000000000010001110001100110;
assign LUT_3[26407] = 32'b00000000000000011000011101000011;
assign LUT_3[26408] = 32'b00000000000000010111110101010010;
assign LUT_3[26409] = 32'b00000000000000011110100000101111;
assign LUT_3[26410] = 32'b00000000000000011001111100110110;
assign LUT_3[26411] = 32'b00000000000000100000101000010011;
assign LUT_3[26412] = 32'b00000000000000010101000011001000;
assign LUT_3[26413] = 32'b00000000000000011011101110100101;
assign LUT_3[26414] = 32'b00000000000000010111001010101100;
assign LUT_3[26415] = 32'b00000000000000011101110110001001;
assign LUT_3[26416] = 32'b00000000000000010101101111001111;
assign LUT_3[26417] = 32'b00000000000000011100011010101100;
assign LUT_3[26418] = 32'b00000000000000010111110110110011;
assign LUT_3[26419] = 32'b00000000000000011110100010010000;
assign LUT_3[26420] = 32'b00000000000000010010111101000101;
assign LUT_3[26421] = 32'b00000000000000011001101000100010;
assign LUT_3[26422] = 32'b00000000000000010101000100101001;
assign LUT_3[26423] = 32'b00000000000000011011110000000110;
assign LUT_3[26424] = 32'b00000000000000011011001000010101;
assign LUT_3[26425] = 32'b00000000000000100001110011110010;
assign LUT_3[26426] = 32'b00000000000000011101001111111001;
assign LUT_3[26427] = 32'b00000000000000100011111011010110;
assign LUT_3[26428] = 32'b00000000000000011000010110001011;
assign LUT_3[26429] = 32'b00000000000000011111000001101000;
assign LUT_3[26430] = 32'b00000000000000011010011101101111;
assign LUT_3[26431] = 32'b00000000000000100001001001001100;
assign LUT_3[26432] = 32'b00000000000000010001000110010111;
assign LUT_3[26433] = 32'b00000000000000010111110001110100;
assign LUT_3[26434] = 32'b00000000000000010011001101111011;
assign LUT_3[26435] = 32'b00000000000000011001111001011000;
assign LUT_3[26436] = 32'b00000000000000001110010100001101;
assign LUT_3[26437] = 32'b00000000000000010100111111101010;
assign LUT_3[26438] = 32'b00000000000000010000011011110001;
assign LUT_3[26439] = 32'b00000000000000010111000111001110;
assign LUT_3[26440] = 32'b00000000000000010110011111011101;
assign LUT_3[26441] = 32'b00000000000000011101001010111010;
assign LUT_3[26442] = 32'b00000000000000011000100111000001;
assign LUT_3[26443] = 32'b00000000000000011111010010011110;
assign LUT_3[26444] = 32'b00000000000000010011101101010011;
assign LUT_3[26445] = 32'b00000000000000011010011000110000;
assign LUT_3[26446] = 32'b00000000000000010101110100110111;
assign LUT_3[26447] = 32'b00000000000000011100100000010100;
assign LUT_3[26448] = 32'b00000000000000010100011001011010;
assign LUT_3[26449] = 32'b00000000000000011011000100110111;
assign LUT_3[26450] = 32'b00000000000000010110100000111110;
assign LUT_3[26451] = 32'b00000000000000011101001100011011;
assign LUT_3[26452] = 32'b00000000000000010001100111010000;
assign LUT_3[26453] = 32'b00000000000000011000010010101101;
assign LUT_3[26454] = 32'b00000000000000010011101110110100;
assign LUT_3[26455] = 32'b00000000000000011010011010010001;
assign LUT_3[26456] = 32'b00000000000000011001110010100000;
assign LUT_3[26457] = 32'b00000000000000100000011101111101;
assign LUT_3[26458] = 32'b00000000000000011011111010000100;
assign LUT_3[26459] = 32'b00000000000000100010100101100001;
assign LUT_3[26460] = 32'b00000000000000010111000000010110;
assign LUT_3[26461] = 32'b00000000000000011101101011110011;
assign LUT_3[26462] = 32'b00000000000000011001000111111010;
assign LUT_3[26463] = 32'b00000000000000011111110011010111;
assign LUT_3[26464] = 32'b00000000000000010010010100110111;
assign LUT_3[26465] = 32'b00000000000000011001000000010100;
assign LUT_3[26466] = 32'b00000000000000010100011100011011;
assign LUT_3[26467] = 32'b00000000000000011011000111111000;
assign LUT_3[26468] = 32'b00000000000000001111100010101101;
assign LUT_3[26469] = 32'b00000000000000010110001110001010;
assign LUT_3[26470] = 32'b00000000000000010001101010010001;
assign LUT_3[26471] = 32'b00000000000000011000010101101110;
assign LUT_3[26472] = 32'b00000000000000010111101101111101;
assign LUT_3[26473] = 32'b00000000000000011110011001011010;
assign LUT_3[26474] = 32'b00000000000000011001110101100001;
assign LUT_3[26475] = 32'b00000000000000100000100000111110;
assign LUT_3[26476] = 32'b00000000000000010100111011110011;
assign LUT_3[26477] = 32'b00000000000000011011100111010000;
assign LUT_3[26478] = 32'b00000000000000010111000011010111;
assign LUT_3[26479] = 32'b00000000000000011101101110110100;
assign LUT_3[26480] = 32'b00000000000000010101100111111010;
assign LUT_3[26481] = 32'b00000000000000011100010011010111;
assign LUT_3[26482] = 32'b00000000000000010111101111011110;
assign LUT_3[26483] = 32'b00000000000000011110011010111011;
assign LUT_3[26484] = 32'b00000000000000010010110101110000;
assign LUT_3[26485] = 32'b00000000000000011001100001001101;
assign LUT_3[26486] = 32'b00000000000000010100111101010100;
assign LUT_3[26487] = 32'b00000000000000011011101000110001;
assign LUT_3[26488] = 32'b00000000000000011011000001000000;
assign LUT_3[26489] = 32'b00000000000000100001101100011101;
assign LUT_3[26490] = 32'b00000000000000011101001000100100;
assign LUT_3[26491] = 32'b00000000000000100011110100000001;
assign LUT_3[26492] = 32'b00000000000000011000001110110110;
assign LUT_3[26493] = 32'b00000000000000011110111010010011;
assign LUT_3[26494] = 32'b00000000000000011010010110011010;
assign LUT_3[26495] = 32'b00000000000000100001000001110111;
assign LUT_3[26496] = 32'b00000000000000010011011000101010;
assign LUT_3[26497] = 32'b00000000000000011010000100000111;
assign LUT_3[26498] = 32'b00000000000000010101100000001110;
assign LUT_3[26499] = 32'b00000000000000011100001011101011;
assign LUT_3[26500] = 32'b00000000000000010000100110100000;
assign LUT_3[26501] = 32'b00000000000000010111010001111101;
assign LUT_3[26502] = 32'b00000000000000010010101110000100;
assign LUT_3[26503] = 32'b00000000000000011001011001100001;
assign LUT_3[26504] = 32'b00000000000000011000110001110000;
assign LUT_3[26505] = 32'b00000000000000011111011101001101;
assign LUT_3[26506] = 32'b00000000000000011010111001010100;
assign LUT_3[26507] = 32'b00000000000000100001100100110001;
assign LUT_3[26508] = 32'b00000000000000010101111111100110;
assign LUT_3[26509] = 32'b00000000000000011100101011000011;
assign LUT_3[26510] = 32'b00000000000000011000000111001010;
assign LUT_3[26511] = 32'b00000000000000011110110010100111;
assign LUT_3[26512] = 32'b00000000000000010110101011101101;
assign LUT_3[26513] = 32'b00000000000000011101010111001010;
assign LUT_3[26514] = 32'b00000000000000011000110011010001;
assign LUT_3[26515] = 32'b00000000000000011111011110101110;
assign LUT_3[26516] = 32'b00000000000000010011111001100011;
assign LUT_3[26517] = 32'b00000000000000011010100101000000;
assign LUT_3[26518] = 32'b00000000000000010110000001000111;
assign LUT_3[26519] = 32'b00000000000000011100101100100100;
assign LUT_3[26520] = 32'b00000000000000011100000100110011;
assign LUT_3[26521] = 32'b00000000000000100010110000010000;
assign LUT_3[26522] = 32'b00000000000000011110001100010111;
assign LUT_3[26523] = 32'b00000000000000100100110111110100;
assign LUT_3[26524] = 32'b00000000000000011001010010101001;
assign LUT_3[26525] = 32'b00000000000000011111111110000110;
assign LUT_3[26526] = 32'b00000000000000011011011010001101;
assign LUT_3[26527] = 32'b00000000000000100010000101101010;
assign LUT_3[26528] = 32'b00000000000000010100100111001010;
assign LUT_3[26529] = 32'b00000000000000011011010010100111;
assign LUT_3[26530] = 32'b00000000000000010110101110101110;
assign LUT_3[26531] = 32'b00000000000000011101011010001011;
assign LUT_3[26532] = 32'b00000000000000010001110101000000;
assign LUT_3[26533] = 32'b00000000000000011000100000011101;
assign LUT_3[26534] = 32'b00000000000000010011111100100100;
assign LUT_3[26535] = 32'b00000000000000011010101000000001;
assign LUT_3[26536] = 32'b00000000000000011010000000010000;
assign LUT_3[26537] = 32'b00000000000000100000101011101101;
assign LUT_3[26538] = 32'b00000000000000011100000111110100;
assign LUT_3[26539] = 32'b00000000000000100010110011010001;
assign LUT_3[26540] = 32'b00000000000000010111001110000110;
assign LUT_3[26541] = 32'b00000000000000011101111001100011;
assign LUT_3[26542] = 32'b00000000000000011001010101101010;
assign LUT_3[26543] = 32'b00000000000000100000000001000111;
assign LUT_3[26544] = 32'b00000000000000010111111010001101;
assign LUT_3[26545] = 32'b00000000000000011110100101101010;
assign LUT_3[26546] = 32'b00000000000000011010000001110001;
assign LUT_3[26547] = 32'b00000000000000100000101101001110;
assign LUT_3[26548] = 32'b00000000000000010101001000000011;
assign LUT_3[26549] = 32'b00000000000000011011110011100000;
assign LUT_3[26550] = 32'b00000000000000010111001111100111;
assign LUT_3[26551] = 32'b00000000000000011101111011000100;
assign LUT_3[26552] = 32'b00000000000000011101010011010011;
assign LUT_3[26553] = 32'b00000000000000100011111110110000;
assign LUT_3[26554] = 32'b00000000000000011111011010110111;
assign LUT_3[26555] = 32'b00000000000000100110000110010100;
assign LUT_3[26556] = 32'b00000000000000011010100001001001;
assign LUT_3[26557] = 32'b00000000000000100001001100100110;
assign LUT_3[26558] = 32'b00000000000000011100101000101101;
assign LUT_3[26559] = 32'b00000000000000100011010100001010;
assign LUT_3[26560] = 32'b00000000000000010011010001010101;
assign LUT_3[26561] = 32'b00000000000000011001111100110010;
assign LUT_3[26562] = 32'b00000000000000010101011000111001;
assign LUT_3[26563] = 32'b00000000000000011100000100010110;
assign LUT_3[26564] = 32'b00000000000000010000011111001011;
assign LUT_3[26565] = 32'b00000000000000010111001010101000;
assign LUT_3[26566] = 32'b00000000000000010010100110101111;
assign LUT_3[26567] = 32'b00000000000000011001010010001100;
assign LUT_3[26568] = 32'b00000000000000011000101010011011;
assign LUT_3[26569] = 32'b00000000000000011111010101111000;
assign LUT_3[26570] = 32'b00000000000000011010110001111111;
assign LUT_3[26571] = 32'b00000000000000100001011101011100;
assign LUT_3[26572] = 32'b00000000000000010101111000010001;
assign LUT_3[26573] = 32'b00000000000000011100100011101110;
assign LUT_3[26574] = 32'b00000000000000010111111111110101;
assign LUT_3[26575] = 32'b00000000000000011110101011010010;
assign LUT_3[26576] = 32'b00000000000000010110100100011000;
assign LUT_3[26577] = 32'b00000000000000011101001111110101;
assign LUT_3[26578] = 32'b00000000000000011000101011111100;
assign LUT_3[26579] = 32'b00000000000000011111010111011001;
assign LUT_3[26580] = 32'b00000000000000010011110010001110;
assign LUT_3[26581] = 32'b00000000000000011010011101101011;
assign LUT_3[26582] = 32'b00000000000000010101111001110010;
assign LUT_3[26583] = 32'b00000000000000011100100101001111;
assign LUT_3[26584] = 32'b00000000000000011011111101011110;
assign LUT_3[26585] = 32'b00000000000000100010101000111011;
assign LUT_3[26586] = 32'b00000000000000011110000101000010;
assign LUT_3[26587] = 32'b00000000000000100100110000011111;
assign LUT_3[26588] = 32'b00000000000000011001001011010100;
assign LUT_3[26589] = 32'b00000000000000011111110110110001;
assign LUT_3[26590] = 32'b00000000000000011011010010111000;
assign LUT_3[26591] = 32'b00000000000000100001111110010101;
assign LUT_3[26592] = 32'b00000000000000010100011111110101;
assign LUT_3[26593] = 32'b00000000000000011011001011010010;
assign LUT_3[26594] = 32'b00000000000000010110100111011001;
assign LUT_3[26595] = 32'b00000000000000011101010010110110;
assign LUT_3[26596] = 32'b00000000000000010001101101101011;
assign LUT_3[26597] = 32'b00000000000000011000011001001000;
assign LUT_3[26598] = 32'b00000000000000010011110101001111;
assign LUT_3[26599] = 32'b00000000000000011010100000101100;
assign LUT_3[26600] = 32'b00000000000000011001111000111011;
assign LUT_3[26601] = 32'b00000000000000100000100100011000;
assign LUT_3[26602] = 32'b00000000000000011100000000011111;
assign LUT_3[26603] = 32'b00000000000000100010101011111100;
assign LUT_3[26604] = 32'b00000000000000010111000110110001;
assign LUT_3[26605] = 32'b00000000000000011101110010001110;
assign LUT_3[26606] = 32'b00000000000000011001001110010101;
assign LUT_3[26607] = 32'b00000000000000011111111001110010;
assign LUT_3[26608] = 32'b00000000000000010111110010111000;
assign LUT_3[26609] = 32'b00000000000000011110011110010101;
assign LUT_3[26610] = 32'b00000000000000011001111010011100;
assign LUT_3[26611] = 32'b00000000000000100000100101111001;
assign LUT_3[26612] = 32'b00000000000000010101000000101110;
assign LUT_3[26613] = 32'b00000000000000011011101100001011;
assign LUT_3[26614] = 32'b00000000000000010111001000010010;
assign LUT_3[26615] = 32'b00000000000000011101110011101111;
assign LUT_3[26616] = 32'b00000000000000011101001011111110;
assign LUT_3[26617] = 32'b00000000000000100011110111011011;
assign LUT_3[26618] = 32'b00000000000000011111010011100010;
assign LUT_3[26619] = 32'b00000000000000100101111110111111;
assign LUT_3[26620] = 32'b00000000000000011010011001110100;
assign LUT_3[26621] = 32'b00000000000000100001000101010001;
assign LUT_3[26622] = 32'b00000000000000011100100001011000;
assign LUT_3[26623] = 32'b00000000000000100011001100110101;
assign LUT_3[26624] = 32'b00000000000000001100111010010000;
assign LUT_3[26625] = 32'b00000000000000010011100101101101;
assign LUT_3[26626] = 32'b00000000000000001111000001110100;
assign LUT_3[26627] = 32'b00000000000000010101101101010001;
assign LUT_3[26628] = 32'b00000000000000001010001000000110;
assign LUT_3[26629] = 32'b00000000000000010000110011100011;
assign LUT_3[26630] = 32'b00000000000000001100001111101010;
assign LUT_3[26631] = 32'b00000000000000010010111011000111;
assign LUT_3[26632] = 32'b00000000000000010010010011010110;
assign LUT_3[26633] = 32'b00000000000000011000111110110011;
assign LUT_3[26634] = 32'b00000000000000010100011010111010;
assign LUT_3[26635] = 32'b00000000000000011011000110010111;
assign LUT_3[26636] = 32'b00000000000000001111100001001100;
assign LUT_3[26637] = 32'b00000000000000010110001100101001;
assign LUT_3[26638] = 32'b00000000000000010001101000110000;
assign LUT_3[26639] = 32'b00000000000000011000010100001101;
assign LUT_3[26640] = 32'b00000000000000010000001101010011;
assign LUT_3[26641] = 32'b00000000000000010110111000110000;
assign LUT_3[26642] = 32'b00000000000000010010010100110111;
assign LUT_3[26643] = 32'b00000000000000011001000000010100;
assign LUT_3[26644] = 32'b00000000000000001101011011001001;
assign LUT_3[26645] = 32'b00000000000000010100000110100110;
assign LUT_3[26646] = 32'b00000000000000001111100010101101;
assign LUT_3[26647] = 32'b00000000000000010110001110001010;
assign LUT_3[26648] = 32'b00000000000000010101100110011001;
assign LUT_3[26649] = 32'b00000000000000011100010001110110;
assign LUT_3[26650] = 32'b00000000000000010111101101111101;
assign LUT_3[26651] = 32'b00000000000000011110011001011010;
assign LUT_3[26652] = 32'b00000000000000010010110100001111;
assign LUT_3[26653] = 32'b00000000000000011001011111101100;
assign LUT_3[26654] = 32'b00000000000000010100111011110011;
assign LUT_3[26655] = 32'b00000000000000011011100111010000;
assign LUT_3[26656] = 32'b00000000000000001110001000110000;
assign LUT_3[26657] = 32'b00000000000000010100110100001101;
assign LUT_3[26658] = 32'b00000000000000010000010000010100;
assign LUT_3[26659] = 32'b00000000000000010110111011110001;
assign LUT_3[26660] = 32'b00000000000000001011010110100110;
assign LUT_3[26661] = 32'b00000000000000010010000010000011;
assign LUT_3[26662] = 32'b00000000000000001101011110001010;
assign LUT_3[26663] = 32'b00000000000000010100001001100111;
assign LUT_3[26664] = 32'b00000000000000010011100001110110;
assign LUT_3[26665] = 32'b00000000000000011010001101010011;
assign LUT_3[26666] = 32'b00000000000000010101101001011010;
assign LUT_3[26667] = 32'b00000000000000011100010100110111;
assign LUT_3[26668] = 32'b00000000000000010000101111101100;
assign LUT_3[26669] = 32'b00000000000000010111011011001001;
assign LUT_3[26670] = 32'b00000000000000010010110111010000;
assign LUT_3[26671] = 32'b00000000000000011001100010101101;
assign LUT_3[26672] = 32'b00000000000000010001011011110011;
assign LUT_3[26673] = 32'b00000000000000011000000111010000;
assign LUT_3[26674] = 32'b00000000000000010011100011010111;
assign LUT_3[26675] = 32'b00000000000000011010001110110100;
assign LUT_3[26676] = 32'b00000000000000001110101001101001;
assign LUT_3[26677] = 32'b00000000000000010101010101000110;
assign LUT_3[26678] = 32'b00000000000000010000110001001101;
assign LUT_3[26679] = 32'b00000000000000010111011100101010;
assign LUT_3[26680] = 32'b00000000000000010110110100111001;
assign LUT_3[26681] = 32'b00000000000000011101100000010110;
assign LUT_3[26682] = 32'b00000000000000011000111100011101;
assign LUT_3[26683] = 32'b00000000000000011111100111111010;
assign LUT_3[26684] = 32'b00000000000000010100000010101111;
assign LUT_3[26685] = 32'b00000000000000011010101110001100;
assign LUT_3[26686] = 32'b00000000000000010110001010010011;
assign LUT_3[26687] = 32'b00000000000000011100110101110000;
assign LUT_3[26688] = 32'b00000000000000001100110010111011;
assign LUT_3[26689] = 32'b00000000000000010011011110011000;
assign LUT_3[26690] = 32'b00000000000000001110111010011111;
assign LUT_3[26691] = 32'b00000000000000010101100101111100;
assign LUT_3[26692] = 32'b00000000000000001010000000110001;
assign LUT_3[26693] = 32'b00000000000000010000101100001110;
assign LUT_3[26694] = 32'b00000000000000001100001000010101;
assign LUT_3[26695] = 32'b00000000000000010010110011110010;
assign LUT_3[26696] = 32'b00000000000000010010001100000001;
assign LUT_3[26697] = 32'b00000000000000011000110111011110;
assign LUT_3[26698] = 32'b00000000000000010100010011100101;
assign LUT_3[26699] = 32'b00000000000000011010111111000010;
assign LUT_3[26700] = 32'b00000000000000001111011001110111;
assign LUT_3[26701] = 32'b00000000000000010110000101010100;
assign LUT_3[26702] = 32'b00000000000000010001100001011011;
assign LUT_3[26703] = 32'b00000000000000011000001100111000;
assign LUT_3[26704] = 32'b00000000000000010000000101111110;
assign LUT_3[26705] = 32'b00000000000000010110110001011011;
assign LUT_3[26706] = 32'b00000000000000010010001101100010;
assign LUT_3[26707] = 32'b00000000000000011000111000111111;
assign LUT_3[26708] = 32'b00000000000000001101010011110100;
assign LUT_3[26709] = 32'b00000000000000010011111111010001;
assign LUT_3[26710] = 32'b00000000000000001111011011011000;
assign LUT_3[26711] = 32'b00000000000000010110000110110101;
assign LUT_3[26712] = 32'b00000000000000010101011111000100;
assign LUT_3[26713] = 32'b00000000000000011100001010100001;
assign LUT_3[26714] = 32'b00000000000000010111100110101000;
assign LUT_3[26715] = 32'b00000000000000011110010010000101;
assign LUT_3[26716] = 32'b00000000000000010010101100111010;
assign LUT_3[26717] = 32'b00000000000000011001011000010111;
assign LUT_3[26718] = 32'b00000000000000010100110100011110;
assign LUT_3[26719] = 32'b00000000000000011011011111111011;
assign LUT_3[26720] = 32'b00000000000000001110000001011011;
assign LUT_3[26721] = 32'b00000000000000010100101100111000;
assign LUT_3[26722] = 32'b00000000000000010000001000111111;
assign LUT_3[26723] = 32'b00000000000000010110110100011100;
assign LUT_3[26724] = 32'b00000000000000001011001111010001;
assign LUT_3[26725] = 32'b00000000000000010001111010101110;
assign LUT_3[26726] = 32'b00000000000000001101010110110101;
assign LUT_3[26727] = 32'b00000000000000010100000010010010;
assign LUT_3[26728] = 32'b00000000000000010011011010100001;
assign LUT_3[26729] = 32'b00000000000000011010000101111110;
assign LUT_3[26730] = 32'b00000000000000010101100010000101;
assign LUT_3[26731] = 32'b00000000000000011100001101100010;
assign LUT_3[26732] = 32'b00000000000000010000101000010111;
assign LUT_3[26733] = 32'b00000000000000010111010011110100;
assign LUT_3[26734] = 32'b00000000000000010010101111111011;
assign LUT_3[26735] = 32'b00000000000000011001011011011000;
assign LUT_3[26736] = 32'b00000000000000010001010100011110;
assign LUT_3[26737] = 32'b00000000000000010111111111111011;
assign LUT_3[26738] = 32'b00000000000000010011011100000010;
assign LUT_3[26739] = 32'b00000000000000011010000111011111;
assign LUT_3[26740] = 32'b00000000000000001110100010010100;
assign LUT_3[26741] = 32'b00000000000000010101001101110001;
assign LUT_3[26742] = 32'b00000000000000010000101001111000;
assign LUT_3[26743] = 32'b00000000000000010111010101010101;
assign LUT_3[26744] = 32'b00000000000000010110101101100100;
assign LUT_3[26745] = 32'b00000000000000011101011001000001;
assign LUT_3[26746] = 32'b00000000000000011000110101001000;
assign LUT_3[26747] = 32'b00000000000000011111100000100101;
assign LUT_3[26748] = 32'b00000000000000010011111011011010;
assign LUT_3[26749] = 32'b00000000000000011010100110110111;
assign LUT_3[26750] = 32'b00000000000000010110000010111110;
assign LUT_3[26751] = 32'b00000000000000011100101110011011;
assign LUT_3[26752] = 32'b00000000000000001111000101001110;
assign LUT_3[26753] = 32'b00000000000000010101110000101011;
assign LUT_3[26754] = 32'b00000000000000010001001100110010;
assign LUT_3[26755] = 32'b00000000000000010111111000001111;
assign LUT_3[26756] = 32'b00000000000000001100010011000100;
assign LUT_3[26757] = 32'b00000000000000010010111110100001;
assign LUT_3[26758] = 32'b00000000000000001110011010101000;
assign LUT_3[26759] = 32'b00000000000000010101000110000101;
assign LUT_3[26760] = 32'b00000000000000010100011110010100;
assign LUT_3[26761] = 32'b00000000000000011011001001110001;
assign LUT_3[26762] = 32'b00000000000000010110100101111000;
assign LUT_3[26763] = 32'b00000000000000011101010001010101;
assign LUT_3[26764] = 32'b00000000000000010001101100001010;
assign LUT_3[26765] = 32'b00000000000000011000010111100111;
assign LUT_3[26766] = 32'b00000000000000010011110011101110;
assign LUT_3[26767] = 32'b00000000000000011010011111001011;
assign LUT_3[26768] = 32'b00000000000000010010011000010001;
assign LUT_3[26769] = 32'b00000000000000011001000011101110;
assign LUT_3[26770] = 32'b00000000000000010100011111110101;
assign LUT_3[26771] = 32'b00000000000000011011001011010010;
assign LUT_3[26772] = 32'b00000000000000001111100110000111;
assign LUT_3[26773] = 32'b00000000000000010110010001100100;
assign LUT_3[26774] = 32'b00000000000000010001101101101011;
assign LUT_3[26775] = 32'b00000000000000011000011001001000;
assign LUT_3[26776] = 32'b00000000000000010111110001010111;
assign LUT_3[26777] = 32'b00000000000000011110011100110100;
assign LUT_3[26778] = 32'b00000000000000011001111000111011;
assign LUT_3[26779] = 32'b00000000000000100000100100011000;
assign LUT_3[26780] = 32'b00000000000000010100111111001101;
assign LUT_3[26781] = 32'b00000000000000011011101010101010;
assign LUT_3[26782] = 32'b00000000000000010111000110110001;
assign LUT_3[26783] = 32'b00000000000000011101110010001110;
assign LUT_3[26784] = 32'b00000000000000010000010011101110;
assign LUT_3[26785] = 32'b00000000000000010110111111001011;
assign LUT_3[26786] = 32'b00000000000000010010011011010010;
assign LUT_3[26787] = 32'b00000000000000011001000110101111;
assign LUT_3[26788] = 32'b00000000000000001101100001100100;
assign LUT_3[26789] = 32'b00000000000000010100001101000001;
assign LUT_3[26790] = 32'b00000000000000001111101001001000;
assign LUT_3[26791] = 32'b00000000000000010110010100100101;
assign LUT_3[26792] = 32'b00000000000000010101101100110100;
assign LUT_3[26793] = 32'b00000000000000011100011000010001;
assign LUT_3[26794] = 32'b00000000000000010111110100011000;
assign LUT_3[26795] = 32'b00000000000000011110011111110101;
assign LUT_3[26796] = 32'b00000000000000010010111010101010;
assign LUT_3[26797] = 32'b00000000000000011001100110000111;
assign LUT_3[26798] = 32'b00000000000000010101000010001110;
assign LUT_3[26799] = 32'b00000000000000011011101101101011;
assign LUT_3[26800] = 32'b00000000000000010011100110110001;
assign LUT_3[26801] = 32'b00000000000000011010010010001110;
assign LUT_3[26802] = 32'b00000000000000010101101110010101;
assign LUT_3[26803] = 32'b00000000000000011100011001110010;
assign LUT_3[26804] = 32'b00000000000000010000110100100111;
assign LUT_3[26805] = 32'b00000000000000010111100000000100;
assign LUT_3[26806] = 32'b00000000000000010010111100001011;
assign LUT_3[26807] = 32'b00000000000000011001100111101000;
assign LUT_3[26808] = 32'b00000000000000011000111111110111;
assign LUT_3[26809] = 32'b00000000000000011111101011010100;
assign LUT_3[26810] = 32'b00000000000000011011000111011011;
assign LUT_3[26811] = 32'b00000000000000100001110010111000;
assign LUT_3[26812] = 32'b00000000000000010110001101101101;
assign LUT_3[26813] = 32'b00000000000000011100111001001010;
assign LUT_3[26814] = 32'b00000000000000011000010101010001;
assign LUT_3[26815] = 32'b00000000000000011111000000101110;
assign LUT_3[26816] = 32'b00000000000000001110111101111001;
assign LUT_3[26817] = 32'b00000000000000010101101001010110;
assign LUT_3[26818] = 32'b00000000000000010001000101011101;
assign LUT_3[26819] = 32'b00000000000000010111110000111010;
assign LUT_3[26820] = 32'b00000000000000001100001011101111;
assign LUT_3[26821] = 32'b00000000000000010010110111001100;
assign LUT_3[26822] = 32'b00000000000000001110010011010011;
assign LUT_3[26823] = 32'b00000000000000010100111110110000;
assign LUT_3[26824] = 32'b00000000000000010100010110111111;
assign LUT_3[26825] = 32'b00000000000000011011000010011100;
assign LUT_3[26826] = 32'b00000000000000010110011110100011;
assign LUT_3[26827] = 32'b00000000000000011101001010000000;
assign LUT_3[26828] = 32'b00000000000000010001100100110101;
assign LUT_3[26829] = 32'b00000000000000011000010000010010;
assign LUT_3[26830] = 32'b00000000000000010011101100011001;
assign LUT_3[26831] = 32'b00000000000000011010010111110110;
assign LUT_3[26832] = 32'b00000000000000010010010000111100;
assign LUT_3[26833] = 32'b00000000000000011000111100011001;
assign LUT_3[26834] = 32'b00000000000000010100011000100000;
assign LUT_3[26835] = 32'b00000000000000011011000011111101;
assign LUT_3[26836] = 32'b00000000000000001111011110110010;
assign LUT_3[26837] = 32'b00000000000000010110001010001111;
assign LUT_3[26838] = 32'b00000000000000010001100110010110;
assign LUT_3[26839] = 32'b00000000000000011000010001110011;
assign LUT_3[26840] = 32'b00000000000000010111101010000010;
assign LUT_3[26841] = 32'b00000000000000011110010101011111;
assign LUT_3[26842] = 32'b00000000000000011001110001100110;
assign LUT_3[26843] = 32'b00000000000000100000011101000011;
assign LUT_3[26844] = 32'b00000000000000010100110111111000;
assign LUT_3[26845] = 32'b00000000000000011011100011010101;
assign LUT_3[26846] = 32'b00000000000000010110111111011100;
assign LUT_3[26847] = 32'b00000000000000011101101010111001;
assign LUT_3[26848] = 32'b00000000000000010000001100011001;
assign LUT_3[26849] = 32'b00000000000000010110110111110110;
assign LUT_3[26850] = 32'b00000000000000010010010011111101;
assign LUT_3[26851] = 32'b00000000000000011000111111011010;
assign LUT_3[26852] = 32'b00000000000000001101011010001111;
assign LUT_3[26853] = 32'b00000000000000010100000101101100;
assign LUT_3[26854] = 32'b00000000000000001111100001110011;
assign LUT_3[26855] = 32'b00000000000000010110001101010000;
assign LUT_3[26856] = 32'b00000000000000010101100101011111;
assign LUT_3[26857] = 32'b00000000000000011100010000111100;
assign LUT_3[26858] = 32'b00000000000000010111101101000011;
assign LUT_3[26859] = 32'b00000000000000011110011000100000;
assign LUT_3[26860] = 32'b00000000000000010010110011010101;
assign LUT_3[26861] = 32'b00000000000000011001011110110010;
assign LUT_3[26862] = 32'b00000000000000010100111010111001;
assign LUT_3[26863] = 32'b00000000000000011011100110010110;
assign LUT_3[26864] = 32'b00000000000000010011011111011100;
assign LUT_3[26865] = 32'b00000000000000011010001010111001;
assign LUT_3[26866] = 32'b00000000000000010101100111000000;
assign LUT_3[26867] = 32'b00000000000000011100010010011101;
assign LUT_3[26868] = 32'b00000000000000010000101101010010;
assign LUT_3[26869] = 32'b00000000000000010111011000101111;
assign LUT_3[26870] = 32'b00000000000000010010110100110110;
assign LUT_3[26871] = 32'b00000000000000011001100000010011;
assign LUT_3[26872] = 32'b00000000000000011000111000100010;
assign LUT_3[26873] = 32'b00000000000000011111100011111111;
assign LUT_3[26874] = 32'b00000000000000011011000000000110;
assign LUT_3[26875] = 32'b00000000000000100001101011100011;
assign LUT_3[26876] = 32'b00000000000000010110000110011000;
assign LUT_3[26877] = 32'b00000000000000011100110001110101;
assign LUT_3[26878] = 32'b00000000000000011000001101111100;
assign LUT_3[26879] = 32'b00000000000000011110111001011001;
assign LUT_3[26880] = 32'b00000000000000001001001001110001;
assign LUT_3[26881] = 32'b00000000000000001111110101001110;
assign LUT_3[26882] = 32'b00000000000000001011010001010101;
assign LUT_3[26883] = 32'b00000000000000010001111100110010;
assign LUT_3[26884] = 32'b00000000000000000110010111100111;
assign LUT_3[26885] = 32'b00000000000000001101000011000100;
assign LUT_3[26886] = 32'b00000000000000001000011111001011;
assign LUT_3[26887] = 32'b00000000000000001111001010101000;
assign LUT_3[26888] = 32'b00000000000000001110100010110111;
assign LUT_3[26889] = 32'b00000000000000010101001110010100;
assign LUT_3[26890] = 32'b00000000000000010000101010011011;
assign LUT_3[26891] = 32'b00000000000000010111010101111000;
assign LUT_3[26892] = 32'b00000000000000001011110000101101;
assign LUT_3[26893] = 32'b00000000000000010010011100001010;
assign LUT_3[26894] = 32'b00000000000000001101111000010001;
assign LUT_3[26895] = 32'b00000000000000010100100011101110;
assign LUT_3[26896] = 32'b00000000000000001100011100110100;
assign LUT_3[26897] = 32'b00000000000000010011001000010001;
assign LUT_3[26898] = 32'b00000000000000001110100100011000;
assign LUT_3[26899] = 32'b00000000000000010101001111110101;
assign LUT_3[26900] = 32'b00000000000000001001101010101010;
assign LUT_3[26901] = 32'b00000000000000010000010110000111;
assign LUT_3[26902] = 32'b00000000000000001011110010001110;
assign LUT_3[26903] = 32'b00000000000000010010011101101011;
assign LUT_3[26904] = 32'b00000000000000010001110101111010;
assign LUT_3[26905] = 32'b00000000000000011000100001010111;
assign LUT_3[26906] = 32'b00000000000000010011111101011110;
assign LUT_3[26907] = 32'b00000000000000011010101000111011;
assign LUT_3[26908] = 32'b00000000000000001111000011110000;
assign LUT_3[26909] = 32'b00000000000000010101101111001101;
assign LUT_3[26910] = 32'b00000000000000010001001011010100;
assign LUT_3[26911] = 32'b00000000000000010111110110110001;
assign LUT_3[26912] = 32'b00000000000000001010011000010001;
assign LUT_3[26913] = 32'b00000000000000010001000011101110;
assign LUT_3[26914] = 32'b00000000000000001100011111110101;
assign LUT_3[26915] = 32'b00000000000000010011001011010010;
assign LUT_3[26916] = 32'b00000000000000000111100110000111;
assign LUT_3[26917] = 32'b00000000000000001110010001100100;
assign LUT_3[26918] = 32'b00000000000000001001101101101011;
assign LUT_3[26919] = 32'b00000000000000010000011001001000;
assign LUT_3[26920] = 32'b00000000000000001111110001010111;
assign LUT_3[26921] = 32'b00000000000000010110011100110100;
assign LUT_3[26922] = 32'b00000000000000010001111000111011;
assign LUT_3[26923] = 32'b00000000000000011000100100011000;
assign LUT_3[26924] = 32'b00000000000000001100111111001101;
assign LUT_3[26925] = 32'b00000000000000010011101010101010;
assign LUT_3[26926] = 32'b00000000000000001111000110110001;
assign LUT_3[26927] = 32'b00000000000000010101110010001110;
assign LUT_3[26928] = 32'b00000000000000001101101011010100;
assign LUT_3[26929] = 32'b00000000000000010100010110110001;
assign LUT_3[26930] = 32'b00000000000000001111110010111000;
assign LUT_3[26931] = 32'b00000000000000010110011110010101;
assign LUT_3[26932] = 32'b00000000000000001010111001001010;
assign LUT_3[26933] = 32'b00000000000000010001100100100111;
assign LUT_3[26934] = 32'b00000000000000001101000000101110;
assign LUT_3[26935] = 32'b00000000000000010011101100001011;
assign LUT_3[26936] = 32'b00000000000000010011000100011010;
assign LUT_3[26937] = 32'b00000000000000011001101111110111;
assign LUT_3[26938] = 32'b00000000000000010101001011111110;
assign LUT_3[26939] = 32'b00000000000000011011110111011011;
assign LUT_3[26940] = 32'b00000000000000010000010010010000;
assign LUT_3[26941] = 32'b00000000000000010110111101101101;
assign LUT_3[26942] = 32'b00000000000000010010011001110100;
assign LUT_3[26943] = 32'b00000000000000011001000101010001;
assign LUT_3[26944] = 32'b00000000000000001001000010011100;
assign LUT_3[26945] = 32'b00000000000000001111101101111001;
assign LUT_3[26946] = 32'b00000000000000001011001010000000;
assign LUT_3[26947] = 32'b00000000000000010001110101011101;
assign LUT_3[26948] = 32'b00000000000000000110010000010010;
assign LUT_3[26949] = 32'b00000000000000001100111011101111;
assign LUT_3[26950] = 32'b00000000000000001000010111110110;
assign LUT_3[26951] = 32'b00000000000000001111000011010011;
assign LUT_3[26952] = 32'b00000000000000001110011011100010;
assign LUT_3[26953] = 32'b00000000000000010101000110111111;
assign LUT_3[26954] = 32'b00000000000000010000100011000110;
assign LUT_3[26955] = 32'b00000000000000010111001110100011;
assign LUT_3[26956] = 32'b00000000000000001011101001011000;
assign LUT_3[26957] = 32'b00000000000000010010010100110101;
assign LUT_3[26958] = 32'b00000000000000001101110000111100;
assign LUT_3[26959] = 32'b00000000000000010100011100011001;
assign LUT_3[26960] = 32'b00000000000000001100010101011111;
assign LUT_3[26961] = 32'b00000000000000010011000000111100;
assign LUT_3[26962] = 32'b00000000000000001110011101000011;
assign LUT_3[26963] = 32'b00000000000000010101001000100000;
assign LUT_3[26964] = 32'b00000000000000001001100011010101;
assign LUT_3[26965] = 32'b00000000000000010000001110110010;
assign LUT_3[26966] = 32'b00000000000000001011101010111001;
assign LUT_3[26967] = 32'b00000000000000010010010110010110;
assign LUT_3[26968] = 32'b00000000000000010001101110100101;
assign LUT_3[26969] = 32'b00000000000000011000011010000010;
assign LUT_3[26970] = 32'b00000000000000010011110110001001;
assign LUT_3[26971] = 32'b00000000000000011010100001100110;
assign LUT_3[26972] = 32'b00000000000000001110111100011011;
assign LUT_3[26973] = 32'b00000000000000010101100111111000;
assign LUT_3[26974] = 32'b00000000000000010001000011111111;
assign LUT_3[26975] = 32'b00000000000000010111101111011100;
assign LUT_3[26976] = 32'b00000000000000001010010000111100;
assign LUT_3[26977] = 32'b00000000000000010000111100011001;
assign LUT_3[26978] = 32'b00000000000000001100011000100000;
assign LUT_3[26979] = 32'b00000000000000010011000011111101;
assign LUT_3[26980] = 32'b00000000000000000111011110110010;
assign LUT_3[26981] = 32'b00000000000000001110001010001111;
assign LUT_3[26982] = 32'b00000000000000001001100110010110;
assign LUT_3[26983] = 32'b00000000000000010000010001110011;
assign LUT_3[26984] = 32'b00000000000000001111101010000010;
assign LUT_3[26985] = 32'b00000000000000010110010101011111;
assign LUT_3[26986] = 32'b00000000000000010001110001100110;
assign LUT_3[26987] = 32'b00000000000000011000011101000011;
assign LUT_3[26988] = 32'b00000000000000001100110111111000;
assign LUT_3[26989] = 32'b00000000000000010011100011010101;
assign LUT_3[26990] = 32'b00000000000000001110111111011100;
assign LUT_3[26991] = 32'b00000000000000010101101010111001;
assign LUT_3[26992] = 32'b00000000000000001101100011111111;
assign LUT_3[26993] = 32'b00000000000000010100001111011100;
assign LUT_3[26994] = 32'b00000000000000001111101011100011;
assign LUT_3[26995] = 32'b00000000000000010110010111000000;
assign LUT_3[26996] = 32'b00000000000000001010110001110101;
assign LUT_3[26997] = 32'b00000000000000010001011101010010;
assign LUT_3[26998] = 32'b00000000000000001100111001011001;
assign LUT_3[26999] = 32'b00000000000000010011100100110110;
assign LUT_3[27000] = 32'b00000000000000010010111101000101;
assign LUT_3[27001] = 32'b00000000000000011001101000100010;
assign LUT_3[27002] = 32'b00000000000000010101000100101001;
assign LUT_3[27003] = 32'b00000000000000011011110000000110;
assign LUT_3[27004] = 32'b00000000000000010000001010111011;
assign LUT_3[27005] = 32'b00000000000000010110110110011000;
assign LUT_3[27006] = 32'b00000000000000010010010010011111;
assign LUT_3[27007] = 32'b00000000000000011000111101111100;
assign LUT_3[27008] = 32'b00000000000000001011010100101111;
assign LUT_3[27009] = 32'b00000000000000010010000000001100;
assign LUT_3[27010] = 32'b00000000000000001101011100010011;
assign LUT_3[27011] = 32'b00000000000000010100000111110000;
assign LUT_3[27012] = 32'b00000000000000001000100010100101;
assign LUT_3[27013] = 32'b00000000000000001111001110000010;
assign LUT_3[27014] = 32'b00000000000000001010101010001001;
assign LUT_3[27015] = 32'b00000000000000010001010101100110;
assign LUT_3[27016] = 32'b00000000000000010000101101110101;
assign LUT_3[27017] = 32'b00000000000000010111011001010010;
assign LUT_3[27018] = 32'b00000000000000010010110101011001;
assign LUT_3[27019] = 32'b00000000000000011001100000110110;
assign LUT_3[27020] = 32'b00000000000000001101111011101011;
assign LUT_3[27021] = 32'b00000000000000010100100111001000;
assign LUT_3[27022] = 32'b00000000000000010000000011001111;
assign LUT_3[27023] = 32'b00000000000000010110101110101100;
assign LUT_3[27024] = 32'b00000000000000001110100111110010;
assign LUT_3[27025] = 32'b00000000000000010101010011001111;
assign LUT_3[27026] = 32'b00000000000000010000101111010110;
assign LUT_3[27027] = 32'b00000000000000010111011010110011;
assign LUT_3[27028] = 32'b00000000000000001011110101101000;
assign LUT_3[27029] = 32'b00000000000000010010100001000101;
assign LUT_3[27030] = 32'b00000000000000001101111101001100;
assign LUT_3[27031] = 32'b00000000000000010100101000101001;
assign LUT_3[27032] = 32'b00000000000000010100000000111000;
assign LUT_3[27033] = 32'b00000000000000011010101100010101;
assign LUT_3[27034] = 32'b00000000000000010110001000011100;
assign LUT_3[27035] = 32'b00000000000000011100110011111001;
assign LUT_3[27036] = 32'b00000000000000010001001110101110;
assign LUT_3[27037] = 32'b00000000000000010111111010001011;
assign LUT_3[27038] = 32'b00000000000000010011010110010010;
assign LUT_3[27039] = 32'b00000000000000011010000001101111;
assign LUT_3[27040] = 32'b00000000000000001100100011001111;
assign LUT_3[27041] = 32'b00000000000000010011001110101100;
assign LUT_3[27042] = 32'b00000000000000001110101010110011;
assign LUT_3[27043] = 32'b00000000000000010101010110010000;
assign LUT_3[27044] = 32'b00000000000000001001110001000101;
assign LUT_3[27045] = 32'b00000000000000010000011100100010;
assign LUT_3[27046] = 32'b00000000000000001011111000101001;
assign LUT_3[27047] = 32'b00000000000000010010100100000110;
assign LUT_3[27048] = 32'b00000000000000010001111100010101;
assign LUT_3[27049] = 32'b00000000000000011000100111110010;
assign LUT_3[27050] = 32'b00000000000000010100000011111001;
assign LUT_3[27051] = 32'b00000000000000011010101111010110;
assign LUT_3[27052] = 32'b00000000000000001111001010001011;
assign LUT_3[27053] = 32'b00000000000000010101110101101000;
assign LUT_3[27054] = 32'b00000000000000010001010001101111;
assign LUT_3[27055] = 32'b00000000000000010111111101001100;
assign LUT_3[27056] = 32'b00000000000000001111110110010010;
assign LUT_3[27057] = 32'b00000000000000010110100001101111;
assign LUT_3[27058] = 32'b00000000000000010001111101110110;
assign LUT_3[27059] = 32'b00000000000000011000101001010011;
assign LUT_3[27060] = 32'b00000000000000001101000100001000;
assign LUT_3[27061] = 32'b00000000000000010011101111100101;
assign LUT_3[27062] = 32'b00000000000000001111001011101100;
assign LUT_3[27063] = 32'b00000000000000010101110111001001;
assign LUT_3[27064] = 32'b00000000000000010101001111011000;
assign LUT_3[27065] = 32'b00000000000000011011111010110101;
assign LUT_3[27066] = 32'b00000000000000010111010110111100;
assign LUT_3[27067] = 32'b00000000000000011110000010011001;
assign LUT_3[27068] = 32'b00000000000000010010011101001110;
assign LUT_3[27069] = 32'b00000000000000011001001000101011;
assign LUT_3[27070] = 32'b00000000000000010100100100110010;
assign LUT_3[27071] = 32'b00000000000000011011010000001111;
assign LUT_3[27072] = 32'b00000000000000001011001101011010;
assign LUT_3[27073] = 32'b00000000000000010001111000110111;
assign LUT_3[27074] = 32'b00000000000000001101010100111110;
assign LUT_3[27075] = 32'b00000000000000010100000000011011;
assign LUT_3[27076] = 32'b00000000000000001000011011010000;
assign LUT_3[27077] = 32'b00000000000000001111000110101101;
assign LUT_3[27078] = 32'b00000000000000001010100010110100;
assign LUT_3[27079] = 32'b00000000000000010001001110010001;
assign LUT_3[27080] = 32'b00000000000000010000100110100000;
assign LUT_3[27081] = 32'b00000000000000010111010001111101;
assign LUT_3[27082] = 32'b00000000000000010010101110000100;
assign LUT_3[27083] = 32'b00000000000000011001011001100001;
assign LUT_3[27084] = 32'b00000000000000001101110100010110;
assign LUT_3[27085] = 32'b00000000000000010100011111110011;
assign LUT_3[27086] = 32'b00000000000000001111111011111010;
assign LUT_3[27087] = 32'b00000000000000010110100111010111;
assign LUT_3[27088] = 32'b00000000000000001110100000011101;
assign LUT_3[27089] = 32'b00000000000000010101001011111010;
assign LUT_3[27090] = 32'b00000000000000010000101000000001;
assign LUT_3[27091] = 32'b00000000000000010111010011011110;
assign LUT_3[27092] = 32'b00000000000000001011101110010011;
assign LUT_3[27093] = 32'b00000000000000010010011001110000;
assign LUT_3[27094] = 32'b00000000000000001101110101110111;
assign LUT_3[27095] = 32'b00000000000000010100100001010100;
assign LUT_3[27096] = 32'b00000000000000010011111001100011;
assign LUT_3[27097] = 32'b00000000000000011010100101000000;
assign LUT_3[27098] = 32'b00000000000000010110000001000111;
assign LUT_3[27099] = 32'b00000000000000011100101100100100;
assign LUT_3[27100] = 32'b00000000000000010001000111011001;
assign LUT_3[27101] = 32'b00000000000000010111110010110110;
assign LUT_3[27102] = 32'b00000000000000010011001110111101;
assign LUT_3[27103] = 32'b00000000000000011001111010011010;
assign LUT_3[27104] = 32'b00000000000000001100011011111010;
assign LUT_3[27105] = 32'b00000000000000010011000111010111;
assign LUT_3[27106] = 32'b00000000000000001110100011011110;
assign LUT_3[27107] = 32'b00000000000000010101001110111011;
assign LUT_3[27108] = 32'b00000000000000001001101001110000;
assign LUT_3[27109] = 32'b00000000000000010000010101001101;
assign LUT_3[27110] = 32'b00000000000000001011110001010100;
assign LUT_3[27111] = 32'b00000000000000010010011100110001;
assign LUT_3[27112] = 32'b00000000000000010001110101000000;
assign LUT_3[27113] = 32'b00000000000000011000100000011101;
assign LUT_3[27114] = 32'b00000000000000010011111100100100;
assign LUT_3[27115] = 32'b00000000000000011010101000000001;
assign LUT_3[27116] = 32'b00000000000000001111000010110110;
assign LUT_3[27117] = 32'b00000000000000010101101110010011;
assign LUT_3[27118] = 32'b00000000000000010001001010011010;
assign LUT_3[27119] = 32'b00000000000000010111110101110111;
assign LUT_3[27120] = 32'b00000000000000001111101110111101;
assign LUT_3[27121] = 32'b00000000000000010110011010011010;
assign LUT_3[27122] = 32'b00000000000000010001110110100001;
assign LUT_3[27123] = 32'b00000000000000011000100001111110;
assign LUT_3[27124] = 32'b00000000000000001100111100110011;
assign LUT_3[27125] = 32'b00000000000000010011101000010000;
assign LUT_3[27126] = 32'b00000000000000001111000100010111;
assign LUT_3[27127] = 32'b00000000000000010101101111110100;
assign LUT_3[27128] = 32'b00000000000000010101001000000011;
assign LUT_3[27129] = 32'b00000000000000011011110011100000;
assign LUT_3[27130] = 32'b00000000000000010111001111100111;
assign LUT_3[27131] = 32'b00000000000000011101111011000100;
assign LUT_3[27132] = 32'b00000000000000010010010101111001;
assign LUT_3[27133] = 32'b00000000000000011001000001010110;
assign LUT_3[27134] = 32'b00000000000000010100011101011101;
assign LUT_3[27135] = 32'b00000000000000011011001000111010;
assign LUT_3[27136] = 32'b00000000000000010000001111011100;
assign LUT_3[27137] = 32'b00000000000000010110111010111001;
assign LUT_3[27138] = 32'b00000000000000010010010111000000;
assign LUT_3[27139] = 32'b00000000000000011001000010011101;
assign LUT_3[27140] = 32'b00000000000000001101011101010010;
assign LUT_3[27141] = 32'b00000000000000010100001000101111;
assign LUT_3[27142] = 32'b00000000000000001111100100110110;
assign LUT_3[27143] = 32'b00000000000000010110010000010011;
assign LUT_3[27144] = 32'b00000000000000010101101000100010;
assign LUT_3[27145] = 32'b00000000000000011100010011111111;
assign LUT_3[27146] = 32'b00000000000000010111110000000110;
assign LUT_3[27147] = 32'b00000000000000011110011011100011;
assign LUT_3[27148] = 32'b00000000000000010010110110011000;
assign LUT_3[27149] = 32'b00000000000000011001100001110101;
assign LUT_3[27150] = 32'b00000000000000010100111101111100;
assign LUT_3[27151] = 32'b00000000000000011011101001011001;
assign LUT_3[27152] = 32'b00000000000000010011100010011111;
assign LUT_3[27153] = 32'b00000000000000011010001101111100;
assign LUT_3[27154] = 32'b00000000000000010101101010000011;
assign LUT_3[27155] = 32'b00000000000000011100010101100000;
assign LUT_3[27156] = 32'b00000000000000010000110000010101;
assign LUT_3[27157] = 32'b00000000000000010111011011110010;
assign LUT_3[27158] = 32'b00000000000000010010110111111001;
assign LUT_3[27159] = 32'b00000000000000011001100011010110;
assign LUT_3[27160] = 32'b00000000000000011000111011100101;
assign LUT_3[27161] = 32'b00000000000000011111100111000010;
assign LUT_3[27162] = 32'b00000000000000011011000011001001;
assign LUT_3[27163] = 32'b00000000000000100001101110100110;
assign LUT_3[27164] = 32'b00000000000000010110001001011011;
assign LUT_3[27165] = 32'b00000000000000011100110100111000;
assign LUT_3[27166] = 32'b00000000000000011000010000111111;
assign LUT_3[27167] = 32'b00000000000000011110111100011100;
assign LUT_3[27168] = 32'b00000000000000010001011101111100;
assign LUT_3[27169] = 32'b00000000000000011000001001011001;
assign LUT_3[27170] = 32'b00000000000000010011100101100000;
assign LUT_3[27171] = 32'b00000000000000011010010000111101;
assign LUT_3[27172] = 32'b00000000000000001110101011110010;
assign LUT_3[27173] = 32'b00000000000000010101010111001111;
assign LUT_3[27174] = 32'b00000000000000010000110011010110;
assign LUT_3[27175] = 32'b00000000000000010111011110110011;
assign LUT_3[27176] = 32'b00000000000000010110110111000010;
assign LUT_3[27177] = 32'b00000000000000011101100010011111;
assign LUT_3[27178] = 32'b00000000000000011000111110100110;
assign LUT_3[27179] = 32'b00000000000000011111101010000011;
assign LUT_3[27180] = 32'b00000000000000010100000100111000;
assign LUT_3[27181] = 32'b00000000000000011010110000010101;
assign LUT_3[27182] = 32'b00000000000000010110001100011100;
assign LUT_3[27183] = 32'b00000000000000011100110111111001;
assign LUT_3[27184] = 32'b00000000000000010100110000111111;
assign LUT_3[27185] = 32'b00000000000000011011011100011100;
assign LUT_3[27186] = 32'b00000000000000010110111000100011;
assign LUT_3[27187] = 32'b00000000000000011101100100000000;
assign LUT_3[27188] = 32'b00000000000000010001111110110101;
assign LUT_3[27189] = 32'b00000000000000011000101010010010;
assign LUT_3[27190] = 32'b00000000000000010100000110011001;
assign LUT_3[27191] = 32'b00000000000000011010110001110110;
assign LUT_3[27192] = 32'b00000000000000011010001010000101;
assign LUT_3[27193] = 32'b00000000000000100000110101100010;
assign LUT_3[27194] = 32'b00000000000000011100010001101001;
assign LUT_3[27195] = 32'b00000000000000100010111101000110;
assign LUT_3[27196] = 32'b00000000000000010111010111111011;
assign LUT_3[27197] = 32'b00000000000000011110000011011000;
assign LUT_3[27198] = 32'b00000000000000011001011111011111;
assign LUT_3[27199] = 32'b00000000000000100000001010111100;
assign LUT_3[27200] = 32'b00000000000000010000001000000111;
assign LUT_3[27201] = 32'b00000000000000010110110011100100;
assign LUT_3[27202] = 32'b00000000000000010010001111101011;
assign LUT_3[27203] = 32'b00000000000000011000111011001000;
assign LUT_3[27204] = 32'b00000000000000001101010101111101;
assign LUT_3[27205] = 32'b00000000000000010100000001011010;
assign LUT_3[27206] = 32'b00000000000000001111011101100001;
assign LUT_3[27207] = 32'b00000000000000010110001000111110;
assign LUT_3[27208] = 32'b00000000000000010101100001001101;
assign LUT_3[27209] = 32'b00000000000000011100001100101010;
assign LUT_3[27210] = 32'b00000000000000010111101000110001;
assign LUT_3[27211] = 32'b00000000000000011110010100001110;
assign LUT_3[27212] = 32'b00000000000000010010101111000011;
assign LUT_3[27213] = 32'b00000000000000011001011010100000;
assign LUT_3[27214] = 32'b00000000000000010100110110100111;
assign LUT_3[27215] = 32'b00000000000000011011100010000100;
assign LUT_3[27216] = 32'b00000000000000010011011011001010;
assign LUT_3[27217] = 32'b00000000000000011010000110100111;
assign LUT_3[27218] = 32'b00000000000000010101100010101110;
assign LUT_3[27219] = 32'b00000000000000011100001110001011;
assign LUT_3[27220] = 32'b00000000000000010000101001000000;
assign LUT_3[27221] = 32'b00000000000000010111010100011101;
assign LUT_3[27222] = 32'b00000000000000010010110000100100;
assign LUT_3[27223] = 32'b00000000000000011001011100000001;
assign LUT_3[27224] = 32'b00000000000000011000110100010000;
assign LUT_3[27225] = 32'b00000000000000011111011111101101;
assign LUT_3[27226] = 32'b00000000000000011010111011110100;
assign LUT_3[27227] = 32'b00000000000000100001100111010001;
assign LUT_3[27228] = 32'b00000000000000010110000010000110;
assign LUT_3[27229] = 32'b00000000000000011100101101100011;
assign LUT_3[27230] = 32'b00000000000000011000001001101010;
assign LUT_3[27231] = 32'b00000000000000011110110101000111;
assign LUT_3[27232] = 32'b00000000000000010001010110100111;
assign LUT_3[27233] = 32'b00000000000000011000000010000100;
assign LUT_3[27234] = 32'b00000000000000010011011110001011;
assign LUT_3[27235] = 32'b00000000000000011010001001101000;
assign LUT_3[27236] = 32'b00000000000000001110100100011101;
assign LUT_3[27237] = 32'b00000000000000010101001111111010;
assign LUT_3[27238] = 32'b00000000000000010000101100000001;
assign LUT_3[27239] = 32'b00000000000000010111010111011110;
assign LUT_3[27240] = 32'b00000000000000010110101111101101;
assign LUT_3[27241] = 32'b00000000000000011101011011001010;
assign LUT_3[27242] = 32'b00000000000000011000110111010001;
assign LUT_3[27243] = 32'b00000000000000011111100010101110;
assign LUT_3[27244] = 32'b00000000000000010011111101100011;
assign LUT_3[27245] = 32'b00000000000000011010101001000000;
assign LUT_3[27246] = 32'b00000000000000010110000101000111;
assign LUT_3[27247] = 32'b00000000000000011100110000100100;
assign LUT_3[27248] = 32'b00000000000000010100101001101010;
assign LUT_3[27249] = 32'b00000000000000011011010101000111;
assign LUT_3[27250] = 32'b00000000000000010110110001001110;
assign LUT_3[27251] = 32'b00000000000000011101011100101011;
assign LUT_3[27252] = 32'b00000000000000010001110111100000;
assign LUT_3[27253] = 32'b00000000000000011000100010111101;
assign LUT_3[27254] = 32'b00000000000000010011111111000100;
assign LUT_3[27255] = 32'b00000000000000011010101010100001;
assign LUT_3[27256] = 32'b00000000000000011010000010110000;
assign LUT_3[27257] = 32'b00000000000000100000101110001101;
assign LUT_3[27258] = 32'b00000000000000011100001010010100;
assign LUT_3[27259] = 32'b00000000000000100010110101110001;
assign LUT_3[27260] = 32'b00000000000000010111010000100110;
assign LUT_3[27261] = 32'b00000000000000011101111100000011;
assign LUT_3[27262] = 32'b00000000000000011001011000001010;
assign LUT_3[27263] = 32'b00000000000000100000000011100111;
assign LUT_3[27264] = 32'b00000000000000010010011010011010;
assign LUT_3[27265] = 32'b00000000000000011001000101110111;
assign LUT_3[27266] = 32'b00000000000000010100100001111110;
assign LUT_3[27267] = 32'b00000000000000011011001101011011;
assign LUT_3[27268] = 32'b00000000000000001111101000010000;
assign LUT_3[27269] = 32'b00000000000000010110010011101101;
assign LUT_3[27270] = 32'b00000000000000010001101111110100;
assign LUT_3[27271] = 32'b00000000000000011000011011010001;
assign LUT_3[27272] = 32'b00000000000000010111110011100000;
assign LUT_3[27273] = 32'b00000000000000011110011110111101;
assign LUT_3[27274] = 32'b00000000000000011001111011000100;
assign LUT_3[27275] = 32'b00000000000000100000100110100001;
assign LUT_3[27276] = 32'b00000000000000010101000001010110;
assign LUT_3[27277] = 32'b00000000000000011011101100110011;
assign LUT_3[27278] = 32'b00000000000000010111001000111010;
assign LUT_3[27279] = 32'b00000000000000011101110100010111;
assign LUT_3[27280] = 32'b00000000000000010101101101011101;
assign LUT_3[27281] = 32'b00000000000000011100011000111010;
assign LUT_3[27282] = 32'b00000000000000010111110101000001;
assign LUT_3[27283] = 32'b00000000000000011110100000011110;
assign LUT_3[27284] = 32'b00000000000000010010111011010011;
assign LUT_3[27285] = 32'b00000000000000011001100110110000;
assign LUT_3[27286] = 32'b00000000000000010101000010110111;
assign LUT_3[27287] = 32'b00000000000000011011101110010100;
assign LUT_3[27288] = 32'b00000000000000011011000110100011;
assign LUT_3[27289] = 32'b00000000000000100001110010000000;
assign LUT_3[27290] = 32'b00000000000000011101001110000111;
assign LUT_3[27291] = 32'b00000000000000100011111001100100;
assign LUT_3[27292] = 32'b00000000000000011000010100011001;
assign LUT_3[27293] = 32'b00000000000000011110111111110110;
assign LUT_3[27294] = 32'b00000000000000011010011011111101;
assign LUT_3[27295] = 32'b00000000000000100001000111011010;
assign LUT_3[27296] = 32'b00000000000000010011101000111010;
assign LUT_3[27297] = 32'b00000000000000011010010100010111;
assign LUT_3[27298] = 32'b00000000000000010101110000011110;
assign LUT_3[27299] = 32'b00000000000000011100011011111011;
assign LUT_3[27300] = 32'b00000000000000010000110110110000;
assign LUT_3[27301] = 32'b00000000000000010111100010001101;
assign LUT_3[27302] = 32'b00000000000000010010111110010100;
assign LUT_3[27303] = 32'b00000000000000011001101001110001;
assign LUT_3[27304] = 32'b00000000000000011001000010000000;
assign LUT_3[27305] = 32'b00000000000000011111101101011101;
assign LUT_3[27306] = 32'b00000000000000011011001001100100;
assign LUT_3[27307] = 32'b00000000000000100001110101000001;
assign LUT_3[27308] = 32'b00000000000000010110001111110110;
assign LUT_3[27309] = 32'b00000000000000011100111011010011;
assign LUT_3[27310] = 32'b00000000000000011000010111011010;
assign LUT_3[27311] = 32'b00000000000000011111000010110111;
assign LUT_3[27312] = 32'b00000000000000010110111011111101;
assign LUT_3[27313] = 32'b00000000000000011101100111011010;
assign LUT_3[27314] = 32'b00000000000000011001000011100001;
assign LUT_3[27315] = 32'b00000000000000011111101110111110;
assign LUT_3[27316] = 32'b00000000000000010100001001110011;
assign LUT_3[27317] = 32'b00000000000000011010110101010000;
assign LUT_3[27318] = 32'b00000000000000010110010001010111;
assign LUT_3[27319] = 32'b00000000000000011100111100110100;
assign LUT_3[27320] = 32'b00000000000000011100010101000011;
assign LUT_3[27321] = 32'b00000000000000100011000000100000;
assign LUT_3[27322] = 32'b00000000000000011110011100100111;
assign LUT_3[27323] = 32'b00000000000000100101001000000100;
assign LUT_3[27324] = 32'b00000000000000011001100010111001;
assign LUT_3[27325] = 32'b00000000000000100000001110010110;
assign LUT_3[27326] = 32'b00000000000000011011101010011101;
assign LUT_3[27327] = 32'b00000000000000100010010101111010;
assign LUT_3[27328] = 32'b00000000000000010010010011000101;
assign LUT_3[27329] = 32'b00000000000000011000111110100010;
assign LUT_3[27330] = 32'b00000000000000010100011010101001;
assign LUT_3[27331] = 32'b00000000000000011011000110000110;
assign LUT_3[27332] = 32'b00000000000000001111100000111011;
assign LUT_3[27333] = 32'b00000000000000010110001100011000;
assign LUT_3[27334] = 32'b00000000000000010001101000011111;
assign LUT_3[27335] = 32'b00000000000000011000010011111100;
assign LUT_3[27336] = 32'b00000000000000010111101100001011;
assign LUT_3[27337] = 32'b00000000000000011110010111101000;
assign LUT_3[27338] = 32'b00000000000000011001110011101111;
assign LUT_3[27339] = 32'b00000000000000100000011111001100;
assign LUT_3[27340] = 32'b00000000000000010100111010000001;
assign LUT_3[27341] = 32'b00000000000000011011100101011110;
assign LUT_3[27342] = 32'b00000000000000010111000001100101;
assign LUT_3[27343] = 32'b00000000000000011101101101000010;
assign LUT_3[27344] = 32'b00000000000000010101100110001000;
assign LUT_3[27345] = 32'b00000000000000011100010001100101;
assign LUT_3[27346] = 32'b00000000000000010111101101101100;
assign LUT_3[27347] = 32'b00000000000000011110011001001001;
assign LUT_3[27348] = 32'b00000000000000010010110011111110;
assign LUT_3[27349] = 32'b00000000000000011001011111011011;
assign LUT_3[27350] = 32'b00000000000000010100111011100010;
assign LUT_3[27351] = 32'b00000000000000011011100110111111;
assign LUT_3[27352] = 32'b00000000000000011010111111001110;
assign LUT_3[27353] = 32'b00000000000000100001101010101011;
assign LUT_3[27354] = 32'b00000000000000011101000110110010;
assign LUT_3[27355] = 32'b00000000000000100011110010001111;
assign LUT_3[27356] = 32'b00000000000000011000001101000100;
assign LUT_3[27357] = 32'b00000000000000011110111000100001;
assign LUT_3[27358] = 32'b00000000000000011010010100101000;
assign LUT_3[27359] = 32'b00000000000000100001000000000101;
assign LUT_3[27360] = 32'b00000000000000010011100001100101;
assign LUT_3[27361] = 32'b00000000000000011010001101000010;
assign LUT_3[27362] = 32'b00000000000000010101101001001001;
assign LUT_3[27363] = 32'b00000000000000011100010100100110;
assign LUT_3[27364] = 32'b00000000000000010000101111011011;
assign LUT_3[27365] = 32'b00000000000000010111011010111000;
assign LUT_3[27366] = 32'b00000000000000010010110110111111;
assign LUT_3[27367] = 32'b00000000000000011001100010011100;
assign LUT_3[27368] = 32'b00000000000000011000111010101011;
assign LUT_3[27369] = 32'b00000000000000011111100110001000;
assign LUT_3[27370] = 32'b00000000000000011011000010001111;
assign LUT_3[27371] = 32'b00000000000000100001101101101100;
assign LUT_3[27372] = 32'b00000000000000010110001000100001;
assign LUT_3[27373] = 32'b00000000000000011100110011111110;
assign LUT_3[27374] = 32'b00000000000000011000010000000101;
assign LUT_3[27375] = 32'b00000000000000011110111011100010;
assign LUT_3[27376] = 32'b00000000000000010110110100101000;
assign LUT_3[27377] = 32'b00000000000000011101100000000101;
assign LUT_3[27378] = 32'b00000000000000011000111100001100;
assign LUT_3[27379] = 32'b00000000000000011111100111101001;
assign LUT_3[27380] = 32'b00000000000000010100000010011110;
assign LUT_3[27381] = 32'b00000000000000011010101101111011;
assign LUT_3[27382] = 32'b00000000000000010110001010000010;
assign LUT_3[27383] = 32'b00000000000000011100110101011111;
assign LUT_3[27384] = 32'b00000000000000011100001101101110;
assign LUT_3[27385] = 32'b00000000000000100010111001001011;
assign LUT_3[27386] = 32'b00000000000000011110010101010010;
assign LUT_3[27387] = 32'b00000000000000100101000000101111;
assign LUT_3[27388] = 32'b00000000000000011001011011100100;
assign LUT_3[27389] = 32'b00000000000000100000000111000001;
assign LUT_3[27390] = 32'b00000000000000011011100011001000;
assign LUT_3[27391] = 32'b00000000000000100010001110100101;
assign LUT_3[27392] = 32'b00000000000000001100011110111101;
assign LUT_3[27393] = 32'b00000000000000010011001010011010;
assign LUT_3[27394] = 32'b00000000000000001110100110100001;
assign LUT_3[27395] = 32'b00000000000000010101010001111110;
assign LUT_3[27396] = 32'b00000000000000001001101100110011;
assign LUT_3[27397] = 32'b00000000000000010000011000010000;
assign LUT_3[27398] = 32'b00000000000000001011110100010111;
assign LUT_3[27399] = 32'b00000000000000010010011111110100;
assign LUT_3[27400] = 32'b00000000000000010001111000000011;
assign LUT_3[27401] = 32'b00000000000000011000100011100000;
assign LUT_3[27402] = 32'b00000000000000010011111111100111;
assign LUT_3[27403] = 32'b00000000000000011010101011000100;
assign LUT_3[27404] = 32'b00000000000000001111000101111001;
assign LUT_3[27405] = 32'b00000000000000010101110001010110;
assign LUT_3[27406] = 32'b00000000000000010001001101011101;
assign LUT_3[27407] = 32'b00000000000000010111111000111010;
assign LUT_3[27408] = 32'b00000000000000001111110010000000;
assign LUT_3[27409] = 32'b00000000000000010110011101011101;
assign LUT_3[27410] = 32'b00000000000000010001111001100100;
assign LUT_3[27411] = 32'b00000000000000011000100101000001;
assign LUT_3[27412] = 32'b00000000000000001100111111110110;
assign LUT_3[27413] = 32'b00000000000000010011101011010011;
assign LUT_3[27414] = 32'b00000000000000001111000111011010;
assign LUT_3[27415] = 32'b00000000000000010101110010110111;
assign LUT_3[27416] = 32'b00000000000000010101001011000110;
assign LUT_3[27417] = 32'b00000000000000011011110110100011;
assign LUT_3[27418] = 32'b00000000000000010111010010101010;
assign LUT_3[27419] = 32'b00000000000000011101111110000111;
assign LUT_3[27420] = 32'b00000000000000010010011000111100;
assign LUT_3[27421] = 32'b00000000000000011001000100011001;
assign LUT_3[27422] = 32'b00000000000000010100100000100000;
assign LUT_3[27423] = 32'b00000000000000011011001011111101;
assign LUT_3[27424] = 32'b00000000000000001101101101011101;
assign LUT_3[27425] = 32'b00000000000000010100011000111010;
assign LUT_3[27426] = 32'b00000000000000001111110101000001;
assign LUT_3[27427] = 32'b00000000000000010110100000011110;
assign LUT_3[27428] = 32'b00000000000000001010111011010011;
assign LUT_3[27429] = 32'b00000000000000010001100110110000;
assign LUT_3[27430] = 32'b00000000000000001101000010110111;
assign LUT_3[27431] = 32'b00000000000000010011101110010100;
assign LUT_3[27432] = 32'b00000000000000010011000110100011;
assign LUT_3[27433] = 32'b00000000000000011001110010000000;
assign LUT_3[27434] = 32'b00000000000000010101001110000111;
assign LUT_3[27435] = 32'b00000000000000011011111001100100;
assign LUT_3[27436] = 32'b00000000000000010000010100011001;
assign LUT_3[27437] = 32'b00000000000000010110111111110110;
assign LUT_3[27438] = 32'b00000000000000010010011011111101;
assign LUT_3[27439] = 32'b00000000000000011001000111011010;
assign LUT_3[27440] = 32'b00000000000000010001000000100000;
assign LUT_3[27441] = 32'b00000000000000010111101011111101;
assign LUT_3[27442] = 32'b00000000000000010011001000000100;
assign LUT_3[27443] = 32'b00000000000000011001110011100001;
assign LUT_3[27444] = 32'b00000000000000001110001110010110;
assign LUT_3[27445] = 32'b00000000000000010100111001110011;
assign LUT_3[27446] = 32'b00000000000000010000010101111010;
assign LUT_3[27447] = 32'b00000000000000010111000001010111;
assign LUT_3[27448] = 32'b00000000000000010110011001100110;
assign LUT_3[27449] = 32'b00000000000000011101000101000011;
assign LUT_3[27450] = 32'b00000000000000011000100001001010;
assign LUT_3[27451] = 32'b00000000000000011111001100100111;
assign LUT_3[27452] = 32'b00000000000000010011100111011100;
assign LUT_3[27453] = 32'b00000000000000011010010010111001;
assign LUT_3[27454] = 32'b00000000000000010101101111000000;
assign LUT_3[27455] = 32'b00000000000000011100011010011101;
assign LUT_3[27456] = 32'b00000000000000001100010111101000;
assign LUT_3[27457] = 32'b00000000000000010011000011000101;
assign LUT_3[27458] = 32'b00000000000000001110011111001100;
assign LUT_3[27459] = 32'b00000000000000010101001010101001;
assign LUT_3[27460] = 32'b00000000000000001001100101011110;
assign LUT_3[27461] = 32'b00000000000000010000010000111011;
assign LUT_3[27462] = 32'b00000000000000001011101101000010;
assign LUT_3[27463] = 32'b00000000000000010010011000011111;
assign LUT_3[27464] = 32'b00000000000000010001110000101110;
assign LUT_3[27465] = 32'b00000000000000011000011100001011;
assign LUT_3[27466] = 32'b00000000000000010011111000010010;
assign LUT_3[27467] = 32'b00000000000000011010100011101111;
assign LUT_3[27468] = 32'b00000000000000001110111110100100;
assign LUT_3[27469] = 32'b00000000000000010101101010000001;
assign LUT_3[27470] = 32'b00000000000000010001000110001000;
assign LUT_3[27471] = 32'b00000000000000010111110001100101;
assign LUT_3[27472] = 32'b00000000000000001111101010101011;
assign LUT_3[27473] = 32'b00000000000000010110010110001000;
assign LUT_3[27474] = 32'b00000000000000010001110010001111;
assign LUT_3[27475] = 32'b00000000000000011000011101101100;
assign LUT_3[27476] = 32'b00000000000000001100111000100001;
assign LUT_3[27477] = 32'b00000000000000010011100011111110;
assign LUT_3[27478] = 32'b00000000000000001111000000000101;
assign LUT_3[27479] = 32'b00000000000000010101101011100010;
assign LUT_3[27480] = 32'b00000000000000010101000011110001;
assign LUT_3[27481] = 32'b00000000000000011011101111001110;
assign LUT_3[27482] = 32'b00000000000000010111001011010101;
assign LUT_3[27483] = 32'b00000000000000011101110110110010;
assign LUT_3[27484] = 32'b00000000000000010010010001100111;
assign LUT_3[27485] = 32'b00000000000000011000111101000100;
assign LUT_3[27486] = 32'b00000000000000010100011001001011;
assign LUT_3[27487] = 32'b00000000000000011011000100101000;
assign LUT_3[27488] = 32'b00000000000000001101100110001000;
assign LUT_3[27489] = 32'b00000000000000010100010001100101;
assign LUT_3[27490] = 32'b00000000000000001111101101101100;
assign LUT_3[27491] = 32'b00000000000000010110011001001001;
assign LUT_3[27492] = 32'b00000000000000001010110011111110;
assign LUT_3[27493] = 32'b00000000000000010001011111011011;
assign LUT_3[27494] = 32'b00000000000000001100111011100010;
assign LUT_3[27495] = 32'b00000000000000010011100110111111;
assign LUT_3[27496] = 32'b00000000000000010010111111001110;
assign LUT_3[27497] = 32'b00000000000000011001101010101011;
assign LUT_3[27498] = 32'b00000000000000010101000110110010;
assign LUT_3[27499] = 32'b00000000000000011011110010001111;
assign LUT_3[27500] = 32'b00000000000000010000001101000100;
assign LUT_3[27501] = 32'b00000000000000010110111000100001;
assign LUT_3[27502] = 32'b00000000000000010010010100101000;
assign LUT_3[27503] = 32'b00000000000000011001000000000101;
assign LUT_3[27504] = 32'b00000000000000010000111001001011;
assign LUT_3[27505] = 32'b00000000000000010111100100101000;
assign LUT_3[27506] = 32'b00000000000000010011000000101111;
assign LUT_3[27507] = 32'b00000000000000011001101100001100;
assign LUT_3[27508] = 32'b00000000000000001110000111000001;
assign LUT_3[27509] = 32'b00000000000000010100110010011110;
assign LUT_3[27510] = 32'b00000000000000010000001110100101;
assign LUT_3[27511] = 32'b00000000000000010110111010000010;
assign LUT_3[27512] = 32'b00000000000000010110010010010001;
assign LUT_3[27513] = 32'b00000000000000011100111101101110;
assign LUT_3[27514] = 32'b00000000000000011000011001110101;
assign LUT_3[27515] = 32'b00000000000000011111000101010010;
assign LUT_3[27516] = 32'b00000000000000010011100000000111;
assign LUT_3[27517] = 32'b00000000000000011010001011100100;
assign LUT_3[27518] = 32'b00000000000000010101100111101011;
assign LUT_3[27519] = 32'b00000000000000011100010011001000;
assign LUT_3[27520] = 32'b00000000000000001110101001111011;
assign LUT_3[27521] = 32'b00000000000000010101010101011000;
assign LUT_3[27522] = 32'b00000000000000010000110001011111;
assign LUT_3[27523] = 32'b00000000000000010111011100111100;
assign LUT_3[27524] = 32'b00000000000000001011110111110001;
assign LUT_3[27525] = 32'b00000000000000010010100011001110;
assign LUT_3[27526] = 32'b00000000000000001101111111010101;
assign LUT_3[27527] = 32'b00000000000000010100101010110010;
assign LUT_3[27528] = 32'b00000000000000010100000011000001;
assign LUT_3[27529] = 32'b00000000000000011010101110011110;
assign LUT_3[27530] = 32'b00000000000000010110001010100101;
assign LUT_3[27531] = 32'b00000000000000011100110110000010;
assign LUT_3[27532] = 32'b00000000000000010001010000110111;
assign LUT_3[27533] = 32'b00000000000000010111111100010100;
assign LUT_3[27534] = 32'b00000000000000010011011000011011;
assign LUT_3[27535] = 32'b00000000000000011010000011111000;
assign LUT_3[27536] = 32'b00000000000000010001111100111110;
assign LUT_3[27537] = 32'b00000000000000011000101000011011;
assign LUT_3[27538] = 32'b00000000000000010100000100100010;
assign LUT_3[27539] = 32'b00000000000000011010101111111111;
assign LUT_3[27540] = 32'b00000000000000001111001010110100;
assign LUT_3[27541] = 32'b00000000000000010101110110010001;
assign LUT_3[27542] = 32'b00000000000000010001010010011000;
assign LUT_3[27543] = 32'b00000000000000010111111101110101;
assign LUT_3[27544] = 32'b00000000000000010111010110000100;
assign LUT_3[27545] = 32'b00000000000000011110000001100001;
assign LUT_3[27546] = 32'b00000000000000011001011101101000;
assign LUT_3[27547] = 32'b00000000000000100000001001000101;
assign LUT_3[27548] = 32'b00000000000000010100100011111010;
assign LUT_3[27549] = 32'b00000000000000011011001111010111;
assign LUT_3[27550] = 32'b00000000000000010110101011011110;
assign LUT_3[27551] = 32'b00000000000000011101010110111011;
assign LUT_3[27552] = 32'b00000000000000001111111000011011;
assign LUT_3[27553] = 32'b00000000000000010110100011111000;
assign LUT_3[27554] = 32'b00000000000000010001111111111111;
assign LUT_3[27555] = 32'b00000000000000011000101011011100;
assign LUT_3[27556] = 32'b00000000000000001101000110010001;
assign LUT_3[27557] = 32'b00000000000000010011110001101110;
assign LUT_3[27558] = 32'b00000000000000001111001101110101;
assign LUT_3[27559] = 32'b00000000000000010101111001010010;
assign LUT_3[27560] = 32'b00000000000000010101010001100001;
assign LUT_3[27561] = 32'b00000000000000011011111100111110;
assign LUT_3[27562] = 32'b00000000000000010111011001000101;
assign LUT_3[27563] = 32'b00000000000000011110000100100010;
assign LUT_3[27564] = 32'b00000000000000010010011111010111;
assign LUT_3[27565] = 32'b00000000000000011001001010110100;
assign LUT_3[27566] = 32'b00000000000000010100100110111011;
assign LUT_3[27567] = 32'b00000000000000011011010010011000;
assign LUT_3[27568] = 32'b00000000000000010011001011011110;
assign LUT_3[27569] = 32'b00000000000000011001110110111011;
assign LUT_3[27570] = 32'b00000000000000010101010011000010;
assign LUT_3[27571] = 32'b00000000000000011011111110011111;
assign LUT_3[27572] = 32'b00000000000000010000011001010100;
assign LUT_3[27573] = 32'b00000000000000010111000100110001;
assign LUT_3[27574] = 32'b00000000000000010010100000111000;
assign LUT_3[27575] = 32'b00000000000000011001001100010101;
assign LUT_3[27576] = 32'b00000000000000011000100100100100;
assign LUT_3[27577] = 32'b00000000000000011111010000000001;
assign LUT_3[27578] = 32'b00000000000000011010101100001000;
assign LUT_3[27579] = 32'b00000000000000100001010111100101;
assign LUT_3[27580] = 32'b00000000000000010101110010011010;
assign LUT_3[27581] = 32'b00000000000000011100011101110111;
assign LUT_3[27582] = 32'b00000000000000010111111001111110;
assign LUT_3[27583] = 32'b00000000000000011110100101011011;
assign LUT_3[27584] = 32'b00000000000000001110100010100110;
assign LUT_3[27585] = 32'b00000000000000010101001110000011;
assign LUT_3[27586] = 32'b00000000000000010000101010001010;
assign LUT_3[27587] = 32'b00000000000000010111010101100111;
assign LUT_3[27588] = 32'b00000000000000001011110000011100;
assign LUT_3[27589] = 32'b00000000000000010010011011111001;
assign LUT_3[27590] = 32'b00000000000000001101111000000000;
assign LUT_3[27591] = 32'b00000000000000010100100011011101;
assign LUT_3[27592] = 32'b00000000000000010011111011101100;
assign LUT_3[27593] = 32'b00000000000000011010100111001001;
assign LUT_3[27594] = 32'b00000000000000010110000011010000;
assign LUT_3[27595] = 32'b00000000000000011100101110101101;
assign LUT_3[27596] = 32'b00000000000000010001001001100010;
assign LUT_3[27597] = 32'b00000000000000010111110100111111;
assign LUT_3[27598] = 32'b00000000000000010011010001000110;
assign LUT_3[27599] = 32'b00000000000000011001111100100011;
assign LUT_3[27600] = 32'b00000000000000010001110101101001;
assign LUT_3[27601] = 32'b00000000000000011000100001000110;
assign LUT_3[27602] = 32'b00000000000000010011111101001101;
assign LUT_3[27603] = 32'b00000000000000011010101000101010;
assign LUT_3[27604] = 32'b00000000000000001111000011011111;
assign LUT_3[27605] = 32'b00000000000000010101101110111100;
assign LUT_3[27606] = 32'b00000000000000010001001011000011;
assign LUT_3[27607] = 32'b00000000000000010111110110100000;
assign LUT_3[27608] = 32'b00000000000000010111001110101111;
assign LUT_3[27609] = 32'b00000000000000011101111010001100;
assign LUT_3[27610] = 32'b00000000000000011001010110010011;
assign LUT_3[27611] = 32'b00000000000000100000000001110000;
assign LUT_3[27612] = 32'b00000000000000010100011100100101;
assign LUT_3[27613] = 32'b00000000000000011011001000000010;
assign LUT_3[27614] = 32'b00000000000000010110100100001001;
assign LUT_3[27615] = 32'b00000000000000011101001111100110;
assign LUT_3[27616] = 32'b00000000000000001111110001000110;
assign LUT_3[27617] = 32'b00000000000000010110011100100011;
assign LUT_3[27618] = 32'b00000000000000010001111000101010;
assign LUT_3[27619] = 32'b00000000000000011000100100000111;
assign LUT_3[27620] = 32'b00000000000000001100111110111100;
assign LUT_3[27621] = 32'b00000000000000010011101010011001;
assign LUT_3[27622] = 32'b00000000000000001111000110100000;
assign LUT_3[27623] = 32'b00000000000000010101110001111101;
assign LUT_3[27624] = 32'b00000000000000010101001010001100;
assign LUT_3[27625] = 32'b00000000000000011011110101101001;
assign LUT_3[27626] = 32'b00000000000000010111010001110000;
assign LUT_3[27627] = 32'b00000000000000011101111101001101;
assign LUT_3[27628] = 32'b00000000000000010010011000000010;
assign LUT_3[27629] = 32'b00000000000000011001000011011111;
assign LUT_3[27630] = 32'b00000000000000010100011111100110;
assign LUT_3[27631] = 32'b00000000000000011011001011000011;
assign LUT_3[27632] = 32'b00000000000000010011000100001001;
assign LUT_3[27633] = 32'b00000000000000011001101111100110;
assign LUT_3[27634] = 32'b00000000000000010101001011101101;
assign LUT_3[27635] = 32'b00000000000000011011110111001010;
assign LUT_3[27636] = 32'b00000000000000010000010001111111;
assign LUT_3[27637] = 32'b00000000000000010110111101011100;
assign LUT_3[27638] = 32'b00000000000000010010011001100011;
assign LUT_3[27639] = 32'b00000000000000011001000101000000;
assign LUT_3[27640] = 32'b00000000000000011000011101001111;
assign LUT_3[27641] = 32'b00000000000000011111001000101100;
assign LUT_3[27642] = 32'b00000000000000011010100100110011;
assign LUT_3[27643] = 32'b00000000000000100001010000010000;
assign LUT_3[27644] = 32'b00000000000000010101101011000101;
assign LUT_3[27645] = 32'b00000000000000011100010110100010;
assign LUT_3[27646] = 32'b00000000000000010111110010101001;
assign LUT_3[27647] = 32'b00000000000000011110011110000110;
assign LUT_3[27648] = 32'b00000000000000010011011111001101;
assign LUT_3[27649] = 32'b00000000000000011010001010101010;
assign LUT_3[27650] = 32'b00000000000000010101100110110001;
assign LUT_3[27651] = 32'b00000000000000011100010010001110;
assign LUT_3[27652] = 32'b00000000000000010000101101000011;
assign LUT_3[27653] = 32'b00000000000000010111011000100000;
assign LUT_3[27654] = 32'b00000000000000010010110100100111;
assign LUT_3[27655] = 32'b00000000000000011001100000000100;
assign LUT_3[27656] = 32'b00000000000000011000111000010011;
assign LUT_3[27657] = 32'b00000000000000011111100011110000;
assign LUT_3[27658] = 32'b00000000000000011010111111110111;
assign LUT_3[27659] = 32'b00000000000000100001101011010100;
assign LUT_3[27660] = 32'b00000000000000010110000110001001;
assign LUT_3[27661] = 32'b00000000000000011100110001100110;
assign LUT_3[27662] = 32'b00000000000000011000001101101101;
assign LUT_3[27663] = 32'b00000000000000011110111001001010;
assign LUT_3[27664] = 32'b00000000000000010110110010010000;
assign LUT_3[27665] = 32'b00000000000000011101011101101101;
assign LUT_3[27666] = 32'b00000000000000011000111001110100;
assign LUT_3[27667] = 32'b00000000000000011111100101010001;
assign LUT_3[27668] = 32'b00000000000000010100000000000110;
assign LUT_3[27669] = 32'b00000000000000011010101011100011;
assign LUT_3[27670] = 32'b00000000000000010110000111101010;
assign LUT_3[27671] = 32'b00000000000000011100110011000111;
assign LUT_3[27672] = 32'b00000000000000011100001011010110;
assign LUT_3[27673] = 32'b00000000000000100010110110110011;
assign LUT_3[27674] = 32'b00000000000000011110010010111010;
assign LUT_3[27675] = 32'b00000000000000100100111110010111;
assign LUT_3[27676] = 32'b00000000000000011001011001001100;
assign LUT_3[27677] = 32'b00000000000000100000000100101001;
assign LUT_3[27678] = 32'b00000000000000011011100000110000;
assign LUT_3[27679] = 32'b00000000000000100010001100001101;
assign LUT_3[27680] = 32'b00000000000000010100101101101101;
assign LUT_3[27681] = 32'b00000000000000011011011001001010;
assign LUT_3[27682] = 32'b00000000000000010110110101010001;
assign LUT_3[27683] = 32'b00000000000000011101100000101110;
assign LUT_3[27684] = 32'b00000000000000010001111011100011;
assign LUT_3[27685] = 32'b00000000000000011000100111000000;
assign LUT_3[27686] = 32'b00000000000000010100000011000111;
assign LUT_3[27687] = 32'b00000000000000011010101110100100;
assign LUT_3[27688] = 32'b00000000000000011010000110110011;
assign LUT_3[27689] = 32'b00000000000000100000110010010000;
assign LUT_3[27690] = 32'b00000000000000011100001110010111;
assign LUT_3[27691] = 32'b00000000000000100010111001110100;
assign LUT_3[27692] = 32'b00000000000000010111010100101001;
assign LUT_3[27693] = 32'b00000000000000011110000000000110;
assign LUT_3[27694] = 32'b00000000000000011001011100001101;
assign LUT_3[27695] = 32'b00000000000000100000000111101010;
assign LUT_3[27696] = 32'b00000000000000011000000000110000;
assign LUT_3[27697] = 32'b00000000000000011110101100001101;
assign LUT_3[27698] = 32'b00000000000000011010001000010100;
assign LUT_3[27699] = 32'b00000000000000100000110011110001;
assign LUT_3[27700] = 32'b00000000000000010101001110100110;
assign LUT_3[27701] = 32'b00000000000000011011111010000011;
assign LUT_3[27702] = 32'b00000000000000010111010110001010;
assign LUT_3[27703] = 32'b00000000000000011110000001100111;
assign LUT_3[27704] = 32'b00000000000000011101011001110110;
assign LUT_3[27705] = 32'b00000000000000100100000101010011;
assign LUT_3[27706] = 32'b00000000000000011111100001011010;
assign LUT_3[27707] = 32'b00000000000000100110001100110111;
assign LUT_3[27708] = 32'b00000000000000011010100111101100;
assign LUT_3[27709] = 32'b00000000000000100001010011001001;
assign LUT_3[27710] = 32'b00000000000000011100101111010000;
assign LUT_3[27711] = 32'b00000000000000100011011010101101;
assign LUT_3[27712] = 32'b00000000000000010011010111111000;
assign LUT_3[27713] = 32'b00000000000000011010000011010101;
assign LUT_3[27714] = 32'b00000000000000010101011111011100;
assign LUT_3[27715] = 32'b00000000000000011100001010111001;
assign LUT_3[27716] = 32'b00000000000000010000100101101110;
assign LUT_3[27717] = 32'b00000000000000010111010001001011;
assign LUT_3[27718] = 32'b00000000000000010010101101010010;
assign LUT_3[27719] = 32'b00000000000000011001011000101111;
assign LUT_3[27720] = 32'b00000000000000011000110000111110;
assign LUT_3[27721] = 32'b00000000000000011111011100011011;
assign LUT_3[27722] = 32'b00000000000000011010111000100010;
assign LUT_3[27723] = 32'b00000000000000100001100011111111;
assign LUT_3[27724] = 32'b00000000000000010101111110110100;
assign LUT_3[27725] = 32'b00000000000000011100101010010001;
assign LUT_3[27726] = 32'b00000000000000011000000110011000;
assign LUT_3[27727] = 32'b00000000000000011110110001110101;
assign LUT_3[27728] = 32'b00000000000000010110101010111011;
assign LUT_3[27729] = 32'b00000000000000011101010110011000;
assign LUT_3[27730] = 32'b00000000000000011000110010011111;
assign LUT_3[27731] = 32'b00000000000000011111011101111100;
assign LUT_3[27732] = 32'b00000000000000010011111000110001;
assign LUT_3[27733] = 32'b00000000000000011010100100001110;
assign LUT_3[27734] = 32'b00000000000000010110000000010101;
assign LUT_3[27735] = 32'b00000000000000011100101011110010;
assign LUT_3[27736] = 32'b00000000000000011100000100000001;
assign LUT_3[27737] = 32'b00000000000000100010101111011110;
assign LUT_3[27738] = 32'b00000000000000011110001011100101;
assign LUT_3[27739] = 32'b00000000000000100100110111000010;
assign LUT_3[27740] = 32'b00000000000000011001010001110111;
assign LUT_3[27741] = 32'b00000000000000011111111101010100;
assign LUT_3[27742] = 32'b00000000000000011011011001011011;
assign LUT_3[27743] = 32'b00000000000000100010000100111000;
assign LUT_3[27744] = 32'b00000000000000010100100110011000;
assign LUT_3[27745] = 32'b00000000000000011011010001110101;
assign LUT_3[27746] = 32'b00000000000000010110101101111100;
assign LUT_3[27747] = 32'b00000000000000011101011001011001;
assign LUT_3[27748] = 32'b00000000000000010001110100001110;
assign LUT_3[27749] = 32'b00000000000000011000011111101011;
assign LUT_3[27750] = 32'b00000000000000010011111011110010;
assign LUT_3[27751] = 32'b00000000000000011010100111001111;
assign LUT_3[27752] = 32'b00000000000000011001111111011110;
assign LUT_3[27753] = 32'b00000000000000100000101010111011;
assign LUT_3[27754] = 32'b00000000000000011100000111000010;
assign LUT_3[27755] = 32'b00000000000000100010110010011111;
assign LUT_3[27756] = 32'b00000000000000010111001101010100;
assign LUT_3[27757] = 32'b00000000000000011101111000110001;
assign LUT_3[27758] = 32'b00000000000000011001010100111000;
assign LUT_3[27759] = 32'b00000000000000100000000000010101;
assign LUT_3[27760] = 32'b00000000000000010111111001011011;
assign LUT_3[27761] = 32'b00000000000000011110100100111000;
assign LUT_3[27762] = 32'b00000000000000011010000000111111;
assign LUT_3[27763] = 32'b00000000000000100000101100011100;
assign LUT_3[27764] = 32'b00000000000000010101000111010001;
assign LUT_3[27765] = 32'b00000000000000011011110010101110;
assign LUT_3[27766] = 32'b00000000000000010111001110110101;
assign LUT_3[27767] = 32'b00000000000000011101111010010010;
assign LUT_3[27768] = 32'b00000000000000011101010010100001;
assign LUT_3[27769] = 32'b00000000000000100011111101111110;
assign LUT_3[27770] = 32'b00000000000000011111011010000101;
assign LUT_3[27771] = 32'b00000000000000100110000101100010;
assign LUT_3[27772] = 32'b00000000000000011010100000010111;
assign LUT_3[27773] = 32'b00000000000000100001001011110100;
assign LUT_3[27774] = 32'b00000000000000011100100111111011;
assign LUT_3[27775] = 32'b00000000000000100011010011011000;
assign LUT_3[27776] = 32'b00000000000000010101101010001011;
assign LUT_3[27777] = 32'b00000000000000011100010101101000;
assign LUT_3[27778] = 32'b00000000000000010111110001101111;
assign LUT_3[27779] = 32'b00000000000000011110011101001100;
assign LUT_3[27780] = 32'b00000000000000010010111000000001;
assign LUT_3[27781] = 32'b00000000000000011001100011011110;
assign LUT_3[27782] = 32'b00000000000000010100111111100101;
assign LUT_3[27783] = 32'b00000000000000011011101011000010;
assign LUT_3[27784] = 32'b00000000000000011011000011010001;
assign LUT_3[27785] = 32'b00000000000000100001101110101110;
assign LUT_3[27786] = 32'b00000000000000011101001010110101;
assign LUT_3[27787] = 32'b00000000000000100011110110010010;
assign LUT_3[27788] = 32'b00000000000000011000010001000111;
assign LUT_3[27789] = 32'b00000000000000011110111100100100;
assign LUT_3[27790] = 32'b00000000000000011010011000101011;
assign LUT_3[27791] = 32'b00000000000000100001000100001000;
assign LUT_3[27792] = 32'b00000000000000011000111101001110;
assign LUT_3[27793] = 32'b00000000000000011111101000101011;
assign LUT_3[27794] = 32'b00000000000000011011000100110010;
assign LUT_3[27795] = 32'b00000000000000100001110000001111;
assign LUT_3[27796] = 32'b00000000000000010110001011000100;
assign LUT_3[27797] = 32'b00000000000000011100110110100001;
assign LUT_3[27798] = 32'b00000000000000011000010010101000;
assign LUT_3[27799] = 32'b00000000000000011110111110000101;
assign LUT_3[27800] = 32'b00000000000000011110010110010100;
assign LUT_3[27801] = 32'b00000000000000100101000001110001;
assign LUT_3[27802] = 32'b00000000000000100000011101111000;
assign LUT_3[27803] = 32'b00000000000000100111001001010101;
assign LUT_3[27804] = 32'b00000000000000011011100100001010;
assign LUT_3[27805] = 32'b00000000000000100010001111100111;
assign LUT_3[27806] = 32'b00000000000000011101101011101110;
assign LUT_3[27807] = 32'b00000000000000100100010111001011;
assign LUT_3[27808] = 32'b00000000000000010110111000101011;
assign LUT_3[27809] = 32'b00000000000000011101100100001000;
assign LUT_3[27810] = 32'b00000000000000011001000000001111;
assign LUT_3[27811] = 32'b00000000000000011111101011101100;
assign LUT_3[27812] = 32'b00000000000000010100000110100001;
assign LUT_3[27813] = 32'b00000000000000011010110001111110;
assign LUT_3[27814] = 32'b00000000000000010110001110000101;
assign LUT_3[27815] = 32'b00000000000000011100111001100010;
assign LUT_3[27816] = 32'b00000000000000011100010001110001;
assign LUT_3[27817] = 32'b00000000000000100010111101001110;
assign LUT_3[27818] = 32'b00000000000000011110011001010101;
assign LUT_3[27819] = 32'b00000000000000100101000100110010;
assign LUT_3[27820] = 32'b00000000000000011001011111100111;
assign LUT_3[27821] = 32'b00000000000000100000001011000100;
assign LUT_3[27822] = 32'b00000000000000011011100111001011;
assign LUT_3[27823] = 32'b00000000000000100010010010101000;
assign LUT_3[27824] = 32'b00000000000000011010001011101110;
assign LUT_3[27825] = 32'b00000000000000100000110111001011;
assign LUT_3[27826] = 32'b00000000000000011100010011010010;
assign LUT_3[27827] = 32'b00000000000000100010111110101111;
assign LUT_3[27828] = 32'b00000000000000010111011001100100;
assign LUT_3[27829] = 32'b00000000000000011110000101000001;
assign LUT_3[27830] = 32'b00000000000000011001100001001000;
assign LUT_3[27831] = 32'b00000000000000100000001100100101;
assign LUT_3[27832] = 32'b00000000000000011111100100110100;
assign LUT_3[27833] = 32'b00000000000000100110010000010001;
assign LUT_3[27834] = 32'b00000000000000100001101100011000;
assign LUT_3[27835] = 32'b00000000000000101000010111110101;
assign LUT_3[27836] = 32'b00000000000000011100110010101010;
assign LUT_3[27837] = 32'b00000000000000100011011110000111;
assign LUT_3[27838] = 32'b00000000000000011110111010001110;
assign LUT_3[27839] = 32'b00000000000000100101100101101011;
assign LUT_3[27840] = 32'b00000000000000010101100010110110;
assign LUT_3[27841] = 32'b00000000000000011100001110010011;
assign LUT_3[27842] = 32'b00000000000000010111101010011010;
assign LUT_3[27843] = 32'b00000000000000011110010101110111;
assign LUT_3[27844] = 32'b00000000000000010010110000101100;
assign LUT_3[27845] = 32'b00000000000000011001011100001001;
assign LUT_3[27846] = 32'b00000000000000010100111000010000;
assign LUT_3[27847] = 32'b00000000000000011011100011101101;
assign LUT_3[27848] = 32'b00000000000000011010111011111100;
assign LUT_3[27849] = 32'b00000000000000100001100111011001;
assign LUT_3[27850] = 32'b00000000000000011101000011100000;
assign LUT_3[27851] = 32'b00000000000000100011101110111101;
assign LUT_3[27852] = 32'b00000000000000011000001001110010;
assign LUT_3[27853] = 32'b00000000000000011110110101001111;
assign LUT_3[27854] = 32'b00000000000000011010010001010110;
assign LUT_3[27855] = 32'b00000000000000100000111100110011;
assign LUT_3[27856] = 32'b00000000000000011000110101111001;
assign LUT_3[27857] = 32'b00000000000000011111100001010110;
assign LUT_3[27858] = 32'b00000000000000011010111101011101;
assign LUT_3[27859] = 32'b00000000000000100001101000111010;
assign LUT_3[27860] = 32'b00000000000000010110000011101111;
assign LUT_3[27861] = 32'b00000000000000011100101111001100;
assign LUT_3[27862] = 32'b00000000000000011000001011010011;
assign LUT_3[27863] = 32'b00000000000000011110110110110000;
assign LUT_3[27864] = 32'b00000000000000011110001110111111;
assign LUT_3[27865] = 32'b00000000000000100100111010011100;
assign LUT_3[27866] = 32'b00000000000000100000010110100011;
assign LUT_3[27867] = 32'b00000000000000100111000010000000;
assign LUT_3[27868] = 32'b00000000000000011011011100110101;
assign LUT_3[27869] = 32'b00000000000000100010001000010010;
assign LUT_3[27870] = 32'b00000000000000011101100100011001;
assign LUT_3[27871] = 32'b00000000000000100100001111110110;
assign LUT_3[27872] = 32'b00000000000000010110110001010110;
assign LUT_3[27873] = 32'b00000000000000011101011100110011;
assign LUT_3[27874] = 32'b00000000000000011000111000111010;
assign LUT_3[27875] = 32'b00000000000000011111100100010111;
assign LUT_3[27876] = 32'b00000000000000010011111111001100;
assign LUT_3[27877] = 32'b00000000000000011010101010101001;
assign LUT_3[27878] = 32'b00000000000000010110000110110000;
assign LUT_3[27879] = 32'b00000000000000011100110010001101;
assign LUT_3[27880] = 32'b00000000000000011100001010011100;
assign LUT_3[27881] = 32'b00000000000000100010110101111001;
assign LUT_3[27882] = 32'b00000000000000011110010010000000;
assign LUT_3[27883] = 32'b00000000000000100100111101011101;
assign LUT_3[27884] = 32'b00000000000000011001011000010010;
assign LUT_3[27885] = 32'b00000000000000100000000011101111;
assign LUT_3[27886] = 32'b00000000000000011011011111110110;
assign LUT_3[27887] = 32'b00000000000000100010001011010011;
assign LUT_3[27888] = 32'b00000000000000011010000100011001;
assign LUT_3[27889] = 32'b00000000000000100000101111110110;
assign LUT_3[27890] = 32'b00000000000000011100001011111101;
assign LUT_3[27891] = 32'b00000000000000100010110111011010;
assign LUT_3[27892] = 32'b00000000000000010111010010001111;
assign LUT_3[27893] = 32'b00000000000000011101111101101100;
assign LUT_3[27894] = 32'b00000000000000011001011001110011;
assign LUT_3[27895] = 32'b00000000000000100000000101010000;
assign LUT_3[27896] = 32'b00000000000000011111011101011111;
assign LUT_3[27897] = 32'b00000000000000100110001000111100;
assign LUT_3[27898] = 32'b00000000000000100001100101000011;
assign LUT_3[27899] = 32'b00000000000000101000010000100000;
assign LUT_3[27900] = 32'b00000000000000011100101011010101;
assign LUT_3[27901] = 32'b00000000000000100011010110110010;
assign LUT_3[27902] = 32'b00000000000000011110110010111001;
assign LUT_3[27903] = 32'b00000000000000100101011110010110;
assign LUT_3[27904] = 32'b00000000000000001111101110101110;
assign LUT_3[27905] = 32'b00000000000000010110011010001011;
assign LUT_3[27906] = 32'b00000000000000010001110110010010;
assign LUT_3[27907] = 32'b00000000000000011000100001101111;
assign LUT_3[27908] = 32'b00000000000000001100111100100100;
assign LUT_3[27909] = 32'b00000000000000010011101000000001;
assign LUT_3[27910] = 32'b00000000000000001111000100001000;
assign LUT_3[27911] = 32'b00000000000000010101101111100101;
assign LUT_3[27912] = 32'b00000000000000010101000111110100;
assign LUT_3[27913] = 32'b00000000000000011011110011010001;
assign LUT_3[27914] = 32'b00000000000000010111001111011000;
assign LUT_3[27915] = 32'b00000000000000011101111010110101;
assign LUT_3[27916] = 32'b00000000000000010010010101101010;
assign LUT_3[27917] = 32'b00000000000000011001000001000111;
assign LUT_3[27918] = 32'b00000000000000010100011101001110;
assign LUT_3[27919] = 32'b00000000000000011011001000101011;
assign LUT_3[27920] = 32'b00000000000000010011000001110001;
assign LUT_3[27921] = 32'b00000000000000011001101101001110;
assign LUT_3[27922] = 32'b00000000000000010101001001010101;
assign LUT_3[27923] = 32'b00000000000000011011110100110010;
assign LUT_3[27924] = 32'b00000000000000010000001111100111;
assign LUT_3[27925] = 32'b00000000000000010110111011000100;
assign LUT_3[27926] = 32'b00000000000000010010010111001011;
assign LUT_3[27927] = 32'b00000000000000011001000010101000;
assign LUT_3[27928] = 32'b00000000000000011000011010110111;
assign LUT_3[27929] = 32'b00000000000000011111000110010100;
assign LUT_3[27930] = 32'b00000000000000011010100010011011;
assign LUT_3[27931] = 32'b00000000000000100001001101111000;
assign LUT_3[27932] = 32'b00000000000000010101101000101101;
assign LUT_3[27933] = 32'b00000000000000011100010100001010;
assign LUT_3[27934] = 32'b00000000000000010111110000010001;
assign LUT_3[27935] = 32'b00000000000000011110011011101110;
assign LUT_3[27936] = 32'b00000000000000010000111101001110;
assign LUT_3[27937] = 32'b00000000000000010111101000101011;
assign LUT_3[27938] = 32'b00000000000000010011000100110010;
assign LUT_3[27939] = 32'b00000000000000011001110000001111;
assign LUT_3[27940] = 32'b00000000000000001110001011000100;
assign LUT_3[27941] = 32'b00000000000000010100110110100001;
assign LUT_3[27942] = 32'b00000000000000010000010010101000;
assign LUT_3[27943] = 32'b00000000000000010110111110000101;
assign LUT_3[27944] = 32'b00000000000000010110010110010100;
assign LUT_3[27945] = 32'b00000000000000011101000001110001;
assign LUT_3[27946] = 32'b00000000000000011000011101111000;
assign LUT_3[27947] = 32'b00000000000000011111001001010101;
assign LUT_3[27948] = 32'b00000000000000010011100100001010;
assign LUT_3[27949] = 32'b00000000000000011010001111100111;
assign LUT_3[27950] = 32'b00000000000000010101101011101110;
assign LUT_3[27951] = 32'b00000000000000011100010111001011;
assign LUT_3[27952] = 32'b00000000000000010100010000010001;
assign LUT_3[27953] = 32'b00000000000000011010111011101110;
assign LUT_3[27954] = 32'b00000000000000010110010111110101;
assign LUT_3[27955] = 32'b00000000000000011101000011010010;
assign LUT_3[27956] = 32'b00000000000000010001011110000111;
assign LUT_3[27957] = 32'b00000000000000011000001001100100;
assign LUT_3[27958] = 32'b00000000000000010011100101101011;
assign LUT_3[27959] = 32'b00000000000000011010010001001000;
assign LUT_3[27960] = 32'b00000000000000011001101001010111;
assign LUT_3[27961] = 32'b00000000000000100000010100110100;
assign LUT_3[27962] = 32'b00000000000000011011110000111011;
assign LUT_3[27963] = 32'b00000000000000100010011100011000;
assign LUT_3[27964] = 32'b00000000000000010110110111001101;
assign LUT_3[27965] = 32'b00000000000000011101100010101010;
assign LUT_3[27966] = 32'b00000000000000011000111110110001;
assign LUT_3[27967] = 32'b00000000000000011111101010001110;
assign LUT_3[27968] = 32'b00000000000000001111100111011001;
assign LUT_3[27969] = 32'b00000000000000010110010010110110;
assign LUT_3[27970] = 32'b00000000000000010001101110111101;
assign LUT_3[27971] = 32'b00000000000000011000011010011010;
assign LUT_3[27972] = 32'b00000000000000001100110101001111;
assign LUT_3[27973] = 32'b00000000000000010011100000101100;
assign LUT_3[27974] = 32'b00000000000000001110111100110011;
assign LUT_3[27975] = 32'b00000000000000010101101000010000;
assign LUT_3[27976] = 32'b00000000000000010101000000011111;
assign LUT_3[27977] = 32'b00000000000000011011101011111100;
assign LUT_3[27978] = 32'b00000000000000010111001000000011;
assign LUT_3[27979] = 32'b00000000000000011101110011100000;
assign LUT_3[27980] = 32'b00000000000000010010001110010101;
assign LUT_3[27981] = 32'b00000000000000011000111001110010;
assign LUT_3[27982] = 32'b00000000000000010100010101111001;
assign LUT_3[27983] = 32'b00000000000000011011000001010110;
assign LUT_3[27984] = 32'b00000000000000010010111010011100;
assign LUT_3[27985] = 32'b00000000000000011001100101111001;
assign LUT_3[27986] = 32'b00000000000000010101000010000000;
assign LUT_3[27987] = 32'b00000000000000011011101101011101;
assign LUT_3[27988] = 32'b00000000000000010000001000010010;
assign LUT_3[27989] = 32'b00000000000000010110110011101111;
assign LUT_3[27990] = 32'b00000000000000010010001111110110;
assign LUT_3[27991] = 32'b00000000000000011000111011010011;
assign LUT_3[27992] = 32'b00000000000000011000010011100010;
assign LUT_3[27993] = 32'b00000000000000011110111110111111;
assign LUT_3[27994] = 32'b00000000000000011010011011000110;
assign LUT_3[27995] = 32'b00000000000000100001000110100011;
assign LUT_3[27996] = 32'b00000000000000010101100001011000;
assign LUT_3[27997] = 32'b00000000000000011100001100110101;
assign LUT_3[27998] = 32'b00000000000000010111101000111100;
assign LUT_3[27999] = 32'b00000000000000011110010100011001;
assign LUT_3[28000] = 32'b00000000000000010000110101111001;
assign LUT_3[28001] = 32'b00000000000000010111100001010110;
assign LUT_3[28002] = 32'b00000000000000010010111101011101;
assign LUT_3[28003] = 32'b00000000000000011001101000111010;
assign LUT_3[28004] = 32'b00000000000000001110000011101111;
assign LUT_3[28005] = 32'b00000000000000010100101111001100;
assign LUT_3[28006] = 32'b00000000000000010000001011010011;
assign LUT_3[28007] = 32'b00000000000000010110110110110000;
assign LUT_3[28008] = 32'b00000000000000010110001110111111;
assign LUT_3[28009] = 32'b00000000000000011100111010011100;
assign LUT_3[28010] = 32'b00000000000000011000010110100011;
assign LUT_3[28011] = 32'b00000000000000011111000010000000;
assign LUT_3[28012] = 32'b00000000000000010011011100110101;
assign LUT_3[28013] = 32'b00000000000000011010001000010010;
assign LUT_3[28014] = 32'b00000000000000010101100100011001;
assign LUT_3[28015] = 32'b00000000000000011100001111110110;
assign LUT_3[28016] = 32'b00000000000000010100001000111100;
assign LUT_3[28017] = 32'b00000000000000011010110100011001;
assign LUT_3[28018] = 32'b00000000000000010110010000100000;
assign LUT_3[28019] = 32'b00000000000000011100111011111101;
assign LUT_3[28020] = 32'b00000000000000010001010110110010;
assign LUT_3[28021] = 32'b00000000000000011000000010001111;
assign LUT_3[28022] = 32'b00000000000000010011011110010110;
assign LUT_3[28023] = 32'b00000000000000011010001001110011;
assign LUT_3[28024] = 32'b00000000000000011001100010000010;
assign LUT_3[28025] = 32'b00000000000000100000001101011111;
assign LUT_3[28026] = 32'b00000000000000011011101001100110;
assign LUT_3[28027] = 32'b00000000000000100010010101000011;
assign LUT_3[28028] = 32'b00000000000000010110101111111000;
assign LUT_3[28029] = 32'b00000000000000011101011011010101;
assign LUT_3[28030] = 32'b00000000000000011000110111011100;
assign LUT_3[28031] = 32'b00000000000000011111100010111001;
assign LUT_3[28032] = 32'b00000000000000010001111001101100;
assign LUT_3[28033] = 32'b00000000000000011000100101001001;
assign LUT_3[28034] = 32'b00000000000000010100000001010000;
assign LUT_3[28035] = 32'b00000000000000011010101100101101;
assign LUT_3[28036] = 32'b00000000000000001111000111100010;
assign LUT_3[28037] = 32'b00000000000000010101110010111111;
assign LUT_3[28038] = 32'b00000000000000010001001111000110;
assign LUT_3[28039] = 32'b00000000000000010111111010100011;
assign LUT_3[28040] = 32'b00000000000000010111010010110010;
assign LUT_3[28041] = 32'b00000000000000011101111110001111;
assign LUT_3[28042] = 32'b00000000000000011001011010010110;
assign LUT_3[28043] = 32'b00000000000000100000000101110011;
assign LUT_3[28044] = 32'b00000000000000010100100000101000;
assign LUT_3[28045] = 32'b00000000000000011011001100000101;
assign LUT_3[28046] = 32'b00000000000000010110101000001100;
assign LUT_3[28047] = 32'b00000000000000011101010011101001;
assign LUT_3[28048] = 32'b00000000000000010101001100101111;
assign LUT_3[28049] = 32'b00000000000000011011111000001100;
assign LUT_3[28050] = 32'b00000000000000010111010100010011;
assign LUT_3[28051] = 32'b00000000000000011101111111110000;
assign LUT_3[28052] = 32'b00000000000000010010011010100101;
assign LUT_3[28053] = 32'b00000000000000011001000110000010;
assign LUT_3[28054] = 32'b00000000000000010100100010001001;
assign LUT_3[28055] = 32'b00000000000000011011001101100110;
assign LUT_3[28056] = 32'b00000000000000011010100101110101;
assign LUT_3[28057] = 32'b00000000000000100001010001010010;
assign LUT_3[28058] = 32'b00000000000000011100101101011001;
assign LUT_3[28059] = 32'b00000000000000100011011000110110;
assign LUT_3[28060] = 32'b00000000000000010111110011101011;
assign LUT_3[28061] = 32'b00000000000000011110011111001000;
assign LUT_3[28062] = 32'b00000000000000011001111011001111;
assign LUT_3[28063] = 32'b00000000000000100000100110101100;
assign LUT_3[28064] = 32'b00000000000000010011001000001100;
assign LUT_3[28065] = 32'b00000000000000011001110011101001;
assign LUT_3[28066] = 32'b00000000000000010101001111110000;
assign LUT_3[28067] = 32'b00000000000000011011111011001101;
assign LUT_3[28068] = 32'b00000000000000010000010110000010;
assign LUT_3[28069] = 32'b00000000000000010111000001011111;
assign LUT_3[28070] = 32'b00000000000000010010011101100110;
assign LUT_3[28071] = 32'b00000000000000011001001001000011;
assign LUT_3[28072] = 32'b00000000000000011000100001010010;
assign LUT_3[28073] = 32'b00000000000000011111001100101111;
assign LUT_3[28074] = 32'b00000000000000011010101000110110;
assign LUT_3[28075] = 32'b00000000000000100001010100010011;
assign LUT_3[28076] = 32'b00000000000000010101101111001000;
assign LUT_3[28077] = 32'b00000000000000011100011010100101;
assign LUT_3[28078] = 32'b00000000000000010111110110101100;
assign LUT_3[28079] = 32'b00000000000000011110100010001001;
assign LUT_3[28080] = 32'b00000000000000010110011011001111;
assign LUT_3[28081] = 32'b00000000000000011101000110101100;
assign LUT_3[28082] = 32'b00000000000000011000100010110011;
assign LUT_3[28083] = 32'b00000000000000011111001110010000;
assign LUT_3[28084] = 32'b00000000000000010011101001000101;
assign LUT_3[28085] = 32'b00000000000000011010010100100010;
assign LUT_3[28086] = 32'b00000000000000010101110000101001;
assign LUT_3[28087] = 32'b00000000000000011100011100000110;
assign LUT_3[28088] = 32'b00000000000000011011110100010101;
assign LUT_3[28089] = 32'b00000000000000100010011111110010;
assign LUT_3[28090] = 32'b00000000000000011101111011111001;
assign LUT_3[28091] = 32'b00000000000000100100100111010110;
assign LUT_3[28092] = 32'b00000000000000011001000010001011;
assign LUT_3[28093] = 32'b00000000000000011111101101101000;
assign LUT_3[28094] = 32'b00000000000000011011001001101111;
assign LUT_3[28095] = 32'b00000000000000100001110101001100;
assign LUT_3[28096] = 32'b00000000000000010001110010010111;
assign LUT_3[28097] = 32'b00000000000000011000011101110100;
assign LUT_3[28098] = 32'b00000000000000010011111001111011;
assign LUT_3[28099] = 32'b00000000000000011010100101011000;
assign LUT_3[28100] = 32'b00000000000000001111000000001101;
assign LUT_3[28101] = 32'b00000000000000010101101011101010;
assign LUT_3[28102] = 32'b00000000000000010001000111110001;
assign LUT_3[28103] = 32'b00000000000000010111110011001110;
assign LUT_3[28104] = 32'b00000000000000010111001011011101;
assign LUT_3[28105] = 32'b00000000000000011101110110111010;
assign LUT_3[28106] = 32'b00000000000000011001010011000001;
assign LUT_3[28107] = 32'b00000000000000011111111110011110;
assign LUT_3[28108] = 32'b00000000000000010100011001010011;
assign LUT_3[28109] = 32'b00000000000000011011000100110000;
assign LUT_3[28110] = 32'b00000000000000010110100000110111;
assign LUT_3[28111] = 32'b00000000000000011101001100010100;
assign LUT_3[28112] = 32'b00000000000000010101000101011010;
assign LUT_3[28113] = 32'b00000000000000011011110000110111;
assign LUT_3[28114] = 32'b00000000000000010111001100111110;
assign LUT_3[28115] = 32'b00000000000000011101111000011011;
assign LUT_3[28116] = 32'b00000000000000010010010011010000;
assign LUT_3[28117] = 32'b00000000000000011000111110101101;
assign LUT_3[28118] = 32'b00000000000000010100011010110100;
assign LUT_3[28119] = 32'b00000000000000011011000110010001;
assign LUT_3[28120] = 32'b00000000000000011010011110100000;
assign LUT_3[28121] = 32'b00000000000000100001001001111101;
assign LUT_3[28122] = 32'b00000000000000011100100110000100;
assign LUT_3[28123] = 32'b00000000000000100011010001100001;
assign LUT_3[28124] = 32'b00000000000000010111101100010110;
assign LUT_3[28125] = 32'b00000000000000011110010111110011;
assign LUT_3[28126] = 32'b00000000000000011001110011111010;
assign LUT_3[28127] = 32'b00000000000000100000011111010111;
assign LUT_3[28128] = 32'b00000000000000010011000000110111;
assign LUT_3[28129] = 32'b00000000000000011001101100010100;
assign LUT_3[28130] = 32'b00000000000000010101001000011011;
assign LUT_3[28131] = 32'b00000000000000011011110011111000;
assign LUT_3[28132] = 32'b00000000000000010000001110101101;
assign LUT_3[28133] = 32'b00000000000000010110111010001010;
assign LUT_3[28134] = 32'b00000000000000010010010110010001;
assign LUT_3[28135] = 32'b00000000000000011001000001101110;
assign LUT_3[28136] = 32'b00000000000000011000011001111101;
assign LUT_3[28137] = 32'b00000000000000011111000101011010;
assign LUT_3[28138] = 32'b00000000000000011010100001100001;
assign LUT_3[28139] = 32'b00000000000000100001001100111110;
assign LUT_3[28140] = 32'b00000000000000010101100111110011;
assign LUT_3[28141] = 32'b00000000000000011100010011010000;
assign LUT_3[28142] = 32'b00000000000000010111101111010111;
assign LUT_3[28143] = 32'b00000000000000011110011010110100;
assign LUT_3[28144] = 32'b00000000000000010110010011111010;
assign LUT_3[28145] = 32'b00000000000000011100111111010111;
assign LUT_3[28146] = 32'b00000000000000011000011011011110;
assign LUT_3[28147] = 32'b00000000000000011111000110111011;
assign LUT_3[28148] = 32'b00000000000000010011100001110000;
assign LUT_3[28149] = 32'b00000000000000011010001101001101;
assign LUT_3[28150] = 32'b00000000000000010101101001010100;
assign LUT_3[28151] = 32'b00000000000000011100010100110001;
assign LUT_3[28152] = 32'b00000000000000011011101101000000;
assign LUT_3[28153] = 32'b00000000000000100010011000011101;
assign LUT_3[28154] = 32'b00000000000000011101110100100100;
assign LUT_3[28155] = 32'b00000000000000100100100000000001;
assign LUT_3[28156] = 32'b00000000000000011000111010110110;
assign LUT_3[28157] = 32'b00000000000000011111100110010011;
assign LUT_3[28158] = 32'b00000000000000011011000010011010;
assign LUT_3[28159] = 32'b00000000000000100001101101110111;
assign LUT_3[28160] = 32'b00000000000000010110110100011001;
assign LUT_3[28161] = 32'b00000000000000011101011111110110;
assign LUT_3[28162] = 32'b00000000000000011000111011111101;
assign LUT_3[28163] = 32'b00000000000000011111100111011010;
assign LUT_3[28164] = 32'b00000000000000010100000010001111;
assign LUT_3[28165] = 32'b00000000000000011010101101101100;
assign LUT_3[28166] = 32'b00000000000000010110001001110011;
assign LUT_3[28167] = 32'b00000000000000011100110101010000;
assign LUT_3[28168] = 32'b00000000000000011100001101011111;
assign LUT_3[28169] = 32'b00000000000000100010111000111100;
assign LUT_3[28170] = 32'b00000000000000011110010101000011;
assign LUT_3[28171] = 32'b00000000000000100101000000100000;
assign LUT_3[28172] = 32'b00000000000000011001011011010101;
assign LUT_3[28173] = 32'b00000000000000100000000110110010;
assign LUT_3[28174] = 32'b00000000000000011011100010111001;
assign LUT_3[28175] = 32'b00000000000000100010001110010110;
assign LUT_3[28176] = 32'b00000000000000011010000111011100;
assign LUT_3[28177] = 32'b00000000000000100000110010111001;
assign LUT_3[28178] = 32'b00000000000000011100001111000000;
assign LUT_3[28179] = 32'b00000000000000100010111010011101;
assign LUT_3[28180] = 32'b00000000000000010111010101010010;
assign LUT_3[28181] = 32'b00000000000000011110000000101111;
assign LUT_3[28182] = 32'b00000000000000011001011100110110;
assign LUT_3[28183] = 32'b00000000000000100000001000010011;
assign LUT_3[28184] = 32'b00000000000000011111100000100010;
assign LUT_3[28185] = 32'b00000000000000100110001011111111;
assign LUT_3[28186] = 32'b00000000000000100001101000000110;
assign LUT_3[28187] = 32'b00000000000000101000010011100011;
assign LUT_3[28188] = 32'b00000000000000011100101110011000;
assign LUT_3[28189] = 32'b00000000000000100011011001110101;
assign LUT_3[28190] = 32'b00000000000000011110110101111100;
assign LUT_3[28191] = 32'b00000000000000100101100001011001;
assign LUT_3[28192] = 32'b00000000000000011000000010111001;
assign LUT_3[28193] = 32'b00000000000000011110101110010110;
assign LUT_3[28194] = 32'b00000000000000011010001010011101;
assign LUT_3[28195] = 32'b00000000000000100000110101111010;
assign LUT_3[28196] = 32'b00000000000000010101010000101111;
assign LUT_3[28197] = 32'b00000000000000011011111100001100;
assign LUT_3[28198] = 32'b00000000000000010111011000010011;
assign LUT_3[28199] = 32'b00000000000000011110000011110000;
assign LUT_3[28200] = 32'b00000000000000011101011011111111;
assign LUT_3[28201] = 32'b00000000000000100100000111011100;
assign LUT_3[28202] = 32'b00000000000000011111100011100011;
assign LUT_3[28203] = 32'b00000000000000100110001111000000;
assign LUT_3[28204] = 32'b00000000000000011010101001110101;
assign LUT_3[28205] = 32'b00000000000000100001010101010010;
assign LUT_3[28206] = 32'b00000000000000011100110001011001;
assign LUT_3[28207] = 32'b00000000000000100011011100110110;
assign LUT_3[28208] = 32'b00000000000000011011010101111100;
assign LUT_3[28209] = 32'b00000000000000100010000001011001;
assign LUT_3[28210] = 32'b00000000000000011101011101100000;
assign LUT_3[28211] = 32'b00000000000000100100001000111101;
assign LUT_3[28212] = 32'b00000000000000011000100011110010;
assign LUT_3[28213] = 32'b00000000000000011111001111001111;
assign LUT_3[28214] = 32'b00000000000000011010101011010110;
assign LUT_3[28215] = 32'b00000000000000100001010110110011;
assign LUT_3[28216] = 32'b00000000000000100000101111000010;
assign LUT_3[28217] = 32'b00000000000000100111011010011111;
assign LUT_3[28218] = 32'b00000000000000100010110110100110;
assign LUT_3[28219] = 32'b00000000000000101001100010000011;
assign LUT_3[28220] = 32'b00000000000000011101111100111000;
assign LUT_3[28221] = 32'b00000000000000100100101000010101;
assign LUT_3[28222] = 32'b00000000000000100000000100011100;
assign LUT_3[28223] = 32'b00000000000000100110101111111001;
assign LUT_3[28224] = 32'b00000000000000010110101101000100;
assign LUT_3[28225] = 32'b00000000000000011101011000100001;
assign LUT_3[28226] = 32'b00000000000000011000110100101000;
assign LUT_3[28227] = 32'b00000000000000011111100000000101;
assign LUT_3[28228] = 32'b00000000000000010011111010111010;
assign LUT_3[28229] = 32'b00000000000000011010100110010111;
assign LUT_3[28230] = 32'b00000000000000010110000010011110;
assign LUT_3[28231] = 32'b00000000000000011100101101111011;
assign LUT_3[28232] = 32'b00000000000000011100000110001010;
assign LUT_3[28233] = 32'b00000000000000100010110001100111;
assign LUT_3[28234] = 32'b00000000000000011110001101101110;
assign LUT_3[28235] = 32'b00000000000000100100111001001011;
assign LUT_3[28236] = 32'b00000000000000011001010100000000;
assign LUT_3[28237] = 32'b00000000000000011111111111011101;
assign LUT_3[28238] = 32'b00000000000000011011011011100100;
assign LUT_3[28239] = 32'b00000000000000100010000111000001;
assign LUT_3[28240] = 32'b00000000000000011010000000000111;
assign LUT_3[28241] = 32'b00000000000000100000101011100100;
assign LUT_3[28242] = 32'b00000000000000011100000111101011;
assign LUT_3[28243] = 32'b00000000000000100010110011001000;
assign LUT_3[28244] = 32'b00000000000000010111001101111101;
assign LUT_3[28245] = 32'b00000000000000011101111001011010;
assign LUT_3[28246] = 32'b00000000000000011001010101100001;
assign LUT_3[28247] = 32'b00000000000000100000000000111110;
assign LUT_3[28248] = 32'b00000000000000011111011001001101;
assign LUT_3[28249] = 32'b00000000000000100110000100101010;
assign LUT_3[28250] = 32'b00000000000000100001100000110001;
assign LUT_3[28251] = 32'b00000000000000101000001100001110;
assign LUT_3[28252] = 32'b00000000000000011100100111000011;
assign LUT_3[28253] = 32'b00000000000000100011010010100000;
assign LUT_3[28254] = 32'b00000000000000011110101110100111;
assign LUT_3[28255] = 32'b00000000000000100101011010000100;
assign LUT_3[28256] = 32'b00000000000000010111111011100100;
assign LUT_3[28257] = 32'b00000000000000011110100111000001;
assign LUT_3[28258] = 32'b00000000000000011010000011001000;
assign LUT_3[28259] = 32'b00000000000000100000101110100101;
assign LUT_3[28260] = 32'b00000000000000010101001001011010;
assign LUT_3[28261] = 32'b00000000000000011011110100110111;
assign LUT_3[28262] = 32'b00000000000000010111010000111110;
assign LUT_3[28263] = 32'b00000000000000011101111100011011;
assign LUT_3[28264] = 32'b00000000000000011101010100101010;
assign LUT_3[28265] = 32'b00000000000000100100000000000111;
assign LUT_3[28266] = 32'b00000000000000011111011100001110;
assign LUT_3[28267] = 32'b00000000000000100110000111101011;
assign LUT_3[28268] = 32'b00000000000000011010100010100000;
assign LUT_3[28269] = 32'b00000000000000100001001101111101;
assign LUT_3[28270] = 32'b00000000000000011100101010000100;
assign LUT_3[28271] = 32'b00000000000000100011010101100001;
assign LUT_3[28272] = 32'b00000000000000011011001110100111;
assign LUT_3[28273] = 32'b00000000000000100001111010000100;
assign LUT_3[28274] = 32'b00000000000000011101010110001011;
assign LUT_3[28275] = 32'b00000000000000100100000001101000;
assign LUT_3[28276] = 32'b00000000000000011000011100011101;
assign LUT_3[28277] = 32'b00000000000000011111000111111010;
assign LUT_3[28278] = 32'b00000000000000011010100100000001;
assign LUT_3[28279] = 32'b00000000000000100001001111011110;
assign LUT_3[28280] = 32'b00000000000000100000100111101101;
assign LUT_3[28281] = 32'b00000000000000100111010011001010;
assign LUT_3[28282] = 32'b00000000000000100010101111010001;
assign LUT_3[28283] = 32'b00000000000000101001011010101110;
assign LUT_3[28284] = 32'b00000000000000011101110101100011;
assign LUT_3[28285] = 32'b00000000000000100100100001000000;
assign LUT_3[28286] = 32'b00000000000000011111111101000111;
assign LUT_3[28287] = 32'b00000000000000100110101000100100;
assign LUT_3[28288] = 32'b00000000000000011000111111010111;
assign LUT_3[28289] = 32'b00000000000000011111101010110100;
assign LUT_3[28290] = 32'b00000000000000011011000110111011;
assign LUT_3[28291] = 32'b00000000000000100001110010011000;
assign LUT_3[28292] = 32'b00000000000000010110001101001101;
assign LUT_3[28293] = 32'b00000000000000011100111000101010;
assign LUT_3[28294] = 32'b00000000000000011000010100110001;
assign LUT_3[28295] = 32'b00000000000000011111000000001110;
assign LUT_3[28296] = 32'b00000000000000011110011000011101;
assign LUT_3[28297] = 32'b00000000000000100101000011111010;
assign LUT_3[28298] = 32'b00000000000000100000100000000001;
assign LUT_3[28299] = 32'b00000000000000100111001011011110;
assign LUT_3[28300] = 32'b00000000000000011011100110010011;
assign LUT_3[28301] = 32'b00000000000000100010010001110000;
assign LUT_3[28302] = 32'b00000000000000011101101101110111;
assign LUT_3[28303] = 32'b00000000000000100100011001010100;
assign LUT_3[28304] = 32'b00000000000000011100010010011010;
assign LUT_3[28305] = 32'b00000000000000100010111101110111;
assign LUT_3[28306] = 32'b00000000000000011110011001111110;
assign LUT_3[28307] = 32'b00000000000000100101000101011011;
assign LUT_3[28308] = 32'b00000000000000011001100000010000;
assign LUT_3[28309] = 32'b00000000000000100000001011101101;
assign LUT_3[28310] = 32'b00000000000000011011100111110100;
assign LUT_3[28311] = 32'b00000000000000100010010011010001;
assign LUT_3[28312] = 32'b00000000000000100001101011100000;
assign LUT_3[28313] = 32'b00000000000000101000010110111101;
assign LUT_3[28314] = 32'b00000000000000100011110011000100;
assign LUT_3[28315] = 32'b00000000000000101010011110100001;
assign LUT_3[28316] = 32'b00000000000000011110111001010110;
assign LUT_3[28317] = 32'b00000000000000100101100100110011;
assign LUT_3[28318] = 32'b00000000000000100001000000111010;
assign LUT_3[28319] = 32'b00000000000000100111101100010111;
assign LUT_3[28320] = 32'b00000000000000011010001101110111;
assign LUT_3[28321] = 32'b00000000000000100000111001010100;
assign LUT_3[28322] = 32'b00000000000000011100010101011011;
assign LUT_3[28323] = 32'b00000000000000100011000000111000;
assign LUT_3[28324] = 32'b00000000000000010111011011101101;
assign LUT_3[28325] = 32'b00000000000000011110000111001010;
assign LUT_3[28326] = 32'b00000000000000011001100011010001;
assign LUT_3[28327] = 32'b00000000000000100000001110101110;
assign LUT_3[28328] = 32'b00000000000000011111100110111101;
assign LUT_3[28329] = 32'b00000000000000100110010010011010;
assign LUT_3[28330] = 32'b00000000000000100001101110100001;
assign LUT_3[28331] = 32'b00000000000000101000011001111110;
assign LUT_3[28332] = 32'b00000000000000011100110100110011;
assign LUT_3[28333] = 32'b00000000000000100011100000010000;
assign LUT_3[28334] = 32'b00000000000000011110111100010111;
assign LUT_3[28335] = 32'b00000000000000100101100111110100;
assign LUT_3[28336] = 32'b00000000000000011101100000111010;
assign LUT_3[28337] = 32'b00000000000000100100001100010111;
assign LUT_3[28338] = 32'b00000000000000011111101000011110;
assign LUT_3[28339] = 32'b00000000000000100110010011111011;
assign LUT_3[28340] = 32'b00000000000000011010101110110000;
assign LUT_3[28341] = 32'b00000000000000100001011010001101;
assign LUT_3[28342] = 32'b00000000000000011100110110010100;
assign LUT_3[28343] = 32'b00000000000000100011100001110001;
assign LUT_3[28344] = 32'b00000000000000100010111010000000;
assign LUT_3[28345] = 32'b00000000000000101001100101011101;
assign LUT_3[28346] = 32'b00000000000000100101000001100100;
assign LUT_3[28347] = 32'b00000000000000101011101101000001;
assign LUT_3[28348] = 32'b00000000000000100000000111110110;
assign LUT_3[28349] = 32'b00000000000000100110110011010011;
assign LUT_3[28350] = 32'b00000000000000100010001111011010;
assign LUT_3[28351] = 32'b00000000000000101000111010110111;
assign LUT_3[28352] = 32'b00000000000000011000111000000010;
assign LUT_3[28353] = 32'b00000000000000011111100011011111;
assign LUT_3[28354] = 32'b00000000000000011010111111100110;
assign LUT_3[28355] = 32'b00000000000000100001101011000011;
assign LUT_3[28356] = 32'b00000000000000010110000101111000;
assign LUT_3[28357] = 32'b00000000000000011100110001010101;
assign LUT_3[28358] = 32'b00000000000000011000001101011100;
assign LUT_3[28359] = 32'b00000000000000011110111000111001;
assign LUT_3[28360] = 32'b00000000000000011110010001001000;
assign LUT_3[28361] = 32'b00000000000000100100111100100101;
assign LUT_3[28362] = 32'b00000000000000100000011000101100;
assign LUT_3[28363] = 32'b00000000000000100111000100001001;
assign LUT_3[28364] = 32'b00000000000000011011011110111110;
assign LUT_3[28365] = 32'b00000000000000100010001010011011;
assign LUT_3[28366] = 32'b00000000000000011101100110100010;
assign LUT_3[28367] = 32'b00000000000000100100010001111111;
assign LUT_3[28368] = 32'b00000000000000011100001011000101;
assign LUT_3[28369] = 32'b00000000000000100010110110100010;
assign LUT_3[28370] = 32'b00000000000000011110010010101001;
assign LUT_3[28371] = 32'b00000000000000100100111110000110;
assign LUT_3[28372] = 32'b00000000000000011001011000111011;
assign LUT_3[28373] = 32'b00000000000000100000000100011000;
assign LUT_3[28374] = 32'b00000000000000011011100000011111;
assign LUT_3[28375] = 32'b00000000000000100010001011111100;
assign LUT_3[28376] = 32'b00000000000000100001100100001011;
assign LUT_3[28377] = 32'b00000000000000101000001111101000;
assign LUT_3[28378] = 32'b00000000000000100011101011101111;
assign LUT_3[28379] = 32'b00000000000000101010010111001100;
assign LUT_3[28380] = 32'b00000000000000011110110010000001;
assign LUT_3[28381] = 32'b00000000000000100101011101011110;
assign LUT_3[28382] = 32'b00000000000000100000111001100101;
assign LUT_3[28383] = 32'b00000000000000100111100101000010;
assign LUT_3[28384] = 32'b00000000000000011010000110100010;
assign LUT_3[28385] = 32'b00000000000000100000110001111111;
assign LUT_3[28386] = 32'b00000000000000011100001110000110;
assign LUT_3[28387] = 32'b00000000000000100010111001100011;
assign LUT_3[28388] = 32'b00000000000000010111010100011000;
assign LUT_3[28389] = 32'b00000000000000011101111111110101;
assign LUT_3[28390] = 32'b00000000000000011001011011111100;
assign LUT_3[28391] = 32'b00000000000000100000000111011001;
assign LUT_3[28392] = 32'b00000000000000011111011111101000;
assign LUT_3[28393] = 32'b00000000000000100110001011000101;
assign LUT_3[28394] = 32'b00000000000000100001100111001100;
assign LUT_3[28395] = 32'b00000000000000101000010010101001;
assign LUT_3[28396] = 32'b00000000000000011100101101011110;
assign LUT_3[28397] = 32'b00000000000000100011011000111011;
assign LUT_3[28398] = 32'b00000000000000011110110101000010;
assign LUT_3[28399] = 32'b00000000000000100101100000011111;
assign LUT_3[28400] = 32'b00000000000000011101011001100101;
assign LUT_3[28401] = 32'b00000000000000100100000101000010;
assign LUT_3[28402] = 32'b00000000000000011111100001001001;
assign LUT_3[28403] = 32'b00000000000000100110001100100110;
assign LUT_3[28404] = 32'b00000000000000011010100111011011;
assign LUT_3[28405] = 32'b00000000000000100001010010111000;
assign LUT_3[28406] = 32'b00000000000000011100101110111111;
assign LUT_3[28407] = 32'b00000000000000100011011010011100;
assign LUT_3[28408] = 32'b00000000000000100010110010101011;
assign LUT_3[28409] = 32'b00000000000000101001011110001000;
assign LUT_3[28410] = 32'b00000000000000100100111010001111;
assign LUT_3[28411] = 32'b00000000000000101011100101101100;
assign LUT_3[28412] = 32'b00000000000000100000000000100001;
assign LUT_3[28413] = 32'b00000000000000100110101011111110;
assign LUT_3[28414] = 32'b00000000000000100010001000000101;
assign LUT_3[28415] = 32'b00000000000000101000110011100010;
assign LUT_3[28416] = 32'b00000000000000010011000011111010;
assign LUT_3[28417] = 32'b00000000000000011001101111010111;
assign LUT_3[28418] = 32'b00000000000000010101001011011110;
assign LUT_3[28419] = 32'b00000000000000011011110110111011;
assign LUT_3[28420] = 32'b00000000000000010000010001110000;
assign LUT_3[28421] = 32'b00000000000000010110111101001101;
assign LUT_3[28422] = 32'b00000000000000010010011001010100;
assign LUT_3[28423] = 32'b00000000000000011001000100110001;
assign LUT_3[28424] = 32'b00000000000000011000011101000000;
assign LUT_3[28425] = 32'b00000000000000011111001000011101;
assign LUT_3[28426] = 32'b00000000000000011010100100100100;
assign LUT_3[28427] = 32'b00000000000000100001010000000001;
assign LUT_3[28428] = 32'b00000000000000010101101010110110;
assign LUT_3[28429] = 32'b00000000000000011100010110010011;
assign LUT_3[28430] = 32'b00000000000000010111110010011010;
assign LUT_3[28431] = 32'b00000000000000011110011101110111;
assign LUT_3[28432] = 32'b00000000000000010110010110111101;
assign LUT_3[28433] = 32'b00000000000000011101000010011010;
assign LUT_3[28434] = 32'b00000000000000011000011110100001;
assign LUT_3[28435] = 32'b00000000000000011111001001111110;
assign LUT_3[28436] = 32'b00000000000000010011100100110011;
assign LUT_3[28437] = 32'b00000000000000011010010000010000;
assign LUT_3[28438] = 32'b00000000000000010101101100010111;
assign LUT_3[28439] = 32'b00000000000000011100010111110100;
assign LUT_3[28440] = 32'b00000000000000011011110000000011;
assign LUT_3[28441] = 32'b00000000000000100010011011100000;
assign LUT_3[28442] = 32'b00000000000000011101110111100111;
assign LUT_3[28443] = 32'b00000000000000100100100011000100;
assign LUT_3[28444] = 32'b00000000000000011000111101111001;
assign LUT_3[28445] = 32'b00000000000000011111101001010110;
assign LUT_3[28446] = 32'b00000000000000011011000101011101;
assign LUT_3[28447] = 32'b00000000000000100001110000111010;
assign LUT_3[28448] = 32'b00000000000000010100010010011010;
assign LUT_3[28449] = 32'b00000000000000011010111101110111;
assign LUT_3[28450] = 32'b00000000000000010110011001111110;
assign LUT_3[28451] = 32'b00000000000000011101000101011011;
assign LUT_3[28452] = 32'b00000000000000010001100000010000;
assign LUT_3[28453] = 32'b00000000000000011000001011101101;
assign LUT_3[28454] = 32'b00000000000000010011100111110100;
assign LUT_3[28455] = 32'b00000000000000011010010011010001;
assign LUT_3[28456] = 32'b00000000000000011001101011100000;
assign LUT_3[28457] = 32'b00000000000000100000010110111101;
assign LUT_3[28458] = 32'b00000000000000011011110011000100;
assign LUT_3[28459] = 32'b00000000000000100010011110100001;
assign LUT_3[28460] = 32'b00000000000000010110111001010110;
assign LUT_3[28461] = 32'b00000000000000011101100100110011;
assign LUT_3[28462] = 32'b00000000000000011001000000111010;
assign LUT_3[28463] = 32'b00000000000000011111101100010111;
assign LUT_3[28464] = 32'b00000000000000010111100101011101;
assign LUT_3[28465] = 32'b00000000000000011110010000111010;
assign LUT_3[28466] = 32'b00000000000000011001101101000001;
assign LUT_3[28467] = 32'b00000000000000100000011000011110;
assign LUT_3[28468] = 32'b00000000000000010100110011010011;
assign LUT_3[28469] = 32'b00000000000000011011011110110000;
assign LUT_3[28470] = 32'b00000000000000010110111010110111;
assign LUT_3[28471] = 32'b00000000000000011101100110010100;
assign LUT_3[28472] = 32'b00000000000000011100111110100011;
assign LUT_3[28473] = 32'b00000000000000100011101010000000;
assign LUT_3[28474] = 32'b00000000000000011111000110000111;
assign LUT_3[28475] = 32'b00000000000000100101110001100100;
assign LUT_3[28476] = 32'b00000000000000011010001100011001;
assign LUT_3[28477] = 32'b00000000000000100000110111110110;
assign LUT_3[28478] = 32'b00000000000000011100010011111101;
assign LUT_3[28479] = 32'b00000000000000100010111111011010;
assign LUT_3[28480] = 32'b00000000000000010010111100100101;
assign LUT_3[28481] = 32'b00000000000000011001101000000010;
assign LUT_3[28482] = 32'b00000000000000010101000100001001;
assign LUT_3[28483] = 32'b00000000000000011011101111100110;
assign LUT_3[28484] = 32'b00000000000000010000001010011011;
assign LUT_3[28485] = 32'b00000000000000010110110101111000;
assign LUT_3[28486] = 32'b00000000000000010010010001111111;
assign LUT_3[28487] = 32'b00000000000000011000111101011100;
assign LUT_3[28488] = 32'b00000000000000011000010101101011;
assign LUT_3[28489] = 32'b00000000000000011111000001001000;
assign LUT_3[28490] = 32'b00000000000000011010011101001111;
assign LUT_3[28491] = 32'b00000000000000100001001000101100;
assign LUT_3[28492] = 32'b00000000000000010101100011100001;
assign LUT_3[28493] = 32'b00000000000000011100001110111110;
assign LUT_3[28494] = 32'b00000000000000010111101011000101;
assign LUT_3[28495] = 32'b00000000000000011110010110100010;
assign LUT_3[28496] = 32'b00000000000000010110001111101000;
assign LUT_3[28497] = 32'b00000000000000011100111011000101;
assign LUT_3[28498] = 32'b00000000000000011000010111001100;
assign LUT_3[28499] = 32'b00000000000000011111000010101001;
assign LUT_3[28500] = 32'b00000000000000010011011101011110;
assign LUT_3[28501] = 32'b00000000000000011010001000111011;
assign LUT_3[28502] = 32'b00000000000000010101100101000010;
assign LUT_3[28503] = 32'b00000000000000011100010000011111;
assign LUT_3[28504] = 32'b00000000000000011011101000101110;
assign LUT_3[28505] = 32'b00000000000000100010010100001011;
assign LUT_3[28506] = 32'b00000000000000011101110000010010;
assign LUT_3[28507] = 32'b00000000000000100100011011101111;
assign LUT_3[28508] = 32'b00000000000000011000110110100100;
assign LUT_3[28509] = 32'b00000000000000011111100010000001;
assign LUT_3[28510] = 32'b00000000000000011010111110001000;
assign LUT_3[28511] = 32'b00000000000000100001101001100101;
assign LUT_3[28512] = 32'b00000000000000010100001011000101;
assign LUT_3[28513] = 32'b00000000000000011010110110100010;
assign LUT_3[28514] = 32'b00000000000000010110010010101001;
assign LUT_3[28515] = 32'b00000000000000011100111110000110;
assign LUT_3[28516] = 32'b00000000000000010001011000111011;
assign LUT_3[28517] = 32'b00000000000000011000000100011000;
assign LUT_3[28518] = 32'b00000000000000010011100000011111;
assign LUT_3[28519] = 32'b00000000000000011010001011111100;
assign LUT_3[28520] = 32'b00000000000000011001100100001011;
assign LUT_3[28521] = 32'b00000000000000100000001111101000;
assign LUT_3[28522] = 32'b00000000000000011011101011101111;
assign LUT_3[28523] = 32'b00000000000000100010010111001100;
assign LUT_3[28524] = 32'b00000000000000010110110010000001;
assign LUT_3[28525] = 32'b00000000000000011101011101011110;
assign LUT_3[28526] = 32'b00000000000000011000111001100101;
assign LUT_3[28527] = 32'b00000000000000011111100101000010;
assign LUT_3[28528] = 32'b00000000000000010111011110001000;
assign LUT_3[28529] = 32'b00000000000000011110001001100101;
assign LUT_3[28530] = 32'b00000000000000011001100101101100;
assign LUT_3[28531] = 32'b00000000000000100000010001001001;
assign LUT_3[28532] = 32'b00000000000000010100101011111110;
assign LUT_3[28533] = 32'b00000000000000011011010111011011;
assign LUT_3[28534] = 32'b00000000000000010110110011100010;
assign LUT_3[28535] = 32'b00000000000000011101011110111111;
assign LUT_3[28536] = 32'b00000000000000011100110111001110;
assign LUT_3[28537] = 32'b00000000000000100011100010101011;
assign LUT_3[28538] = 32'b00000000000000011110111110110010;
assign LUT_3[28539] = 32'b00000000000000100101101010001111;
assign LUT_3[28540] = 32'b00000000000000011010000101000100;
assign LUT_3[28541] = 32'b00000000000000100000110000100001;
assign LUT_3[28542] = 32'b00000000000000011100001100101000;
assign LUT_3[28543] = 32'b00000000000000100010111000000101;
assign LUT_3[28544] = 32'b00000000000000010101001110111000;
assign LUT_3[28545] = 32'b00000000000000011011111010010101;
assign LUT_3[28546] = 32'b00000000000000010111010110011100;
assign LUT_3[28547] = 32'b00000000000000011110000001111001;
assign LUT_3[28548] = 32'b00000000000000010010011100101110;
assign LUT_3[28549] = 32'b00000000000000011001001000001011;
assign LUT_3[28550] = 32'b00000000000000010100100100010010;
assign LUT_3[28551] = 32'b00000000000000011011001111101111;
assign LUT_3[28552] = 32'b00000000000000011010100111111110;
assign LUT_3[28553] = 32'b00000000000000100001010011011011;
assign LUT_3[28554] = 32'b00000000000000011100101111100010;
assign LUT_3[28555] = 32'b00000000000000100011011010111111;
assign LUT_3[28556] = 32'b00000000000000010111110101110100;
assign LUT_3[28557] = 32'b00000000000000011110100001010001;
assign LUT_3[28558] = 32'b00000000000000011001111101011000;
assign LUT_3[28559] = 32'b00000000000000100000101000110101;
assign LUT_3[28560] = 32'b00000000000000011000100001111011;
assign LUT_3[28561] = 32'b00000000000000011111001101011000;
assign LUT_3[28562] = 32'b00000000000000011010101001011111;
assign LUT_3[28563] = 32'b00000000000000100001010100111100;
assign LUT_3[28564] = 32'b00000000000000010101101111110001;
assign LUT_3[28565] = 32'b00000000000000011100011011001110;
assign LUT_3[28566] = 32'b00000000000000010111110111010101;
assign LUT_3[28567] = 32'b00000000000000011110100010110010;
assign LUT_3[28568] = 32'b00000000000000011101111011000001;
assign LUT_3[28569] = 32'b00000000000000100100100110011110;
assign LUT_3[28570] = 32'b00000000000000100000000010100101;
assign LUT_3[28571] = 32'b00000000000000100110101110000010;
assign LUT_3[28572] = 32'b00000000000000011011001000110111;
assign LUT_3[28573] = 32'b00000000000000100001110100010100;
assign LUT_3[28574] = 32'b00000000000000011101010000011011;
assign LUT_3[28575] = 32'b00000000000000100011111011111000;
assign LUT_3[28576] = 32'b00000000000000010110011101011000;
assign LUT_3[28577] = 32'b00000000000000011101001000110101;
assign LUT_3[28578] = 32'b00000000000000011000100100111100;
assign LUT_3[28579] = 32'b00000000000000011111010000011001;
assign LUT_3[28580] = 32'b00000000000000010011101011001110;
assign LUT_3[28581] = 32'b00000000000000011010010110101011;
assign LUT_3[28582] = 32'b00000000000000010101110010110010;
assign LUT_3[28583] = 32'b00000000000000011100011110001111;
assign LUT_3[28584] = 32'b00000000000000011011110110011110;
assign LUT_3[28585] = 32'b00000000000000100010100001111011;
assign LUT_3[28586] = 32'b00000000000000011101111110000010;
assign LUT_3[28587] = 32'b00000000000000100100101001011111;
assign LUT_3[28588] = 32'b00000000000000011001000100010100;
assign LUT_3[28589] = 32'b00000000000000011111101111110001;
assign LUT_3[28590] = 32'b00000000000000011011001011111000;
assign LUT_3[28591] = 32'b00000000000000100001110111010101;
assign LUT_3[28592] = 32'b00000000000000011001110000011011;
assign LUT_3[28593] = 32'b00000000000000100000011011111000;
assign LUT_3[28594] = 32'b00000000000000011011110111111111;
assign LUT_3[28595] = 32'b00000000000000100010100011011100;
assign LUT_3[28596] = 32'b00000000000000010110111110010001;
assign LUT_3[28597] = 32'b00000000000000011101101001101110;
assign LUT_3[28598] = 32'b00000000000000011001000101110101;
assign LUT_3[28599] = 32'b00000000000000011111110001010010;
assign LUT_3[28600] = 32'b00000000000000011111001001100001;
assign LUT_3[28601] = 32'b00000000000000100101110100111110;
assign LUT_3[28602] = 32'b00000000000000100001010001000101;
assign LUT_3[28603] = 32'b00000000000000100111111100100010;
assign LUT_3[28604] = 32'b00000000000000011100010111010111;
assign LUT_3[28605] = 32'b00000000000000100011000010110100;
assign LUT_3[28606] = 32'b00000000000000011110011110111011;
assign LUT_3[28607] = 32'b00000000000000100101001010011000;
assign LUT_3[28608] = 32'b00000000000000010101000111100011;
assign LUT_3[28609] = 32'b00000000000000011011110011000000;
assign LUT_3[28610] = 32'b00000000000000010111001111000111;
assign LUT_3[28611] = 32'b00000000000000011101111010100100;
assign LUT_3[28612] = 32'b00000000000000010010010101011001;
assign LUT_3[28613] = 32'b00000000000000011001000000110110;
assign LUT_3[28614] = 32'b00000000000000010100011100111101;
assign LUT_3[28615] = 32'b00000000000000011011001000011010;
assign LUT_3[28616] = 32'b00000000000000011010100000101001;
assign LUT_3[28617] = 32'b00000000000000100001001100000110;
assign LUT_3[28618] = 32'b00000000000000011100101000001101;
assign LUT_3[28619] = 32'b00000000000000100011010011101010;
assign LUT_3[28620] = 32'b00000000000000010111101110011111;
assign LUT_3[28621] = 32'b00000000000000011110011001111100;
assign LUT_3[28622] = 32'b00000000000000011001110110000011;
assign LUT_3[28623] = 32'b00000000000000100000100001100000;
assign LUT_3[28624] = 32'b00000000000000011000011010100110;
assign LUT_3[28625] = 32'b00000000000000011111000110000011;
assign LUT_3[28626] = 32'b00000000000000011010100010001010;
assign LUT_3[28627] = 32'b00000000000000100001001101100111;
assign LUT_3[28628] = 32'b00000000000000010101101000011100;
assign LUT_3[28629] = 32'b00000000000000011100010011111001;
assign LUT_3[28630] = 32'b00000000000000010111110000000000;
assign LUT_3[28631] = 32'b00000000000000011110011011011101;
assign LUT_3[28632] = 32'b00000000000000011101110011101100;
assign LUT_3[28633] = 32'b00000000000000100100011111001001;
assign LUT_3[28634] = 32'b00000000000000011111111011010000;
assign LUT_3[28635] = 32'b00000000000000100110100110101101;
assign LUT_3[28636] = 32'b00000000000000011011000001100010;
assign LUT_3[28637] = 32'b00000000000000100001101100111111;
assign LUT_3[28638] = 32'b00000000000000011101001001000110;
assign LUT_3[28639] = 32'b00000000000000100011110100100011;
assign LUT_3[28640] = 32'b00000000000000010110010110000011;
assign LUT_3[28641] = 32'b00000000000000011101000001100000;
assign LUT_3[28642] = 32'b00000000000000011000011101100111;
assign LUT_3[28643] = 32'b00000000000000011111001001000100;
assign LUT_3[28644] = 32'b00000000000000010011100011111001;
assign LUT_3[28645] = 32'b00000000000000011010001111010110;
assign LUT_3[28646] = 32'b00000000000000010101101011011101;
assign LUT_3[28647] = 32'b00000000000000011100010110111010;
assign LUT_3[28648] = 32'b00000000000000011011101111001001;
assign LUT_3[28649] = 32'b00000000000000100010011010100110;
assign LUT_3[28650] = 32'b00000000000000011101110110101101;
assign LUT_3[28651] = 32'b00000000000000100100100010001010;
assign LUT_3[28652] = 32'b00000000000000011000111100111111;
assign LUT_3[28653] = 32'b00000000000000011111101000011100;
assign LUT_3[28654] = 32'b00000000000000011011000100100011;
assign LUT_3[28655] = 32'b00000000000000100001110000000000;
assign LUT_3[28656] = 32'b00000000000000011001101001000110;
assign LUT_3[28657] = 32'b00000000000000100000010100100011;
assign LUT_3[28658] = 32'b00000000000000011011110000101010;
assign LUT_3[28659] = 32'b00000000000000100010011100000111;
assign LUT_3[28660] = 32'b00000000000000010110110110111100;
assign LUT_3[28661] = 32'b00000000000000011101100010011001;
assign LUT_3[28662] = 32'b00000000000000011000111110100000;
assign LUT_3[28663] = 32'b00000000000000011111101001111101;
assign LUT_3[28664] = 32'b00000000000000011111000010001100;
assign LUT_3[28665] = 32'b00000000000000100101101101101001;
assign LUT_3[28666] = 32'b00000000000000100001001001110000;
assign LUT_3[28667] = 32'b00000000000000100111110101001101;
assign LUT_3[28668] = 32'b00000000000000011100010000000010;
assign LUT_3[28669] = 32'b00000000000000100010111011011111;
assign LUT_3[28670] = 32'b00000000000000011110010111100110;
assign LUT_3[28671] = 32'b00000000000000100101000011000011;
assign LUT_3[28672] = 32'b00000000000000001111010101011101;
assign LUT_3[28673] = 32'b00000000000000010110000000111010;
assign LUT_3[28674] = 32'b00000000000000010001011101000001;
assign LUT_3[28675] = 32'b00000000000000011000001000011110;
assign LUT_3[28676] = 32'b00000000000000001100100011010011;
assign LUT_3[28677] = 32'b00000000000000010011001110110000;
assign LUT_3[28678] = 32'b00000000000000001110101010110111;
assign LUT_3[28679] = 32'b00000000000000010101010110010100;
assign LUT_3[28680] = 32'b00000000000000010100101110100011;
assign LUT_3[28681] = 32'b00000000000000011011011010000000;
assign LUT_3[28682] = 32'b00000000000000010110110110000111;
assign LUT_3[28683] = 32'b00000000000000011101100001100100;
assign LUT_3[28684] = 32'b00000000000000010001111100011001;
assign LUT_3[28685] = 32'b00000000000000011000100111110110;
assign LUT_3[28686] = 32'b00000000000000010100000011111101;
assign LUT_3[28687] = 32'b00000000000000011010101111011010;
assign LUT_3[28688] = 32'b00000000000000010010101000100000;
assign LUT_3[28689] = 32'b00000000000000011001010011111101;
assign LUT_3[28690] = 32'b00000000000000010100110000000100;
assign LUT_3[28691] = 32'b00000000000000011011011011100001;
assign LUT_3[28692] = 32'b00000000000000001111110110010110;
assign LUT_3[28693] = 32'b00000000000000010110100001110011;
assign LUT_3[28694] = 32'b00000000000000010001111101111010;
assign LUT_3[28695] = 32'b00000000000000011000101001010111;
assign LUT_3[28696] = 32'b00000000000000011000000001100110;
assign LUT_3[28697] = 32'b00000000000000011110101101000011;
assign LUT_3[28698] = 32'b00000000000000011010001001001010;
assign LUT_3[28699] = 32'b00000000000000100000110100100111;
assign LUT_3[28700] = 32'b00000000000000010101001111011100;
assign LUT_3[28701] = 32'b00000000000000011011111010111001;
assign LUT_3[28702] = 32'b00000000000000010111010111000000;
assign LUT_3[28703] = 32'b00000000000000011110000010011101;
assign LUT_3[28704] = 32'b00000000000000010000100011111101;
assign LUT_3[28705] = 32'b00000000000000010111001111011010;
assign LUT_3[28706] = 32'b00000000000000010010101011100001;
assign LUT_3[28707] = 32'b00000000000000011001010110111110;
assign LUT_3[28708] = 32'b00000000000000001101110001110011;
assign LUT_3[28709] = 32'b00000000000000010100011101010000;
assign LUT_3[28710] = 32'b00000000000000001111111001010111;
assign LUT_3[28711] = 32'b00000000000000010110100100110100;
assign LUT_3[28712] = 32'b00000000000000010101111101000011;
assign LUT_3[28713] = 32'b00000000000000011100101000100000;
assign LUT_3[28714] = 32'b00000000000000011000000100100111;
assign LUT_3[28715] = 32'b00000000000000011110110000000100;
assign LUT_3[28716] = 32'b00000000000000010011001010111001;
assign LUT_3[28717] = 32'b00000000000000011001110110010110;
assign LUT_3[28718] = 32'b00000000000000010101010010011101;
assign LUT_3[28719] = 32'b00000000000000011011111101111010;
assign LUT_3[28720] = 32'b00000000000000010011110111000000;
assign LUT_3[28721] = 32'b00000000000000011010100010011101;
assign LUT_3[28722] = 32'b00000000000000010101111110100100;
assign LUT_3[28723] = 32'b00000000000000011100101010000001;
assign LUT_3[28724] = 32'b00000000000000010001000100110110;
assign LUT_3[28725] = 32'b00000000000000010111110000010011;
assign LUT_3[28726] = 32'b00000000000000010011001100011010;
assign LUT_3[28727] = 32'b00000000000000011001110111110111;
assign LUT_3[28728] = 32'b00000000000000011001010000000110;
assign LUT_3[28729] = 32'b00000000000000011111111011100011;
assign LUT_3[28730] = 32'b00000000000000011011010111101010;
assign LUT_3[28731] = 32'b00000000000000100010000011000111;
assign LUT_3[28732] = 32'b00000000000000010110011101111100;
assign LUT_3[28733] = 32'b00000000000000011101001001011001;
assign LUT_3[28734] = 32'b00000000000000011000100101100000;
assign LUT_3[28735] = 32'b00000000000000011111010000111101;
assign LUT_3[28736] = 32'b00000000000000001111001110001000;
assign LUT_3[28737] = 32'b00000000000000010101111001100101;
assign LUT_3[28738] = 32'b00000000000000010001010101101100;
assign LUT_3[28739] = 32'b00000000000000011000000001001001;
assign LUT_3[28740] = 32'b00000000000000001100011011111110;
assign LUT_3[28741] = 32'b00000000000000010011000111011011;
assign LUT_3[28742] = 32'b00000000000000001110100011100010;
assign LUT_3[28743] = 32'b00000000000000010101001110111111;
assign LUT_3[28744] = 32'b00000000000000010100100111001110;
assign LUT_3[28745] = 32'b00000000000000011011010010101011;
assign LUT_3[28746] = 32'b00000000000000010110101110110010;
assign LUT_3[28747] = 32'b00000000000000011101011010001111;
assign LUT_3[28748] = 32'b00000000000000010001110101000100;
assign LUT_3[28749] = 32'b00000000000000011000100000100001;
assign LUT_3[28750] = 32'b00000000000000010011111100101000;
assign LUT_3[28751] = 32'b00000000000000011010101000000101;
assign LUT_3[28752] = 32'b00000000000000010010100001001011;
assign LUT_3[28753] = 32'b00000000000000011001001100101000;
assign LUT_3[28754] = 32'b00000000000000010100101000101111;
assign LUT_3[28755] = 32'b00000000000000011011010100001100;
assign LUT_3[28756] = 32'b00000000000000001111101111000001;
assign LUT_3[28757] = 32'b00000000000000010110011010011110;
assign LUT_3[28758] = 32'b00000000000000010001110110100101;
assign LUT_3[28759] = 32'b00000000000000011000100010000010;
assign LUT_3[28760] = 32'b00000000000000010111111010010001;
assign LUT_3[28761] = 32'b00000000000000011110100101101110;
assign LUT_3[28762] = 32'b00000000000000011010000001110101;
assign LUT_3[28763] = 32'b00000000000000100000101101010010;
assign LUT_3[28764] = 32'b00000000000000010101001000000111;
assign LUT_3[28765] = 32'b00000000000000011011110011100100;
assign LUT_3[28766] = 32'b00000000000000010111001111101011;
assign LUT_3[28767] = 32'b00000000000000011101111011001000;
assign LUT_3[28768] = 32'b00000000000000010000011100101000;
assign LUT_3[28769] = 32'b00000000000000010111001000000101;
assign LUT_3[28770] = 32'b00000000000000010010100100001100;
assign LUT_3[28771] = 32'b00000000000000011001001111101001;
assign LUT_3[28772] = 32'b00000000000000001101101010011110;
assign LUT_3[28773] = 32'b00000000000000010100010101111011;
assign LUT_3[28774] = 32'b00000000000000001111110010000010;
assign LUT_3[28775] = 32'b00000000000000010110011101011111;
assign LUT_3[28776] = 32'b00000000000000010101110101101110;
assign LUT_3[28777] = 32'b00000000000000011100100001001011;
assign LUT_3[28778] = 32'b00000000000000010111111101010010;
assign LUT_3[28779] = 32'b00000000000000011110101000101111;
assign LUT_3[28780] = 32'b00000000000000010011000011100100;
assign LUT_3[28781] = 32'b00000000000000011001101111000001;
assign LUT_3[28782] = 32'b00000000000000010101001011001000;
assign LUT_3[28783] = 32'b00000000000000011011110110100101;
assign LUT_3[28784] = 32'b00000000000000010011101111101011;
assign LUT_3[28785] = 32'b00000000000000011010011011001000;
assign LUT_3[28786] = 32'b00000000000000010101110111001111;
assign LUT_3[28787] = 32'b00000000000000011100100010101100;
assign LUT_3[28788] = 32'b00000000000000010000111101100001;
assign LUT_3[28789] = 32'b00000000000000010111101000111110;
assign LUT_3[28790] = 32'b00000000000000010011000101000101;
assign LUT_3[28791] = 32'b00000000000000011001110000100010;
assign LUT_3[28792] = 32'b00000000000000011001001000110001;
assign LUT_3[28793] = 32'b00000000000000011111110100001110;
assign LUT_3[28794] = 32'b00000000000000011011010000010101;
assign LUT_3[28795] = 32'b00000000000000100001111011110010;
assign LUT_3[28796] = 32'b00000000000000010110010110100111;
assign LUT_3[28797] = 32'b00000000000000011101000010000100;
assign LUT_3[28798] = 32'b00000000000000011000011110001011;
assign LUT_3[28799] = 32'b00000000000000011111001001101000;
assign LUT_3[28800] = 32'b00000000000000010001100000011011;
assign LUT_3[28801] = 32'b00000000000000011000001011111000;
assign LUT_3[28802] = 32'b00000000000000010011100111111111;
assign LUT_3[28803] = 32'b00000000000000011010010011011100;
assign LUT_3[28804] = 32'b00000000000000001110101110010001;
assign LUT_3[28805] = 32'b00000000000000010101011001101110;
assign LUT_3[28806] = 32'b00000000000000010000110101110101;
assign LUT_3[28807] = 32'b00000000000000010111100001010010;
assign LUT_3[28808] = 32'b00000000000000010110111001100001;
assign LUT_3[28809] = 32'b00000000000000011101100100111110;
assign LUT_3[28810] = 32'b00000000000000011001000001000101;
assign LUT_3[28811] = 32'b00000000000000011111101100100010;
assign LUT_3[28812] = 32'b00000000000000010100000111010111;
assign LUT_3[28813] = 32'b00000000000000011010110010110100;
assign LUT_3[28814] = 32'b00000000000000010110001110111011;
assign LUT_3[28815] = 32'b00000000000000011100111010011000;
assign LUT_3[28816] = 32'b00000000000000010100110011011110;
assign LUT_3[28817] = 32'b00000000000000011011011110111011;
assign LUT_3[28818] = 32'b00000000000000010110111011000010;
assign LUT_3[28819] = 32'b00000000000000011101100110011111;
assign LUT_3[28820] = 32'b00000000000000010010000001010100;
assign LUT_3[28821] = 32'b00000000000000011000101100110001;
assign LUT_3[28822] = 32'b00000000000000010100001000111000;
assign LUT_3[28823] = 32'b00000000000000011010110100010101;
assign LUT_3[28824] = 32'b00000000000000011010001100100100;
assign LUT_3[28825] = 32'b00000000000000100000111000000001;
assign LUT_3[28826] = 32'b00000000000000011100010100001000;
assign LUT_3[28827] = 32'b00000000000000100010111111100101;
assign LUT_3[28828] = 32'b00000000000000010111011010011010;
assign LUT_3[28829] = 32'b00000000000000011110000101110111;
assign LUT_3[28830] = 32'b00000000000000011001100001111110;
assign LUT_3[28831] = 32'b00000000000000100000001101011011;
assign LUT_3[28832] = 32'b00000000000000010010101110111011;
assign LUT_3[28833] = 32'b00000000000000011001011010011000;
assign LUT_3[28834] = 32'b00000000000000010100110110011111;
assign LUT_3[28835] = 32'b00000000000000011011100001111100;
assign LUT_3[28836] = 32'b00000000000000001111111100110001;
assign LUT_3[28837] = 32'b00000000000000010110101000001110;
assign LUT_3[28838] = 32'b00000000000000010010000100010101;
assign LUT_3[28839] = 32'b00000000000000011000101111110010;
assign LUT_3[28840] = 32'b00000000000000011000001000000001;
assign LUT_3[28841] = 32'b00000000000000011110110011011110;
assign LUT_3[28842] = 32'b00000000000000011010001111100101;
assign LUT_3[28843] = 32'b00000000000000100000111011000010;
assign LUT_3[28844] = 32'b00000000000000010101010101110111;
assign LUT_3[28845] = 32'b00000000000000011100000001010100;
assign LUT_3[28846] = 32'b00000000000000010111011101011011;
assign LUT_3[28847] = 32'b00000000000000011110001000111000;
assign LUT_3[28848] = 32'b00000000000000010110000001111110;
assign LUT_3[28849] = 32'b00000000000000011100101101011011;
assign LUT_3[28850] = 32'b00000000000000011000001001100010;
assign LUT_3[28851] = 32'b00000000000000011110110100111111;
assign LUT_3[28852] = 32'b00000000000000010011001111110100;
assign LUT_3[28853] = 32'b00000000000000011001111011010001;
assign LUT_3[28854] = 32'b00000000000000010101010111011000;
assign LUT_3[28855] = 32'b00000000000000011100000010110101;
assign LUT_3[28856] = 32'b00000000000000011011011011000100;
assign LUT_3[28857] = 32'b00000000000000100010000110100001;
assign LUT_3[28858] = 32'b00000000000000011101100010101000;
assign LUT_3[28859] = 32'b00000000000000100100001110000101;
assign LUT_3[28860] = 32'b00000000000000011000101000111010;
assign LUT_3[28861] = 32'b00000000000000011111010100010111;
assign LUT_3[28862] = 32'b00000000000000011010110000011110;
assign LUT_3[28863] = 32'b00000000000000100001011011111011;
assign LUT_3[28864] = 32'b00000000000000010001011001000110;
assign LUT_3[28865] = 32'b00000000000000011000000100100011;
assign LUT_3[28866] = 32'b00000000000000010011100000101010;
assign LUT_3[28867] = 32'b00000000000000011010001100000111;
assign LUT_3[28868] = 32'b00000000000000001110100110111100;
assign LUT_3[28869] = 32'b00000000000000010101010010011001;
assign LUT_3[28870] = 32'b00000000000000010000101110100000;
assign LUT_3[28871] = 32'b00000000000000010111011001111101;
assign LUT_3[28872] = 32'b00000000000000010110110010001100;
assign LUT_3[28873] = 32'b00000000000000011101011101101001;
assign LUT_3[28874] = 32'b00000000000000011000111001110000;
assign LUT_3[28875] = 32'b00000000000000011111100101001101;
assign LUT_3[28876] = 32'b00000000000000010100000000000010;
assign LUT_3[28877] = 32'b00000000000000011010101011011111;
assign LUT_3[28878] = 32'b00000000000000010110000111100110;
assign LUT_3[28879] = 32'b00000000000000011100110011000011;
assign LUT_3[28880] = 32'b00000000000000010100101100001001;
assign LUT_3[28881] = 32'b00000000000000011011010111100110;
assign LUT_3[28882] = 32'b00000000000000010110110011101101;
assign LUT_3[28883] = 32'b00000000000000011101011111001010;
assign LUT_3[28884] = 32'b00000000000000010001111001111111;
assign LUT_3[28885] = 32'b00000000000000011000100101011100;
assign LUT_3[28886] = 32'b00000000000000010100000001100011;
assign LUT_3[28887] = 32'b00000000000000011010101101000000;
assign LUT_3[28888] = 32'b00000000000000011010000101001111;
assign LUT_3[28889] = 32'b00000000000000100000110000101100;
assign LUT_3[28890] = 32'b00000000000000011100001100110011;
assign LUT_3[28891] = 32'b00000000000000100010111000010000;
assign LUT_3[28892] = 32'b00000000000000010111010011000101;
assign LUT_3[28893] = 32'b00000000000000011101111110100010;
assign LUT_3[28894] = 32'b00000000000000011001011010101001;
assign LUT_3[28895] = 32'b00000000000000100000000110000110;
assign LUT_3[28896] = 32'b00000000000000010010100111100110;
assign LUT_3[28897] = 32'b00000000000000011001010011000011;
assign LUT_3[28898] = 32'b00000000000000010100101111001010;
assign LUT_3[28899] = 32'b00000000000000011011011010100111;
assign LUT_3[28900] = 32'b00000000000000001111110101011100;
assign LUT_3[28901] = 32'b00000000000000010110100000111001;
assign LUT_3[28902] = 32'b00000000000000010001111101000000;
assign LUT_3[28903] = 32'b00000000000000011000101000011101;
assign LUT_3[28904] = 32'b00000000000000011000000000101100;
assign LUT_3[28905] = 32'b00000000000000011110101100001001;
assign LUT_3[28906] = 32'b00000000000000011010001000010000;
assign LUT_3[28907] = 32'b00000000000000100000110011101101;
assign LUT_3[28908] = 32'b00000000000000010101001110100010;
assign LUT_3[28909] = 32'b00000000000000011011111001111111;
assign LUT_3[28910] = 32'b00000000000000010111010110000110;
assign LUT_3[28911] = 32'b00000000000000011110000001100011;
assign LUT_3[28912] = 32'b00000000000000010101111010101001;
assign LUT_3[28913] = 32'b00000000000000011100100110000110;
assign LUT_3[28914] = 32'b00000000000000011000000010001101;
assign LUT_3[28915] = 32'b00000000000000011110101101101010;
assign LUT_3[28916] = 32'b00000000000000010011001000011111;
assign LUT_3[28917] = 32'b00000000000000011001110011111100;
assign LUT_3[28918] = 32'b00000000000000010101010000000011;
assign LUT_3[28919] = 32'b00000000000000011011111011100000;
assign LUT_3[28920] = 32'b00000000000000011011010011101111;
assign LUT_3[28921] = 32'b00000000000000100001111111001100;
assign LUT_3[28922] = 32'b00000000000000011101011011010011;
assign LUT_3[28923] = 32'b00000000000000100100000110110000;
assign LUT_3[28924] = 32'b00000000000000011000100001100101;
assign LUT_3[28925] = 32'b00000000000000011111001101000010;
assign LUT_3[28926] = 32'b00000000000000011010101001001001;
assign LUT_3[28927] = 32'b00000000000000100001010100100110;
assign LUT_3[28928] = 32'b00000000000000001011100100111110;
assign LUT_3[28929] = 32'b00000000000000010010010000011011;
assign LUT_3[28930] = 32'b00000000000000001101101100100010;
assign LUT_3[28931] = 32'b00000000000000010100010111111111;
assign LUT_3[28932] = 32'b00000000000000001000110010110100;
assign LUT_3[28933] = 32'b00000000000000001111011110010001;
assign LUT_3[28934] = 32'b00000000000000001010111010011000;
assign LUT_3[28935] = 32'b00000000000000010001100101110101;
assign LUT_3[28936] = 32'b00000000000000010000111110000100;
assign LUT_3[28937] = 32'b00000000000000010111101001100001;
assign LUT_3[28938] = 32'b00000000000000010011000101101000;
assign LUT_3[28939] = 32'b00000000000000011001110001000101;
assign LUT_3[28940] = 32'b00000000000000001110001011111010;
assign LUT_3[28941] = 32'b00000000000000010100110111010111;
assign LUT_3[28942] = 32'b00000000000000010000010011011110;
assign LUT_3[28943] = 32'b00000000000000010110111110111011;
assign LUT_3[28944] = 32'b00000000000000001110111000000001;
assign LUT_3[28945] = 32'b00000000000000010101100011011110;
assign LUT_3[28946] = 32'b00000000000000010000111111100101;
assign LUT_3[28947] = 32'b00000000000000010111101011000010;
assign LUT_3[28948] = 32'b00000000000000001100000101110111;
assign LUT_3[28949] = 32'b00000000000000010010110001010100;
assign LUT_3[28950] = 32'b00000000000000001110001101011011;
assign LUT_3[28951] = 32'b00000000000000010100111000111000;
assign LUT_3[28952] = 32'b00000000000000010100010001000111;
assign LUT_3[28953] = 32'b00000000000000011010111100100100;
assign LUT_3[28954] = 32'b00000000000000010110011000101011;
assign LUT_3[28955] = 32'b00000000000000011101000100001000;
assign LUT_3[28956] = 32'b00000000000000010001011110111101;
assign LUT_3[28957] = 32'b00000000000000011000001010011010;
assign LUT_3[28958] = 32'b00000000000000010011100110100001;
assign LUT_3[28959] = 32'b00000000000000011010010001111110;
assign LUT_3[28960] = 32'b00000000000000001100110011011110;
assign LUT_3[28961] = 32'b00000000000000010011011110111011;
assign LUT_3[28962] = 32'b00000000000000001110111011000010;
assign LUT_3[28963] = 32'b00000000000000010101100110011111;
assign LUT_3[28964] = 32'b00000000000000001010000001010100;
assign LUT_3[28965] = 32'b00000000000000010000101100110001;
assign LUT_3[28966] = 32'b00000000000000001100001000111000;
assign LUT_3[28967] = 32'b00000000000000010010110100010101;
assign LUT_3[28968] = 32'b00000000000000010010001100100100;
assign LUT_3[28969] = 32'b00000000000000011000111000000001;
assign LUT_3[28970] = 32'b00000000000000010100010100001000;
assign LUT_3[28971] = 32'b00000000000000011010111111100101;
assign LUT_3[28972] = 32'b00000000000000001111011010011010;
assign LUT_3[28973] = 32'b00000000000000010110000101110111;
assign LUT_3[28974] = 32'b00000000000000010001100001111110;
assign LUT_3[28975] = 32'b00000000000000011000001101011011;
assign LUT_3[28976] = 32'b00000000000000010000000110100001;
assign LUT_3[28977] = 32'b00000000000000010110110001111110;
assign LUT_3[28978] = 32'b00000000000000010010001110000101;
assign LUT_3[28979] = 32'b00000000000000011000111001100010;
assign LUT_3[28980] = 32'b00000000000000001101010100010111;
assign LUT_3[28981] = 32'b00000000000000010011111111110100;
assign LUT_3[28982] = 32'b00000000000000001111011011111011;
assign LUT_3[28983] = 32'b00000000000000010110000111011000;
assign LUT_3[28984] = 32'b00000000000000010101011111100111;
assign LUT_3[28985] = 32'b00000000000000011100001011000100;
assign LUT_3[28986] = 32'b00000000000000010111100111001011;
assign LUT_3[28987] = 32'b00000000000000011110010010101000;
assign LUT_3[28988] = 32'b00000000000000010010101101011101;
assign LUT_3[28989] = 32'b00000000000000011001011000111010;
assign LUT_3[28990] = 32'b00000000000000010100110101000001;
assign LUT_3[28991] = 32'b00000000000000011011100000011110;
assign LUT_3[28992] = 32'b00000000000000001011011101101001;
assign LUT_3[28993] = 32'b00000000000000010010001001000110;
assign LUT_3[28994] = 32'b00000000000000001101100101001101;
assign LUT_3[28995] = 32'b00000000000000010100010000101010;
assign LUT_3[28996] = 32'b00000000000000001000101011011111;
assign LUT_3[28997] = 32'b00000000000000001111010110111100;
assign LUT_3[28998] = 32'b00000000000000001010110011000011;
assign LUT_3[28999] = 32'b00000000000000010001011110100000;
assign LUT_3[29000] = 32'b00000000000000010000110110101111;
assign LUT_3[29001] = 32'b00000000000000010111100010001100;
assign LUT_3[29002] = 32'b00000000000000010010111110010011;
assign LUT_3[29003] = 32'b00000000000000011001101001110000;
assign LUT_3[29004] = 32'b00000000000000001110000100100101;
assign LUT_3[29005] = 32'b00000000000000010100110000000010;
assign LUT_3[29006] = 32'b00000000000000010000001100001001;
assign LUT_3[29007] = 32'b00000000000000010110110111100110;
assign LUT_3[29008] = 32'b00000000000000001110110000101100;
assign LUT_3[29009] = 32'b00000000000000010101011100001001;
assign LUT_3[29010] = 32'b00000000000000010000111000010000;
assign LUT_3[29011] = 32'b00000000000000010111100011101101;
assign LUT_3[29012] = 32'b00000000000000001011111110100010;
assign LUT_3[29013] = 32'b00000000000000010010101001111111;
assign LUT_3[29014] = 32'b00000000000000001110000110000110;
assign LUT_3[29015] = 32'b00000000000000010100110001100011;
assign LUT_3[29016] = 32'b00000000000000010100001001110010;
assign LUT_3[29017] = 32'b00000000000000011010110101001111;
assign LUT_3[29018] = 32'b00000000000000010110010001010110;
assign LUT_3[29019] = 32'b00000000000000011100111100110011;
assign LUT_3[29020] = 32'b00000000000000010001010111101000;
assign LUT_3[29021] = 32'b00000000000000011000000011000101;
assign LUT_3[29022] = 32'b00000000000000010011011111001100;
assign LUT_3[29023] = 32'b00000000000000011010001010101001;
assign LUT_3[29024] = 32'b00000000000000001100101100001001;
assign LUT_3[29025] = 32'b00000000000000010011010111100110;
assign LUT_3[29026] = 32'b00000000000000001110110011101101;
assign LUT_3[29027] = 32'b00000000000000010101011111001010;
assign LUT_3[29028] = 32'b00000000000000001001111001111111;
assign LUT_3[29029] = 32'b00000000000000010000100101011100;
assign LUT_3[29030] = 32'b00000000000000001100000001100011;
assign LUT_3[29031] = 32'b00000000000000010010101101000000;
assign LUT_3[29032] = 32'b00000000000000010010000101001111;
assign LUT_3[29033] = 32'b00000000000000011000110000101100;
assign LUT_3[29034] = 32'b00000000000000010100001100110011;
assign LUT_3[29035] = 32'b00000000000000011010111000010000;
assign LUT_3[29036] = 32'b00000000000000001111010011000101;
assign LUT_3[29037] = 32'b00000000000000010101111110100010;
assign LUT_3[29038] = 32'b00000000000000010001011010101001;
assign LUT_3[29039] = 32'b00000000000000011000000110000110;
assign LUT_3[29040] = 32'b00000000000000001111111111001100;
assign LUT_3[29041] = 32'b00000000000000010110101010101001;
assign LUT_3[29042] = 32'b00000000000000010010000110110000;
assign LUT_3[29043] = 32'b00000000000000011000110010001101;
assign LUT_3[29044] = 32'b00000000000000001101001101000010;
assign LUT_3[29045] = 32'b00000000000000010011111000011111;
assign LUT_3[29046] = 32'b00000000000000001111010100100110;
assign LUT_3[29047] = 32'b00000000000000010110000000000011;
assign LUT_3[29048] = 32'b00000000000000010101011000010010;
assign LUT_3[29049] = 32'b00000000000000011100000011101111;
assign LUT_3[29050] = 32'b00000000000000010111011111110110;
assign LUT_3[29051] = 32'b00000000000000011110001011010011;
assign LUT_3[29052] = 32'b00000000000000010010100110001000;
assign LUT_3[29053] = 32'b00000000000000011001010001100101;
assign LUT_3[29054] = 32'b00000000000000010100101101101100;
assign LUT_3[29055] = 32'b00000000000000011011011001001001;
assign LUT_3[29056] = 32'b00000000000000001101101111111100;
assign LUT_3[29057] = 32'b00000000000000010100011011011001;
assign LUT_3[29058] = 32'b00000000000000001111110111100000;
assign LUT_3[29059] = 32'b00000000000000010110100010111101;
assign LUT_3[29060] = 32'b00000000000000001010111101110010;
assign LUT_3[29061] = 32'b00000000000000010001101001001111;
assign LUT_3[29062] = 32'b00000000000000001101000101010110;
assign LUT_3[29063] = 32'b00000000000000010011110000110011;
assign LUT_3[29064] = 32'b00000000000000010011001001000010;
assign LUT_3[29065] = 32'b00000000000000011001110100011111;
assign LUT_3[29066] = 32'b00000000000000010101010000100110;
assign LUT_3[29067] = 32'b00000000000000011011111100000011;
assign LUT_3[29068] = 32'b00000000000000010000010110111000;
assign LUT_3[29069] = 32'b00000000000000010111000010010101;
assign LUT_3[29070] = 32'b00000000000000010010011110011100;
assign LUT_3[29071] = 32'b00000000000000011001001001111001;
assign LUT_3[29072] = 32'b00000000000000010001000010111111;
assign LUT_3[29073] = 32'b00000000000000010111101110011100;
assign LUT_3[29074] = 32'b00000000000000010011001010100011;
assign LUT_3[29075] = 32'b00000000000000011001110110000000;
assign LUT_3[29076] = 32'b00000000000000001110010000110101;
assign LUT_3[29077] = 32'b00000000000000010100111100010010;
assign LUT_3[29078] = 32'b00000000000000010000011000011001;
assign LUT_3[29079] = 32'b00000000000000010111000011110110;
assign LUT_3[29080] = 32'b00000000000000010110011100000101;
assign LUT_3[29081] = 32'b00000000000000011101000111100010;
assign LUT_3[29082] = 32'b00000000000000011000100011101001;
assign LUT_3[29083] = 32'b00000000000000011111001111000110;
assign LUT_3[29084] = 32'b00000000000000010011101001111011;
assign LUT_3[29085] = 32'b00000000000000011010010101011000;
assign LUT_3[29086] = 32'b00000000000000010101110001011111;
assign LUT_3[29087] = 32'b00000000000000011100011100111100;
assign LUT_3[29088] = 32'b00000000000000001110111110011100;
assign LUT_3[29089] = 32'b00000000000000010101101001111001;
assign LUT_3[29090] = 32'b00000000000000010001000110000000;
assign LUT_3[29091] = 32'b00000000000000010111110001011101;
assign LUT_3[29092] = 32'b00000000000000001100001100010010;
assign LUT_3[29093] = 32'b00000000000000010010110111101111;
assign LUT_3[29094] = 32'b00000000000000001110010011110110;
assign LUT_3[29095] = 32'b00000000000000010100111111010011;
assign LUT_3[29096] = 32'b00000000000000010100010111100010;
assign LUT_3[29097] = 32'b00000000000000011011000010111111;
assign LUT_3[29098] = 32'b00000000000000010110011111000110;
assign LUT_3[29099] = 32'b00000000000000011101001010100011;
assign LUT_3[29100] = 32'b00000000000000010001100101011000;
assign LUT_3[29101] = 32'b00000000000000011000010000110101;
assign LUT_3[29102] = 32'b00000000000000010011101100111100;
assign LUT_3[29103] = 32'b00000000000000011010011000011001;
assign LUT_3[29104] = 32'b00000000000000010010010001011111;
assign LUT_3[29105] = 32'b00000000000000011000111100111100;
assign LUT_3[29106] = 32'b00000000000000010100011001000011;
assign LUT_3[29107] = 32'b00000000000000011011000100100000;
assign LUT_3[29108] = 32'b00000000000000001111011111010101;
assign LUT_3[29109] = 32'b00000000000000010110001010110010;
assign LUT_3[29110] = 32'b00000000000000010001100110111001;
assign LUT_3[29111] = 32'b00000000000000011000010010010110;
assign LUT_3[29112] = 32'b00000000000000010111101010100101;
assign LUT_3[29113] = 32'b00000000000000011110010110000010;
assign LUT_3[29114] = 32'b00000000000000011001110010001001;
assign LUT_3[29115] = 32'b00000000000000100000011101100110;
assign LUT_3[29116] = 32'b00000000000000010100111000011011;
assign LUT_3[29117] = 32'b00000000000000011011100011111000;
assign LUT_3[29118] = 32'b00000000000000010110111111111111;
assign LUT_3[29119] = 32'b00000000000000011101101011011100;
assign LUT_3[29120] = 32'b00000000000000001101101000100111;
assign LUT_3[29121] = 32'b00000000000000010100010100000100;
assign LUT_3[29122] = 32'b00000000000000001111110000001011;
assign LUT_3[29123] = 32'b00000000000000010110011011101000;
assign LUT_3[29124] = 32'b00000000000000001010110110011101;
assign LUT_3[29125] = 32'b00000000000000010001100001111010;
assign LUT_3[29126] = 32'b00000000000000001100111110000001;
assign LUT_3[29127] = 32'b00000000000000010011101001011110;
assign LUT_3[29128] = 32'b00000000000000010011000001101101;
assign LUT_3[29129] = 32'b00000000000000011001101101001010;
assign LUT_3[29130] = 32'b00000000000000010101001001010001;
assign LUT_3[29131] = 32'b00000000000000011011110100101110;
assign LUT_3[29132] = 32'b00000000000000010000001111100011;
assign LUT_3[29133] = 32'b00000000000000010110111011000000;
assign LUT_3[29134] = 32'b00000000000000010010010111000111;
assign LUT_3[29135] = 32'b00000000000000011001000010100100;
assign LUT_3[29136] = 32'b00000000000000010000111011101010;
assign LUT_3[29137] = 32'b00000000000000010111100111000111;
assign LUT_3[29138] = 32'b00000000000000010011000011001110;
assign LUT_3[29139] = 32'b00000000000000011001101110101011;
assign LUT_3[29140] = 32'b00000000000000001110001001100000;
assign LUT_3[29141] = 32'b00000000000000010100110100111101;
assign LUT_3[29142] = 32'b00000000000000010000010001000100;
assign LUT_3[29143] = 32'b00000000000000010110111100100001;
assign LUT_3[29144] = 32'b00000000000000010110010100110000;
assign LUT_3[29145] = 32'b00000000000000011101000000001101;
assign LUT_3[29146] = 32'b00000000000000011000011100010100;
assign LUT_3[29147] = 32'b00000000000000011111000111110001;
assign LUT_3[29148] = 32'b00000000000000010011100010100110;
assign LUT_3[29149] = 32'b00000000000000011010001110000011;
assign LUT_3[29150] = 32'b00000000000000010101101010001010;
assign LUT_3[29151] = 32'b00000000000000011100010101100111;
assign LUT_3[29152] = 32'b00000000000000001110110111000111;
assign LUT_3[29153] = 32'b00000000000000010101100010100100;
assign LUT_3[29154] = 32'b00000000000000010000111110101011;
assign LUT_3[29155] = 32'b00000000000000010111101010001000;
assign LUT_3[29156] = 32'b00000000000000001100000100111101;
assign LUT_3[29157] = 32'b00000000000000010010110000011010;
assign LUT_3[29158] = 32'b00000000000000001110001100100001;
assign LUT_3[29159] = 32'b00000000000000010100110111111110;
assign LUT_3[29160] = 32'b00000000000000010100010000001101;
assign LUT_3[29161] = 32'b00000000000000011010111011101010;
assign LUT_3[29162] = 32'b00000000000000010110010111110001;
assign LUT_3[29163] = 32'b00000000000000011101000011001110;
assign LUT_3[29164] = 32'b00000000000000010001011110000011;
assign LUT_3[29165] = 32'b00000000000000011000001001100000;
assign LUT_3[29166] = 32'b00000000000000010011100101100111;
assign LUT_3[29167] = 32'b00000000000000011010010001000100;
assign LUT_3[29168] = 32'b00000000000000010010001010001010;
assign LUT_3[29169] = 32'b00000000000000011000110101100111;
assign LUT_3[29170] = 32'b00000000000000010100010001101110;
assign LUT_3[29171] = 32'b00000000000000011010111101001011;
assign LUT_3[29172] = 32'b00000000000000001111011000000000;
assign LUT_3[29173] = 32'b00000000000000010110000011011101;
assign LUT_3[29174] = 32'b00000000000000010001011111100100;
assign LUT_3[29175] = 32'b00000000000000011000001011000001;
assign LUT_3[29176] = 32'b00000000000000010111100011010000;
assign LUT_3[29177] = 32'b00000000000000011110001110101101;
assign LUT_3[29178] = 32'b00000000000000011001101010110100;
assign LUT_3[29179] = 32'b00000000000000100000010110010001;
assign LUT_3[29180] = 32'b00000000000000010100110001000110;
assign LUT_3[29181] = 32'b00000000000000011011011100100011;
assign LUT_3[29182] = 32'b00000000000000010110111000101010;
assign LUT_3[29183] = 32'b00000000000000011101100100000111;
assign LUT_3[29184] = 32'b00000000000000010010101010101001;
assign LUT_3[29185] = 32'b00000000000000011001010110000110;
assign LUT_3[29186] = 32'b00000000000000010100110010001101;
assign LUT_3[29187] = 32'b00000000000000011011011101101010;
assign LUT_3[29188] = 32'b00000000000000001111111000011111;
assign LUT_3[29189] = 32'b00000000000000010110100011111100;
assign LUT_3[29190] = 32'b00000000000000010010000000000011;
assign LUT_3[29191] = 32'b00000000000000011000101011100000;
assign LUT_3[29192] = 32'b00000000000000011000000011101111;
assign LUT_3[29193] = 32'b00000000000000011110101111001100;
assign LUT_3[29194] = 32'b00000000000000011010001011010011;
assign LUT_3[29195] = 32'b00000000000000100000110110110000;
assign LUT_3[29196] = 32'b00000000000000010101010001100101;
assign LUT_3[29197] = 32'b00000000000000011011111101000010;
assign LUT_3[29198] = 32'b00000000000000010111011001001001;
assign LUT_3[29199] = 32'b00000000000000011110000100100110;
assign LUT_3[29200] = 32'b00000000000000010101111101101100;
assign LUT_3[29201] = 32'b00000000000000011100101001001001;
assign LUT_3[29202] = 32'b00000000000000011000000101010000;
assign LUT_3[29203] = 32'b00000000000000011110110000101101;
assign LUT_3[29204] = 32'b00000000000000010011001011100010;
assign LUT_3[29205] = 32'b00000000000000011001110110111111;
assign LUT_3[29206] = 32'b00000000000000010101010011000110;
assign LUT_3[29207] = 32'b00000000000000011011111110100011;
assign LUT_3[29208] = 32'b00000000000000011011010110110010;
assign LUT_3[29209] = 32'b00000000000000100010000010001111;
assign LUT_3[29210] = 32'b00000000000000011101011110010110;
assign LUT_3[29211] = 32'b00000000000000100100001001110011;
assign LUT_3[29212] = 32'b00000000000000011000100100101000;
assign LUT_3[29213] = 32'b00000000000000011111010000000101;
assign LUT_3[29214] = 32'b00000000000000011010101100001100;
assign LUT_3[29215] = 32'b00000000000000100001010111101001;
assign LUT_3[29216] = 32'b00000000000000010011111001001001;
assign LUT_3[29217] = 32'b00000000000000011010100100100110;
assign LUT_3[29218] = 32'b00000000000000010110000000101101;
assign LUT_3[29219] = 32'b00000000000000011100101100001010;
assign LUT_3[29220] = 32'b00000000000000010001000110111111;
assign LUT_3[29221] = 32'b00000000000000010111110010011100;
assign LUT_3[29222] = 32'b00000000000000010011001110100011;
assign LUT_3[29223] = 32'b00000000000000011001111010000000;
assign LUT_3[29224] = 32'b00000000000000011001010010001111;
assign LUT_3[29225] = 32'b00000000000000011111111101101100;
assign LUT_3[29226] = 32'b00000000000000011011011001110011;
assign LUT_3[29227] = 32'b00000000000000100010000101010000;
assign LUT_3[29228] = 32'b00000000000000010110100000000101;
assign LUT_3[29229] = 32'b00000000000000011101001011100010;
assign LUT_3[29230] = 32'b00000000000000011000100111101001;
assign LUT_3[29231] = 32'b00000000000000011111010011000110;
assign LUT_3[29232] = 32'b00000000000000010111001100001100;
assign LUT_3[29233] = 32'b00000000000000011101110111101001;
assign LUT_3[29234] = 32'b00000000000000011001010011110000;
assign LUT_3[29235] = 32'b00000000000000011111111111001101;
assign LUT_3[29236] = 32'b00000000000000010100011010000010;
assign LUT_3[29237] = 32'b00000000000000011011000101011111;
assign LUT_3[29238] = 32'b00000000000000010110100001100110;
assign LUT_3[29239] = 32'b00000000000000011101001101000011;
assign LUT_3[29240] = 32'b00000000000000011100100101010010;
assign LUT_3[29241] = 32'b00000000000000100011010000101111;
assign LUT_3[29242] = 32'b00000000000000011110101100110110;
assign LUT_3[29243] = 32'b00000000000000100101011000010011;
assign LUT_3[29244] = 32'b00000000000000011001110011001000;
assign LUT_3[29245] = 32'b00000000000000100000011110100101;
assign LUT_3[29246] = 32'b00000000000000011011111010101100;
assign LUT_3[29247] = 32'b00000000000000100010100110001001;
assign LUT_3[29248] = 32'b00000000000000010010100011010100;
assign LUT_3[29249] = 32'b00000000000000011001001110110001;
assign LUT_3[29250] = 32'b00000000000000010100101010111000;
assign LUT_3[29251] = 32'b00000000000000011011010110010101;
assign LUT_3[29252] = 32'b00000000000000001111110001001010;
assign LUT_3[29253] = 32'b00000000000000010110011100100111;
assign LUT_3[29254] = 32'b00000000000000010001111000101110;
assign LUT_3[29255] = 32'b00000000000000011000100100001011;
assign LUT_3[29256] = 32'b00000000000000010111111100011010;
assign LUT_3[29257] = 32'b00000000000000011110100111110111;
assign LUT_3[29258] = 32'b00000000000000011010000011111110;
assign LUT_3[29259] = 32'b00000000000000100000101111011011;
assign LUT_3[29260] = 32'b00000000000000010101001010010000;
assign LUT_3[29261] = 32'b00000000000000011011110101101101;
assign LUT_3[29262] = 32'b00000000000000010111010001110100;
assign LUT_3[29263] = 32'b00000000000000011101111101010001;
assign LUT_3[29264] = 32'b00000000000000010101110110010111;
assign LUT_3[29265] = 32'b00000000000000011100100001110100;
assign LUT_3[29266] = 32'b00000000000000010111111101111011;
assign LUT_3[29267] = 32'b00000000000000011110101001011000;
assign LUT_3[29268] = 32'b00000000000000010011000100001101;
assign LUT_3[29269] = 32'b00000000000000011001101111101010;
assign LUT_3[29270] = 32'b00000000000000010101001011110001;
assign LUT_3[29271] = 32'b00000000000000011011110111001110;
assign LUT_3[29272] = 32'b00000000000000011011001111011101;
assign LUT_3[29273] = 32'b00000000000000100001111010111010;
assign LUT_3[29274] = 32'b00000000000000011101010111000001;
assign LUT_3[29275] = 32'b00000000000000100100000010011110;
assign LUT_3[29276] = 32'b00000000000000011000011101010011;
assign LUT_3[29277] = 32'b00000000000000011111001000110000;
assign LUT_3[29278] = 32'b00000000000000011010100100110111;
assign LUT_3[29279] = 32'b00000000000000100001010000010100;
assign LUT_3[29280] = 32'b00000000000000010011110001110100;
assign LUT_3[29281] = 32'b00000000000000011010011101010001;
assign LUT_3[29282] = 32'b00000000000000010101111001011000;
assign LUT_3[29283] = 32'b00000000000000011100100100110101;
assign LUT_3[29284] = 32'b00000000000000010000111111101010;
assign LUT_3[29285] = 32'b00000000000000010111101011000111;
assign LUT_3[29286] = 32'b00000000000000010011000111001110;
assign LUT_3[29287] = 32'b00000000000000011001110010101011;
assign LUT_3[29288] = 32'b00000000000000011001001010111010;
assign LUT_3[29289] = 32'b00000000000000011111110110010111;
assign LUT_3[29290] = 32'b00000000000000011011010010011110;
assign LUT_3[29291] = 32'b00000000000000100001111101111011;
assign LUT_3[29292] = 32'b00000000000000010110011000110000;
assign LUT_3[29293] = 32'b00000000000000011101000100001101;
assign LUT_3[29294] = 32'b00000000000000011000100000010100;
assign LUT_3[29295] = 32'b00000000000000011111001011110001;
assign LUT_3[29296] = 32'b00000000000000010111000100110111;
assign LUT_3[29297] = 32'b00000000000000011101110000010100;
assign LUT_3[29298] = 32'b00000000000000011001001100011011;
assign LUT_3[29299] = 32'b00000000000000011111110111111000;
assign LUT_3[29300] = 32'b00000000000000010100010010101101;
assign LUT_3[29301] = 32'b00000000000000011010111110001010;
assign LUT_3[29302] = 32'b00000000000000010110011010010001;
assign LUT_3[29303] = 32'b00000000000000011101000101101110;
assign LUT_3[29304] = 32'b00000000000000011100011101111101;
assign LUT_3[29305] = 32'b00000000000000100011001001011010;
assign LUT_3[29306] = 32'b00000000000000011110100101100001;
assign LUT_3[29307] = 32'b00000000000000100101010000111110;
assign LUT_3[29308] = 32'b00000000000000011001101011110011;
assign LUT_3[29309] = 32'b00000000000000100000010111010000;
assign LUT_3[29310] = 32'b00000000000000011011110011010111;
assign LUT_3[29311] = 32'b00000000000000100010011110110100;
assign LUT_3[29312] = 32'b00000000000000010100110101100111;
assign LUT_3[29313] = 32'b00000000000000011011100001000100;
assign LUT_3[29314] = 32'b00000000000000010110111101001011;
assign LUT_3[29315] = 32'b00000000000000011101101000101000;
assign LUT_3[29316] = 32'b00000000000000010010000011011101;
assign LUT_3[29317] = 32'b00000000000000011000101110111010;
assign LUT_3[29318] = 32'b00000000000000010100001011000001;
assign LUT_3[29319] = 32'b00000000000000011010110110011110;
assign LUT_3[29320] = 32'b00000000000000011010001110101101;
assign LUT_3[29321] = 32'b00000000000000100000111010001010;
assign LUT_3[29322] = 32'b00000000000000011100010110010001;
assign LUT_3[29323] = 32'b00000000000000100011000001101110;
assign LUT_3[29324] = 32'b00000000000000010111011100100011;
assign LUT_3[29325] = 32'b00000000000000011110001000000000;
assign LUT_3[29326] = 32'b00000000000000011001100100000111;
assign LUT_3[29327] = 32'b00000000000000100000001111100100;
assign LUT_3[29328] = 32'b00000000000000011000001000101010;
assign LUT_3[29329] = 32'b00000000000000011110110100000111;
assign LUT_3[29330] = 32'b00000000000000011010010000001110;
assign LUT_3[29331] = 32'b00000000000000100000111011101011;
assign LUT_3[29332] = 32'b00000000000000010101010110100000;
assign LUT_3[29333] = 32'b00000000000000011100000001111101;
assign LUT_3[29334] = 32'b00000000000000010111011110000100;
assign LUT_3[29335] = 32'b00000000000000011110001001100001;
assign LUT_3[29336] = 32'b00000000000000011101100001110000;
assign LUT_3[29337] = 32'b00000000000000100100001101001101;
assign LUT_3[29338] = 32'b00000000000000011111101001010100;
assign LUT_3[29339] = 32'b00000000000000100110010100110001;
assign LUT_3[29340] = 32'b00000000000000011010101111100110;
assign LUT_3[29341] = 32'b00000000000000100001011011000011;
assign LUT_3[29342] = 32'b00000000000000011100110111001010;
assign LUT_3[29343] = 32'b00000000000000100011100010100111;
assign LUT_3[29344] = 32'b00000000000000010110000100000111;
assign LUT_3[29345] = 32'b00000000000000011100101111100100;
assign LUT_3[29346] = 32'b00000000000000011000001011101011;
assign LUT_3[29347] = 32'b00000000000000011110110111001000;
assign LUT_3[29348] = 32'b00000000000000010011010001111101;
assign LUT_3[29349] = 32'b00000000000000011001111101011010;
assign LUT_3[29350] = 32'b00000000000000010101011001100001;
assign LUT_3[29351] = 32'b00000000000000011100000100111110;
assign LUT_3[29352] = 32'b00000000000000011011011101001101;
assign LUT_3[29353] = 32'b00000000000000100010001000101010;
assign LUT_3[29354] = 32'b00000000000000011101100100110001;
assign LUT_3[29355] = 32'b00000000000000100100010000001110;
assign LUT_3[29356] = 32'b00000000000000011000101011000011;
assign LUT_3[29357] = 32'b00000000000000011111010110100000;
assign LUT_3[29358] = 32'b00000000000000011010110010100111;
assign LUT_3[29359] = 32'b00000000000000100001011110000100;
assign LUT_3[29360] = 32'b00000000000000011001010111001010;
assign LUT_3[29361] = 32'b00000000000000100000000010100111;
assign LUT_3[29362] = 32'b00000000000000011011011110101110;
assign LUT_3[29363] = 32'b00000000000000100010001010001011;
assign LUT_3[29364] = 32'b00000000000000010110100101000000;
assign LUT_3[29365] = 32'b00000000000000011101010000011101;
assign LUT_3[29366] = 32'b00000000000000011000101100100100;
assign LUT_3[29367] = 32'b00000000000000011111011000000001;
assign LUT_3[29368] = 32'b00000000000000011110110000010000;
assign LUT_3[29369] = 32'b00000000000000100101011011101101;
assign LUT_3[29370] = 32'b00000000000000100000110111110100;
assign LUT_3[29371] = 32'b00000000000000100111100011010001;
assign LUT_3[29372] = 32'b00000000000000011011111110000110;
assign LUT_3[29373] = 32'b00000000000000100010101001100011;
assign LUT_3[29374] = 32'b00000000000000011110000101101010;
assign LUT_3[29375] = 32'b00000000000000100100110001000111;
assign LUT_3[29376] = 32'b00000000000000010100101110010010;
assign LUT_3[29377] = 32'b00000000000000011011011001101111;
assign LUT_3[29378] = 32'b00000000000000010110110101110110;
assign LUT_3[29379] = 32'b00000000000000011101100001010011;
assign LUT_3[29380] = 32'b00000000000000010001111100001000;
assign LUT_3[29381] = 32'b00000000000000011000100111100101;
assign LUT_3[29382] = 32'b00000000000000010100000011101100;
assign LUT_3[29383] = 32'b00000000000000011010101111001001;
assign LUT_3[29384] = 32'b00000000000000011010000111011000;
assign LUT_3[29385] = 32'b00000000000000100000110010110101;
assign LUT_3[29386] = 32'b00000000000000011100001110111100;
assign LUT_3[29387] = 32'b00000000000000100010111010011001;
assign LUT_3[29388] = 32'b00000000000000010111010101001110;
assign LUT_3[29389] = 32'b00000000000000011110000000101011;
assign LUT_3[29390] = 32'b00000000000000011001011100110010;
assign LUT_3[29391] = 32'b00000000000000100000001000001111;
assign LUT_3[29392] = 32'b00000000000000011000000001010101;
assign LUT_3[29393] = 32'b00000000000000011110101100110010;
assign LUT_3[29394] = 32'b00000000000000011010001000111001;
assign LUT_3[29395] = 32'b00000000000000100000110100010110;
assign LUT_3[29396] = 32'b00000000000000010101001111001011;
assign LUT_3[29397] = 32'b00000000000000011011111010101000;
assign LUT_3[29398] = 32'b00000000000000010111010110101111;
assign LUT_3[29399] = 32'b00000000000000011110000010001100;
assign LUT_3[29400] = 32'b00000000000000011101011010011011;
assign LUT_3[29401] = 32'b00000000000000100100000101111000;
assign LUT_3[29402] = 32'b00000000000000011111100001111111;
assign LUT_3[29403] = 32'b00000000000000100110001101011100;
assign LUT_3[29404] = 32'b00000000000000011010101000010001;
assign LUT_3[29405] = 32'b00000000000000100001010011101110;
assign LUT_3[29406] = 32'b00000000000000011100101111110101;
assign LUT_3[29407] = 32'b00000000000000100011011011010010;
assign LUT_3[29408] = 32'b00000000000000010101111100110010;
assign LUT_3[29409] = 32'b00000000000000011100101000001111;
assign LUT_3[29410] = 32'b00000000000000011000000100010110;
assign LUT_3[29411] = 32'b00000000000000011110101111110011;
assign LUT_3[29412] = 32'b00000000000000010011001010101000;
assign LUT_3[29413] = 32'b00000000000000011001110110000101;
assign LUT_3[29414] = 32'b00000000000000010101010010001100;
assign LUT_3[29415] = 32'b00000000000000011011111101101001;
assign LUT_3[29416] = 32'b00000000000000011011010101111000;
assign LUT_3[29417] = 32'b00000000000000100010000001010101;
assign LUT_3[29418] = 32'b00000000000000011101011101011100;
assign LUT_3[29419] = 32'b00000000000000100100001000111001;
assign LUT_3[29420] = 32'b00000000000000011000100011101110;
assign LUT_3[29421] = 32'b00000000000000011111001111001011;
assign LUT_3[29422] = 32'b00000000000000011010101011010010;
assign LUT_3[29423] = 32'b00000000000000100001010110101111;
assign LUT_3[29424] = 32'b00000000000000011001001111110101;
assign LUT_3[29425] = 32'b00000000000000011111111011010010;
assign LUT_3[29426] = 32'b00000000000000011011010111011001;
assign LUT_3[29427] = 32'b00000000000000100010000010110110;
assign LUT_3[29428] = 32'b00000000000000010110011101101011;
assign LUT_3[29429] = 32'b00000000000000011101001001001000;
assign LUT_3[29430] = 32'b00000000000000011000100101001111;
assign LUT_3[29431] = 32'b00000000000000011111010000101100;
assign LUT_3[29432] = 32'b00000000000000011110101000111011;
assign LUT_3[29433] = 32'b00000000000000100101010100011000;
assign LUT_3[29434] = 32'b00000000000000100000110000011111;
assign LUT_3[29435] = 32'b00000000000000100111011011111100;
assign LUT_3[29436] = 32'b00000000000000011011110110110001;
assign LUT_3[29437] = 32'b00000000000000100010100010001110;
assign LUT_3[29438] = 32'b00000000000000011101111110010101;
assign LUT_3[29439] = 32'b00000000000000100100101001110010;
assign LUT_3[29440] = 32'b00000000000000001110111010001010;
assign LUT_3[29441] = 32'b00000000000000010101100101100111;
assign LUT_3[29442] = 32'b00000000000000010001000001101110;
assign LUT_3[29443] = 32'b00000000000000010111101101001011;
assign LUT_3[29444] = 32'b00000000000000001100001000000000;
assign LUT_3[29445] = 32'b00000000000000010010110011011101;
assign LUT_3[29446] = 32'b00000000000000001110001111100100;
assign LUT_3[29447] = 32'b00000000000000010100111011000001;
assign LUT_3[29448] = 32'b00000000000000010100010011010000;
assign LUT_3[29449] = 32'b00000000000000011010111110101101;
assign LUT_3[29450] = 32'b00000000000000010110011010110100;
assign LUT_3[29451] = 32'b00000000000000011101000110010001;
assign LUT_3[29452] = 32'b00000000000000010001100001000110;
assign LUT_3[29453] = 32'b00000000000000011000001100100011;
assign LUT_3[29454] = 32'b00000000000000010011101000101010;
assign LUT_3[29455] = 32'b00000000000000011010010100000111;
assign LUT_3[29456] = 32'b00000000000000010010001101001101;
assign LUT_3[29457] = 32'b00000000000000011000111000101010;
assign LUT_3[29458] = 32'b00000000000000010100010100110001;
assign LUT_3[29459] = 32'b00000000000000011011000000001110;
assign LUT_3[29460] = 32'b00000000000000001111011011000011;
assign LUT_3[29461] = 32'b00000000000000010110000110100000;
assign LUT_3[29462] = 32'b00000000000000010001100010100111;
assign LUT_3[29463] = 32'b00000000000000011000001110000100;
assign LUT_3[29464] = 32'b00000000000000010111100110010011;
assign LUT_3[29465] = 32'b00000000000000011110010001110000;
assign LUT_3[29466] = 32'b00000000000000011001101101110111;
assign LUT_3[29467] = 32'b00000000000000100000011001010100;
assign LUT_3[29468] = 32'b00000000000000010100110100001001;
assign LUT_3[29469] = 32'b00000000000000011011011111100110;
assign LUT_3[29470] = 32'b00000000000000010110111011101101;
assign LUT_3[29471] = 32'b00000000000000011101100111001010;
assign LUT_3[29472] = 32'b00000000000000010000001000101010;
assign LUT_3[29473] = 32'b00000000000000010110110100000111;
assign LUT_3[29474] = 32'b00000000000000010010010000001110;
assign LUT_3[29475] = 32'b00000000000000011000111011101011;
assign LUT_3[29476] = 32'b00000000000000001101010110100000;
assign LUT_3[29477] = 32'b00000000000000010100000001111101;
assign LUT_3[29478] = 32'b00000000000000001111011110000100;
assign LUT_3[29479] = 32'b00000000000000010110001001100001;
assign LUT_3[29480] = 32'b00000000000000010101100001110000;
assign LUT_3[29481] = 32'b00000000000000011100001101001101;
assign LUT_3[29482] = 32'b00000000000000010111101001010100;
assign LUT_3[29483] = 32'b00000000000000011110010100110001;
assign LUT_3[29484] = 32'b00000000000000010010101111100110;
assign LUT_3[29485] = 32'b00000000000000011001011011000011;
assign LUT_3[29486] = 32'b00000000000000010100110111001010;
assign LUT_3[29487] = 32'b00000000000000011011100010100111;
assign LUT_3[29488] = 32'b00000000000000010011011011101101;
assign LUT_3[29489] = 32'b00000000000000011010000111001010;
assign LUT_3[29490] = 32'b00000000000000010101100011010001;
assign LUT_3[29491] = 32'b00000000000000011100001110101110;
assign LUT_3[29492] = 32'b00000000000000010000101001100011;
assign LUT_3[29493] = 32'b00000000000000010111010101000000;
assign LUT_3[29494] = 32'b00000000000000010010110001000111;
assign LUT_3[29495] = 32'b00000000000000011001011100100100;
assign LUT_3[29496] = 32'b00000000000000011000110100110011;
assign LUT_3[29497] = 32'b00000000000000011111100000010000;
assign LUT_3[29498] = 32'b00000000000000011010111100010111;
assign LUT_3[29499] = 32'b00000000000000100001100111110100;
assign LUT_3[29500] = 32'b00000000000000010110000010101001;
assign LUT_3[29501] = 32'b00000000000000011100101110000110;
assign LUT_3[29502] = 32'b00000000000000011000001010001101;
assign LUT_3[29503] = 32'b00000000000000011110110101101010;
assign LUT_3[29504] = 32'b00000000000000001110110010110101;
assign LUT_3[29505] = 32'b00000000000000010101011110010010;
assign LUT_3[29506] = 32'b00000000000000010000111010011001;
assign LUT_3[29507] = 32'b00000000000000010111100101110110;
assign LUT_3[29508] = 32'b00000000000000001100000000101011;
assign LUT_3[29509] = 32'b00000000000000010010101100001000;
assign LUT_3[29510] = 32'b00000000000000001110001000001111;
assign LUT_3[29511] = 32'b00000000000000010100110011101100;
assign LUT_3[29512] = 32'b00000000000000010100001011111011;
assign LUT_3[29513] = 32'b00000000000000011010110111011000;
assign LUT_3[29514] = 32'b00000000000000010110010011011111;
assign LUT_3[29515] = 32'b00000000000000011100111110111100;
assign LUT_3[29516] = 32'b00000000000000010001011001110001;
assign LUT_3[29517] = 32'b00000000000000011000000101001110;
assign LUT_3[29518] = 32'b00000000000000010011100001010101;
assign LUT_3[29519] = 32'b00000000000000011010001100110010;
assign LUT_3[29520] = 32'b00000000000000010010000101111000;
assign LUT_3[29521] = 32'b00000000000000011000110001010101;
assign LUT_3[29522] = 32'b00000000000000010100001101011100;
assign LUT_3[29523] = 32'b00000000000000011010111000111001;
assign LUT_3[29524] = 32'b00000000000000001111010011101110;
assign LUT_3[29525] = 32'b00000000000000010101111111001011;
assign LUT_3[29526] = 32'b00000000000000010001011011010010;
assign LUT_3[29527] = 32'b00000000000000011000000110101111;
assign LUT_3[29528] = 32'b00000000000000010111011110111110;
assign LUT_3[29529] = 32'b00000000000000011110001010011011;
assign LUT_3[29530] = 32'b00000000000000011001100110100010;
assign LUT_3[29531] = 32'b00000000000000100000010001111111;
assign LUT_3[29532] = 32'b00000000000000010100101100110100;
assign LUT_3[29533] = 32'b00000000000000011011011000010001;
assign LUT_3[29534] = 32'b00000000000000010110110100011000;
assign LUT_3[29535] = 32'b00000000000000011101011111110101;
assign LUT_3[29536] = 32'b00000000000000010000000001010101;
assign LUT_3[29537] = 32'b00000000000000010110101100110010;
assign LUT_3[29538] = 32'b00000000000000010010001000111001;
assign LUT_3[29539] = 32'b00000000000000011000110100010110;
assign LUT_3[29540] = 32'b00000000000000001101001111001011;
assign LUT_3[29541] = 32'b00000000000000010011111010101000;
assign LUT_3[29542] = 32'b00000000000000001111010110101111;
assign LUT_3[29543] = 32'b00000000000000010110000010001100;
assign LUT_3[29544] = 32'b00000000000000010101011010011011;
assign LUT_3[29545] = 32'b00000000000000011100000101111000;
assign LUT_3[29546] = 32'b00000000000000010111100001111111;
assign LUT_3[29547] = 32'b00000000000000011110001101011100;
assign LUT_3[29548] = 32'b00000000000000010010101000010001;
assign LUT_3[29549] = 32'b00000000000000011001010011101110;
assign LUT_3[29550] = 32'b00000000000000010100101111110101;
assign LUT_3[29551] = 32'b00000000000000011011011011010010;
assign LUT_3[29552] = 32'b00000000000000010011010100011000;
assign LUT_3[29553] = 32'b00000000000000011001111111110101;
assign LUT_3[29554] = 32'b00000000000000010101011011111100;
assign LUT_3[29555] = 32'b00000000000000011100000111011001;
assign LUT_3[29556] = 32'b00000000000000010000100010001110;
assign LUT_3[29557] = 32'b00000000000000010111001101101011;
assign LUT_3[29558] = 32'b00000000000000010010101001110010;
assign LUT_3[29559] = 32'b00000000000000011001010101001111;
assign LUT_3[29560] = 32'b00000000000000011000101101011110;
assign LUT_3[29561] = 32'b00000000000000011111011000111011;
assign LUT_3[29562] = 32'b00000000000000011010110101000010;
assign LUT_3[29563] = 32'b00000000000000100001100000011111;
assign LUT_3[29564] = 32'b00000000000000010101111011010100;
assign LUT_3[29565] = 32'b00000000000000011100100110110001;
assign LUT_3[29566] = 32'b00000000000000011000000010111000;
assign LUT_3[29567] = 32'b00000000000000011110101110010101;
assign LUT_3[29568] = 32'b00000000000000010001000101001000;
assign LUT_3[29569] = 32'b00000000000000010111110000100101;
assign LUT_3[29570] = 32'b00000000000000010011001100101100;
assign LUT_3[29571] = 32'b00000000000000011001111000001001;
assign LUT_3[29572] = 32'b00000000000000001110010010111110;
assign LUT_3[29573] = 32'b00000000000000010100111110011011;
assign LUT_3[29574] = 32'b00000000000000010000011010100010;
assign LUT_3[29575] = 32'b00000000000000010111000101111111;
assign LUT_3[29576] = 32'b00000000000000010110011110001110;
assign LUT_3[29577] = 32'b00000000000000011101001001101011;
assign LUT_3[29578] = 32'b00000000000000011000100101110010;
assign LUT_3[29579] = 32'b00000000000000011111010001001111;
assign LUT_3[29580] = 32'b00000000000000010011101100000100;
assign LUT_3[29581] = 32'b00000000000000011010010111100001;
assign LUT_3[29582] = 32'b00000000000000010101110011101000;
assign LUT_3[29583] = 32'b00000000000000011100011111000101;
assign LUT_3[29584] = 32'b00000000000000010100011000001011;
assign LUT_3[29585] = 32'b00000000000000011011000011101000;
assign LUT_3[29586] = 32'b00000000000000010110011111101111;
assign LUT_3[29587] = 32'b00000000000000011101001011001100;
assign LUT_3[29588] = 32'b00000000000000010001100110000001;
assign LUT_3[29589] = 32'b00000000000000011000010001011110;
assign LUT_3[29590] = 32'b00000000000000010011101101100101;
assign LUT_3[29591] = 32'b00000000000000011010011001000010;
assign LUT_3[29592] = 32'b00000000000000011001110001010001;
assign LUT_3[29593] = 32'b00000000000000100000011100101110;
assign LUT_3[29594] = 32'b00000000000000011011111000110101;
assign LUT_3[29595] = 32'b00000000000000100010100100010010;
assign LUT_3[29596] = 32'b00000000000000010110111111000111;
assign LUT_3[29597] = 32'b00000000000000011101101010100100;
assign LUT_3[29598] = 32'b00000000000000011001000110101011;
assign LUT_3[29599] = 32'b00000000000000011111110010001000;
assign LUT_3[29600] = 32'b00000000000000010010010011101000;
assign LUT_3[29601] = 32'b00000000000000011000111111000101;
assign LUT_3[29602] = 32'b00000000000000010100011011001100;
assign LUT_3[29603] = 32'b00000000000000011011000110101001;
assign LUT_3[29604] = 32'b00000000000000001111100001011110;
assign LUT_3[29605] = 32'b00000000000000010110001100111011;
assign LUT_3[29606] = 32'b00000000000000010001101001000010;
assign LUT_3[29607] = 32'b00000000000000011000010100011111;
assign LUT_3[29608] = 32'b00000000000000010111101100101110;
assign LUT_3[29609] = 32'b00000000000000011110011000001011;
assign LUT_3[29610] = 32'b00000000000000011001110100010010;
assign LUT_3[29611] = 32'b00000000000000100000011111101111;
assign LUT_3[29612] = 32'b00000000000000010100111010100100;
assign LUT_3[29613] = 32'b00000000000000011011100110000001;
assign LUT_3[29614] = 32'b00000000000000010111000010001000;
assign LUT_3[29615] = 32'b00000000000000011101101101100101;
assign LUT_3[29616] = 32'b00000000000000010101100110101011;
assign LUT_3[29617] = 32'b00000000000000011100010010001000;
assign LUT_3[29618] = 32'b00000000000000010111101110001111;
assign LUT_3[29619] = 32'b00000000000000011110011001101100;
assign LUT_3[29620] = 32'b00000000000000010010110100100001;
assign LUT_3[29621] = 32'b00000000000000011001011111111110;
assign LUT_3[29622] = 32'b00000000000000010100111100000101;
assign LUT_3[29623] = 32'b00000000000000011011100111100010;
assign LUT_3[29624] = 32'b00000000000000011010111111110001;
assign LUT_3[29625] = 32'b00000000000000100001101011001110;
assign LUT_3[29626] = 32'b00000000000000011101000111010101;
assign LUT_3[29627] = 32'b00000000000000100011110010110010;
assign LUT_3[29628] = 32'b00000000000000011000001101100111;
assign LUT_3[29629] = 32'b00000000000000011110111001000100;
assign LUT_3[29630] = 32'b00000000000000011010010101001011;
assign LUT_3[29631] = 32'b00000000000000100001000000101000;
assign LUT_3[29632] = 32'b00000000000000010000111101110011;
assign LUT_3[29633] = 32'b00000000000000010111101001010000;
assign LUT_3[29634] = 32'b00000000000000010011000101010111;
assign LUT_3[29635] = 32'b00000000000000011001110000110100;
assign LUT_3[29636] = 32'b00000000000000001110001011101001;
assign LUT_3[29637] = 32'b00000000000000010100110111000110;
assign LUT_3[29638] = 32'b00000000000000010000010011001101;
assign LUT_3[29639] = 32'b00000000000000010110111110101010;
assign LUT_3[29640] = 32'b00000000000000010110010110111001;
assign LUT_3[29641] = 32'b00000000000000011101000010010110;
assign LUT_3[29642] = 32'b00000000000000011000011110011101;
assign LUT_3[29643] = 32'b00000000000000011111001001111010;
assign LUT_3[29644] = 32'b00000000000000010011100100101111;
assign LUT_3[29645] = 32'b00000000000000011010010000001100;
assign LUT_3[29646] = 32'b00000000000000010101101100010011;
assign LUT_3[29647] = 32'b00000000000000011100010111110000;
assign LUT_3[29648] = 32'b00000000000000010100010000110110;
assign LUT_3[29649] = 32'b00000000000000011010111100010011;
assign LUT_3[29650] = 32'b00000000000000010110011000011010;
assign LUT_3[29651] = 32'b00000000000000011101000011110111;
assign LUT_3[29652] = 32'b00000000000000010001011110101100;
assign LUT_3[29653] = 32'b00000000000000011000001010001001;
assign LUT_3[29654] = 32'b00000000000000010011100110010000;
assign LUT_3[29655] = 32'b00000000000000011010010001101101;
assign LUT_3[29656] = 32'b00000000000000011001101001111100;
assign LUT_3[29657] = 32'b00000000000000100000010101011001;
assign LUT_3[29658] = 32'b00000000000000011011110001100000;
assign LUT_3[29659] = 32'b00000000000000100010011100111101;
assign LUT_3[29660] = 32'b00000000000000010110110111110010;
assign LUT_3[29661] = 32'b00000000000000011101100011001111;
assign LUT_3[29662] = 32'b00000000000000011000111111010110;
assign LUT_3[29663] = 32'b00000000000000011111101010110011;
assign LUT_3[29664] = 32'b00000000000000010010001100010011;
assign LUT_3[29665] = 32'b00000000000000011000110111110000;
assign LUT_3[29666] = 32'b00000000000000010100010011110111;
assign LUT_3[29667] = 32'b00000000000000011010111111010100;
assign LUT_3[29668] = 32'b00000000000000001111011010001001;
assign LUT_3[29669] = 32'b00000000000000010110000101100110;
assign LUT_3[29670] = 32'b00000000000000010001100001101101;
assign LUT_3[29671] = 32'b00000000000000011000001101001010;
assign LUT_3[29672] = 32'b00000000000000010111100101011001;
assign LUT_3[29673] = 32'b00000000000000011110010000110110;
assign LUT_3[29674] = 32'b00000000000000011001101100111101;
assign LUT_3[29675] = 32'b00000000000000100000011000011010;
assign LUT_3[29676] = 32'b00000000000000010100110011001111;
assign LUT_3[29677] = 32'b00000000000000011011011110101100;
assign LUT_3[29678] = 32'b00000000000000010110111010110011;
assign LUT_3[29679] = 32'b00000000000000011101100110010000;
assign LUT_3[29680] = 32'b00000000000000010101011111010110;
assign LUT_3[29681] = 32'b00000000000000011100001010110011;
assign LUT_3[29682] = 32'b00000000000000010111100110111010;
assign LUT_3[29683] = 32'b00000000000000011110010010010111;
assign LUT_3[29684] = 32'b00000000000000010010101101001100;
assign LUT_3[29685] = 32'b00000000000000011001011000101001;
assign LUT_3[29686] = 32'b00000000000000010100110100110000;
assign LUT_3[29687] = 32'b00000000000000011011100000001101;
assign LUT_3[29688] = 32'b00000000000000011010111000011100;
assign LUT_3[29689] = 32'b00000000000000100001100011111001;
assign LUT_3[29690] = 32'b00000000000000011101000000000000;
assign LUT_3[29691] = 32'b00000000000000100011101011011101;
assign LUT_3[29692] = 32'b00000000000000011000000110010010;
assign LUT_3[29693] = 32'b00000000000000011110110001101111;
assign LUT_3[29694] = 32'b00000000000000011010001101110110;
assign LUT_3[29695] = 32'b00000000000000100000111001010011;
assign LUT_3[29696] = 32'b00000000000000010101111010011010;
assign LUT_3[29697] = 32'b00000000000000011100100101110111;
assign LUT_3[29698] = 32'b00000000000000011000000001111110;
assign LUT_3[29699] = 32'b00000000000000011110101101011011;
assign LUT_3[29700] = 32'b00000000000000010011001000010000;
assign LUT_3[29701] = 32'b00000000000000011001110011101101;
assign LUT_3[29702] = 32'b00000000000000010101001111110100;
assign LUT_3[29703] = 32'b00000000000000011011111011010001;
assign LUT_3[29704] = 32'b00000000000000011011010011100000;
assign LUT_3[29705] = 32'b00000000000000100001111110111101;
assign LUT_3[29706] = 32'b00000000000000011101011011000100;
assign LUT_3[29707] = 32'b00000000000000100100000110100001;
assign LUT_3[29708] = 32'b00000000000000011000100001010110;
assign LUT_3[29709] = 32'b00000000000000011111001100110011;
assign LUT_3[29710] = 32'b00000000000000011010101000111010;
assign LUT_3[29711] = 32'b00000000000000100001010100010111;
assign LUT_3[29712] = 32'b00000000000000011001001101011101;
assign LUT_3[29713] = 32'b00000000000000011111111000111010;
assign LUT_3[29714] = 32'b00000000000000011011010101000001;
assign LUT_3[29715] = 32'b00000000000000100010000000011110;
assign LUT_3[29716] = 32'b00000000000000010110011011010011;
assign LUT_3[29717] = 32'b00000000000000011101000110110000;
assign LUT_3[29718] = 32'b00000000000000011000100010110111;
assign LUT_3[29719] = 32'b00000000000000011111001110010100;
assign LUT_3[29720] = 32'b00000000000000011110100110100011;
assign LUT_3[29721] = 32'b00000000000000100101010010000000;
assign LUT_3[29722] = 32'b00000000000000100000101110000111;
assign LUT_3[29723] = 32'b00000000000000100111011001100100;
assign LUT_3[29724] = 32'b00000000000000011011110100011001;
assign LUT_3[29725] = 32'b00000000000000100010011111110110;
assign LUT_3[29726] = 32'b00000000000000011101111011111101;
assign LUT_3[29727] = 32'b00000000000000100100100111011010;
assign LUT_3[29728] = 32'b00000000000000010111001000111010;
assign LUT_3[29729] = 32'b00000000000000011101110100010111;
assign LUT_3[29730] = 32'b00000000000000011001010000011110;
assign LUT_3[29731] = 32'b00000000000000011111111011111011;
assign LUT_3[29732] = 32'b00000000000000010100010110110000;
assign LUT_3[29733] = 32'b00000000000000011011000010001101;
assign LUT_3[29734] = 32'b00000000000000010110011110010100;
assign LUT_3[29735] = 32'b00000000000000011101001001110001;
assign LUT_3[29736] = 32'b00000000000000011100100010000000;
assign LUT_3[29737] = 32'b00000000000000100011001101011101;
assign LUT_3[29738] = 32'b00000000000000011110101001100100;
assign LUT_3[29739] = 32'b00000000000000100101010101000001;
assign LUT_3[29740] = 32'b00000000000000011001101111110110;
assign LUT_3[29741] = 32'b00000000000000100000011011010011;
assign LUT_3[29742] = 32'b00000000000000011011110111011010;
assign LUT_3[29743] = 32'b00000000000000100010100010110111;
assign LUT_3[29744] = 32'b00000000000000011010011011111101;
assign LUT_3[29745] = 32'b00000000000000100001000111011010;
assign LUT_3[29746] = 32'b00000000000000011100100011100001;
assign LUT_3[29747] = 32'b00000000000000100011001110111110;
assign LUT_3[29748] = 32'b00000000000000010111101001110011;
assign LUT_3[29749] = 32'b00000000000000011110010101010000;
assign LUT_3[29750] = 32'b00000000000000011001110001010111;
assign LUT_3[29751] = 32'b00000000000000100000011100110100;
assign LUT_3[29752] = 32'b00000000000000011111110101000011;
assign LUT_3[29753] = 32'b00000000000000100110100000100000;
assign LUT_3[29754] = 32'b00000000000000100001111100100111;
assign LUT_3[29755] = 32'b00000000000000101000101000000100;
assign LUT_3[29756] = 32'b00000000000000011101000010111001;
assign LUT_3[29757] = 32'b00000000000000100011101110010110;
assign LUT_3[29758] = 32'b00000000000000011111001010011101;
assign LUT_3[29759] = 32'b00000000000000100101110101111010;
assign LUT_3[29760] = 32'b00000000000000010101110011000101;
assign LUT_3[29761] = 32'b00000000000000011100011110100010;
assign LUT_3[29762] = 32'b00000000000000010111111010101001;
assign LUT_3[29763] = 32'b00000000000000011110100110000110;
assign LUT_3[29764] = 32'b00000000000000010011000000111011;
assign LUT_3[29765] = 32'b00000000000000011001101100011000;
assign LUT_3[29766] = 32'b00000000000000010101001000011111;
assign LUT_3[29767] = 32'b00000000000000011011110011111100;
assign LUT_3[29768] = 32'b00000000000000011011001100001011;
assign LUT_3[29769] = 32'b00000000000000100001110111101000;
assign LUT_3[29770] = 32'b00000000000000011101010011101111;
assign LUT_3[29771] = 32'b00000000000000100011111111001100;
assign LUT_3[29772] = 32'b00000000000000011000011010000001;
assign LUT_3[29773] = 32'b00000000000000011111000101011110;
assign LUT_3[29774] = 32'b00000000000000011010100001100101;
assign LUT_3[29775] = 32'b00000000000000100001001101000010;
assign LUT_3[29776] = 32'b00000000000000011001000110001000;
assign LUT_3[29777] = 32'b00000000000000011111110001100101;
assign LUT_3[29778] = 32'b00000000000000011011001101101100;
assign LUT_3[29779] = 32'b00000000000000100001111001001001;
assign LUT_3[29780] = 32'b00000000000000010110010011111110;
assign LUT_3[29781] = 32'b00000000000000011100111111011011;
assign LUT_3[29782] = 32'b00000000000000011000011011100010;
assign LUT_3[29783] = 32'b00000000000000011111000110111111;
assign LUT_3[29784] = 32'b00000000000000011110011111001110;
assign LUT_3[29785] = 32'b00000000000000100101001010101011;
assign LUT_3[29786] = 32'b00000000000000100000100110110010;
assign LUT_3[29787] = 32'b00000000000000100111010010001111;
assign LUT_3[29788] = 32'b00000000000000011011101101000100;
assign LUT_3[29789] = 32'b00000000000000100010011000100001;
assign LUT_3[29790] = 32'b00000000000000011101110100101000;
assign LUT_3[29791] = 32'b00000000000000100100100000000101;
assign LUT_3[29792] = 32'b00000000000000010111000001100101;
assign LUT_3[29793] = 32'b00000000000000011101101101000010;
assign LUT_3[29794] = 32'b00000000000000011001001001001001;
assign LUT_3[29795] = 32'b00000000000000011111110100100110;
assign LUT_3[29796] = 32'b00000000000000010100001111011011;
assign LUT_3[29797] = 32'b00000000000000011010111010111000;
assign LUT_3[29798] = 32'b00000000000000010110010110111111;
assign LUT_3[29799] = 32'b00000000000000011101000010011100;
assign LUT_3[29800] = 32'b00000000000000011100011010101011;
assign LUT_3[29801] = 32'b00000000000000100011000110001000;
assign LUT_3[29802] = 32'b00000000000000011110100010001111;
assign LUT_3[29803] = 32'b00000000000000100101001101101100;
assign LUT_3[29804] = 32'b00000000000000011001101000100001;
assign LUT_3[29805] = 32'b00000000000000100000010011111110;
assign LUT_3[29806] = 32'b00000000000000011011110000000101;
assign LUT_3[29807] = 32'b00000000000000100010011011100010;
assign LUT_3[29808] = 32'b00000000000000011010010100101000;
assign LUT_3[29809] = 32'b00000000000000100001000000000101;
assign LUT_3[29810] = 32'b00000000000000011100011100001100;
assign LUT_3[29811] = 32'b00000000000000100011000111101001;
assign LUT_3[29812] = 32'b00000000000000010111100010011110;
assign LUT_3[29813] = 32'b00000000000000011110001101111011;
assign LUT_3[29814] = 32'b00000000000000011001101010000010;
assign LUT_3[29815] = 32'b00000000000000100000010101011111;
assign LUT_3[29816] = 32'b00000000000000011111101101101110;
assign LUT_3[29817] = 32'b00000000000000100110011001001011;
assign LUT_3[29818] = 32'b00000000000000100001110101010010;
assign LUT_3[29819] = 32'b00000000000000101000100000101111;
assign LUT_3[29820] = 32'b00000000000000011100111011100100;
assign LUT_3[29821] = 32'b00000000000000100011100111000001;
assign LUT_3[29822] = 32'b00000000000000011111000011001000;
assign LUT_3[29823] = 32'b00000000000000100101101110100101;
assign LUT_3[29824] = 32'b00000000000000011000000101011000;
assign LUT_3[29825] = 32'b00000000000000011110110000110101;
assign LUT_3[29826] = 32'b00000000000000011010001100111100;
assign LUT_3[29827] = 32'b00000000000000100000111000011001;
assign LUT_3[29828] = 32'b00000000000000010101010011001110;
assign LUT_3[29829] = 32'b00000000000000011011111110101011;
assign LUT_3[29830] = 32'b00000000000000010111011010110010;
assign LUT_3[29831] = 32'b00000000000000011110000110001111;
assign LUT_3[29832] = 32'b00000000000000011101011110011110;
assign LUT_3[29833] = 32'b00000000000000100100001001111011;
assign LUT_3[29834] = 32'b00000000000000011111100110000010;
assign LUT_3[29835] = 32'b00000000000000100110010001011111;
assign LUT_3[29836] = 32'b00000000000000011010101100010100;
assign LUT_3[29837] = 32'b00000000000000100001010111110001;
assign LUT_3[29838] = 32'b00000000000000011100110011111000;
assign LUT_3[29839] = 32'b00000000000000100011011111010101;
assign LUT_3[29840] = 32'b00000000000000011011011000011011;
assign LUT_3[29841] = 32'b00000000000000100010000011111000;
assign LUT_3[29842] = 32'b00000000000000011101011111111111;
assign LUT_3[29843] = 32'b00000000000000100100001011011100;
assign LUT_3[29844] = 32'b00000000000000011000100110010001;
assign LUT_3[29845] = 32'b00000000000000011111010001101110;
assign LUT_3[29846] = 32'b00000000000000011010101101110101;
assign LUT_3[29847] = 32'b00000000000000100001011001010010;
assign LUT_3[29848] = 32'b00000000000000100000110001100001;
assign LUT_3[29849] = 32'b00000000000000100111011100111110;
assign LUT_3[29850] = 32'b00000000000000100010111001000101;
assign LUT_3[29851] = 32'b00000000000000101001100100100010;
assign LUT_3[29852] = 32'b00000000000000011101111111010111;
assign LUT_3[29853] = 32'b00000000000000100100101010110100;
assign LUT_3[29854] = 32'b00000000000000100000000110111011;
assign LUT_3[29855] = 32'b00000000000000100110110010011000;
assign LUT_3[29856] = 32'b00000000000000011001010011111000;
assign LUT_3[29857] = 32'b00000000000000011111111111010101;
assign LUT_3[29858] = 32'b00000000000000011011011011011100;
assign LUT_3[29859] = 32'b00000000000000100010000110111001;
assign LUT_3[29860] = 32'b00000000000000010110100001101110;
assign LUT_3[29861] = 32'b00000000000000011101001101001011;
assign LUT_3[29862] = 32'b00000000000000011000101001010010;
assign LUT_3[29863] = 32'b00000000000000011111010100101111;
assign LUT_3[29864] = 32'b00000000000000011110101100111110;
assign LUT_3[29865] = 32'b00000000000000100101011000011011;
assign LUT_3[29866] = 32'b00000000000000100000110100100010;
assign LUT_3[29867] = 32'b00000000000000100111011111111111;
assign LUT_3[29868] = 32'b00000000000000011011111010110100;
assign LUT_3[29869] = 32'b00000000000000100010100110010001;
assign LUT_3[29870] = 32'b00000000000000011110000010011000;
assign LUT_3[29871] = 32'b00000000000000100100101101110101;
assign LUT_3[29872] = 32'b00000000000000011100100110111011;
assign LUT_3[29873] = 32'b00000000000000100011010010011000;
assign LUT_3[29874] = 32'b00000000000000011110101110011111;
assign LUT_3[29875] = 32'b00000000000000100101011001111100;
assign LUT_3[29876] = 32'b00000000000000011001110100110001;
assign LUT_3[29877] = 32'b00000000000000100000100000001110;
assign LUT_3[29878] = 32'b00000000000000011011111100010101;
assign LUT_3[29879] = 32'b00000000000000100010100111110010;
assign LUT_3[29880] = 32'b00000000000000100010000000000001;
assign LUT_3[29881] = 32'b00000000000000101000101011011110;
assign LUT_3[29882] = 32'b00000000000000100100000111100101;
assign LUT_3[29883] = 32'b00000000000000101010110011000010;
assign LUT_3[29884] = 32'b00000000000000011111001101110111;
assign LUT_3[29885] = 32'b00000000000000100101111001010100;
assign LUT_3[29886] = 32'b00000000000000100001010101011011;
assign LUT_3[29887] = 32'b00000000000000101000000000111000;
assign LUT_3[29888] = 32'b00000000000000010111111110000011;
assign LUT_3[29889] = 32'b00000000000000011110101001100000;
assign LUT_3[29890] = 32'b00000000000000011010000101100111;
assign LUT_3[29891] = 32'b00000000000000100000110001000100;
assign LUT_3[29892] = 32'b00000000000000010101001011111001;
assign LUT_3[29893] = 32'b00000000000000011011110111010110;
assign LUT_3[29894] = 32'b00000000000000010111010011011101;
assign LUT_3[29895] = 32'b00000000000000011101111110111010;
assign LUT_3[29896] = 32'b00000000000000011101010111001001;
assign LUT_3[29897] = 32'b00000000000000100100000010100110;
assign LUT_3[29898] = 32'b00000000000000011111011110101101;
assign LUT_3[29899] = 32'b00000000000000100110001010001010;
assign LUT_3[29900] = 32'b00000000000000011010100100111111;
assign LUT_3[29901] = 32'b00000000000000100001010000011100;
assign LUT_3[29902] = 32'b00000000000000011100101100100011;
assign LUT_3[29903] = 32'b00000000000000100011011000000000;
assign LUT_3[29904] = 32'b00000000000000011011010001000110;
assign LUT_3[29905] = 32'b00000000000000100001111100100011;
assign LUT_3[29906] = 32'b00000000000000011101011000101010;
assign LUT_3[29907] = 32'b00000000000000100100000100000111;
assign LUT_3[29908] = 32'b00000000000000011000011110111100;
assign LUT_3[29909] = 32'b00000000000000011111001010011001;
assign LUT_3[29910] = 32'b00000000000000011010100110100000;
assign LUT_3[29911] = 32'b00000000000000100001010001111101;
assign LUT_3[29912] = 32'b00000000000000100000101010001100;
assign LUT_3[29913] = 32'b00000000000000100111010101101001;
assign LUT_3[29914] = 32'b00000000000000100010110001110000;
assign LUT_3[29915] = 32'b00000000000000101001011101001101;
assign LUT_3[29916] = 32'b00000000000000011101111000000010;
assign LUT_3[29917] = 32'b00000000000000100100100011011111;
assign LUT_3[29918] = 32'b00000000000000011111111111100110;
assign LUT_3[29919] = 32'b00000000000000100110101011000011;
assign LUT_3[29920] = 32'b00000000000000011001001100100011;
assign LUT_3[29921] = 32'b00000000000000011111111000000000;
assign LUT_3[29922] = 32'b00000000000000011011010100000111;
assign LUT_3[29923] = 32'b00000000000000100001111111100100;
assign LUT_3[29924] = 32'b00000000000000010110011010011001;
assign LUT_3[29925] = 32'b00000000000000011101000101110110;
assign LUT_3[29926] = 32'b00000000000000011000100001111101;
assign LUT_3[29927] = 32'b00000000000000011111001101011010;
assign LUT_3[29928] = 32'b00000000000000011110100101101001;
assign LUT_3[29929] = 32'b00000000000000100101010001000110;
assign LUT_3[29930] = 32'b00000000000000100000101101001101;
assign LUT_3[29931] = 32'b00000000000000100111011000101010;
assign LUT_3[29932] = 32'b00000000000000011011110011011111;
assign LUT_3[29933] = 32'b00000000000000100010011110111100;
assign LUT_3[29934] = 32'b00000000000000011101111011000011;
assign LUT_3[29935] = 32'b00000000000000100100100110100000;
assign LUT_3[29936] = 32'b00000000000000011100011111100110;
assign LUT_3[29937] = 32'b00000000000000100011001011000011;
assign LUT_3[29938] = 32'b00000000000000011110100111001010;
assign LUT_3[29939] = 32'b00000000000000100101010010100111;
assign LUT_3[29940] = 32'b00000000000000011001101101011100;
assign LUT_3[29941] = 32'b00000000000000100000011000111001;
assign LUT_3[29942] = 32'b00000000000000011011110101000000;
assign LUT_3[29943] = 32'b00000000000000100010100000011101;
assign LUT_3[29944] = 32'b00000000000000100001111000101100;
assign LUT_3[29945] = 32'b00000000000000101000100100001001;
assign LUT_3[29946] = 32'b00000000000000100100000000010000;
assign LUT_3[29947] = 32'b00000000000000101010101011101101;
assign LUT_3[29948] = 32'b00000000000000011111000110100010;
assign LUT_3[29949] = 32'b00000000000000100101110001111111;
assign LUT_3[29950] = 32'b00000000000000100001001110000110;
assign LUT_3[29951] = 32'b00000000000000100111111001100011;
assign LUT_3[29952] = 32'b00000000000000010010001001111011;
assign LUT_3[29953] = 32'b00000000000000011000110101011000;
assign LUT_3[29954] = 32'b00000000000000010100010001011111;
assign LUT_3[29955] = 32'b00000000000000011010111100111100;
assign LUT_3[29956] = 32'b00000000000000001111010111110001;
assign LUT_3[29957] = 32'b00000000000000010110000011001110;
assign LUT_3[29958] = 32'b00000000000000010001011111010101;
assign LUT_3[29959] = 32'b00000000000000011000001010110010;
assign LUT_3[29960] = 32'b00000000000000010111100011000001;
assign LUT_3[29961] = 32'b00000000000000011110001110011110;
assign LUT_3[29962] = 32'b00000000000000011001101010100101;
assign LUT_3[29963] = 32'b00000000000000100000010110000010;
assign LUT_3[29964] = 32'b00000000000000010100110000110111;
assign LUT_3[29965] = 32'b00000000000000011011011100010100;
assign LUT_3[29966] = 32'b00000000000000010110111000011011;
assign LUT_3[29967] = 32'b00000000000000011101100011111000;
assign LUT_3[29968] = 32'b00000000000000010101011100111110;
assign LUT_3[29969] = 32'b00000000000000011100001000011011;
assign LUT_3[29970] = 32'b00000000000000010111100100100010;
assign LUT_3[29971] = 32'b00000000000000011110001111111111;
assign LUT_3[29972] = 32'b00000000000000010010101010110100;
assign LUT_3[29973] = 32'b00000000000000011001010110010001;
assign LUT_3[29974] = 32'b00000000000000010100110010011000;
assign LUT_3[29975] = 32'b00000000000000011011011101110101;
assign LUT_3[29976] = 32'b00000000000000011010110110000100;
assign LUT_3[29977] = 32'b00000000000000100001100001100001;
assign LUT_3[29978] = 32'b00000000000000011100111101101000;
assign LUT_3[29979] = 32'b00000000000000100011101001000101;
assign LUT_3[29980] = 32'b00000000000000011000000011111010;
assign LUT_3[29981] = 32'b00000000000000011110101111010111;
assign LUT_3[29982] = 32'b00000000000000011010001011011110;
assign LUT_3[29983] = 32'b00000000000000100000110110111011;
assign LUT_3[29984] = 32'b00000000000000010011011000011011;
assign LUT_3[29985] = 32'b00000000000000011010000011111000;
assign LUT_3[29986] = 32'b00000000000000010101011111111111;
assign LUT_3[29987] = 32'b00000000000000011100001011011100;
assign LUT_3[29988] = 32'b00000000000000010000100110010001;
assign LUT_3[29989] = 32'b00000000000000010111010001101110;
assign LUT_3[29990] = 32'b00000000000000010010101101110101;
assign LUT_3[29991] = 32'b00000000000000011001011001010010;
assign LUT_3[29992] = 32'b00000000000000011000110001100001;
assign LUT_3[29993] = 32'b00000000000000011111011100111110;
assign LUT_3[29994] = 32'b00000000000000011010111001000101;
assign LUT_3[29995] = 32'b00000000000000100001100100100010;
assign LUT_3[29996] = 32'b00000000000000010101111111010111;
assign LUT_3[29997] = 32'b00000000000000011100101010110100;
assign LUT_3[29998] = 32'b00000000000000011000000110111011;
assign LUT_3[29999] = 32'b00000000000000011110110010011000;
assign LUT_3[30000] = 32'b00000000000000010110101011011110;
assign LUT_3[30001] = 32'b00000000000000011101010110111011;
assign LUT_3[30002] = 32'b00000000000000011000110011000010;
assign LUT_3[30003] = 32'b00000000000000011111011110011111;
assign LUT_3[30004] = 32'b00000000000000010011111001010100;
assign LUT_3[30005] = 32'b00000000000000011010100100110001;
assign LUT_3[30006] = 32'b00000000000000010110000000111000;
assign LUT_3[30007] = 32'b00000000000000011100101100010101;
assign LUT_3[30008] = 32'b00000000000000011100000100100100;
assign LUT_3[30009] = 32'b00000000000000100010110000000001;
assign LUT_3[30010] = 32'b00000000000000011110001100001000;
assign LUT_3[30011] = 32'b00000000000000100100110111100101;
assign LUT_3[30012] = 32'b00000000000000011001010010011010;
assign LUT_3[30013] = 32'b00000000000000011111111101110111;
assign LUT_3[30014] = 32'b00000000000000011011011001111110;
assign LUT_3[30015] = 32'b00000000000000100010000101011011;
assign LUT_3[30016] = 32'b00000000000000010010000010100110;
assign LUT_3[30017] = 32'b00000000000000011000101110000011;
assign LUT_3[30018] = 32'b00000000000000010100001010001010;
assign LUT_3[30019] = 32'b00000000000000011010110101100111;
assign LUT_3[30020] = 32'b00000000000000001111010000011100;
assign LUT_3[30021] = 32'b00000000000000010101111011111001;
assign LUT_3[30022] = 32'b00000000000000010001011000000000;
assign LUT_3[30023] = 32'b00000000000000011000000011011101;
assign LUT_3[30024] = 32'b00000000000000010111011011101100;
assign LUT_3[30025] = 32'b00000000000000011110000111001001;
assign LUT_3[30026] = 32'b00000000000000011001100011010000;
assign LUT_3[30027] = 32'b00000000000000100000001110101101;
assign LUT_3[30028] = 32'b00000000000000010100101001100010;
assign LUT_3[30029] = 32'b00000000000000011011010100111111;
assign LUT_3[30030] = 32'b00000000000000010110110001000110;
assign LUT_3[30031] = 32'b00000000000000011101011100100011;
assign LUT_3[30032] = 32'b00000000000000010101010101101001;
assign LUT_3[30033] = 32'b00000000000000011100000001000110;
assign LUT_3[30034] = 32'b00000000000000010111011101001101;
assign LUT_3[30035] = 32'b00000000000000011110001000101010;
assign LUT_3[30036] = 32'b00000000000000010010100011011111;
assign LUT_3[30037] = 32'b00000000000000011001001110111100;
assign LUT_3[30038] = 32'b00000000000000010100101011000011;
assign LUT_3[30039] = 32'b00000000000000011011010110100000;
assign LUT_3[30040] = 32'b00000000000000011010101110101111;
assign LUT_3[30041] = 32'b00000000000000100001011010001100;
assign LUT_3[30042] = 32'b00000000000000011100110110010011;
assign LUT_3[30043] = 32'b00000000000000100011100001110000;
assign LUT_3[30044] = 32'b00000000000000010111111100100101;
assign LUT_3[30045] = 32'b00000000000000011110101000000010;
assign LUT_3[30046] = 32'b00000000000000011010000100001001;
assign LUT_3[30047] = 32'b00000000000000100000101111100110;
assign LUT_3[30048] = 32'b00000000000000010011010001000110;
assign LUT_3[30049] = 32'b00000000000000011001111100100011;
assign LUT_3[30050] = 32'b00000000000000010101011000101010;
assign LUT_3[30051] = 32'b00000000000000011100000100000111;
assign LUT_3[30052] = 32'b00000000000000010000011110111100;
assign LUT_3[30053] = 32'b00000000000000010111001010011001;
assign LUT_3[30054] = 32'b00000000000000010010100110100000;
assign LUT_3[30055] = 32'b00000000000000011001010001111101;
assign LUT_3[30056] = 32'b00000000000000011000101010001100;
assign LUT_3[30057] = 32'b00000000000000011111010101101001;
assign LUT_3[30058] = 32'b00000000000000011010110001110000;
assign LUT_3[30059] = 32'b00000000000000100001011101001101;
assign LUT_3[30060] = 32'b00000000000000010101111000000010;
assign LUT_3[30061] = 32'b00000000000000011100100011011111;
assign LUT_3[30062] = 32'b00000000000000010111111111100110;
assign LUT_3[30063] = 32'b00000000000000011110101011000011;
assign LUT_3[30064] = 32'b00000000000000010110100100001001;
assign LUT_3[30065] = 32'b00000000000000011101001111100110;
assign LUT_3[30066] = 32'b00000000000000011000101011101101;
assign LUT_3[30067] = 32'b00000000000000011111010111001010;
assign LUT_3[30068] = 32'b00000000000000010011110001111111;
assign LUT_3[30069] = 32'b00000000000000011010011101011100;
assign LUT_3[30070] = 32'b00000000000000010101111001100011;
assign LUT_3[30071] = 32'b00000000000000011100100101000000;
assign LUT_3[30072] = 32'b00000000000000011011111101001111;
assign LUT_3[30073] = 32'b00000000000000100010101000101100;
assign LUT_3[30074] = 32'b00000000000000011110000100110011;
assign LUT_3[30075] = 32'b00000000000000100100110000010000;
assign LUT_3[30076] = 32'b00000000000000011001001011000101;
assign LUT_3[30077] = 32'b00000000000000011111110110100010;
assign LUT_3[30078] = 32'b00000000000000011011010010101001;
assign LUT_3[30079] = 32'b00000000000000100001111110000110;
assign LUT_3[30080] = 32'b00000000000000010100010100111001;
assign LUT_3[30081] = 32'b00000000000000011011000000010110;
assign LUT_3[30082] = 32'b00000000000000010110011100011101;
assign LUT_3[30083] = 32'b00000000000000011101000111111010;
assign LUT_3[30084] = 32'b00000000000000010001100010101111;
assign LUT_3[30085] = 32'b00000000000000011000001110001100;
assign LUT_3[30086] = 32'b00000000000000010011101010010011;
assign LUT_3[30087] = 32'b00000000000000011010010101110000;
assign LUT_3[30088] = 32'b00000000000000011001101101111111;
assign LUT_3[30089] = 32'b00000000000000100000011001011100;
assign LUT_3[30090] = 32'b00000000000000011011110101100011;
assign LUT_3[30091] = 32'b00000000000000100010100001000000;
assign LUT_3[30092] = 32'b00000000000000010110111011110101;
assign LUT_3[30093] = 32'b00000000000000011101100111010010;
assign LUT_3[30094] = 32'b00000000000000011001000011011001;
assign LUT_3[30095] = 32'b00000000000000011111101110110110;
assign LUT_3[30096] = 32'b00000000000000010111100111111100;
assign LUT_3[30097] = 32'b00000000000000011110010011011001;
assign LUT_3[30098] = 32'b00000000000000011001101111100000;
assign LUT_3[30099] = 32'b00000000000000100000011010111101;
assign LUT_3[30100] = 32'b00000000000000010100110101110010;
assign LUT_3[30101] = 32'b00000000000000011011100001001111;
assign LUT_3[30102] = 32'b00000000000000010110111101010110;
assign LUT_3[30103] = 32'b00000000000000011101101000110011;
assign LUT_3[30104] = 32'b00000000000000011101000001000010;
assign LUT_3[30105] = 32'b00000000000000100011101100011111;
assign LUT_3[30106] = 32'b00000000000000011111001000100110;
assign LUT_3[30107] = 32'b00000000000000100101110100000011;
assign LUT_3[30108] = 32'b00000000000000011010001110111000;
assign LUT_3[30109] = 32'b00000000000000100000111010010101;
assign LUT_3[30110] = 32'b00000000000000011100010110011100;
assign LUT_3[30111] = 32'b00000000000000100011000001111001;
assign LUT_3[30112] = 32'b00000000000000010101100011011001;
assign LUT_3[30113] = 32'b00000000000000011100001110110110;
assign LUT_3[30114] = 32'b00000000000000010111101010111101;
assign LUT_3[30115] = 32'b00000000000000011110010110011010;
assign LUT_3[30116] = 32'b00000000000000010010110001001111;
assign LUT_3[30117] = 32'b00000000000000011001011100101100;
assign LUT_3[30118] = 32'b00000000000000010100111000110011;
assign LUT_3[30119] = 32'b00000000000000011011100100010000;
assign LUT_3[30120] = 32'b00000000000000011010111100011111;
assign LUT_3[30121] = 32'b00000000000000100001100111111100;
assign LUT_3[30122] = 32'b00000000000000011101000100000011;
assign LUT_3[30123] = 32'b00000000000000100011101111100000;
assign LUT_3[30124] = 32'b00000000000000011000001010010101;
assign LUT_3[30125] = 32'b00000000000000011110110101110010;
assign LUT_3[30126] = 32'b00000000000000011010010001111001;
assign LUT_3[30127] = 32'b00000000000000100000111101010110;
assign LUT_3[30128] = 32'b00000000000000011000110110011100;
assign LUT_3[30129] = 32'b00000000000000011111100001111001;
assign LUT_3[30130] = 32'b00000000000000011010111110000000;
assign LUT_3[30131] = 32'b00000000000000100001101001011101;
assign LUT_3[30132] = 32'b00000000000000010110000100010010;
assign LUT_3[30133] = 32'b00000000000000011100101111101111;
assign LUT_3[30134] = 32'b00000000000000011000001011110110;
assign LUT_3[30135] = 32'b00000000000000011110110111010011;
assign LUT_3[30136] = 32'b00000000000000011110001111100010;
assign LUT_3[30137] = 32'b00000000000000100100111010111111;
assign LUT_3[30138] = 32'b00000000000000100000010111000110;
assign LUT_3[30139] = 32'b00000000000000100111000010100011;
assign LUT_3[30140] = 32'b00000000000000011011011101011000;
assign LUT_3[30141] = 32'b00000000000000100010001000110101;
assign LUT_3[30142] = 32'b00000000000000011101100100111100;
assign LUT_3[30143] = 32'b00000000000000100100010000011001;
assign LUT_3[30144] = 32'b00000000000000010100001101100100;
assign LUT_3[30145] = 32'b00000000000000011010111001000001;
assign LUT_3[30146] = 32'b00000000000000010110010101001000;
assign LUT_3[30147] = 32'b00000000000000011101000000100101;
assign LUT_3[30148] = 32'b00000000000000010001011011011010;
assign LUT_3[30149] = 32'b00000000000000011000000110110111;
assign LUT_3[30150] = 32'b00000000000000010011100010111110;
assign LUT_3[30151] = 32'b00000000000000011010001110011011;
assign LUT_3[30152] = 32'b00000000000000011001100110101010;
assign LUT_3[30153] = 32'b00000000000000100000010010000111;
assign LUT_3[30154] = 32'b00000000000000011011101110001110;
assign LUT_3[30155] = 32'b00000000000000100010011001101011;
assign LUT_3[30156] = 32'b00000000000000010110110100100000;
assign LUT_3[30157] = 32'b00000000000000011101011111111101;
assign LUT_3[30158] = 32'b00000000000000011000111100000100;
assign LUT_3[30159] = 32'b00000000000000011111100111100001;
assign LUT_3[30160] = 32'b00000000000000010111100000100111;
assign LUT_3[30161] = 32'b00000000000000011110001100000100;
assign LUT_3[30162] = 32'b00000000000000011001101000001011;
assign LUT_3[30163] = 32'b00000000000000100000010011101000;
assign LUT_3[30164] = 32'b00000000000000010100101110011101;
assign LUT_3[30165] = 32'b00000000000000011011011001111010;
assign LUT_3[30166] = 32'b00000000000000010110110110000001;
assign LUT_3[30167] = 32'b00000000000000011101100001011110;
assign LUT_3[30168] = 32'b00000000000000011100111001101101;
assign LUT_3[30169] = 32'b00000000000000100011100101001010;
assign LUT_3[30170] = 32'b00000000000000011111000001010001;
assign LUT_3[30171] = 32'b00000000000000100101101100101110;
assign LUT_3[30172] = 32'b00000000000000011010000111100011;
assign LUT_3[30173] = 32'b00000000000000100000110011000000;
assign LUT_3[30174] = 32'b00000000000000011100001111000111;
assign LUT_3[30175] = 32'b00000000000000100010111010100100;
assign LUT_3[30176] = 32'b00000000000000010101011100000100;
assign LUT_3[30177] = 32'b00000000000000011100000111100001;
assign LUT_3[30178] = 32'b00000000000000010111100011101000;
assign LUT_3[30179] = 32'b00000000000000011110001111000101;
assign LUT_3[30180] = 32'b00000000000000010010101001111010;
assign LUT_3[30181] = 32'b00000000000000011001010101010111;
assign LUT_3[30182] = 32'b00000000000000010100110001011110;
assign LUT_3[30183] = 32'b00000000000000011011011100111011;
assign LUT_3[30184] = 32'b00000000000000011010110101001010;
assign LUT_3[30185] = 32'b00000000000000100001100000100111;
assign LUT_3[30186] = 32'b00000000000000011100111100101110;
assign LUT_3[30187] = 32'b00000000000000100011101000001011;
assign LUT_3[30188] = 32'b00000000000000011000000011000000;
assign LUT_3[30189] = 32'b00000000000000011110101110011101;
assign LUT_3[30190] = 32'b00000000000000011010001010100100;
assign LUT_3[30191] = 32'b00000000000000100000110110000001;
assign LUT_3[30192] = 32'b00000000000000011000101111000111;
assign LUT_3[30193] = 32'b00000000000000011111011010100100;
assign LUT_3[30194] = 32'b00000000000000011010110110101011;
assign LUT_3[30195] = 32'b00000000000000100001100010001000;
assign LUT_3[30196] = 32'b00000000000000010101111100111101;
assign LUT_3[30197] = 32'b00000000000000011100101000011010;
assign LUT_3[30198] = 32'b00000000000000011000000100100001;
assign LUT_3[30199] = 32'b00000000000000011110101111111110;
assign LUT_3[30200] = 32'b00000000000000011110001000001101;
assign LUT_3[30201] = 32'b00000000000000100100110011101010;
assign LUT_3[30202] = 32'b00000000000000100000001111110001;
assign LUT_3[30203] = 32'b00000000000000100110111011001110;
assign LUT_3[30204] = 32'b00000000000000011011010110000011;
assign LUT_3[30205] = 32'b00000000000000100010000001100000;
assign LUT_3[30206] = 32'b00000000000000011101011101100111;
assign LUT_3[30207] = 32'b00000000000000100100001001000100;
assign LUT_3[30208] = 32'b00000000000000011001001111100110;
assign LUT_3[30209] = 32'b00000000000000011111111011000011;
assign LUT_3[30210] = 32'b00000000000000011011010111001010;
assign LUT_3[30211] = 32'b00000000000000100010000010100111;
assign LUT_3[30212] = 32'b00000000000000010110011101011100;
assign LUT_3[30213] = 32'b00000000000000011101001000111001;
assign LUT_3[30214] = 32'b00000000000000011000100101000000;
assign LUT_3[30215] = 32'b00000000000000011111010000011101;
assign LUT_3[30216] = 32'b00000000000000011110101000101100;
assign LUT_3[30217] = 32'b00000000000000100101010100001001;
assign LUT_3[30218] = 32'b00000000000000100000110000010000;
assign LUT_3[30219] = 32'b00000000000000100111011011101101;
assign LUT_3[30220] = 32'b00000000000000011011110110100010;
assign LUT_3[30221] = 32'b00000000000000100010100001111111;
assign LUT_3[30222] = 32'b00000000000000011101111110000110;
assign LUT_3[30223] = 32'b00000000000000100100101001100011;
assign LUT_3[30224] = 32'b00000000000000011100100010101001;
assign LUT_3[30225] = 32'b00000000000000100011001110000110;
assign LUT_3[30226] = 32'b00000000000000011110101010001101;
assign LUT_3[30227] = 32'b00000000000000100101010101101010;
assign LUT_3[30228] = 32'b00000000000000011001110000011111;
assign LUT_3[30229] = 32'b00000000000000100000011011111100;
assign LUT_3[30230] = 32'b00000000000000011011111000000011;
assign LUT_3[30231] = 32'b00000000000000100010100011100000;
assign LUT_3[30232] = 32'b00000000000000100001111011101111;
assign LUT_3[30233] = 32'b00000000000000101000100111001100;
assign LUT_3[30234] = 32'b00000000000000100100000011010011;
assign LUT_3[30235] = 32'b00000000000000101010101110110000;
assign LUT_3[30236] = 32'b00000000000000011111001001100101;
assign LUT_3[30237] = 32'b00000000000000100101110101000010;
assign LUT_3[30238] = 32'b00000000000000100001010001001001;
assign LUT_3[30239] = 32'b00000000000000100111111100100110;
assign LUT_3[30240] = 32'b00000000000000011010011110000110;
assign LUT_3[30241] = 32'b00000000000000100001001001100011;
assign LUT_3[30242] = 32'b00000000000000011100100101101010;
assign LUT_3[30243] = 32'b00000000000000100011010001000111;
assign LUT_3[30244] = 32'b00000000000000010111101011111100;
assign LUT_3[30245] = 32'b00000000000000011110010111011001;
assign LUT_3[30246] = 32'b00000000000000011001110011100000;
assign LUT_3[30247] = 32'b00000000000000100000011110111101;
assign LUT_3[30248] = 32'b00000000000000011111110111001100;
assign LUT_3[30249] = 32'b00000000000000100110100010101001;
assign LUT_3[30250] = 32'b00000000000000100001111110110000;
assign LUT_3[30251] = 32'b00000000000000101000101010001101;
assign LUT_3[30252] = 32'b00000000000000011101000101000010;
assign LUT_3[30253] = 32'b00000000000000100011110000011111;
assign LUT_3[30254] = 32'b00000000000000011111001100100110;
assign LUT_3[30255] = 32'b00000000000000100101111000000011;
assign LUT_3[30256] = 32'b00000000000000011101110001001001;
assign LUT_3[30257] = 32'b00000000000000100100011100100110;
assign LUT_3[30258] = 32'b00000000000000011111111000101101;
assign LUT_3[30259] = 32'b00000000000000100110100100001010;
assign LUT_3[30260] = 32'b00000000000000011010111110111111;
assign LUT_3[30261] = 32'b00000000000000100001101010011100;
assign LUT_3[30262] = 32'b00000000000000011101000110100011;
assign LUT_3[30263] = 32'b00000000000000100011110010000000;
assign LUT_3[30264] = 32'b00000000000000100011001010001111;
assign LUT_3[30265] = 32'b00000000000000101001110101101100;
assign LUT_3[30266] = 32'b00000000000000100101010001110011;
assign LUT_3[30267] = 32'b00000000000000101011111101010000;
assign LUT_3[30268] = 32'b00000000000000100000011000000101;
assign LUT_3[30269] = 32'b00000000000000100111000011100010;
assign LUT_3[30270] = 32'b00000000000000100010011111101001;
assign LUT_3[30271] = 32'b00000000000000101001001011000110;
assign LUT_3[30272] = 32'b00000000000000011001001000010001;
assign LUT_3[30273] = 32'b00000000000000011111110011101110;
assign LUT_3[30274] = 32'b00000000000000011011001111110101;
assign LUT_3[30275] = 32'b00000000000000100001111011010010;
assign LUT_3[30276] = 32'b00000000000000010110010110000111;
assign LUT_3[30277] = 32'b00000000000000011101000001100100;
assign LUT_3[30278] = 32'b00000000000000011000011101101011;
assign LUT_3[30279] = 32'b00000000000000011111001001001000;
assign LUT_3[30280] = 32'b00000000000000011110100001010111;
assign LUT_3[30281] = 32'b00000000000000100101001100110100;
assign LUT_3[30282] = 32'b00000000000000100000101000111011;
assign LUT_3[30283] = 32'b00000000000000100111010100011000;
assign LUT_3[30284] = 32'b00000000000000011011101111001101;
assign LUT_3[30285] = 32'b00000000000000100010011010101010;
assign LUT_3[30286] = 32'b00000000000000011101110110110001;
assign LUT_3[30287] = 32'b00000000000000100100100010001110;
assign LUT_3[30288] = 32'b00000000000000011100011011010100;
assign LUT_3[30289] = 32'b00000000000000100011000110110001;
assign LUT_3[30290] = 32'b00000000000000011110100010111000;
assign LUT_3[30291] = 32'b00000000000000100101001110010101;
assign LUT_3[30292] = 32'b00000000000000011001101001001010;
assign LUT_3[30293] = 32'b00000000000000100000010100100111;
assign LUT_3[30294] = 32'b00000000000000011011110000101110;
assign LUT_3[30295] = 32'b00000000000000100010011100001011;
assign LUT_3[30296] = 32'b00000000000000100001110100011010;
assign LUT_3[30297] = 32'b00000000000000101000011111110111;
assign LUT_3[30298] = 32'b00000000000000100011111011111110;
assign LUT_3[30299] = 32'b00000000000000101010100111011011;
assign LUT_3[30300] = 32'b00000000000000011111000010010000;
assign LUT_3[30301] = 32'b00000000000000100101101101101101;
assign LUT_3[30302] = 32'b00000000000000100001001001110100;
assign LUT_3[30303] = 32'b00000000000000100111110101010001;
assign LUT_3[30304] = 32'b00000000000000011010010110110001;
assign LUT_3[30305] = 32'b00000000000000100001000010001110;
assign LUT_3[30306] = 32'b00000000000000011100011110010101;
assign LUT_3[30307] = 32'b00000000000000100011001001110010;
assign LUT_3[30308] = 32'b00000000000000010111100100100111;
assign LUT_3[30309] = 32'b00000000000000011110010000000100;
assign LUT_3[30310] = 32'b00000000000000011001101100001011;
assign LUT_3[30311] = 32'b00000000000000100000010111101000;
assign LUT_3[30312] = 32'b00000000000000011111101111110111;
assign LUT_3[30313] = 32'b00000000000000100110011011010100;
assign LUT_3[30314] = 32'b00000000000000100001110111011011;
assign LUT_3[30315] = 32'b00000000000000101000100010111000;
assign LUT_3[30316] = 32'b00000000000000011100111101101101;
assign LUT_3[30317] = 32'b00000000000000100011101001001010;
assign LUT_3[30318] = 32'b00000000000000011111000101010001;
assign LUT_3[30319] = 32'b00000000000000100101110000101110;
assign LUT_3[30320] = 32'b00000000000000011101101001110100;
assign LUT_3[30321] = 32'b00000000000000100100010101010001;
assign LUT_3[30322] = 32'b00000000000000011111110001011000;
assign LUT_3[30323] = 32'b00000000000000100110011100110101;
assign LUT_3[30324] = 32'b00000000000000011010110111101010;
assign LUT_3[30325] = 32'b00000000000000100001100011000111;
assign LUT_3[30326] = 32'b00000000000000011100111111001110;
assign LUT_3[30327] = 32'b00000000000000100011101010101011;
assign LUT_3[30328] = 32'b00000000000000100011000010111010;
assign LUT_3[30329] = 32'b00000000000000101001101110010111;
assign LUT_3[30330] = 32'b00000000000000100101001010011110;
assign LUT_3[30331] = 32'b00000000000000101011110101111011;
assign LUT_3[30332] = 32'b00000000000000100000010000110000;
assign LUT_3[30333] = 32'b00000000000000100110111100001101;
assign LUT_3[30334] = 32'b00000000000000100010011000010100;
assign LUT_3[30335] = 32'b00000000000000101001000011110001;
assign LUT_3[30336] = 32'b00000000000000011011011010100100;
assign LUT_3[30337] = 32'b00000000000000100010000110000001;
assign LUT_3[30338] = 32'b00000000000000011101100010001000;
assign LUT_3[30339] = 32'b00000000000000100100001101100101;
assign LUT_3[30340] = 32'b00000000000000011000101000011010;
assign LUT_3[30341] = 32'b00000000000000011111010011110111;
assign LUT_3[30342] = 32'b00000000000000011010101111111110;
assign LUT_3[30343] = 32'b00000000000000100001011011011011;
assign LUT_3[30344] = 32'b00000000000000100000110011101010;
assign LUT_3[30345] = 32'b00000000000000100111011111000111;
assign LUT_3[30346] = 32'b00000000000000100010111011001110;
assign LUT_3[30347] = 32'b00000000000000101001100110101011;
assign LUT_3[30348] = 32'b00000000000000011110000001100000;
assign LUT_3[30349] = 32'b00000000000000100100101100111101;
assign LUT_3[30350] = 32'b00000000000000100000001001000100;
assign LUT_3[30351] = 32'b00000000000000100110110100100001;
assign LUT_3[30352] = 32'b00000000000000011110101101100111;
assign LUT_3[30353] = 32'b00000000000000100101011001000100;
assign LUT_3[30354] = 32'b00000000000000100000110101001011;
assign LUT_3[30355] = 32'b00000000000000100111100000101000;
assign LUT_3[30356] = 32'b00000000000000011011111011011101;
assign LUT_3[30357] = 32'b00000000000000100010100110111010;
assign LUT_3[30358] = 32'b00000000000000011110000011000001;
assign LUT_3[30359] = 32'b00000000000000100100101110011110;
assign LUT_3[30360] = 32'b00000000000000100100000110101101;
assign LUT_3[30361] = 32'b00000000000000101010110010001010;
assign LUT_3[30362] = 32'b00000000000000100110001110010001;
assign LUT_3[30363] = 32'b00000000000000101100111001101110;
assign LUT_3[30364] = 32'b00000000000000100001010100100011;
assign LUT_3[30365] = 32'b00000000000000101000000000000000;
assign LUT_3[30366] = 32'b00000000000000100011011100000111;
assign LUT_3[30367] = 32'b00000000000000101010000111100100;
assign LUT_3[30368] = 32'b00000000000000011100101001000100;
assign LUT_3[30369] = 32'b00000000000000100011010100100001;
assign LUT_3[30370] = 32'b00000000000000011110110000101000;
assign LUT_3[30371] = 32'b00000000000000100101011100000101;
assign LUT_3[30372] = 32'b00000000000000011001110110111010;
assign LUT_3[30373] = 32'b00000000000000100000100010010111;
assign LUT_3[30374] = 32'b00000000000000011011111110011110;
assign LUT_3[30375] = 32'b00000000000000100010101001111011;
assign LUT_3[30376] = 32'b00000000000000100010000010001010;
assign LUT_3[30377] = 32'b00000000000000101000101101100111;
assign LUT_3[30378] = 32'b00000000000000100100001001101110;
assign LUT_3[30379] = 32'b00000000000000101010110101001011;
assign LUT_3[30380] = 32'b00000000000000011111010000000000;
assign LUT_3[30381] = 32'b00000000000000100101111011011101;
assign LUT_3[30382] = 32'b00000000000000100001010111100100;
assign LUT_3[30383] = 32'b00000000000000101000000011000001;
assign LUT_3[30384] = 32'b00000000000000011111111100000111;
assign LUT_3[30385] = 32'b00000000000000100110100111100100;
assign LUT_3[30386] = 32'b00000000000000100010000011101011;
assign LUT_3[30387] = 32'b00000000000000101000101111001000;
assign LUT_3[30388] = 32'b00000000000000011101001001111101;
assign LUT_3[30389] = 32'b00000000000000100011110101011010;
assign LUT_3[30390] = 32'b00000000000000011111010001100001;
assign LUT_3[30391] = 32'b00000000000000100101111100111110;
assign LUT_3[30392] = 32'b00000000000000100101010101001101;
assign LUT_3[30393] = 32'b00000000000000101100000000101010;
assign LUT_3[30394] = 32'b00000000000000100111011100110001;
assign LUT_3[30395] = 32'b00000000000000101110001000001110;
assign LUT_3[30396] = 32'b00000000000000100010100011000011;
assign LUT_3[30397] = 32'b00000000000000101001001110100000;
assign LUT_3[30398] = 32'b00000000000000100100101010100111;
assign LUT_3[30399] = 32'b00000000000000101011010110000100;
assign LUT_3[30400] = 32'b00000000000000011011010011001111;
assign LUT_3[30401] = 32'b00000000000000100001111110101100;
assign LUT_3[30402] = 32'b00000000000000011101011010110011;
assign LUT_3[30403] = 32'b00000000000000100100000110010000;
assign LUT_3[30404] = 32'b00000000000000011000100001000101;
assign LUT_3[30405] = 32'b00000000000000011111001100100010;
assign LUT_3[30406] = 32'b00000000000000011010101000101001;
assign LUT_3[30407] = 32'b00000000000000100001010100000110;
assign LUT_3[30408] = 32'b00000000000000100000101100010101;
assign LUT_3[30409] = 32'b00000000000000100111010111110010;
assign LUT_3[30410] = 32'b00000000000000100010110011111001;
assign LUT_3[30411] = 32'b00000000000000101001011111010110;
assign LUT_3[30412] = 32'b00000000000000011101111010001011;
assign LUT_3[30413] = 32'b00000000000000100100100101101000;
assign LUT_3[30414] = 32'b00000000000000100000000001101111;
assign LUT_3[30415] = 32'b00000000000000100110101101001100;
assign LUT_3[30416] = 32'b00000000000000011110100110010010;
assign LUT_3[30417] = 32'b00000000000000100101010001101111;
assign LUT_3[30418] = 32'b00000000000000100000101101110110;
assign LUT_3[30419] = 32'b00000000000000100111011001010011;
assign LUT_3[30420] = 32'b00000000000000011011110100001000;
assign LUT_3[30421] = 32'b00000000000000100010011111100101;
assign LUT_3[30422] = 32'b00000000000000011101111011101100;
assign LUT_3[30423] = 32'b00000000000000100100100111001001;
assign LUT_3[30424] = 32'b00000000000000100011111111011000;
assign LUT_3[30425] = 32'b00000000000000101010101010110101;
assign LUT_3[30426] = 32'b00000000000000100110000110111100;
assign LUT_3[30427] = 32'b00000000000000101100110010011001;
assign LUT_3[30428] = 32'b00000000000000100001001101001110;
assign LUT_3[30429] = 32'b00000000000000100111111000101011;
assign LUT_3[30430] = 32'b00000000000000100011010100110010;
assign LUT_3[30431] = 32'b00000000000000101010000000001111;
assign LUT_3[30432] = 32'b00000000000000011100100001101111;
assign LUT_3[30433] = 32'b00000000000000100011001101001100;
assign LUT_3[30434] = 32'b00000000000000011110101001010011;
assign LUT_3[30435] = 32'b00000000000000100101010100110000;
assign LUT_3[30436] = 32'b00000000000000011001101111100101;
assign LUT_3[30437] = 32'b00000000000000100000011011000010;
assign LUT_3[30438] = 32'b00000000000000011011110111001001;
assign LUT_3[30439] = 32'b00000000000000100010100010100110;
assign LUT_3[30440] = 32'b00000000000000100001111010110101;
assign LUT_3[30441] = 32'b00000000000000101000100110010010;
assign LUT_3[30442] = 32'b00000000000000100100000010011001;
assign LUT_3[30443] = 32'b00000000000000101010101101110110;
assign LUT_3[30444] = 32'b00000000000000011111001000101011;
assign LUT_3[30445] = 32'b00000000000000100101110100001000;
assign LUT_3[30446] = 32'b00000000000000100001010000001111;
assign LUT_3[30447] = 32'b00000000000000100111111011101100;
assign LUT_3[30448] = 32'b00000000000000011111110100110010;
assign LUT_3[30449] = 32'b00000000000000100110100000001111;
assign LUT_3[30450] = 32'b00000000000000100001111100010110;
assign LUT_3[30451] = 32'b00000000000000101000100111110011;
assign LUT_3[30452] = 32'b00000000000000011101000010101000;
assign LUT_3[30453] = 32'b00000000000000100011101110000101;
assign LUT_3[30454] = 32'b00000000000000011111001010001100;
assign LUT_3[30455] = 32'b00000000000000100101110101101001;
assign LUT_3[30456] = 32'b00000000000000100101001101111000;
assign LUT_3[30457] = 32'b00000000000000101011111001010101;
assign LUT_3[30458] = 32'b00000000000000100111010101011100;
assign LUT_3[30459] = 32'b00000000000000101110000000111001;
assign LUT_3[30460] = 32'b00000000000000100010011011101110;
assign LUT_3[30461] = 32'b00000000000000101001000111001011;
assign LUT_3[30462] = 32'b00000000000000100100100011010010;
assign LUT_3[30463] = 32'b00000000000000101011001110101111;
assign LUT_3[30464] = 32'b00000000000000010101011111000111;
assign LUT_3[30465] = 32'b00000000000000011100001010100100;
assign LUT_3[30466] = 32'b00000000000000010111100110101011;
assign LUT_3[30467] = 32'b00000000000000011110010010001000;
assign LUT_3[30468] = 32'b00000000000000010010101100111101;
assign LUT_3[30469] = 32'b00000000000000011001011000011010;
assign LUT_3[30470] = 32'b00000000000000010100110100100001;
assign LUT_3[30471] = 32'b00000000000000011011011111111110;
assign LUT_3[30472] = 32'b00000000000000011010111000001101;
assign LUT_3[30473] = 32'b00000000000000100001100011101010;
assign LUT_3[30474] = 32'b00000000000000011100111111110001;
assign LUT_3[30475] = 32'b00000000000000100011101011001110;
assign LUT_3[30476] = 32'b00000000000000011000000110000011;
assign LUT_3[30477] = 32'b00000000000000011110110001100000;
assign LUT_3[30478] = 32'b00000000000000011010001101100111;
assign LUT_3[30479] = 32'b00000000000000100000111001000100;
assign LUT_3[30480] = 32'b00000000000000011000110010001010;
assign LUT_3[30481] = 32'b00000000000000011111011101100111;
assign LUT_3[30482] = 32'b00000000000000011010111001101110;
assign LUT_3[30483] = 32'b00000000000000100001100101001011;
assign LUT_3[30484] = 32'b00000000000000010110000000000000;
assign LUT_3[30485] = 32'b00000000000000011100101011011101;
assign LUT_3[30486] = 32'b00000000000000011000000111100100;
assign LUT_3[30487] = 32'b00000000000000011110110011000001;
assign LUT_3[30488] = 32'b00000000000000011110001011010000;
assign LUT_3[30489] = 32'b00000000000000100100110110101101;
assign LUT_3[30490] = 32'b00000000000000100000010010110100;
assign LUT_3[30491] = 32'b00000000000000100110111110010001;
assign LUT_3[30492] = 32'b00000000000000011011011001000110;
assign LUT_3[30493] = 32'b00000000000000100010000100100011;
assign LUT_3[30494] = 32'b00000000000000011101100000101010;
assign LUT_3[30495] = 32'b00000000000000100100001100000111;
assign LUT_3[30496] = 32'b00000000000000010110101101100111;
assign LUT_3[30497] = 32'b00000000000000011101011001000100;
assign LUT_3[30498] = 32'b00000000000000011000110101001011;
assign LUT_3[30499] = 32'b00000000000000011111100000101000;
assign LUT_3[30500] = 32'b00000000000000010011111011011101;
assign LUT_3[30501] = 32'b00000000000000011010100110111010;
assign LUT_3[30502] = 32'b00000000000000010110000011000001;
assign LUT_3[30503] = 32'b00000000000000011100101110011110;
assign LUT_3[30504] = 32'b00000000000000011100000110101101;
assign LUT_3[30505] = 32'b00000000000000100010110010001010;
assign LUT_3[30506] = 32'b00000000000000011110001110010001;
assign LUT_3[30507] = 32'b00000000000000100100111001101110;
assign LUT_3[30508] = 32'b00000000000000011001010100100011;
assign LUT_3[30509] = 32'b00000000000000100000000000000000;
assign LUT_3[30510] = 32'b00000000000000011011011100000111;
assign LUT_3[30511] = 32'b00000000000000100010000111100100;
assign LUT_3[30512] = 32'b00000000000000011010000000101010;
assign LUT_3[30513] = 32'b00000000000000100000101100000111;
assign LUT_3[30514] = 32'b00000000000000011100001000001110;
assign LUT_3[30515] = 32'b00000000000000100010110011101011;
assign LUT_3[30516] = 32'b00000000000000010111001110100000;
assign LUT_3[30517] = 32'b00000000000000011101111001111101;
assign LUT_3[30518] = 32'b00000000000000011001010110000100;
assign LUT_3[30519] = 32'b00000000000000100000000001100001;
assign LUT_3[30520] = 32'b00000000000000011111011001110000;
assign LUT_3[30521] = 32'b00000000000000100110000101001101;
assign LUT_3[30522] = 32'b00000000000000100001100001010100;
assign LUT_3[30523] = 32'b00000000000000101000001100110001;
assign LUT_3[30524] = 32'b00000000000000011100100111100110;
assign LUT_3[30525] = 32'b00000000000000100011010011000011;
assign LUT_3[30526] = 32'b00000000000000011110101111001010;
assign LUT_3[30527] = 32'b00000000000000100101011010100111;
assign LUT_3[30528] = 32'b00000000000000010101010111110010;
assign LUT_3[30529] = 32'b00000000000000011100000011001111;
assign LUT_3[30530] = 32'b00000000000000010111011111010110;
assign LUT_3[30531] = 32'b00000000000000011110001010110011;
assign LUT_3[30532] = 32'b00000000000000010010100101101000;
assign LUT_3[30533] = 32'b00000000000000011001010001000101;
assign LUT_3[30534] = 32'b00000000000000010100101101001100;
assign LUT_3[30535] = 32'b00000000000000011011011000101001;
assign LUT_3[30536] = 32'b00000000000000011010110000111000;
assign LUT_3[30537] = 32'b00000000000000100001011100010101;
assign LUT_3[30538] = 32'b00000000000000011100111000011100;
assign LUT_3[30539] = 32'b00000000000000100011100011111001;
assign LUT_3[30540] = 32'b00000000000000010111111110101110;
assign LUT_3[30541] = 32'b00000000000000011110101010001011;
assign LUT_3[30542] = 32'b00000000000000011010000110010010;
assign LUT_3[30543] = 32'b00000000000000100000110001101111;
assign LUT_3[30544] = 32'b00000000000000011000101010110101;
assign LUT_3[30545] = 32'b00000000000000011111010110010010;
assign LUT_3[30546] = 32'b00000000000000011010110010011001;
assign LUT_3[30547] = 32'b00000000000000100001011101110110;
assign LUT_3[30548] = 32'b00000000000000010101111000101011;
assign LUT_3[30549] = 32'b00000000000000011100100100001000;
assign LUT_3[30550] = 32'b00000000000000011000000000001111;
assign LUT_3[30551] = 32'b00000000000000011110101011101100;
assign LUT_3[30552] = 32'b00000000000000011110000011111011;
assign LUT_3[30553] = 32'b00000000000000100100101111011000;
assign LUT_3[30554] = 32'b00000000000000100000001011011111;
assign LUT_3[30555] = 32'b00000000000000100110110110111100;
assign LUT_3[30556] = 32'b00000000000000011011010001110001;
assign LUT_3[30557] = 32'b00000000000000100001111101001110;
assign LUT_3[30558] = 32'b00000000000000011101011001010101;
assign LUT_3[30559] = 32'b00000000000000100100000100110010;
assign LUT_3[30560] = 32'b00000000000000010110100110010010;
assign LUT_3[30561] = 32'b00000000000000011101010001101111;
assign LUT_3[30562] = 32'b00000000000000011000101101110110;
assign LUT_3[30563] = 32'b00000000000000011111011001010011;
assign LUT_3[30564] = 32'b00000000000000010011110100001000;
assign LUT_3[30565] = 32'b00000000000000011010011111100101;
assign LUT_3[30566] = 32'b00000000000000010101111011101100;
assign LUT_3[30567] = 32'b00000000000000011100100111001001;
assign LUT_3[30568] = 32'b00000000000000011011111111011000;
assign LUT_3[30569] = 32'b00000000000000100010101010110101;
assign LUT_3[30570] = 32'b00000000000000011110000110111100;
assign LUT_3[30571] = 32'b00000000000000100100110010011001;
assign LUT_3[30572] = 32'b00000000000000011001001101001110;
assign LUT_3[30573] = 32'b00000000000000011111111000101011;
assign LUT_3[30574] = 32'b00000000000000011011010100110010;
assign LUT_3[30575] = 32'b00000000000000100010000000001111;
assign LUT_3[30576] = 32'b00000000000000011001111001010101;
assign LUT_3[30577] = 32'b00000000000000100000100100110010;
assign LUT_3[30578] = 32'b00000000000000011100000000111001;
assign LUT_3[30579] = 32'b00000000000000100010101100010110;
assign LUT_3[30580] = 32'b00000000000000010111000111001011;
assign LUT_3[30581] = 32'b00000000000000011101110010101000;
assign LUT_3[30582] = 32'b00000000000000011001001110101111;
assign LUT_3[30583] = 32'b00000000000000011111111010001100;
assign LUT_3[30584] = 32'b00000000000000011111010010011011;
assign LUT_3[30585] = 32'b00000000000000100101111101111000;
assign LUT_3[30586] = 32'b00000000000000100001011001111111;
assign LUT_3[30587] = 32'b00000000000000101000000101011100;
assign LUT_3[30588] = 32'b00000000000000011100100000010001;
assign LUT_3[30589] = 32'b00000000000000100011001011101110;
assign LUT_3[30590] = 32'b00000000000000011110100111110101;
assign LUT_3[30591] = 32'b00000000000000100101010011010010;
assign LUT_3[30592] = 32'b00000000000000010111101010000101;
assign LUT_3[30593] = 32'b00000000000000011110010101100010;
assign LUT_3[30594] = 32'b00000000000000011001110001101001;
assign LUT_3[30595] = 32'b00000000000000100000011101000110;
assign LUT_3[30596] = 32'b00000000000000010100110111111011;
assign LUT_3[30597] = 32'b00000000000000011011100011011000;
assign LUT_3[30598] = 32'b00000000000000010110111111011111;
assign LUT_3[30599] = 32'b00000000000000011101101010111100;
assign LUT_3[30600] = 32'b00000000000000011101000011001011;
assign LUT_3[30601] = 32'b00000000000000100011101110101000;
assign LUT_3[30602] = 32'b00000000000000011111001010101111;
assign LUT_3[30603] = 32'b00000000000000100101110110001100;
assign LUT_3[30604] = 32'b00000000000000011010010001000001;
assign LUT_3[30605] = 32'b00000000000000100000111100011110;
assign LUT_3[30606] = 32'b00000000000000011100011000100101;
assign LUT_3[30607] = 32'b00000000000000100011000100000010;
assign LUT_3[30608] = 32'b00000000000000011010111101001000;
assign LUT_3[30609] = 32'b00000000000000100001101000100101;
assign LUT_3[30610] = 32'b00000000000000011101000100101100;
assign LUT_3[30611] = 32'b00000000000000100011110000001001;
assign LUT_3[30612] = 32'b00000000000000011000001010111110;
assign LUT_3[30613] = 32'b00000000000000011110110110011011;
assign LUT_3[30614] = 32'b00000000000000011010010010100010;
assign LUT_3[30615] = 32'b00000000000000100000111101111111;
assign LUT_3[30616] = 32'b00000000000000100000010110001110;
assign LUT_3[30617] = 32'b00000000000000100111000001101011;
assign LUT_3[30618] = 32'b00000000000000100010011101110010;
assign LUT_3[30619] = 32'b00000000000000101001001001001111;
assign LUT_3[30620] = 32'b00000000000000011101100100000100;
assign LUT_3[30621] = 32'b00000000000000100100001111100001;
assign LUT_3[30622] = 32'b00000000000000011111101011101000;
assign LUT_3[30623] = 32'b00000000000000100110010111000101;
assign LUT_3[30624] = 32'b00000000000000011000111000100101;
assign LUT_3[30625] = 32'b00000000000000011111100100000010;
assign LUT_3[30626] = 32'b00000000000000011011000000001001;
assign LUT_3[30627] = 32'b00000000000000100001101011100110;
assign LUT_3[30628] = 32'b00000000000000010110000110011011;
assign LUT_3[30629] = 32'b00000000000000011100110001111000;
assign LUT_3[30630] = 32'b00000000000000011000001101111111;
assign LUT_3[30631] = 32'b00000000000000011110111001011100;
assign LUT_3[30632] = 32'b00000000000000011110010001101011;
assign LUT_3[30633] = 32'b00000000000000100100111101001000;
assign LUT_3[30634] = 32'b00000000000000100000011001001111;
assign LUT_3[30635] = 32'b00000000000000100111000100101100;
assign LUT_3[30636] = 32'b00000000000000011011011111100001;
assign LUT_3[30637] = 32'b00000000000000100010001010111110;
assign LUT_3[30638] = 32'b00000000000000011101100111000101;
assign LUT_3[30639] = 32'b00000000000000100100010010100010;
assign LUT_3[30640] = 32'b00000000000000011100001011101000;
assign LUT_3[30641] = 32'b00000000000000100010110111000101;
assign LUT_3[30642] = 32'b00000000000000011110010011001100;
assign LUT_3[30643] = 32'b00000000000000100100111110101001;
assign LUT_3[30644] = 32'b00000000000000011001011001011110;
assign LUT_3[30645] = 32'b00000000000000100000000100111011;
assign LUT_3[30646] = 32'b00000000000000011011100001000010;
assign LUT_3[30647] = 32'b00000000000000100010001100011111;
assign LUT_3[30648] = 32'b00000000000000100001100100101110;
assign LUT_3[30649] = 32'b00000000000000101000010000001011;
assign LUT_3[30650] = 32'b00000000000000100011101100010010;
assign LUT_3[30651] = 32'b00000000000000101010010111101111;
assign LUT_3[30652] = 32'b00000000000000011110110010100100;
assign LUT_3[30653] = 32'b00000000000000100101011110000001;
assign LUT_3[30654] = 32'b00000000000000100000111010001000;
assign LUT_3[30655] = 32'b00000000000000100111100101100101;
assign LUT_3[30656] = 32'b00000000000000010111100010110000;
assign LUT_3[30657] = 32'b00000000000000011110001110001101;
assign LUT_3[30658] = 32'b00000000000000011001101010010100;
assign LUT_3[30659] = 32'b00000000000000100000010101110001;
assign LUT_3[30660] = 32'b00000000000000010100110000100110;
assign LUT_3[30661] = 32'b00000000000000011011011100000011;
assign LUT_3[30662] = 32'b00000000000000010110111000001010;
assign LUT_3[30663] = 32'b00000000000000011101100011100111;
assign LUT_3[30664] = 32'b00000000000000011100111011110110;
assign LUT_3[30665] = 32'b00000000000000100011100111010011;
assign LUT_3[30666] = 32'b00000000000000011111000011011010;
assign LUT_3[30667] = 32'b00000000000000100101101110110111;
assign LUT_3[30668] = 32'b00000000000000011010001001101100;
assign LUT_3[30669] = 32'b00000000000000100000110101001001;
assign LUT_3[30670] = 32'b00000000000000011100010001010000;
assign LUT_3[30671] = 32'b00000000000000100010111100101101;
assign LUT_3[30672] = 32'b00000000000000011010110101110011;
assign LUT_3[30673] = 32'b00000000000000100001100001010000;
assign LUT_3[30674] = 32'b00000000000000011100111101010111;
assign LUT_3[30675] = 32'b00000000000000100011101000110100;
assign LUT_3[30676] = 32'b00000000000000011000000011101001;
assign LUT_3[30677] = 32'b00000000000000011110101111000110;
assign LUT_3[30678] = 32'b00000000000000011010001011001101;
assign LUT_3[30679] = 32'b00000000000000100000110110101010;
assign LUT_3[30680] = 32'b00000000000000100000001110111001;
assign LUT_3[30681] = 32'b00000000000000100110111010010110;
assign LUT_3[30682] = 32'b00000000000000100010010110011101;
assign LUT_3[30683] = 32'b00000000000000101001000001111010;
assign LUT_3[30684] = 32'b00000000000000011101011100101111;
assign LUT_3[30685] = 32'b00000000000000100100001000001100;
assign LUT_3[30686] = 32'b00000000000000011111100100010011;
assign LUT_3[30687] = 32'b00000000000000100110001111110000;
assign LUT_3[30688] = 32'b00000000000000011000110001010000;
assign LUT_3[30689] = 32'b00000000000000011111011100101101;
assign LUT_3[30690] = 32'b00000000000000011010111000110100;
assign LUT_3[30691] = 32'b00000000000000100001100100010001;
assign LUT_3[30692] = 32'b00000000000000010101111111000110;
assign LUT_3[30693] = 32'b00000000000000011100101010100011;
assign LUT_3[30694] = 32'b00000000000000011000000110101010;
assign LUT_3[30695] = 32'b00000000000000011110110010000111;
assign LUT_3[30696] = 32'b00000000000000011110001010010110;
assign LUT_3[30697] = 32'b00000000000000100100110101110011;
assign LUT_3[30698] = 32'b00000000000000100000010001111010;
assign LUT_3[30699] = 32'b00000000000000100110111101010111;
assign LUT_3[30700] = 32'b00000000000000011011011000001100;
assign LUT_3[30701] = 32'b00000000000000100010000011101001;
assign LUT_3[30702] = 32'b00000000000000011101011111110000;
assign LUT_3[30703] = 32'b00000000000000100100001011001101;
assign LUT_3[30704] = 32'b00000000000000011100000100010011;
assign LUT_3[30705] = 32'b00000000000000100010101111110000;
assign LUT_3[30706] = 32'b00000000000000011110001011110111;
assign LUT_3[30707] = 32'b00000000000000100100110111010100;
assign LUT_3[30708] = 32'b00000000000000011001010010001001;
assign LUT_3[30709] = 32'b00000000000000011111111101100110;
assign LUT_3[30710] = 32'b00000000000000011011011001101101;
assign LUT_3[30711] = 32'b00000000000000100010000101001010;
assign LUT_3[30712] = 32'b00000000000000100001011101011001;
assign LUT_3[30713] = 32'b00000000000000101000001000110110;
assign LUT_3[30714] = 32'b00000000000000100011100100111101;
assign LUT_3[30715] = 32'b00000000000000101010010000011010;
assign LUT_3[30716] = 32'b00000000000000011110101011001111;
assign LUT_3[30717] = 32'b00000000000000100101010110101100;
assign LUT_3[30718] = 32'b00000000000000100000110010110011;
assign LUT_3[30719] = 32'b00000000000000100111011110010000;
assign LUT_3[30720] = 32'b00000000000000010001001011101011;
assign LUT_3[30721] = 32'b00000000000000010111110111001000;
assign LUT_3[30722] = 32'b00000000000000010011010011001111;
assign LUT_3[30723] = 32'b00000000000000011001111110101100;
assign LUT_3[30724] = 32'b00000000000000001110011001100001;
assign LUT_3[30725] = 32'b00000000000000010101000100111110;
assign LUT_3[30726] = 32'b00000000000000010000100001000101;
assign LUT_3[30727] = 32'b00000000000000010111001100100010;
assign LUT_3[30728] = 32'b00000000000000010110100100110001;
assign LUT_3[30729] = 32'b00000000000000011101010000001110;
assign LUT_3[30730] = 32'b00000000000000011000101100010101;
assign LUT_3[30731] = 32'b00000000000000011111010111110010;
assign LUT_3[30732] = 32'b00000000000000010011110010100111;
assign LUT_3[30733] = 32'b00000000000000011010011110000100;
assign LUT_3[30734] = 32'b00000000000000010101111010001011;
assign LUT_3[30735] = 32'b00000000000000011100100101101000;
assign LUT_3[30736] = 32'b00000000000000010100011110101110;
assign LUT_3[30737] = 32'b00000000000000011011001010001011;
assign LUT_3[30738] = 32'b00000000000000010110100110010010;
assign LUT_3[30739] = 32'b00000000000000011101010001101111;
assign LUT_3[30740] = 32'b00000000000000010001101100100100;
assign LUT_3[30741] = 32'b00000000000000011000011000000001;
assign LUT_3[30742] = 32'b00000000000000010011110100001000;
assign LUT_3[30743] = 32'b00000000000000011010011111100101;
assign LUT_3[30744] = 32'b00000000000000011001110111110100;
assign LUT_3[30745] = 32'b00000000000000100000100011010001;
assign LUT_3[30746] = 32'b00000000000000011011111111011000;
assign LUT_3[30747] = 32'b00000000000000100010101010110101;
assign LUT_3[30748] = 32'b00000000000000010111000101101010;
assign LUT_3[30749] = 32'b00000000000000011101110001000111;
assign LUT_3[30750] = 32'b00000000000000011001001101001110;
assign LUT_3[30751] = 32'b00000000000000011111111000101011;
assign LUT_3[30752] = 32'b00000000000000010010011010001011;
assign LUT_3[30753] = 32'b00000000000000011001000101101000;
assign LUT_3[30754] = 32'b00000000000000010100100001101111;
assign LUT_3[30755] = 32'b00000000000000011011001101001100;
assign LUT_3[30756] = 32'b00000000000000001111101000000001;
assign LUT_3[30757] = 32'b00000000000000010110010011011110;
assign LUT_3[30758] = 32'b00000000000000010001101111100101;
assign LUT_3[30759] = 32'b00000000000000011000011011000010;
assign LUT_3[30760] = 32'b00000000000000010111110011010001;
assign LUT_3[30761] = 32'b00000000000000011110011110101110;
assign LUT_3[30762] = 32'b00000000000000011001111010110101;
assign LUT_3[30763] = 32'b00000000000000100000100110010010;
assign LUT_3[30764] = 32'b00000000000000010101000001000111;
assign LUT_3[30765] = 32'b00000000000000011011101100100100;
assign LUT_3[30766] = 32'b00000000000000010111001000101011;
assign LUT_3[30767] = 32'b00000000000000011101110100001000;
assign LUT_3[30768] = 32'b00000000000000010101101101001110;
assign LUT_3[30769] = 32'b00000000000000011100011000101011;
assign LUT_3[30770] = 32'b00000000000000010111110100110010;
assign LUT_3[30771] = 32'b00000000000000011110100000001111;
assign LUT_3[30772] = 32'b00000000000000010010111011000100;
assign LUT_3[30773] = 32'b00000000000000011001100110100001;
assign LUT_3[30774] = 32'b00000000000000010101000010101000;
assign LUT_3[30775] = 32'b00000000000000011011101110000101;
assign LUT_3[30776] = 32'b00000000000000011011000110010100;
assign LUT_3[30777] = 32'b00000000000000100001110001110001;
assign LUT_3[30778] = 32'b00000000000000011101001101111000;
assign LUT_3[30779] = 32'b00000000000000100011111001010101;
assign LUT_3[30780] = 32'b00000000000000011000010100001010;
assign LUT_3[30781] = 32'b00000000000000011110111111100111;
assign LUT_3[30782] = 32'b00000000000000011010011011101110;
assign LUT_3[30783] = 32'b00000000000000100001000111001011;
assign LUT_3[30784] = 32'b00000000000000010001000100010110;
assign LUT_3[30785] = 32'b00000000000000010111101111110011;
assign LUT_3[30786] = 32'b00000000000000010011001011111010;
assign LUT_3[30787] = 32'b00000000000000011001110111010111;
assign LUT_3[30788] = 32'b00000000000000001110010010001100;
assign LUT_3[30789] = 32'b00000000000000010100111101101001;
assign LUT_3[30790] = 32'b00000000000000010000011001110000;
assign LUT_3[30791] = 32'b00000000000000010111000101001101;
assign LUT_3[30792] = 32'b00000000000000010110011101011100;
assign LUT_3[30793] = 32'b00000000000000011101001000111001;
assign LUT_3[30794] = 32'b00000000000000011000100101000000;
assign LUT_3[30795] = 32'b00000000000000011111010000011101;
assign LUT_3[30796] = 32'b00000000000000010011101011010010;
assign LUT_3[30797] = 32'b00000000000000011010010110101111;
assign LUT_3[30798] = 32'b00000000000000010101110010110110;
assign LUT_3[30799] = 32'b00000000000000011100011110010011;
assign LUT_3[30800] = 32'b00000000000000010100010111011001;
assign LUT_3[30801] = 32'b00000000000000011011000010110110;
assign LUT_3[30802] = 32'b00000000000000010110011110111101;
assign LUT_3[30803] = 32'b00000000000000011101001010011010;
assign LUT_3[30804] = 32'b00000000000000010001100101001111;
assign LUT_3[30805] = 32'b00000000000000011000010000101100;
assign LUT_3[30806] = 32'b00000000000000010011101100110011;
assign LUT_3[30807] = 32'b00000000000000011010011000010000;
assign LUT_3[30808] = 32'b00000000000000011001110000011111;
assign LUT_3[30809] = 32'b00000000000000100000011011111100;
assign LUT_3[30810] = 32'b00000000000000011011111000000011;
assign LUT_3[30811] = 32'b00000000000000100010100011100000;
assign LUT_3[30812] = 32'b00000000000000010110111110010101;
assign LUT_3[30813] = 32'b00000000000000011101101001110010;
assign LUT_3[30814] = 32'b00000000000000011001000101111001;
assign LUT_3[30815] = 32'b00000000000000011111110001010110;
assign LUT_3[30816] = 32'b00000000000000010010010010110110;
assign LUT_3[30817] = 32'b00000000000000011000111110010011;
assign LUT_3[30818] = 32'b00000000000000010100011010011010;
assign LUT_3[30819] = 32'b00000000000000011011000101110111;
assign LUT_3[30820] = 32'b00000000000000001111100000101100;
assign LUT_3[30821] = 32'b00000000000000010110001100001001;
assign LUT_3[30822] = 32'b00000000000000010001101000010000;
assign LUT_3[30823] = 32'b00000000000000011000010011101101;
assign LUT_3[30824] = 32'b00000000000000010111101011111100;
assign LUT_3[30825] = 32'b00000000000000011110010111011001;
assign LUT_3[30826] = 32'b00000000000000011001110011100000;
assign LUT_3[30827] = 32'b00000000000000100000011110111101;
assign LUT_3[30828] = 32'b00000000000000010100111001110010;
assign LUT_3[30829] = 32'b00000000000000011011100101001111;
assign LUT_3[30830] = 32'b00000000000000010111000001010110;
assign LUT_3[30831] = 32'b00000000000000011101101100110011;
assign LUT_3[30832] = 32'b00000000000000010101100101111001;
assign LUT_3[30833] = 32'b00000000000000011100010001010110;
assign LUT_3[30834] = 32'b00000000000000010111101101011101;
assign LUT_3[30835] = 32'b00000000000000011110011000111010;
assign LUT_3[30836] = 32'b00000000000000010010110011101111;
assign LUT_3[30837] = 32'b00000000000000011001011111001100;
assign LUT_3[30838] = 32'b00000000000000010100111011010011;
assign LUT_3[30839] = 32'b00000000000000011011100110110000;
assign LUT_3[30840] = 32'b00000000000000011010111110111111;
assign LUT_3[30841] = 32'b00000000000000100001101010011100;
assign LUT_3[30842] = 32'b00000000000000011101000110100011;
assign LUT_3[30843] = 32'b00000000000000100011110010000000;
assign LUT_3[30844] = 32'b00000000000000011000001100110101;
assign LUT_3[30845] = 32'b00000000000000011110111000010010;
assign LUT_3[30846] = 32'b00000000000000011010010100011001;
assign LUT_3[30847] = 32'b00000000000000100000111111110110;
assign LUT_3[30848] = 32'b00000000000000010011010110101001;
assign LUT_3[30849] = 32'b00000000000000011010000010000110;
assign LUT_3[30850] = 32'b00000000000000010101011110001101;
assign LUT_3[30851] = 32'b00000000000000011100001001101010;
assign LUT_3[30852] = 32'b00000000000000010000100100011111;
assign LUT_3[30853] = 32'b00000000000000010111001111111100;
assign LUT_3[30854] = 32'b00000000000000010010101100000011;
assign LUT_3[30855] = 32'b00000000000000011001010111100000;
assign LUT_3[30856] = 32'b00000000000000011000101111101111;
assign LUT_3[30857] = 32'b00000000000000011111011011001100;
assign LUT_3[30858] = 32'b00000000000000011010110111010011;
assign LUT_3[30859] = 32'b00000000000000100001100010110000;
assign LUT_3[30860] = 32'b00000000000000010101111101100101;
assign LUT_3[30861] = 32'b00000000000000011100101001000010;
assign LUT_3[30862] = 32'b00000000000000011000000101001001;
assign LUT_3[30863] = 32'b00000000000000011110110000100110;
assign LUT_3[30864] = 32'b00000000000000010110101001101100;
assign LUT_3[30865] = 32'b00000000000000011101010101001001;
assign LUT_3[30866] = 32'b00000000000000011000110001010000;
assign LUT_3[30867] = 32'b00000000000000011111011100101101;
assign LUT_3[30868] = 32'b00000000000000010011110111100010;
assign LUT_3[30869] = 32'b00000000000000011010100010111111;
assign LUT_3[30870] = 32'b00000000000000010101111111000110;
assign LUT_3[30871] = 32'b00000000000000011100101010100011;
assign LUT_3[30872] = 32'b00000000000000011100000010110010;
assign LUT_3[30873] = 32'b00000000000000100010101110001111;
assign LUT_3[30874] = 32'b00000000000000011110001010010110;
assign LUT_3[30875] = 32'b00000000000000100100110101110011;
assign LUT_3[30876] = 32'b00000000000000011001010000101000;
assign LUT_3[30877] = 32'b00000000000000011111111100000101;
assign LUT_3[30878] = 32'b00000000000000011011011000001100;
assign LUT_3[30879] = 32'b00000000000000100010000011101001;
assign LUT_3[30880] = 32'b00000000000000010100100101001001;
assign LUT_3[30881] = 32'b00000000000000011011010000100110;
assign LUT_3[30882] = 32'b00000000000000010110101100101101;
assign LUT_3[30883] = 32'b00000000000000011101011000001010;
assign LUT_3[30884] = 32'b00000000000000010001110010111111;
assign LUT_3[30885] = 32'b00000000000000011000011110011100;
assign LUT_3[30886] = 32'b00000000000000010011111010100011;
assign LUT_3[30887] = 32'b00000000000000011010100110000000;
assign LUT_3[30888] = 32'b00000000000000011001111110001111;
assign LUT_3[30889] = 32'b00000000000000100000101001101100;
assign LUT_3[30890] = 32'b00000000000000011100000101110011;
assign LUT_3[30891] = 32'b00000000000000100010110001010000;
assign LUT_3[30892] = 32'b00000000000000010111001100000101;
assign LUT_3[30893] = 32'b00000000000000011101110111100010;
assign LUT_3[30894] = 32'b00000000000000011001010011101001;
assign LUT_3[30895] = 32'b00000000000000011111111111000110;
assign LUT_3[30896] = 32'b00000000000000010111111000001100;
assign LUT_3[30897] = 32'b00000000000000011110100011101001;
assign LUT_3[30898] = 32'b00000000000000011001111111110000;
assign LUT_3[30899] = 32'b00000000000000100000101011001101;
assign LUT_3[30900] = 32'b00000000000000010101000110000010;
assign LUT_3[30901] = 32'b00000000000000011011110001011111;
assign LUT_3[30902] = 32'b00000000000000010111001101100110;
assign LUT_3[30903] = 32'b00000000000000011101111001000011;
assign LUT_3[30904] = 32'b00000000000000011101010001010010;
assign LUT_3[30905] = 32'b00000000000000100011111100101111;
assign LUT_3[30906] = 32'b00000000000000011111011000110110;
assign LUT_3[30907] = 32'b00000000000000100110000100010011;
assign LUT_3[30908] = 32'b00000000000000011010011111001000;
assign LUT_3[30909] = 32'b00000000000000100001001010100101;
assign LUT_3[30910] = 32'b00000000000000011100100110101100;
assign LUT_3[30911] = 32'b00000000000000100011010010001001;
assign LUT_3[30912] = 32'b00000000000000010011001111010100;
assign LUT_3[30913] = 32'b00000000000000011001111010110001;
assign LUT_3[30914] = 32'b00000000000000010101010110111000;
assign LUT_3[30915] = 32'b00000000000000011100000010010101;
assign LUT_3[30916] = 32'b00000000000000010000011101001010;
assign LUT_3[30917] = 32'b00000000000000010111001000100111;
assign LUT_3[30918] = 32'b00000000000000010010100100101110;
assign LUT_3[30919] = 32'b00000000000000011001010000001011;
assign LUT_3[30920] = 32'b00000000000000011000101000011010;
assign LUT_3[30921] = 32'b00000000000000011111010011110111;
assign LUT_3[30922] = 32'b00000000000000011010101111111110;
assign LUT_3[30923] = 32'b00000000000000100001011011011011;
assign LUT_3[30924] = 32'b00000000000000010101110110010000;
assign LUT_3[30925] = 32'b00000000000000011100100001101101;
assign LUT_3[30926] = 32'b00000000000000010111111101110100;
assign LUT_3[30927] = 32'b00000000000000011110101001010001;
assign LUT_3[30928] = 32'b00000000000000010110100010010111;
assign LUT_3[30929] = 32'b00000000000000011101001101110100;
assign LUT_3[30930] = 32'b00000000000000011000101001111011;
assign LUT_3[30931] = 32'b00000000000000011111010101011000;
assign LUT_3[30932] = 32'b00000000000000010011110000001101;
assign LUT_3[30933] = 32'b00000000000000011010011011101010;
assign LUT_3[30934] = 32'b00000000000000010101110111110001;
assign LUT_3[30935] = 32'b00000000000000011100100011001110;
assign LUT_3[30936] = 32'b00000000000000011011111011011101;
assign LUT_3[30937] = 32'b00000000000000100010100110111010;
assign LUT_3[30938] = 32'b00000000000000011110000011000001;
assign LUT_3[30939] = 32'b00000000000000100100101110011110;
assign LUT_3[30940] = 32'b00000000000000011001001001010011;
assign LUT_3[30941] = 32'b00000000000000011111110100110000;
assign LUT_3[30942] = 32'b00000000000000011011010000110111;
assign LUT_3[30943] = 32'b00000000000000100001111100010100;
assign LUT_3[30944] = 32'b00000000000000010100011101110100;
assign LUT_3[30945] = 32'b00000000000000011011001001010001;
assign LUT_3[30946] = 32'b00000000000000010110100101011000;
assign LUT_3[30947] = 32'b00000000000000011101010000110101;
assign LUT_3[30948] = 32'b00000000000000010001101011101010;
assign LUT_3[30949] = 32'b00000000000000011000010111000111;
assign LUT_3[30950] = 32'b00000000000000010011110011001110;
assign LUT_3[30951] = 32'b00000000000000011010011110101011;
assign LUT_3[30952] = 32'b00000000000000011001110110111010;
assign LUT_3[30953] = 32'b00000000000000100000100010010111;
assign LUT_3[30954] = 32'b00000000000000011011111110011110;
assign LUT_3[30955] = 32'b00000000000000100010101001111011;
assign LUT_3[30956] = 32'b00000000000000010111000100110000;
assign LUT_3[30957] = 32'b00000000000000011101110000001101;
assign LUT_3[30958] = 32'b00000000000000011001001100010100;
assign LUT_3[30959] = 32'b00000000000000011111110111110001;
assign LUT_3[30960] = 32'b00000000000000010111110000110111;
assign LUT_3[30961] = 32'b00000000000000011110011100010100;
assign LUT_3[30962] = 32'b00000000000000011001111000011011;
assign LUT_3[30963] = 32'b00000000000000100000100011111000;
assign LUT_3[30964] = 32'b00000000000000010100111110101101;
assign LUT_3[30965] = 32'b00000000000000011011101010001010;
assign LUT_3[30966] = 32'b00000000000000010111000110010001;
assign LUT_3[30967] = 32'b00000000000000011101110001101110;
assign LUT_3[30968] = 32'b00000000000000011101001001111101;
assign LUT_3[30969] = 32'b00000000000000100011110101011010;
assign LUT_3[30970] = 32'b00000000000000011111010001100001;
assign LUT_3[30971] = 32'b00000000000000100101111100111110;
assign LUT_3[30972] = 32'b00000000000000011010010111110011;
assign LUT_3[30973] = 32'b00000000000000100001000011010000;
assign LUT_3[30974] = 32'b00000000000000011100011111010111;
assign LUT_3[30975] = 32'b00000000000000100011001010110100;
assign LUT_3[30976] = 32'b00000000000000001101011011001100;
assign LUT_3[30977] = 32'b00000000000000010100000110101001;
assign LUT_3[30978] = 32'b00000000000000001111100010110000;
assign LUT_3[30979] = 32'b00000000000000010110001110001101;
assign LUT_3[30980] = 32'b00000000000000001010101001000010;
assign LUT_3[30981] = 32'b00000000000000010001010100011111;
assign LUT_3[30982] = 32'b00000000000000001100110000100110;
assign LUT_3[30983] = 32'b00000000000000010011011100000011;
assign LUT_3[30984] = 32'b00000000000000010010110100010010;
assign LUT_3[30985] = 32'b00000000000000011001011111101111;
assign LUT_3[30986] = 32'b00000000000000010100111011110110;
assign LUT_3[30987] = 32'b00000000000000011011100111010011;
assign LUT_3[30988] = 32'b00000000000000010000000010001000;
assign LUT_3[30989] = 32'b00000000000000010110101101100101;
assign LUT_3[30990] = 32'b00000000000000010010001001101100;
assign LUT_3[30991] = 32'b00000000000000011000110101001001;
assign LUT_3[30992] = 32'b00000000000000010000101110001111;
assign LUT_3[30993] = 32'b00000000000000010111011001101100;
assign LUT_3[30994] = 32'b00000000000000010010110101110011;
assign LUT_3[30995] = 32'b00000000000000011001100001010000;
assign LUT_3[30996] = 32'b00000000000000001101111100000101;
assign LUT_3[30997] = 32'b00000000000000010100100111100010;
assign LUT_3[30998] = 32'b00000000000000010000000011101001;
assign LUT_3[30999] = 32'b00000000000000010110101111000110;
assign LUT_3[31000] = 32'b00000000000000010110000111010101;
assign LUT_3[31001] = 32'b00000000000000011100110010110010;
assign LUT_3[31002] = 32'b00000000000000011000001110111001;
assign LUT_3[31003] = 32'b00000000000000011110111010010110;
assign LUT_3[31004] = 32'b00000000000000010011010101001011;
assign LUT_3[31005] = 32'b00000000000000011010000000101000;
assign LUT_3[31006] = 32'b00000000000000010101011100101111;
assign LUT_3[31007] = 32'b00000000000000011100001000001100;
assign LUT_3[31008] = 32'b00000000000000001110101001101100;
assign LUT_3[31009] = 32'b00000000000000010101010101001001;
assign LUT_3[31010] = 32'b00000000000000010000110001010000;
assign LUT_3[31011] = 32'b00000000000000010111011100101101;
assign LUT_3[31012] = 32'b00000000000000001011110111100010;
assign LUT_3[31013] = 32'b00000000000000010010100010111111;
assign LUT_3[31014] = 32'b00000000000000001101111111000110;
assign LUT_3[31015] = 32'b00000000000000010100101010100011;
assign LUT_3[31016] = 32'b00000000000000010100000010110010;
assign LUT_3[31017] = 32'b00000000000000011010101110001111;
assign LUT_3[31018] = 32'b00000000000000010110001010010110;
assign LUT_3[31019] = 32'b00000000000000011100110101110011;
assign LUT_3[31020] = 32'b00000000000000010001010000101000;
assign LUT_3[31021] = 32'b00000000000000010111111100000101;
assign LUT_3[31022] = 32'b00000000000000010011011000001100;
assign LUT_3[31023] = 32'b00000000000000011010000011101001;
assign LUT_3[31024] = 32'b00000000000000010001111100101111;
assign LUT_3[31025] = 32'b00000000000000011000101000001100;
assign LUT_3[31026] = 32'b00000000000000010100000100010011;
assign LUT_3[31027] = 32'b00000000000000011010101111110000;
assign LUT_3[31028] = 32'b00000000000000001111001010100101;
assign LUT_3[31029] = 32'b00000000000000010101110110000010;
assign LUT_3[31030] = 32'b00000000000000010001010010001001;
assign LUT_3[31031] = 32'b00000000000000010111111101100110;
assign LUT_3[31032] = 32'b00000000000000010111010101110101;
assign LUT_3[31033] = 32'b00000000000000011110000001010010;
assign LUT_3[31034] = 32'b00000000000000011001011101011001;
assign LUT_3[31035] = 32'b00000000000000100000001000110110;
assign LUT_3[31036] = 32'b00000000000000010100100011101011;
assign LUT_3[31037] = 32'b00000000000000011011001111001000;
assign LUT_3[31038] = 32'b00000000000000010110101011001111;
assign LUT_3[31039] = 32'b00000000000000011101010110101100;
assign LUT_3[31040] = 32'b00000000000000001101010011110111;
assign LUT_3[31041] = 32'b00000000000000010011111111010100;
assign LUT_3[31042] = 32'b00000000000000001111011011011011;
assign LUT_3[31043] = 32'b00000000000000010110000110111000;
assign LUT_3[31044] = 32'b00000000000000001010100001101101;
assign LUT_3[31045] = 32'b00000000000000010001001101001010;
assign LUT_3[31046] = 32'b00000000000000001100101001010001;
assign LUT_3[31047] = 32'b00000000000000010011010100101110;
assign LUT_3[31048] = 32'b00000000000000010010101100111101;
assign LUT_3[31049] = 32'b00000000000000011001011000011010;
assign LUT_3[31050] = 32'b00000000000000010100110100100001;
assign LUT_3[31051] = 32'b00000000000000011011011111111110;
assign LUT_3[31052] = 32'b00000000000000001111111010110011;
assign LUT_3[31053] = 32'b00000000000000010110100110010000;
assign LUT_3[31054] = 32'b00000000000000010010000010010111;
assign LUT_3[31055] = 32'b00000000000000011000101101110100;
assign LUT_3[31056] = 32'b00000000000000010000100110111010;
assign LUT_3[31057] = 32'b00000000000000010111010010010111;
assign LUT_3[31058] = 32'b00000000000000010010101110011110;
assign LUT_3[31059] = 32'b00000000000000011001011001111011;
assign LUT_3[31060] = 32'b00000000000000001101110100110000;
assign LUT_3[31061] = 32'b00000000000000010100100000001101;
assign LUT_3[31062] = 32'b00000000000000001111111100010100;
assign LUT_3[31063] = 32'b00000000000000010110100111110001;
assign LUT_3[31064] = 32'b00000000000000010110000000000000;
assign LUT_3[31065] = 32'b00000000000000011100101011011101;
assign LUT_3[31066] = 32'b00000000000000011000000111100100;
assign LUT_3[31067] = 32'b00000000000000011110110011000001;
assign LUT_3[31068] = 32'b00000000000000010011001101110110;
assign LUT_3[31069] = 32'b00000000000000011001111001010011;
assign LUT_3[31070] = 32'b00000000000000010101010101011010;
assign LUT_3[31071] = 32'b00000000000000011100000000110111;
assign LUT_3[31072] = 32'b00000000000000001110100010010111;
assign LUT_3[31073] = 32'b00000000000000010101001101110100;
assign LUT_3[31074] = 32'b00000000000000010000101001111011;
assign LUT_3[31075] = 32'b00000000000000010111010101011000;
assign LUT_3[31076] = 32'b00000000000000001011110000001101;
assign LUT_3[31077] = 32'b00000000000000010010011011101010;
assign LUT_3[31078] = 32'b00000000000000001101110111110001;
assign LUT_3[31079] = 32'b00000000000000010100100011001110;
assign LUT_3[31080] = 32'b00000000000000010011111011011101;
assign LUT_3[31081] = 32'b00000000000000011010100110111010;
assign LUT_3[31082] = 32'b00000000000000010110000011000001;
assign LUT_3[31083] = 32'b00000000000000011100101110011110;
assign LUT_3[31084] = 32'b00000000000000010001001001010011;
assign LUT_3[31085] = 32'b00000000000000010111110100110000;
assign LUT_3[31086] = 32'b00000000000000010011010000110111;
assign LUT_3[31087] = 32'b00000000000000011001111100010100;
assign LUT_3[31088] = 32'b00000000000000010001110101011010;
assign LUT_3[31089] = 32'b00000000000000011000100000110111;
assign LUT_3[31090] = 32'b00000000000000010011111100111110;
assign LUT_3[31091] = 32'b00000000000000011010101000011011;
assign LUT_3[31092] = 32'b00000000000000001111000011010000;
assign LUT_3[31093] = 32'b00000000000000010101101110101101;
assign LUT_3[31094] = 32'b00000000000000010001001010110100;
assign LUT_3[31095] = 32'b00000000000000010111110110010001;
assign LUT_3[31096] = 32'b00000000000000010111001110100000;
assign LUT_3[31097] = 32'b00000000000000011101111001111101;
assign LUT_3[31098] = 32'b00000000000000011001010110000100;
assign LUT_3[31099] = 32'b00000000000000100000000001100001;
assign LUT_3[31100] = 32'b00000000000000010100011100010110;
assign LUT_3[31101] = 32'b00000000000000011011000111110011;
assign LUT_3[31102] = 32'b00000000000000010110100011111010;
assign LUT_3[31103] = 32'b00000000000000011101001111010111;
assign LUT_3[31104] = 32'b00000000000000001111100110001010;
assign LUT_3[31105] = 32'b00000000000000010110010001100111;
assign LUT_3[31106] = 32'b00000000000000010001101101101110;
assign LUT_3[31107] = 32'b00000000000000011000011001001011;
assign LUT_3[31108] = 32'b00000000000000001100110100000000;
assign LUT_3[31109] = 32'b00000000000000010011011111011101;
assign LUT_3[31110] = 32'b00000000000000001110111011100100;
assign LUT_3[31111] = 32'b00000000000000010101100111000001;
assign LUT_3[31112] = 32'b00000000000000010100111111010000;
assign LUT_3[31113] = 32'b00000000000000011011101010101101;
assign LUT_3[31114] = 32'b00000000000000010111000110110100;
assign LUT_3[31115] = 32'b00000000000000011101110010010001;
assign LUT_3[31116] = 32'b00000000000000010010001101000110;
assign LUT_3[31117] = 32'b00000000000000011000111000100011;
assign LUT_3[31118] = 32'b00000000000000010100010100101010;
assign LUT_3[31119] = 32'b00000000000000011011000000000111;
assign LUT_3[31120] = 32'b00000000000000010010111001001101;
assign LUT_3[31121] = 32'b00000000000000011001100100101010;
assign LUT_3[31122] = 32'b00000000000000010101000000110001;
assign LUT_3[31123] = 32'b00000000000000011011101100001110;
assign LUT_3[31124] = 32'b00000000000000010000000111000011;
assign LUT_3[31125] = 32'b00000000000000010110110010100000;
assign LUT_3[31126] = 32'b00000000000000010010001110100111;
assign LUT_3[31127] = 32'b00000000000000011000111010000100;
assign LUT_3[31128] = 32'b00000000000000011000010010010011;
assign LUT_3[31129] = 32'b00000000000000011110111101110000;
assign LUT_3[31130] = 32'b00000000000000011010011001110111;
assign LUT_3[31131] = 32'b00000000000000100001000101010100;
assign LUT_3[31132] = 32'b00000000000000010101100000001001;
assign LUT_3[31133] = 32'b00000000000000011100001011100110;
assign LUT_3[31134] = 32'b00000000000000010111100111101101;
assign LUT_3[31135] = 32'b00000000000000011110010011001010;
assign LUT_3[31136] = 32'b00000000000000010000110100101010;
assign LUT_3[31137] = 32'b00000000000000010111100000000111;
assign LUT_3[31138] = 32'b00000000000000010010111100001110;
assign LUT_3[31139] = 32'b00000000000000011001100111101011;
assign LUT_3[31140] = 32'b00000000000000001110000010100000;
assign LUT_3[31141] = 32'b00000000000000010100101101111101;
assign LUT_3[31142] = 32'b00000000000000010000001010000100;
assign LUT_3[31143] = 32'b00000000000000010110110101100001;
assign LUT_3[31144] = 32'b00000000000000010110001101110000;
assign LUT_3[31145] = 32'b00000000000000011100111001001101;
assign LUT_3[31146] = 32'b00000000000000011000010101010100;
assign LUT_3[31147] = 32'b00000000000000011111000000110001;
assign LUT_3[31148] = 32'b00000000000000010011011011100110;
assign LUT_3[31149] = 32'b00000000000000011010000111000011;
assign LUT_3[31150] = 32'b00000000000000010101100011001010;
assign LUT_3[31151] = 32'b00000000000000011100001110100111;
assign LUT_3[31152] = 32'b00000000000000010100000111101101;
assign LUT_3[31153] = 32'b00000000000000011010110011001010;
assign LUT_3[31154] = 32'b00000000000000010110001111010001;
assign LUT_3[31155] = 32'b00000000000000011100111010101110;
assign LUT_3[31156] = 32'b00000000000000010001010101100011;
assign LUT_3[31157] = 32'b00000000000000011000000001000000;
assign LUT_3[31158] = 32'b00000000000000010011011101000111;
assign LUT_3[31159] = 32'b00000000000000011010001000100100;
assign LUT_3[31160] = 32'b00000000000000011001100000110011;
assign LUT_3[31161] = 32'b00000000000000100000001100010000;
assign LUT_3[31162] = 32'b00000000000000011011101000010111;
assign LUT_3[31163] = 32'b00000000000000100010010011110100;
assign LUT_3[31164] = 32'b00000000000000010110101110101001;
assign LUT_3[31165] = 32'b00000000000000011101011010000110;
assign LUT_3[31166] = 32'b00000000000000011000110110001101;
assign LUT_3[31167] = 32'b00000000000000011111100001101010;
assign LUT_3[31168] = 32'b00000000000000001111011110110101;
assign LUT_3[31169] = 32'b00000000000000010110001010010010;
assign LUT_3[31170] = 32'b00000000000000010001100110011001;
assign LUT_3[31171] = 32'b00000000000000011000010001110110;
assign LUT_3[31172] = 32'b00000000000000001100101100101011;
assign LUT_3[31173] = 32'b00000000000000010011011000001000;
assign LUT_3[31174] = 32'b00000000000000001110110100001111;
assign LUT_3[31175] = 32'b00000000000000010101011111101100;
assign LUT_3[31176] = 32'b00000000000000010100110111111011;
assign LUT_3[31177] = 32'b00000000000000011011100011011000;
assign LUT_3[31178] = 32'b00000000000000010110111111011111;
assign LUT_3[31179] = 32'b00000000000000011101101010111100;
assign LUT_3[31180] = 32'b00000000000000010010000101110001;
assign LUT_3[31181] = 32'b00000000000000011000110001001110;
assign LUT_3[31182] = 32'b00000000000000010100001101010101;
assign LUT_3[31183] = 32'b00000000000000011010111000110010;
assign LUT_3[31184] = 32'b00000000000000010010110001111000;
assign LUT_3[31185] = 32'b00000000000000011001011101010101;
assign LUT_3[31186] = 32'b00000000000000010100111001011100;
assign LUT_3[31187] = 32'b00000000000000011011100100111001;
assign LUT_3[31188] = 32'b00000000000000001111111111101110;
assign LUT_3[31189] = 32'b00000000000000010110101011001011;
assign LUT_3[31190] = 32'b00000000000000010010000111010010;
assign LUT_3[31191] = 32'b00000000000000011000110010101111;
assign LUT_3[31192] = 32'b00000000000000011000001010111110;
assign LUT_3[31193] = 32'b00000000000000011110110110011011;
assign LUT_3[31194] = 32'b00000000000000011010010010100010;
assign LUT_3[31195] = 32'b00000000000000100000111101111111;
assign LUT_3[31196] = 32'b00000000000000010101011000110100;
assign LUT_3[31197] = 32'b00000000000000011100000100010001;
assign LUT_3[31198] = 32'b00000000000000010111100000011000;
assign LUT_3[31199] = 32'b00000000000000011110001011110101;
assign LUT_3[31200] = 32'b00000000000000010000101101010101;
assign LUT_3[31201] = 32'b00000000000000010111011000110010;
assign LUT_3[31202] = 32'b00000000000000010010110100111001;
assign LUT_3[31203] = 32'b00000000000000011001100000010110;
assign LUT_3[31204] = 32'b00000000000000001101111011001011;
assign LUT_3[31205] = 32'b00000000000000010100100110101000;
assign LUT_3[31206] = 32'b00000000000000010000000010101111;
assign LUT_3[31207] = 32'b00000000000000010110101110001100;
assign LUT_3[31208] = 32'b00000000000000010110000110011011;
assign LUT_3[31209] = 32'b00000000000000011100110001111000;
assign LUT_3[31210] = 32'b00000000000000011000001101111111;
assign LUT_3[31211] = 32'b00000000000000011110111001011100;
assign LUT_3[31212] = 32'b00000000000000010011010100010001;
assign LUT_3[31213] = 32'b00000000000000011001111111101110;
assign LUT_3[31214] = 32'b00000000000000010101011011110101;
assign LUT_3[31215] = 32'b00000000000000011100000111010010;
assign LUT_3[31216] = 32'b00000000000000010100000000011000;
assign LUT_3[31217] = 32'b00000000000000011010101011110101;
assign LUT_3[31218] = 32'b00000000000000010110000111111100;
assign LUT_3[31219] = 32'b00000000000000011100110011011001;
assign LUT_3[31220] = 32'b00000000000000010001001110001110;
assign LUT_3[31221] = 32'b00000000000000010111111001101011;
assign LUT_3[31222] = 32'b00000000000000010011010101110010;
assign LUT_3[31223] = 32'b00000000000000011010000001001111;
assign LUT_3[31224] = 32'b00000000000000011001011001011110;
assign LUT_3[31225] = 32'b00000000000000100000000100111011;
assign LUT_3[31226] = 32'b00000000000000011011100001000010;
assign LUT_3[31227] = 32'b00000000000000100010001100011111;
assign LUT_3[31228] = 32'b00000000000000010110100111010100;
assign LUT_3[31229] = 32'b00000000000000011101010010110001;
assign LUT_3[31230] = 32'b00000000000000011000101110111000;
assign LUT_3[31231] = 32'b00000000000000011111011010010101;
assign LUT_3[31232] = 32'b00000000000000010100100000110111;
assign LUT_3[31233] = 32'b00000000000000011011001100010100;
assign LUT_3[31234] = 32'b00000000000000010110101000011011;
assign LUT_3[31235] = 32'b00000000000000011101010011111000;
assign LUT_3[31236] = 32'b00000000000000010001101110101101;
assign LUT_3[31237] = 32'b00000000000000011000011010001010;
assign LUT_3[31238] = 32'b00000000000000010011110110010001;
assign LUT_3[31239] = 32'b00000000000000011010100001101110;
assign LUT_3[31240] = 32'b00000000000000011001111001111101;
assign LUT_3[31241] = 32'b00000000000000100000100101011010;
assign LUT_3[31242] = 32'b00000000000000011100000001100001;
assign LUT_3[31243] = 32'b00000000000000100010101100111110;
assign LUT_3[31244] = 32'b00000000000000010111000111110011;
assign LUT_3[31245] = 32'b00000000000000011101110011010000;
assign LUT_3[31246] = 32'b00000000000000011001001111010111;
assign LUT_3[31247] = 32'b00000000000000011111111010110100;
assign LUT_3[31248] = 32'b00000000000000010111110011111010;
assign LUT_3[31249] = 32'b00000000000000011110011111010111;
assign LUT_3[31250] = 32'b00000000000000011001111011011110;
assign LUT_3[31251] = 32'b00000000000000100000100110111011;
assign LUT_3[31252] = 32'b00000000000000010101000001110000;
assign LUT_3[31253] = 32'b00000000000000011011101101001101;
assign LUT_3[31254] = 32'b00000000000000010111001001010100;
assign LUT_3[31255] = 32'b00000000000000011101110100110001;
assign LUT_3[31256] = 32'b00000000000000011101001101000000;
assign LUT_3[31257] = 32'b00000000000000100011111000011101;
assign LUT_3[31258] = 32'b00000000000000011111010100100100;
assign LUT_3[31259] = 32'b00000000000000100110000000000001;
assign LUT_3[31260] = 32'b00000000000000011010011010110110;
assign LUT_3[31261] = 32'b00000000000000100001000110010011;
assign LUT_3[31262] = 32'b00000000000000011100100010011010;
assign LUT_3[31263] = 32'b00000000000000100011001101110111;
assign LUT_3[31264] = 32'b00000000000000010101101111010111;
assign LUT_3[31265] = 32'b00000000000000011100011010110100;
assign LUT_3[31266] = 32'b00000000000000010111110110111011;
assign LUT_3[31267] = 32'b00000000000000011110100010011000;
assign LUT_3[31268] = 32'b00000000000000010010111101001101;
assign LUT_3[31269] = 32'b00000000000000011001101000101010;
assign LUT_3[31270] = 32'b00000000000000010101000100110001;
assign LUT_3[31271] = 32'b00000000000000011011110000001110;
assign LUT_3[31272] = 32'b00000000000000011011001000011101;
assign LUT_3[31273] = 32'b00000000000000100001110011111010;
assign LUT_3[31274] = 32'b00000000000000011101010000000001;
assign LUT_3[31275] = 32'b00000000000000100011111011011110;
assign LUT_3[31276] = 32'b00000000000000011000010110010011;
assign LUT_3[31277] = 32'b00000000000000011111000001110000;
assign LUT_3[31278] = 32'b00000000000000011010011101110111;
assign LUT_3[31279] = 32'b00000000000000100001001001010100;
assign LUT_3[31280] = 32'b00000000000000011001000010011010;
assign LUT_3[31281] = 32'b00000000000000011111101101110111;
assign LUT_3[31282] = 32'b00000000000000011011001001111110;
assign LUT_3[31283] = 32'b00000000000000100001110101011011;
assign LUT_3[31284] = 32'b00000000000000010110010000010000;
assign LUT_3[31285] = 32'b00000000000000011100111011101101;
assign LUT_3[31286] = 32'b00000000000000011000010111110100;
assign LUT_3[31287] = 32'b00000000000000011111000011010001;
assign LUT_3[31288] = 32'b00000000000000011110011011100000;
assign LUT_3[31289] = 32'b00000000000000100101000110111101;
assign LUT_3[31290] = 32'b00000000000000100000100011000100;
assign LUT_3[31291] = 32'b00000000000000100111001110100001;
assign LUT_3[31292] = 32'b00000000000000011011101001010110;
assign LUT_3[31293] = 32'b00000000000000100010010100110011;
assign LUT_3[31294] = 32'b00000000000000011101110000111010;
assign LUT_3[31295] = 32'b00000000000000100100011100010111;
assign LUT_3[31296] = 32'b00000000000000010100011001100010;
assign LUT_3[31297] = 32'b00000000000000011011000100111111;
assign LUT_3[31298] = 32'b00000000000000010110100001000110;
assign LUT_3[31299] = 32'b00000000000000011101001100100011;
assign LUT_3[31300] = 32'b00000000000000010001100111011000;
assign LUT_3[31301] = 32'b00000000000000011000010010110101;
assign LUT_3[31302] = 32'b00000000000000010011101110111100;
assign LUT_3[31303] = 32'b00000000000000011010011010011001;
assign LUT_3[31304] = 32'b00000000000000011001110010101000;
assign LUT_3[31305] = 32'b00000000000000100000011110000101;
assign LUT_3[31306] = 32'b00000000000000011011111010001100;
assign LUT_3[31307] = 32'b00000000000000100010100101101001;
assign LUT_3[31308] = 32'b00000000000000010111000000011110;
assign LUT_3[31309] = 32'b00000000000000011101101011111011;
assign LUT_3[31310] = 32'b00000000000000011001001000000010;
assign LUT_3[31311] = 32'b00000000000000011111110011011111;
assign LUT_3[31312] = 32'b00000000000000010111101100100101;
assign LUT_3[31313] = 32'b00000000000000011110011000000010;
assign LUT_3[31314] = 32'b00000000000000011001110100001001;
assign LUT_3[31315] = 32'b00000000000000100000011111100110;
assign LUT_3[31316] = 32'b00000000000000010100111010011011;
assign LUT_3[31317] = 32'b00000000000000011011100101111000;
assign LUT_3[31318] = 32'b00000000000000010111000001111111;
assign LUT_3[31319] = 32'b00000000000000011101101101011100;
assign LUT_3[31320] = 32'b00000000000000011101000101101011;
assign LUT_3[31321] = 32'b00000000000000100011110001001000;
assign LUT_3[31322] = 32'b00000000000000011111001101001111;
assign LUT_3[31323] = 32'b00000000000000100101111000101100;
assign LUT_3[31324] = 32'b00000000000000011010010011100001;
assign LUT_3[31325] = 32'b00000000000000100000111110111110;
assign LUT_3[31326] = 32'b00000000000000011100011011000101;
assign LUT_3[31327] = 32'b00000000000000100011000110100010;
assign LUT_3[31328] = 32'b00000000000000010101101000000010;
assign LUT_3[31329] = 32'b00000000000000011100010011011111;
assign LUT_3[31330] = 32'b00000000000000010111101111100110;
assign LUT_3[31331] = 32'b00000000000000011110011011000011;
assign LUT_3[31332] = 32'b00000000000000010010110101111000;
assign LUT_3[31333] = 32'b00000000000000011001100001010101;
assign LUT_3[31334] = 32'b00000000000000010100111101011100;
assign LUT_3[31335] = 32'b00000000000000011011101000111001;
assign LUT_3[31336] = 32'b00000000000000011011000001001000;
assign LUT_3[31337] = 32'b00000000000000100001101100100101;
assign LUT_3[31338] = 32'b00000000000000011101001000101100;
assign LUT_3[31339] = 32'b00000000000000100011110100001001;
assign LUT_3[31340] = 32'b00000000000000011000001110111110;
assign LUT_3[31341] = 32'b00000000000000011110111010011011;
assign LUT_3[31342] = 32'b00000000000000011010010110100010;
assign LUT_3[31343] = 32'b00000000000000100001000001111111;
assign LUT_3[31344] = 32'b00000000000000011000111011000101;
assign LUT_3[31345] = 32'b00000000000000011111100110100010;
assign LUT_3[31346] = 32'b00000000000000011011000010101001;
assign LUT_3[31347] = 32'b00000000000000100001101110000110;
assign LUT_3[31348] = 32'b00000000000000010110001000111011;
assign LUT_3[31349] = 32'b00000000000000011100110100011000;
assign LUT_3[31350] = 32'b00000000000000011000010000011111;
assign LUT_3[31351] = 32'b00000000000000011110111011111100;
assign LUT_3[31352] = 32'b00000000000000011110010100001011;
assign LUT_3[31353] = 32'b00000000000000100100111111101000;
assign LUT_3[31354] = 32'b00000000000000100000011011101111;
assign LUT_3[31355] = 32'b00000000000000100111000111001100;
assign LUT_3[31356] = 32'b00000000000000011011100010000001;
assign LUT_3[31357] = 32'b00000000000000100010001101011110;
assign LUT_3[31358] = 32'b00000000000000011101101001100101;
assign LUT_3[31359] = 32'b00000000000000100100010101000010;
assign LUT_3[31360] = 32'b00000000000000010110101011110101;
assign LUT_3[31361] = 32'b00000000000000011101010111010010;
assign LUT_3[31362] = 32'b00000000000000011000110011011001;
assign LUT_3[31363] = 32'b00000000000000011111011110110110;
assign LUT_3[31364] = 32'b00000000000000010011111001101011;
assign LUT_3[31365] = 32'b00000000000000011010100101001000;
assign LUT_3[31366] = 32'b00000000000000010110000001001111;
assign LUT_3[31367] = 32'b00000000000000011100101100101100;
assign LUT_3[31368] = 32'b00000000000000011100000100111011;
assign LUT_3[31369] = 32'b00000000000000100010110000011000;
assign LUT_3[31370] = 32'b00000000000000011110001100011111;
assign LUT_3[31371] = 32'b00000000000000100100110111111100;
assign LUT_3[31372] = 32'b00000000000000011001010010110001;
assign LUT_3[31373] = 32'b00000000000000011111111110001110;
assign LUT_3[31374] = 32'b00000000000000011011011010010101;
assign LUT_3[31375] = 32'b00000000000000100010000101110010;
assign LUT_3[31376] = 32'b00000000000000011001111110111000;
assign LUT_3[31377] = 32'b00000000000000100000101010010101;
assign LUT_3[31378] = 32'b00000000000000011100000110011100;
assign LUT_3[31379] = 32'b00000000000000100010110001111001;
assign LUT_3[31380] = 32'b00000000000000010111001100101110;
assign LUT_3[31381] = 32'b00000000000000011101111000001011;
assign LUT_3[31382] = 32'b00000000000000011001010100010010;
assign LUT_3[31383] = 32'b00000000000000011111111111101111;
assign LUT_3[31384] = 32'b00000000000000011111010111111110;
assign LUT_3[31385] = 32'b00000000000000100110000011011011;
assign LUT_3[31386] = 32'b00000000000000100001011111100010;
assign LUT_3[31387] = 32'b00000000000000101000001010111111;
assign LUT_3[31388] = 32'b00000000000000011100100101110100;
assign LUT_3[31389] = 32'b00000000000000100011010001010001;
assign LUT_3[31390] = 32'b00000000000000011110101101011000;
assign LUT_3[31391] = 32'b00000000000000100101011000110101;
assign LUT_3[31392] = 32'b00000000000000010111111010010101;
assign LUT_3[31393] = 32'b00000000000000011110100101110010;
assign LUT_3[31394] = 32'b00000000000000011010000001111001;
assign LUT_3[31395] = 32'b00000000000000100000101101010110;
assign LUT_3[31396] = 32'b00000000000000010101001000001011;
assign LUT_3[31397] = 32'b00000000000000011011110011101000;
assign LUT_3[31398] = 32'b00000000000000010111001111101111;
assign LUT_3[31399] = 32'b00000000000000011101111011001100;
assign LUT_3[31400] = 32'b00000000000000011101010011011011;
assign LUT_3[31401] = 32'b00000000000000100011111110111000;
assign LUT_3[31402] = 32'b00000000000000011111011010111111;
assign LUT_3[31403] = 32'b00000000000000100110000110011100;
assign LUT_3[31404] = 32'b00000000000000011010100001010001;
assign LUT_3[31405] = 32'b00000000000000100001001100101110;
assign LUT_3[31406] = 32'b00000000000000011100101000110101;
assign LUT_3[31407] = 32'b00000000000000100011010100010010;
assign LUT_3[31408] = 32'b00000000000000011011001101011000;
assign LUT_3[31409] = 32'b00000000000000100001111000110101;
assign LUT_3[31410] = 32'b00000000000000011101010100111100;
assign LUT_3[31411] = 32'b00000000000000100100000000011001;
assign LUT_3[31412] = 32'b00000000000000011000011011001110;
assign LUT_3[31413] = 32'b00000000000000011111000110101011;
assign LUT_3[31414] = 32'b00000000000000011010100010110010;
assign LUT_3[31415] = 32'b00000000000000100001001110001111;
assign LUT_3[31416] = 32'b00000000000000100000100110011110;
assign LUT_3[31417] = 32'b00000000000000100111010001111011;
assign LUT_3[31418] = 32'b00000000000000100010101110000010;
assign LUT_3[31419] = 32'b00000000000000101001011001011111;
assign LUT_3[31420] = 32'b00000000000000011101110100010100;
assign LUT_3[31421] = 32'b00000000000000100100011111110001;
assign LUT_3[31422] = 32'b00000000000000011111111011111000;
assign LUT_3[31423] = 32'b00000000000000100110100111010101;
assign LUT_3[31424] = 32'b00000000000000010110100100100000;
assign LUT_3[31425] = 32'b00000000000000011101001111111101;
assign LUT_3[31426] = 32'b00000000000000011000101100000100;
assign LUT_3[31427] = 32'b00000000000000011111010111100001;
assign LUT_3[31428] = 32'b00000000000000010011110010010110;
assign LUT_3[31429] = 32'b00000000000000011010011101110011;
assign LUT_3[31430] = 32'b00000000000000010101111001111010;
assign LUT_3[31431] = 32'b00000000000000011100100101010111;
assign LUT_3[31432] = 32'b00000000000000011011111101100110;
assign LUT_3[31433] = 32'b00000000000000100010101001000011;
assign LUT_3[31434] = 32'b00000000000000011110000101001010;
assign LUT_3[31435] = 32'b00000000000000100100110000100111;
assign LUT_3[31436] = 32'b00000000000000011001001011011100;
assign LUT_3[31437] = 32'b00000000000000011111110110111001;
assign LUT_3[31438] = 32'b00000000000000011011010011000000;
assign LUT_3[31439] = 32'b00000000000000100001111110011101;
assign LUT_3[31440] = 32'b00000000000000011001110111100011;
assign LUT_3[31441] = 32'b00000000000000100000100011000000;
assign LUT_3[31442] = 32'b00000000000000011011111111000111;
assign LUT_3[31443] = 32'b00000000000000100010101010100100;
assign LUT_3[31444] = 32'b00000000000000010111000101011001;
assign LUT_3[31445] = 32'b00000000000000011101110000110110;
assign LUT_3[31446] = 32'b00000000000000011001001100111101;
assign LUT_3[31447] = 32'b00000000000000011111111000011010;
assign LUT_3[31448] = 32'b00000000000000011111010000101001;
assign LUT_3[31449] = 32'b00000000000000100101111100000110;
assign LUT_3[31450] = 32'b00000000000000100001011000001101;
assign LUT_3[31451] = 32'b00000000000000101000000011101010;
assign LUT_3[31452] = 32'b00000000000000011100011110011111;
assign LUT_3[31453] = 32'b00000000000000100011001001111100;
assign LUT_3[31454] = 32'b00000000000000011110100110000011;
assign LUT_3[31455] = 32'b00000000000000100101010001100000;
assign LUT_3[31456] = 32'b00000000000000010111110011000000;
assign LUT_3[31457] = 32'b00000000000000011110011110011101;
assign LUT_3[31458] = 32'b00000000000000011001111010100100;
assign LUT_3[31459] = 32'b00000000000000100000100110000001;
assign LUT_3[31460] = 32'b00000000000000010101000000110110;
assign LUT_3[31461] = 32'b00000000000000011011101100010011;
assign LUT_3[31462] = 32'b00000000000000010111001000011010;
assign LUT_3[31463] = 32'b00000000000000011101110011110111;
assign LUT_3[31464] = 32'b00000000000000011101001100000110;
assign LUT_3[31465] = 32'b00000000000000100011110111100011;
assign LUT_3[31466] = 32'b00000000000000011111010011101010;
assign LUT_3[31467] = 32'b00000000000000100101111111000111;
assign LUT_3[31468] = 32'b00000000000000011010011001111100;
assign LUT_3[31469] = 32'b00000000000000100001000101011001;
assign LUT_3[31470] = 32'b00000000000000011100100001100000;
assign LUT_3[31471] = 32'b00000000000000100011001100111101;
assign LUT_3[31472] = 32'b00000000000000011011000110000011;
assign LUT_3[31473] = 32'b00000000000000100001110001100000;
assign LUT_3[31474] = 32'b00000000000000011101001101100111;
assign LUT_3[31475] = 32'b00000000000000100011111001000100;
assign LUT_3[31476] = 32'b00000000000000011000010011111001;
assign LUT_3[31477] = 32'b00000000000000011110111111010110;
assign LUT_3[31478] = 32'b00000000000000011010011011011101;
assign LUT_3[31479] = 32'b00000000000000100001000110111010;
assign LUT_3[31480] = 32'b00000000000000100000011111001001;
assign LUT_3[31481] = 32'b00000000000000100111001010100110;
assign LUT_3[31482] = 32'b00000000000000100010100110101101;
assign LUT_3[31483] = 32'b00000000000000101001010010001010;
assign LUT_3[31484] = 32'b00000000000000011101101100111111;
assign LUT_3[31485] = 32'b00000000000000100100011000011100;
assign LUT_3[31486] = 32'b00000000000000011111110100100011;
assign LUT_3[31487] = 32'b00000000000000100110100000000000;
assign LUT_3[31488] = 32'b00000000000000010000110000011000;
assign LUT_3[31489] = 32'b00000000000000010111011011110101;
assign LUT_3[31490] = 32'b00000000000000010010110111111100;
assign LUT_3[31491] = 32'b00000000000000011001100011011001;
assign LUT_3[31492] = 32'b00000000000000001101111110001110;
assign LUT_3[31493] = 32'b00000000000000010100101001101011;
assign LUT_3[31494] = 32'b00000000000000010000000101110010;
assign LUT_3[31495] = 32'b00000000000000010110110001001111;
assign LUT_3[31496] = 32'b00000000000000010110001001011110;
assign LUT_3[31497] = 32'b00000000000000011100110100111011;
assign LUT_3[31498] = 32'b00000000000000011000010001000010;
assign LUT_3[31499] = 32'b00000000000000011110111100011111;
assign LUT_3[31500] = 32'b00000000000000010011010111010100;
assign LUT_3[31501] = 32'b00000000000000011010000010110001;
assign LUT_3[31502] = 32'b00000000000000010101011110111000;
assign LUT_3[31503] = 32'b00000000000000011100001010010101;
assign LUT_3[31504] = 32'b00000000000000010100000011011011;
assign LUT_3[31505] = 32'b00000000000000011010101110111000;
assign LUT_3[31506] = 32'b00000000000000010110001010111111;
assign LUT_3[31507] = 32'b00000000000000011100110110011100;
assign LUT_3[31508] = 32'b00000000000000010001010001010001;
assign LUT_3[31509] = 32'b00000000000000010111111100101110;
assign LUT_3[31510] = 32'b00000000000000010011011000110101;
assign LUT_3[31511] = 32'b00000000000000011010000100010010;
assign LUT_3[31512] = 32'b00000000000000011001011100100001;
assign LUT_3[31513] = 32'b00000000000000100000000111111110;
assign LUT_3[31514] = 32'b00000000000000011011100100000101;
assign LUT_3[31515] = 32'b00000000000000100010001111100010;
assign LUT_3[31516] = 32'b00000000000000010110101010010111;
assign LUT_3[31517] = 32'b00000000000000011101010101110100;
assign LUT_3[31518] = 32'b00000000000000011000110001111011;
assign LUT_3[31519] = 32'b00000000000000011111011101011000;
assign LUT_3[31520] = 32'b00000000000000010001111110111000;
assign LUT_3[31521] = 32'b00000000000000011000101010010101;
assign LUT_3[31522] = 32'b00000000000000010100000110011100;
assign LUT_3[31523] = 32'b00000000000000011010110001111001;
assign LUT_3[31524] = 32'b00000000000000001111001100101110;
assign LUT_3[31525] = 32'b00000000000000010101111000001011;
assign LUT_3[31526] = 32'b00000000000000010001010100010010;
assign LUT_3[31527] = 32'b00000000000000010111111111101111;
assign LUT_3[31528] = 32'b00000000000000010111010111111110;
assign LUT_3[31529] = 32'b00000000000000011110000011011011;
assign LUT_3[31530] = 32'b00000000000000011001011111100010;
assign LUT_3[31531] = 32'b00000000000000100000001010111111;
assign LUT_3[31532] = 32'b00000000000000010100100101110100;
assign LUT_3[31533] = 32'b00000000000000011011010001010001;
assign LUT_3[31534] = 32'b00000000000000010110101101011000;
assign LUT_3[31535] = 32'b00000000000000011101011000110101;
assign LUT_3[31536] = 32'b00000000000000010101010001111011;
assign LUT_3[31537] = 32'b00000000000000011011111101011000;
assign LUT_3[31538] = 32'b00000000000000010111011001011111;
assign LUT_3[31539] = 32'b00000000000000011110000100111100;
assign LUT_3[31540] = 32'b00000000000000010010011111110001;
assign LUT_3[31541] = 32'b00000000000000011001001011001110;
assign LUT_3[31542] = 32'b00000000000000010100100111010101;
assign LUT_3[31543] = 32'b00000000000000011011010010110010;
assign LUT_3[31544] = 32'b00000000000000011010101011000001;
assign LUT_3[31545] = 32'b00000000000000100001010110011110;
assign LUT_3[31546] = 32'b00000000000000011100110010100101;
assign LUT_3[31547] = 32'b00000000000000100011011110000010;
assign LUT_3[31548] = 32'b00000000000000010111111000110111;
assign LUT_3[31549] = 32'b00000000000000011110100100010100;
assign LUT_3[31550] = 32'b00000000000000011010000000011011;
assign LUT_3[31551] = 32'b00000000000000100000101011111000;
assign LUT_3[31552] = 32'b00000000000000010000101001000011;
assign LUT_3[31553] = 32'b00000000000000010111010100100000;
assign LUT_3[31554] = 32'b00000000000000010010110000100111;
assign LUT_3[31555] = 32'b00000000000000011001011100000100;
assign LUT_3[31556] = 32'b00000000000000001101110110111001;
assign LUT_3[31557] = 32'b00000000000000010100100010010110;
assign LUT_3[31558] = 32'b00000000000000001111111110011101;
assign LUT_3[31559] = 32'b00000000000000010110101001111010;
assign LUT_3[31560] = 32'b00000000000000010110000010001001;
assign LUT_3[31561] = 32'b00000000000000011100101101100110;
assign LUT_3[31562] = 32'b00000000000000011000001001101101;
assign LUT_3[31563] = 32'b00000000000000011110110101001010;
assign LUT_3[31564] = 32'b00000000000000010011001111111111;
assign LUT_3[31565] = 32'b00000000000000011001111011011100;
assign LUT_3[31566] = 32'b00000000000000010101010111100011;
assign LUT_3[31567] = 32'b00000000000000011100000011000000;
assign LUT_3[31568] = 32'b00000000000000010011111100000110;
assign LUT_3[31569] = 32'b00000000000000011010100111100011;
assign LUT_3[31570] = 32'b00000000000000010110000011101010;
assign LUT_3[31571] = 32'b00000000000000011100101111000111;
assign LUT_3[31572] = 32'b00000000000000010001001001111100;
assign LUT_3[31573] = 32'b00000000000000010111110101011001;
assign LUT_3[31574] = 32'b00000000000000010011010001100000;
assign LUT_3[31575] = 32'b00000000000000011001111100111101;
assign LUT_3[31576] = 32'b00000000000000011001010101001100;
assign LUT_3[31577] = 32'b00000000000000100000000000101001;
assign LUT_3[31578] = 32'b00000000000000011011011100110000;
assign LUT_3[31579] = 32'b00000000000000100010001000001101;
assign LUT_3[31580] = 32'b00000000000000010110100011000010;
assign LUT_3[31581] = 32'b00000000000000011101001110011111;
assign LUT_3[31582] = 32'b00000000000000011000101010100110;
assign LUT_3[31583] = 32'b00000000000000011111010110000011;
assign LUT_3[31584] = 32'b00000000000000010001110111100011;
assign LUT_3[31585] = 32'b00000000000000011000100011000000;
assign LUT_3[31586] = 32'b00000000000000010011111111000111;
assign LUT_3[31587] = 32'b00000000000000011010101010100100;
assign LUT_3[31588] = 32'b00000000000000001111000101011001;
assign LUT_3[31589] = 32'b00000000000000010101110000110110;
assign LUT_3[31590] = 32'b00000000000000010001001100111101;
assign LUT_3[31591] = 32'b00000000000000010111111000011010;
assign LUT_3[31592] = 32'b00000000000000010111010000101001;
assign LUT_3[31593] = 32'b00000000000000011101111100000110;
assign LUT_3[31594] = 32'b00000000000000011001011000001101;
assign LUT_3[31595] = 32'b00000000000000100000000011101010;
assign LUT_3[31596] = 32'b00000000000000010100011110011111;
assign LUT_3[31597] = 32'b00000000000000011011001001111100;
assign LUT_3[31598] = 32'b00000000000000010110100110000011;
assign LUT_3[31599] = 32'b00000000000000011101010001100000;
assign LUT_3[31600] = 32'b00000000000000010101001010100110;
assign LUT_3[31601] = 32'b00000000000000011011110110000011;
assign LUT_3[31602] = 32'b00000000000000010111010010001010;
assign LUT_3[31603] = 32'b00000000000000011101111101100111;
assign LUT_3[31604] = 32'b00000000000000010010011000011100;
assign LUT_3[31605] = 32'b00000000000000011001000011111001;
assign LUT_3[31606] = 32'b00000000000000010100100000000000;
assign LUT_3[31607] = 32'b00000000000000011011001011011101;
assign LUT_3[31608] = 32'b00000000000000011010100011101100;
assign LUT_3[31609] = 32'b00000000000000100001001111001001;
assign LUT_3[31610] = 32'b00000000000000011100101011010000;
assign LUT_3[31611] = 32'b00000000000000100011010110101101;
assign LUT_3[31612] = 32'b00000000000000010111110001100010;
assign LUT_3[31613] = 32'b00000000000000011110011100111111;
assign LUT_3[31614] = 32'b00000000000000011001111001000110;
assign LUT_3[31615] = 32'b00000000000000100000100100100011;
assign LUT_3[31616] = 32'b00000000000000010010111011010110;
assign LUT_3[31617] = 32'b00000000000000011001100110110011;
assign LUT_3[31618] = 32'b00000000000000010101000010111010;
assign LUT_3[31619] = 32'b00000000000000011011101110010111;
assign LUT_3[31620] = 32'b00000000000000010000001001001100;
assign LUT_3[31621] = 32'b00000000000000010110110100101001;
assign LUT_3[31622] = 32'b00000000000000010010010000110000;
assign LUT_3[31623] = 32'b00000000000000011000111100001101;
assign LUT_3[31624] = 32'b00000000000000011000010100011100;
assign LUT_3[31625] = 32'b00000000000000011110111111111001;
assign LUT_3[31626] = 32'b00000000000000011010011100000000;
assign LUT_3[31627] = 32'b00000000000000100001000111011101;
assign LUT_3[31628] = 32'b00000000000000010101100010010010;
assign LUT_3[31629] = 32'b00000000000000011100001101101111;
assign LUT_3[31630] = 32'b00000000000000010111101001110110;
assign LUT_3[31631] = 32'b00000000000000011110010101010011;
assign LUT_3[31632] = 32'b00000000000000010110001110011001;
assign LUT_3[31633] = 32'b00000000000000011100111001110110;
assign LUT_3[31634] = 32'b00000000000000011000010101111101;
assign LUT_3[31635] = 32'b00000000000000011111000001011010;
assign LUT_3[31636] = 32'b00000000000000010011011100001111;
assign LUT_3[31637] = 32'b00000000000000011010000111101100;
assign LUT_3[31638] = 32'b00000000000000010101100011110011;
assign LUT_3[31639] = 32'b00000000000000011100001111010000;
assign LUT_3[31640] = 32'b00000000000000011011100111011111;
assign LUT_3[31641] = 32'b00000000000000100010010010111100;
assign LUT_3[31642] = 32'b00000000000000011101101111000011;
assign LUT_3[31643] = 32'b00000000000000100100011010100000;
assign LUT_3[31644] = 32'b00000000000000011000110101010101;
assign LUT_3[31645] = 32'b00000000000000011111100000110010;
assign LUT_3[31646] = 32'b00000000000000011010111100111001;
assign LUT_3[31647] = 32'b00000000000000100001101000010110;
assign LUT_3[31648] = 32'b00000000000000010100001001110110;
assign LUT_3[31649] = 32'b00000000000000011010110101010011;
assign LUT_3[31650] = 32'b00000000000000010110010001011010;
assign LUT_3[31651] = 32'b00000000000000011100111100110111;
assign LUT_3[31652] = 32'b00000000000000010001010111101100;
assign LUT_3[31653] = 32'b00000000000000011000000011001001;
assign LUT_3[31654] = 32'b00000000000000010011011111010000;
assign LUT_3[31655] = 32'b00000000000000011010001010101101;
assign LUT_3[31656] = 32'b00000000000000011001100010111100;
assign LUT_3[31657] = 32'b00000000000000100000001110011001;
assign LUT_3[31658] = 32'b00000000000000011011101010100000;
assign LUT_3[31659] = 32'b00000000000000100010010101111101;
assign LUT_3[31660] = 32'b00000000000000010110110000110010;
assign LUT_3[31661] = 32'b00000000000000011101011100001111;
assign LUT_3[31662] = 32'b00000000000000011000111000010110;
assign LUT_3[31663] = 32'b00000000000000011111100011110011;
assign LUT_3[31664] = 32'b00000000000000010111011100111001;
assign LUT_3[31665] = 32'b00000000000000011110001000010110;
assign LUT_3[31666] = 32'b00000000000000011001100100011101;
assign LUT_3[31667] = 32'b00000000000000100000001111111010;
assign LUT_3[31668] = 32'b00000000000000010100101010101111;
assign LUT_3[31669] = 32'b00000000000000011011010110001100;
assign LUT_3[31670] = 32'b00000000000000010110110010010011;
assign LUT_3[31671] = 32'b00000000000000011101011101110000;
assign LUT_3[31672] = 32'b00000000000000011100110101111111;
assign LUT_3[31673] = 32'b00000000000000100011100001011100;
assign LUT_3[31674] = 32'b00000000000000011110111101100011;
assign LUT_3[31675] = 32'b00000000000000100101101001000000;
assign LUT_3[31676] = 32'b00000000000000011010000011110101;
assign LUT_3[31677] = 32'b00000000000000100000101111010010;
assign LUT_3[31678] = 32'b00000000000000011100001011011001;
assign LUT_3[31679] = 32'b00000000000000100010110110110110;
assign LUT_3[31680] = 32'b00000000000000010010110100000001;
assign LUT_3[31681] = 32'b00000000000000011001011111011110;
assign LUT_3[31682] = 32'b00000000000000010100111011100101;
assign LUT_3[31683] = 32'b00000000000000011011100111000010;
assign LUT_3[31684] = 32'b00000000000000010000000001110111;
assign LUT_3[31685] = 32'b00000000000000010110101101010100;
assign LUT_3[31686] = 32'b00000000000000010010001001011011;
assign LUT_3[31687] = 32'b00000000000000011000110100111000;
assign LUT_3[31688] = 32'b00000000000000011000001101000111;
assign LUT_3[31689] = 32'b00000000000000011110111000100100;
assign LUT_3[31690] = 32'b00000000000000011010010100101011;
assign LUT_3[31691] = 32'b00000000000000100001000000001000;
assign LUT_3[31692] = 32'b00000000000000010101011010111101;
assign LUT_3[31693] = 32'b00000000000000011100000110011010;
assign LUT_3[31694] = 32'b00000000000000010111100010100001;
assign LUT_3[31695] = 32'b00000000000000011110001101111110;
assign LUT_3[31696] = 32'b00000000000000010110000111000100;
assign LUT_3[31697] = 32'b00000000000000011100110010100001;
assign LUT_3[31698] = 32'b00000000000000011000001110101000;
assign LUT_3[31699] = 32'b00000000000000011110111010000101;
assign LUT_3[31700] = 32'b00000000000000010011010100111010;
assign LUT_3[31701] = 32'b00000000000000011010000000010111;
assign LUT_3[31702] = 32'b00000000000000010101011100011110;
assign LUT_3[31703] = 32'b00000000000000011100000111111011;
assign LUT_3[31704] = 32'b00000000000000011011100000001010;
assign LUT_3[31705] = 32'b00000000000000100010001011100111;
assign LUT_3[31706] = 32'b00000000000000011101100111101110;
assign LUT_3[31707] = 32'b00000000000000100100010011001011;
assign LUT_3[31708] = 32'b00000000000000011000101110000000;
assign LUT_3[31709] = 32'b00000000000000011111011001011101;
assign LUT_3[31710] = 32'b00000000000000011010110101100100;
assign LUT_3[31711] = 32'b00000000000000100001100001000001;
assign LUT_3[31712] = 32'b00000000000000010100000010100001;
assign LUT_3[31713] = 32'b00000000000000011010101101111110;
assign LUT_3[31714] = 32'b00000000000000010110001010000101;
assign LUT_3[31715] = 32'b00000000000000011100110101100010;
assign LUT_3[31716] = 32'b00000000000000010001010000010111;
assign LUT_3[31717] = 32'b00000000000000010111111011110100;
assign LUT_3[31718] = 32'b00000000000000010011010111111011;
assign LUT_3[31719] = 32'b00000000000000011010000011011000;
assign LUT_3[31720] = 32'b00000000000000011001011011100111;
assign LUT_3[31721] = 32'b00000000000000100000000111000100;
assign LUT_3[31722] = 32'b00000000000000011011100011001011;
assign LUT_3[31723] = 32'b00000000000000100010001110101000;
assign LUT_3[31724] = 32'b00000000000000010110101001011101;
assign LUT_3[31725] = 32'b00000000000000011101010100111010;
assign LUT_3[31726] = 32'b00000000000000011000110001000001;
assign LUT_3[31727] = 32'b00000000000000011111011100011110;
assign LUT_3[31728] = 32'b00000000000000010111010101100100;
assign LUT_3[31729] = 32'b00000000000000011110000001000001;
assign LUT_3[31730] = 32'b00000000000000011001011101001000;
assign LUT_3[31731] = 32'b00000000000000100000001000100101;
assign LUT_3[31732] = 32'b00000000000000010100100011011010;
assign LUT_3[31733] = 32'b00000000000000011011001110110111;
assign LUT_3[31734] = 32'b00000000000000010110101010111110;
assign LUT_3[31735] = 32'b00000000000000011101010110011011;
assign LUT_3[31736] = 32'b00000000000000011100101110101010;
assign LUT_3[31737] = 32'b00000000000000100011011010000111;
assign LUT_3[31738] = 32'b00000000000000011110110110001110;
assign LUT_3[31739] = 32'b00000000000000100101100001101011;
assign LUT_3[31740] = 32'b00000000000000011001111100100000;
assign LUT_3[31741] = 32'b00000000000000100000100111111101;
assign LUT_3[31742] = 32'b00000000000000011100000100000100;
assign LUT_3[31743] = 32'b00000000000000100010101111100001;
assign LUT_3[31744] = 32'b00000000000000010111110000101000;
assign LUT_3[31745] = 32'b00000000000000011110011100000101;
assign LUT_3[31746] = 32'b00000000000000011001111000001100;
assign LUT_3[31747] = 32'b00000000000000100000100011101001;
assign LUT_3[31748] = 32'b00000000000000010100111110011110;
assign LUT_3[31749] = 32'b00000000000000011011101001111011;
assign LUT_3[31750] = 32'b00000000000000010111000110000010;
assign LUT_3[31751] = 32'b00000000000000011101110001011111;
assign LUT_3[31752] = 32'b00000000000000011101001001101110;
assign LUT_3[31753] = 32'b00000000000000100011110101001011;
assign LUT_3[31754] = 32'b00000000000000011111010001010010;
assign LUT_3[31755] = 32'b00000000000000100101111100101111;
assign LUT_3[31756] = 32'b00000000000000011010010111100100;
assign LUT_3[31757] = 32'b00000000000000100001000011000001;
assign LUT_3[31758] = 32'b00000000000000011100011111001000;
assign LUT_3[31759] = 32'b00000000000000100011001010100101;
assign LUT_3[31760] = 32'b00000000000000011011000011101011;
assign LUT_3[31761] = 32'b00000000000000100001101111001000;
assign LUT_3[31762] = 32'b00000000000000011101001011001111;
assign LUT_3[31763] = 32'b00000000000000100011110110101100;
assign LUT_3[31764] = 32'b00000000000000011000010001100001;
assign LUT_3[31765] = 32'b00000000000000011110111100111110;
assign LUT_3[31766] = 32'b00000000000000011010011001000101;
assign LUT_3[31767] = 32'b00000000000000100001000100100010;
assign LUT_3[31768] = 32'b00000000000000100000011100110001;
assign LUT_3[31769] = 32'b00000000000000100111001000001110;
assign LUT_3[31770] = 32'b00000000000000100010100100010101;
assign LUT_3[31771] = 32'b00000000000000101001001111110010;
assign LUT_3[31772] = 32'b00000000000000011101101010100111;
assign LUT_3[31773] = 32'b00000000000000100100010110000100;
assign LUT_3[31774] = 32'b00000000000000011111110010001011;
assign LUT_3[31775] = 32'b00000000000000100110011101101000;
assign LUT_3[31776] = 32'b00000000000000011000111111001000;
assign LUT_3[31777] = 32'b00000000000000011111101010100101;
assign LUT_3[31778] = 32'b00000000000000011011000110101100;
assign LUT_3[31779] = 32'b00000000000000100001110010001001;
assign LUT_3[31780] = 32'b00000000000000010110001100111110;
assign LUT_3[31781] = 32'b00000000000000011100111000011011;
assign LUT_3[31782] = 32'b00000000000000011000010100100010;
assign LUT_3[31783] = 32'b00000000000000011110111111111111;
assign LUT_3[31784] = 32'b00000000000000011110011000001110;
assign LUT_3[31785] = 32'b00000000000000100101000011101011;
assign LUT_3[31786] = 32'b00000000000000100000011111110010;
assign LUT_3[31787] = 32'b00000000000000100111001011001111;
assign LUT_3[31788] = 32'b00000000000000011011100110000100;
assign LUT_3[31789] = 32'b00000000000000100010010001100001;
assign LUT_3[31790] = 32'b00000000000000011101101101101000;
assign LUT_3[31791] = 32'b00000000000000100100011001000101;
assign LUT_3[31792] = 32'b00000000000000011100010010001011;
assign LUT_3[31793] = 32'b00000000000000100010111101101000;
assign LUT_3[31794] = 32'b00000000000000011110011001101111;
assign LUT_3[31795] = 32'b00000000000000100101000101001100;
assign LUT_3[31796] = 32'b00000000000000011001100000000001;
assign LUT_3[31797] = 32'b00000000000000100000001011011110;
assign LUT_3[31798] = 32'b00000000000000011011100111100101;
assign LUT_3[31799] = 32'b00000000000000100010010011000010;
assign LUT_3[31800] = 32'b00000000000000100001101011010001;
assign LUT_3[31801] = 32'b00000000000000101000010110101110;
assign LUT_3[31802] = 32'b00000000000000100011110010110101;
assign LUT_3[31803] = 32'b00000000000000101010011110010010;
assign LUT_3[31804] = 32'b00000000000000011110111001000111;
assign LUT_3[31805] = 32'b00000000000000100101100100100100;
assign LUT_3[31806] = 32'b00000000000000100001000000101011;
assign LUT_3[31807] = 32'b00000000000000100111101100001000;
assign LUT_3[31808] = 32'b00000000000000010111101001010011;
assign LUT_3[31809] = 32'b00000000000000011110010100110000;
assign LUT_3[31810] = 32'b00000000000000011001110000110111;
assign LUT_3[31811] = 32'b00000000000000100000011100010100;
assign LUT_3[31812] = 32'b00000000000000010100110111001001;
assign LUT_3[31813] = 32'b00000000000000011011100010100110;
assign LUT_3[31814] = 32'b00000000000000010110111110101101;
assign LUT_3[31815] = 32'b00000000000000011101101010001010;
assign LUT_3[31816] = 32'b00000000000000011101000010011001;
assign LUT_3[31817] = 32'b00000000000000100011101101110110;
assign LUT_3[31818] = 32'b00000000000000011111001001111101;
assign LUT_3[31819] = 32'b00000000000000100101110101011010;
assign LUT_3[31820] = 32'b00000000000000011010010000001111;
assign LUT_3[31821] = 32'b00000000000000100000111011101100;
assign LUT_3[31822] = 32'b00000000000000011100010111110011;
assign LUT_3[31823] = 32'b00000000000000100011000011010000;
assign LUT_3[31824] = 32'b00000000000000011010111100010110;
assign LUT_3[31825] = 32'b00000000000000100001100111110011;
assign LUT_3[31826] = 32'b00000000000000011101000011111010;
assign LUT_3[31827] = 32'b00000000000000100011101111010111;
assign LUT_3[31828] = 32'b00000000000000011000001010001100;
assign LUT_3[31829] = 32'b00000000000000011110110101101001;
assign LUT_3[31830] = 32'b00000000000000011010010001110000;
assign LUT_3[31831] = 32'b00000000000000100000111101001101;
assign LUT_3[31832] = 32'b00000000000000100000010101011100;
assign LUT_3[31833] = 32'b00000000000000100111000000111001;
assign LUT_3[31834] = 32'b00000000000000100010011101000000;
assign LUT_3[31835] = 32'b00000000000000101001001000011101;
assign LUT_3[31836] = 32'b00000000000000011101100011010010;
assign LUT_3[31837] = 32'b00000000000000100100001110101111;
assign LUT_3[31838] = 32'b00000000000000011111101010110110;
assign LUT_3[31839] = 32'b00000000000000100110010110010011;
assign LUT_3[31840] = 32'b00000000000000011000110111110011;
assign LUT_3[31841] = 32'b00000000000000011111100011010000;
assign LUT_3[31842] = 32'b00000000000000011010111111010111;
assign LUT_3[31843] = 32'b00000000000000100001101010110100;
assign LUT_3[31844] = 32'b00000000000000010110000101101001;
assign LUT_3[31845] = 32'b00000000000000011100110001000110;
assign LUT_3[31846] = 32'b00000000000000011000001101001101;
assign LUT_3[31847] = 32'b00000000000000011110111000101010;
assign LUT_3[31848] = 32'b00000000000000011110010000111001;
assign LUT_3[31849] = 32'b00000000000000100100111100010110;
assign LUT_3[31850] = 32'b00000000000000100000011000011101;
assign LUT_3[31851] = 32'b00000000000000100111000011111010;
assign LUT_3[31852] = 32'b00000000000000011011011110101111;
assign LUT_3[31853] = 32'b00000000000000100010001010001100;
assign LUT_3[31854] = 32'b00000000000000011101100110010011;
assign LUT_3[31855] = 32'b00000000000000100100010001110000;
assign LUT_3[31856] = 32'b00000000000000011100001010110110;
assign LUT_3[31857] = 32'b00000000000000100010110110010011;
assign LUT_3[31858] = 32'b00000000000000011110010010011010;
assign LUT_3[31859] = 32'b00000000000000100100111101110111;
assign LUT_3[31860] = 32'b00000000000000011001011000101100;
assign LUT_3[31861] = 32'b00000000000000100000000100001001;
assign LUT_3[31862] = 32'b00000000000000011011100000010000;
assign LUT_3[31863] = 32'b00000000000000100010001011101101;
assign LUT_3[31864] = 32'b00000000000000100001100011111100;
assign LUT_3[31865] = 32'b00000000000000101000001111011001;
assign LUT_3[31866] = 32'b00000000000000100011101011100000;
assign LUT_3[31867] = 32'b00000000000000101010010110111101;
assign LUT_3[31868] = 32'b00000000000000011110110001110010;
assign LUT_3[31869] = 32'b00000000000000100101011101001111;
assign LUT_3[31870] = 32'b00000000000000100000111001010110;
assign LUT_3[31871] = 32'b00000000000000100111100100110011;
assign LUT_3[31872] = 32'b00000000000000011001111011100110;
assign LUT_3[31873] = 32'b00000000000000100000100111000011;
assign LUT_3[31874] = 32'b00000000000000011100000011001010;
assign LUT_3[31875] = 32'b00000000000000100010101110100111;
assign LUT_3[31876] = 32'b00000000000000010111001001011100;
assign LUT_3[31877] = 32'b00000000000000011101110100111001;
assign LUT_3[31878] = 32'b00000000000000011001010001000000;
assign LUT_3[31879] = 32'b00000000000000011111111100011101;
assign LUT_3[31880] = 32'b00000000000000011111010100101100;
assign LUT_3[31881] = 32'b00000000000000100110000000001001;
assign LUT_3[31882] = 32'b00000000000000100001011100010000;
assign LUT_3[31883] = 32'b00000000000000101000000111101101;
assign LUT_3[31884] = 32'b00000000000000011100100010100010;
assign LUT_3[31885] = 32'b00000000000000100011001101111111;
assign LUT_3[31886] = 32'b00000000000000011110101010000110;
assign LUT_3[31887] = 32'b00000000000000100101010101100011;
assign LUT_3[31888] = 32'b00000000000000011101001110101001;
assign LUT_3[31889] = 32'b00000000000000100011111010000110;
assign LUT_3[31890] = 32'b00000000000000011111010110001101;
assign LUT_3[31891] = 32'b00000000000000100110000001101010;
assign LUT_3[31892] = 32'b00000000000000011010011100011111;
assign LUT_3[31893] = 32'b00000000000000100001000111111100;
assign LUT_3[31894] = 32'b00000000000000011100100100000011;
assign LUT_3[31895] = 32'b00000000000000100011001111100000;
assign LUT_3[31896] = 32'b00000000000000100010100111101111;
assign LUT_3[31897] = 32'b00000000000000101001010011001100;
assign LUT_3[31898] = 32'b00000000000000100100101111010011;
assign LUT_3[31899] = 32'b00000000000000101011011010110000;
assign LUT_3[31900] = 32'b00000000000000011111110101100101;
assign LUT_3[31901] = 32'b00000000000000100110100001000010;
assign LUT_3[31902] = 32'b00000000000000100001111101001001;
assign LUT_3[31903] = 32'b00000000000000101000101000100110;
assign LUT_3[31904] = 32'b00000000000000011011001010000110;
assign LUT_3[31905] = 32'b00000000000000100001110101100011;
assign LUT_3[31906] = 32'b00000000000000011101010001101010;
assign LUT_3[31907] = 32'b00000000000000100011111101000111;
assign LUT_3[31908] = 32'b00000000000000011000010111111100;
assign LUT_3[31909] = 32'b00000000000000011111000011011001;
assign LUT_3[31910] = 32'b00000000000000011010011111100000;
assign LUT_3[31911] = 32'b00000000000000100001001010111101;
assign LUT_3[31912] = 32'b00000000000000100000100011001100;
assign LUT_3[31913] = 32'b00000000000000100111001110101001;
assign LUT_3[31914] = 32'b00000000000000100010101010110000;
assign LUT_3[31915] = 32'b00000000000000101001010110001101;
assign LUT_3[31916] = 32'b00000000000000011101110001000010;
assign LUT_3[31917] = 32'b00000000000000100100011100011111;
assign LUT_3[31918] = 32'b00000000000000011111111000100110;
assign LUT_3[31919] = 32'b00000000000000100110100100000011;
assign LUT_3[31920] = 32'b00000000000000011110011101001001;
assign LUT_3[31921] = 32'b00000000000000100101001000100110;
assign LUT_3[31922] = 32'b00000000000000100000100100101101;
assign LUT_3[31923] = 32'b00000000000000100111010000001010;
assign LUT_3[31924] = 32'b00000000000000011011101010111111;
assign LUT_3[31925] = 32'b00000000000000100010010110011100;
assign LUT_3[31926] = 32'b00000000000000011101110010100011;
assign LUT_3[31927] = 32'b00000000000000100100011110000000;
assign LUT_3[31928] = 32'b00000000000000100011110110001111;
assign LUT_3[31929] = 32'b00000000000000101010100001101100;
assign LUT_3[31930] = 32'b00000000000000100101111101110011;
assign LUT_3[31931] = 32'b00000000000000101100101001010000;
assign LUT_3[31932] = 32'b00000000000000100001000100000101;
assign LUT_3[31933] = 32'b00000000000000100111101111100010;
assign LUT_3[31934] = 32'b00000000000000100011001011101001;
assign LUT_3[31935] = 32'b00000000000000101001110111000110;
assign LUT_3[31936] = 32'b00000000000000011001110100010001;
assign LUT_3[31937] = 32'b00000000000000100000011111101110;
assign LUT_3[31938] = 32'b00000000000000011011111011110101;
assign LUT_3[31939] = 32'b00000000000000100010100111010010;
assign LUT_3[31940] = 32'b00000000000000010111000010000111;
assign LUT_3[31941] = 32'b00000000000000011101101101100100;
assign LUT_3[31942] = 32'b00000000000000011001001001101011;
assign LUT_3[31943] = 32'b00000000000000011111110101001000;
assign LUT_3[31944] = 32'b00000000000000011111001101010111;
assign LUT_3[31945] = 32'b00000000000000100101111000110100;
assign LUT_3[31946] = 32'b00000000000000100001010100111011;
assign LUT_3[31947] = 32'b00000000000000101000000000011000;
assign LUT_3[31948] = 32'b00000000000000011100011011001101;
assign LUT_3[31949] = 32'b00000000000000100011000110101010;
assign LUT_3[31950] = 32'b00000000000000011110100010110001;
assign LUT_3[31951] = 32'b00000000000000100101001110001110;
assign LUT_3[31952] = 32'b00000000000000011101000111010100;
assign LUT_3[31953] = 32'b00000000000000100011110010110001;
assign LUT_3[31954] = 32'b00000000000000011111001110111000;
assign LUT_3[31955] = 32'b00000000000000100101111010010101;
assign LUT_3[31956] = 32'b00000000000000011010010101001010;
assign LUT_3[31957] = 32'b00000000000000100001000000100111;
assign LUT_3[31958] = 32'b00000000000000011100011100101110;
assign LUT_3[31959] = 32'b00000000000000100011001000001011;
assign LUT_3[31960] = 32'b00000000000000100010100000011010;
assign LUT_3[31961] = 32'b00000000000000101001001011110111;
assign LUT_3[31962] = 32'b00000000000000100100100111111110;
assign LUT_3[31963] = 32'b00000000000000101011010011011011;
assign LUT_3[31964] = 32'b00000000000000011111101110010000;
assign LUT_3[31965] = 32'b00000000000000100110011001101101;
assign LUT_3[31966] = 32'b00000000000000100001110101110100;
assign LUT_3[31967] = 32'b00000000000000101000100001010001;
assign LUT_3[31968] = 32'b00000000000000011011000010110001;
assign LUT_3[31969] = 32'b00000000000000100001101110001110;
assign LUT_3[31970] = 32'b00000000000000011101001010010101;
assign LUT_3[31971] = 32'b00000000000000100011110101110010;
assign LUT_3[31972] = 32'b00000000000000011000010000100111;
assign LUT_3[31973] = 32'b00000000000000011110111100000100;
assign LUT_3[31974] = 32'b00000000000000011010011000001011;
assign LUT_3[31975] = 32'b00000000000000100001000011101000;
assign LUT_3[31976] = 32'b00000000000000100000011011110111;
assign LUT_3[31977] = 32'b00000000000000100111000111010100;
assign LUT_3[31978] = 32'b00000000000000100010100011011011;
assign LUT_3[31979] = 32'b00000000000000101001001110111000;
assign LUT_3[31980] = 32'b00000000000000011101101001101101;
assign LUT_3[31981] = 32'b00000000000000100100010101001010;
assign LUT_3[31982] = 32'b00000000000000011111110001010001;
assign LUT_3[31983] = 32'b00000000000000100110011100101110;
assign LUT_3[31984] = 32'b00000000000000011110010101110100;
assign LUT_3[31985] = 32'b00000000000000100101000001010001;
assign LUT_3[31986] = 32'b00000000000000100000011101011000;
assign LUT_3[31987] = 32'b00000000000000100111001000110101;
assign LUT_3[31988] = 32'b00000000000000011011100011101010;
assign LUT_3[31989] = 32'b00000000000000100010001111000111;
assign LUT_3[31990] = 32'b00000000000000011101101011001110;
assign LUT_3[31991] = 32'b00000000000000100100010110101011;
assign LUT_3[31992] = 32'b00000000000000100011101110111010;
assign LUT_3[31993] = 32'b00000000000000101010011010010111;
assign LUT_3[31994] = 32'b00000000000000100101110110011110;
assign LUT_3[31995] = 32'b00000000000000101100100001111011;
assign LUT_3[31996] = 32'b00000000000000100000111100110000;
assign LUT_3[31997] = 32'b00000000000000100111101000001101;
assign LUT_3[31998] = 32'b00000000000000100011000100010100;
assign LUT_3[31999] = 32'b00000000000000101001101111110001;
assign LUT_3[32000] = 32'b00000000000000010100000000001001;
assign LUT_3[32001] = 32'b00000000000000011010101011100110;
assign LUT_3[32002] = 32'b00000000000000010110000111101101;
assign LUT_3[32003] = 32'b00000000000000011100110011001010;
assign LUT_3[32004] = 32'b00000000000000010001001101111111;
assign LUT_3[32005] = 32'b00000000000000010111111001011100;
assign LUT_3[32006] = 32'b00000000000000010011010101100011;
assign LUT_3[32007] = 32'b00000000000000011010000001000000;
assign LUT_3[32008] = 32'b00000000000000011001011001001111;
assign LUT_3[32009] = 32'b00000000000000100000000100101100;
assign LUT_3[32010] = 32'b00000000000000011011100000110011;
assign LUT_3[32011] = 32'b00000000000000100010001100010000;
assign LUT_3[32012] = 32'b00000000000000010110100111000101;
assign LUT_3[32013] = 32'b00000000000000011101010010100010;
assign LUT_3[32014] = 32'b00000000000000011000101110101001;
assign LUT_3[32015] = 32'b00000000000000011111011010000110;
assign LUT_3[32016] = 32'b00000000000000010111010011001100;
assign LUT_3[32017] = 32'b00000000000000011101111110101001;
assign LUT_3[32018] = 32'b00000000000000011001011010110000;
assign LUT_3[32019] = 32'b00000000000000100000000110001101;
assign LUT_3[32020] = 32'b00000000000000010100100001000010;
assign LUT_3[32021] = 32'b00000000000000011011001100011111;
assign LUT_3[32022] = 32'b00000000000000010110101000100110;
assign LUT_3[32023] = 32'b00000000000000011101010100000011;
assign LUT_3[32024] = 32'b00000000000000011100101100010010;
assign LUT_3[32025] = 32'b00000000000000100011010111101111;
assign LUT_3[32026] = 32'b00000000000000011110110011110110;
assign LUT_3[32027] = 32'b00000000000000100101011111010011;
assign LUT_3[32028] = 32'b00000000000000011001111010001000;
assign LUT_3[32029] = 32'b00000000000000100000100101100101;
assign LUT_3[32030] = 32'b00000000000000011100000001101100;
assign LUT_3[32031] = 32'b00000000000000100010101101001001;
assign LUT_3[32032] = 32'b00000000000000010101001110101001;
assign LUT_3[32033] = 32'b00000000000000011011111010000110;
assign LUT_3[32034] = 32'b00000000000000010111010110001101;
assign LUT_3[32035] = 32'b00000000000000011110000001101010;
assign LUT_3[32036] = 32'b00000000000000010010011100011111;
assign LUT_3[32037] = 32'b00000000000000011001000111111100;
assign LUT_3[32038] = 32'b00000000000000010100100100000011;
assign LUT_3[32039] = 32'b00000000000000011011001111100000;
assign LUT_3[32040] = 32'b00000000000000011010100111101111;
assign LUT_3[32041] = 32'b00000000000000100001010011001100;
assign LUT_3[32042] = 32'b00000000000000011100101111010011;
assign LUT_3[32043] = 32'b00000000000000100011011010110000;
assign LUT_3[32044] = 32'b00000000000000010111110101100101;
assign LUT_3[32045] = 32'b00000000000000011110100001000010;
assign LUT_3[32046] = 32'b00000000000000011001111101001001;
assign LUT_3[32047] = 32'b00000000000000100000101000100110;
assign LUT_3[32048] = 32'b00000000000000011000100001101100;
assign LUT_3[32049] = 32'b00000000000000011111001101001001;
assign LUT_3[32050] = 32'b00000000000000011010101001010000;
assign LUT_3[32051] = 32'b00000000000000100001010100101101;
assign LUT_3[32052] = 32'b00000000000000010101101111100010;
assign LUT_3[32053] = 32'b00000000000000011100011010111111;
assign LUT_3[32054] = 32'b00000000000000010111110111000110;
assign LUT_3[32055] = 32'b00000000000000011110100010100011;
assign LUT_3[32056] = 32'b00000000000000011101111010110010;
assign LUT_3[32057] = 32'b00000000000000100100100110001111;
assign LUT_3[32058] = 32'b00000000000000100000000010010110;
assign LUT_3[32059] = 32'b00000000000000100110101101110011;
assign LUT_3[32060] = 32'b00000000000000011011001000101000;
assign LUT_3[32061] = 32'b00000000000000100001110100000101;
assign LUT_3[32062] = 32'b00000000000000011101010000001100;
assign LUT_3[32063] = 32'b00000000000000100011111011101001;
assign LUT_3[32064] = 32'b00000000000000010011111000110100;
assign LUT_3[32065] = 32'b00000000000000011010100100010001;
assign LUT_3[32066] = 32'b00000000000000010110000000011000;
assign LUT_3[32067] = 32'b00000000000000011100101011110101;
assign LUT_3[32068] = 32'b00000000000000010001000110101010;
assign LUT_3[32069] = 32'b00000000000000010111110010000111;
assign LUT_3[32070] = 32'b00000000000000010011001110001110;
assign LUT_3[32071] = 32'b00000000000000011001111001101011;
assign LUT_3[32072] = 32'b00000000000000011001010001111010;
assign LUT_3[32073] = 32'b00000000000000011111111101010111;
assign LUT_3[32074] = 32'b00000000000000011011011001011110;
assign LUT_3[32075] = 32'b00000000000000100010000100111011;
assign LUT_3[32076] = 32'b00000000000000010110011111110000;
assign LUT_3[32077] = 32'b00000000000000011101001011001101;
assign LUT_3[32078] = 32'b00000000000000011000100111010100;
assign LUT_3[32079] = 32'b00000000000000011111010010110001;
assign LUT_3[32080] = 32'b00000000000000010111001011110111;
assign LUT_3[32081] = 32'b00000000000000011101110111010100;
assign LUT_3[32082] = 32'b00000000000000011001010011011011;
assign LUT_3[32083] = 32'b00000000000000011111111110111000;
assign LUT_3[32084] = 32'b00000000000000010100011001101101;
assign LUT_3[32085] = 32'b00000000000000011011000101001010;
assign LUT_3[32086] = 32'b00000000000000010110100001010001;
assign LUT_3[32087] = 32'b00000000000000011101001100101110;
assign LUT_3[32088] = 32'b00000000000000011100100100111101;
assign LUT_3[32089] = 32'b00000000000000100011010000011010;
assign LUT_3[32090] = 32'b00000000000000011110101100100001;
assign LUT_3[32091] = 32'b00000000000000100101010111111110;
assign LUT_3[32092] = 32'b00000000000000011001110010110011;
assign LUT_3[32093] = 32'b00000000000000100000011110010000;
assign LUT_3[32094] = 32'b00000000000000011011111010010111;
assign LUT_3[32095] = 32'b00000000000000100010100101110100;
assign LUT_3[32096] = 32'b00000000000000010101000111010100;
assign LUT_3[32097] = 32'b00000000000000011011110010110001;
assign LUT_3[32098] = 32'b00000000000000010111001110111000;
assign LUT_3[32099] = 32'b00000000000000011101111010010101;
assign LUT_3[32100] = 32'b00000000000000010010010101001010;
assign LUT_3[32101] = 32'b00000000000000011001000000100111;
assign LUT_3[32102] = 32'b00000000000000010100011100101110;
assign LUT_3[32103] = 32'b00000000000000011011001000001011;
assign LUT_3[32104] = 32'b00000000000000011010100000011010;
assign LUT_3[32105] = 32'b00000000000000100001001011110111;
assign LUT_3[32106] = 32'b00000000000000011100100111111110;
assign LUT_3[32107] = 32'b00000000000000100011010011011011;
assign LUT_3[32108] = 32'b00000000000000010111101110010000;
assign LUT_3[32109] = 32'b00000000000000011110011001101101;
assign LUT_3[32110] = 32'b00000000000000011001110101110100;
assign LUT_3[32111] = 32'b00000000000000100000100001010001;
assign LUT_3[32112] = 32'b00000000000000011000011010010111;
assign LUT_3[32113] = 32'b00000000000000011111000101110100;
assign LUT_3[32114] = 32'b00000000000000011010100001111011;
assign LUT_3[32115] = 32'b00000000000000100001001101011000;
assign LUT_3[32116] = 32'b00000000000000010101101000001101;
assign LUT_3[32117] = 32'b00000000000000011100010011101010;
assign LUT_3[32118] = 32'b00000000000000010111101111110001;
assign LUT_3[32119] = 32'b00000000000000011110011011001110;
assign LUT_3[32120] = 32'b00000000000000011101110011011101;
assign LUT_3[32121] = 32'b00000000000000100100011110111010;
assign LUT_3[32122] = 32'b00000000000000011111111011000001;
assign LUT_3[32123] = 32'b00000000000000100110100110011110;
assign LUT_3[32124] = 32'b00000000000000011011000001010011;
assign LUT_3[32125] = 32'b00000000000000100001101100110000;
assign LUT_3[32126] = 32'b00000000000000011101001000110111;
assign LUT_3[32127] = 32'b00000000000000100011110100010100;
assign LUT_3[32128] = 32'b00000000000000010110001011000111;
assign LUT_3[32129] = 32'b00000000000000011100110110100100;
assign LUT_3[32130] = 32'b00000000000000011000010010101011;
assign LUT_3[32131] = 32'b00000000000000011110111110001000;
assign LUT_3[32132] = 32'b00000000000000010011011000111101;
assign LUT_3[32133] = 32'b00000000000000011010000100011010;
assign LUT_3[32134] = 32'b00000000000000010101100000100001;
assign LUT_3[32135] = 32'b00000000000000011100001011111110;
assign LUT_3[32136] = 32'b00000000000000011011100100001101;
assign LUT_3[32137] = 32'b00000000000000100010001111101010;
assign LUT_3[32138] = 32'b00000000000000011101101011110001;
assign LUT_3[32139] = 32'b00000000000000100100010111001110;
assign LUT_3[32140] = 32'b00000000000000011000110010000011;
assign LUT_3[32141] = 32'b00000000000000011111011101100000;
assign LUT_3[32142] = 32'b00000000000000011010111001100111;
assign LUT_3[32143] = 32'b00000000000000100001100101000100;
assign LUT_3[32144] = 32'b00000000000000011001011110001010;
assign LUT_3[32145] = 32'b00000000000000100000001001100111;
assign LUT_3[32146] = 32'b00000000000000011011100101101110;
assign LUT_3[32147] = 32'b00000000000000100010010001001011;
assign LUT_3[32148] = 32'b00000000000000010110101100000000;
assign LUT_3[32149] = 32'b00000000000000011101010111011101;
assign LUT_3[32150] = 32'b00000000000000011000110011100100;
assign LUT_3[32151] = 32'b00000000000000011111011111000001;
assign LUT_3[32152] = 32'b00000000000000011110110111010000;
assign LUT_3[32153] = 32'b00000000000000100101100010101101;
assign LUT_3[32154] = 32'b00000000000000100000111110110100;
assign LUT_3[32155] = 32'b00000000000000100111101010010001;
assign LUT_3[32156] = 32'b00000000000000011100000101000110;
assign LUT_3[32157] = 32'b00000000000000100010110000100011;
assign LUT_3[32158] = 32'b00000000000000011110001100101010;
assign LUT_3[32159] = 32'b00000000000000100100111000000111;
assign LUT_3[32160] = 32'b00000000000000010111011001100111;
assign LUT_3[32161] = 32'b00000000000000011110000101000100;
assign LUT_3[32162] = 32'b00000000000000011001100001001011;
assign LUT_3[32163] = 32'b00000000000000100000001100101000;
assign LUT_3[32164] = 32'b00000000000000010100100111011101;
assign LUT_3[32165] = 32'b00000000000000011011010010111010;
assign LUT_3[32166] = 32'b00000000000000010110101111000001;
assign LUT_3[32167] = 32'b00000000000000011101011010011110;
assign LUT_3[32168] = 32'b00000000000000011100110010101101;
assign LUT_3[32169] = 32'b00000000000000100011011110001010;
assign LUT_3[32170] = 32'b00000000000000011110111010010001;
assign LUT_3[32171] = 32'b00000000000000100101100101101110;
assign LUT_3[32172] = 32'b00000000000000011010000000100011;
assign LUT_3[32173] = 32'b00000000000000100000101100000000;
assign LUT_3[32174] = 32'b00000000000000011100001000000111;
assign LUT_3[32175] = 32'b00000000000000100010110011100100;
assign LUT_3[32176] = 32'b00000000000000011010101100101010;
assign LUT_3[32177] = 32'b00000000000000100001011000000111;
assign LUT_3[32178] = 32'b00000000000000011100110100001110;
assign LUT_3[32179] = 32'b00000000000000100011011111101011;
assign LUT_3[32180] = 32'b00000000000000010111111010100000;
assign LUT_3[32181] = 32'b00000000000000011110100101111101;
assign LUT_3[32182] = 32'b00000000000000011010000010000100;
assign LUT_3[32183] = 32'b00000000000000100000101101100001;
assign LUT_3[32184] = 32'b00000000000000100000000101110000;
assign LUT_3[32185] = 32'b00000000000000100110110001001101;
assign LUT_3[32186] = 32'b00000000000000100010001101010100;
assign LUT_3[32187] = 32'b00000000000000101000111000110001;
assign LUT_3[32188] = 32'b00000000000000011101010011100110;
assign LUT_3[32189] = 32'b00000000000000100011111111000011;
assign LUT_3[32190] = 32'b00000000000000011111011011001010;
assign LUT_3[32191] = 32'b00000000000000100110000110100111;
assign LUT_3[32192] = 32'b00000000000000010110000011110010;
assign LUT_3[32193] = 32'b00000000000000011100101111001111;
assign LUT_3[32194] = 32'b00000000000000011000001011010110;
assign LUT_3[32195] = 32'b00000000000000011110110110110011;
assign LUT_3[32196] = 32'b00000000000000010011010001101000;
assign LUT_3[32197] = 32'b00000000000000011001111101000101;
assign LUT_3[32198] = 32'b00000000000000010101011001001100;
assign LUT_3[32199] = 32'b00000000000000011100000100101001;
assign LUT_3[32200] = 32'b00000000000000011011011100111000;
assign LUT_3[32201] = 32'b00000000000000100010001000010101;
assign LUT_3[32202] = 32'b00000000000000011101100100011100;
assign LUT_3[32203] = 32'b00000000000000100100001111111001;
assign LUT_3[32204] = 32'b00000000000000011000101010101110;
assign LUT_3[32205] = 32'b00000000000000011111010110001011;
assign LUT_3[32206] = 32'b00000000000000011010110010010010;
assign LUT_3[32207] = 32'b00000000000000100001011101101111;
assign LUT_3[32208] = 32'b00000000000000011001010110110101;
assign LUT_3[32209] = 32'b00000000000000100000000010010010;
assign LUT_3[32210] = 32'b00000000000000011011011110011001;
assign LUT_3[32211] = 32'b00000000000000100010001001110110;
assign LUT_3[32212] = 32'b00000000000000010110100100101011;
assign LUT_3[32213] = 32'b00000000000000011101010000001000;
assign LUT_3[32214] = 32'b00000000000000011000101100001111;
assign LUT_3[32215] = 32'b00000000000000011111010111101100;
assign LUT_3[32216] = 32'b00000000000000011110101111111011;
assign LUT_3[32217] = 32'b00000000000000100101011011011000;
assign LUT_3[32218] = 32'b00000000000000100000110111011111;
assign LUT_3[32219] = 32'b00000000000000100111100010111100;
assign LUT_3[32220] = 32'b00000000000000011011111101110001;
assign LUT_3[32221] = 32'b00000000000000100010101001001110;
assign LUT_3[32222] = 32'b00000000000000011110000101010101;
assign LUT_3[32223] = 32'b00000000000000100100110000110010;
assign LUT_3[32224] = 32'b00000000000000010111010010010010;
assign LUT_3[32225] = 32'b00000000000000011101111101101111;
assign LUT_3[32226] = 32'b00000000000000011001011001110110;
assign LUT_3[32227] = 32'b00000000000000100000000101010011;
assign LUT_3[32228] = 32'b00000000000000010100100000001000;
assign LUT_3[32229] = 32'b00000000000000011011001011100101;
assign LUT_3[32230] = 32'b00000000000000010110100111101100;
assign LUT_3[32231] = 32'b00000000000000011101010011001001;
assign LUT_3[32232] = 32'b00000000000000011100101011011000;
assign LUT_3[32233] = 32'b00000000000000100011010110110101;
assign LUT_3[32234] = 32'b00000000000000011110110010111100;
assign LUT_3[32235] = 32'b00000000000000100101011110011001;
assign LUT_3[32236] = 32'b00000000000000011001111001001110;
assign LUT_3[32237] = 32'b00000000000000100000100100101011;
assign LUT_3[32238] = 32'b00000000000000011100000000110010;
assign LUT_3[32239] = 32'b00000000000000100010101100001111;
assign LUT_3[32240] = 32'b00000000000000011010100101010101;
assign LUT_3[32241] = 32'b00000000000000100001010000110010;
assign LUT_3[32242] = 32'b00000000000000011100101100111001;
assign LUT_3[32243] = 32'b00000000000000100011011000010110;
assign LUT_3[32244] = 32'b00000000000000010111110011001011;
assign LUT_3[32245] = 32'b00000000000000011110011110101000;
assign LUT_3[32246] = 32'b00000000000000011001111010101111;
assign LUT_3[32247] = 32'b00000000000000100000100110001100;
assign LUT_3[32248] = 32'b00000000000000011111111110011011;
assign LUT_3[32249] = 32'b00000000000000100110101001111000;
assign LUT_3[32250] = 32'b00000000000000100010000101111111;
assign LUT_3[32251] = 32'b00000000000000101000110001011100;
assign LUT_3[32252] = 32'b00000000000000011101001100010001;
assign LUT_3[32253] = 32'b00000000000000100011110111101110;
assign LUT_3[32254] = 32'b00000000000000011111010011110101;
assign LUT_3[32255] = 32'b00000000000000100101111111010010;
assign LUT_3[32256] = 32'b00000000000000011011000101110100;
assign LUT_3[32257] = 32'b00000000000000100001110001010001;
assign LUT_3[32258] = 32'b00000000000000011101001101011000;
assign LUT_3[32259] = 32'b00000000000000100011111000110101;
assign LUT_3[32260] = 32'b00000000000000011000010011101010;
assign LUT_3[32261] = 32'b00000000000000011110111111000111;
assign LUT_3[32262] = 32'b00000000000000011010011011001110;
assign LUT_3[32263] = 32'b00000000000000100001000110101011;
assign LUT_3[32264] = 32'b00000000000000100000011110111010;
assign LUT_3[32265] = 32'b00000000000000100111001010010111;
assign LUT_3[32266] = 32'b00000000000000100010100110011110;
assign LUT_3[32267] = 32'b00000000000000101001010001111011;
assign LUT_3[32268] = 32'b00000000000000011101101100110000;
assign LUT_3[32269] = 32'b00000000000000100100011000001101;
assign LUT_3[32270] = 32'b00000000000000011111110100010100;
assign LUT_3[32271] = 32'b00000000000000100110011111110001;
assign LUT_3[32272] = 32'b00000000000000011110011000110111;
assign LUT_3[32273] = 32'b00000000000000100101000100010100;
assign LUT_3[32274] = 32'b00000000000000100000100000011011;
assign LUT_3[32275] = 32'b00000000000000100111001011111000;
assign LUT_3[32276] = 32'b00000000000000011011100110101101;
assign LUT_3[32277] = 32'b00000000000000100010010010001010;
assign LUT_3[32278] = 32'b00000000000000011101101110010001;
assign LUT_3[32279] = 32'b00000000000000100100011001101110;
assign LUT_3[32280] = 32'b00000000000000100011110001111101;
assign LUT_3[32281] = 32'b00000000000000101010011101011010;
assign LUT_3[32282] = 32'b00000000000000100101111001100001;
assign LUT_3[32283] = 32'b00000000000000101100100100111110;
assign LUT_3[32284] = 32'b00000000000000100000111111110011;
assign LUT_3[32285] = 32'b00000000000000100111101011010000;
assign LUT_3[32286] = 32'b00000000000000100011000111010111;
assign LUT_3[32287] = 32'b00000000000000101001110010110100;
assign LUT_3[32288] = 32'b00000000000000011100010100010100;
assign LUT_3[32289] = 32'b00000000000000100010111111110001;
assign LUT_3[32290] = 32'b00000000000000011110011011111000;
assign LUT_3[32291] = 32'b00000000000000100101000111010101;
assign LUT_3[32292] = 32'b00000000000000011001100010001010;
assign LUT_3[32293] = 32'b00000000000000100000001101100111;
assign LUT_3[32294] = 32'b00000000000000011011101001101110;
assign LUT_3[32295] = 32'b00000000000000100010010101001011;
assign LUT_3[32296] = 32'b00000000000000100001101101011010;
assign LUT_3[32297] = 32'b00000000000000101000011000110111;
assign LUT_3[32298] = 32'b00000000000000100011110100111110;
assign LUT_3[32299] = 32'b00000000000000101010100000011011;
assign LUT_3[32300] = 32'b00000000000000011110111011010000;
assign LUT_3[32301] = 32'b00000000000000100101100110101101;
assign LUT_3[32302] = 32'b00000000000000100001000010110100;
assign LUT_3[32303] = 32'b00000000000000100111101110010001;
assign LUT_3[32304] = 32'b00000000000000011111100111010111;
assign LUT_3[32305] = 32'b00000000000000100110010010110100;
assign LUT_3[32306] = 32'b00000000000000100001101110111011;
assign LUT_3[32307] = 32'b00000000000000101000011010011000;
assign LUT_3[32308] = 32'b00000000000000011100110101001101;
assign LUT_3[32309] = 32'b00000000000000100011100000101010;
assign LUT_3[32310] = 32'b00000000000000011110111100110001;
assign LUT_3[32311] = 32'b00000000000000100101101000001110;
assign LUT_3[32312] = 32'b00000000000000100101000000011101;
assign LUT_3[32313] = 32'b00000000000000101011101011111010;
assign LUT_3[32314] = 32'b00000000000000100111001000000001;
assign LUT_3[32315] = 32'b00000000000000101101110011011110;
assign LUT_3[32316] = 32'b00000000000000100010001110010011;
assign LUT_3[32317] = 32'b00000000000000101000111001110000;
assign LUT_3[32318] = 32'b00000000000000100100010101110111;
assign LUT_3[32319] = 32'b00000000000000101011000001010100;
assign LUT_3[32320] = 32'b00000000000000011010111110011111;
assign LUT_3[32321] = 32'b00000000000000100001101001111100;
assign LUT_3[32322] = 32'b00000000000000011101000110000011;
assign LUT_3[32323] = 32'b00000000000000100011110001100000;
assign LUT_3[32324] = 32'b00000000000000011000001100010101;
assign LUT_3[32325] = 32'b00000000000000011110110111110010;
assign LUT_3[32326] = 32'b00000000000000011010010011111001;
assign LUT_3[32327] = 32'b00000000000000100000111111010110;
assign LUT_3[32328] = 32'b00000000000000100000010111100101;
assign LUT_3[32329] = 32'b00000000000000100111000011000010;
assign LUT_3[32330] = 32'b00000000000000100010011111001001;
assign LUT_3[32331] = 32'b00000000000000101001001010100110;
assign LUT_3[32332] = 32'b00000000000000011101100101011011;
assign LUT_3[32333] = 32'b00000000000000100100010000111000;
assign LUT_3[32334] = 32'b00000000000000011111101100111111;
assign LUT_3[32335] = 32'b00000000000000100110011000011100;
assign LUT_3[32336] = 32'b00000000000000011110010001100010;
assign LUT_3[32337] = 32'b00000000000000100100111100111111;
assign LUT_3[32338] = 32'b00000000000000100000011001000110;
assign LUT_3[32339] = 32'b00000000000000100111000100100011;
assign LUT_3[32340] = 32'b00000000000000011011011111011000;
assign LUT_3[32341] = 32'b00000000000000100010001010110101;
assign LUT_3[32342] = 32'b00000000000000011101100110111100;
assign LUT_3[32343] = 32'b00000000000000100100010010011001;
assign LUT_3[32344] = 32'b00000000000000100011101010101000;
assign LUT_3[32345] = 32'b00000000000000101010010110000101;
assign LUT_3[32346] = 32'b00000000000000100101110010001100;
assign LUT_3[32347] = 32'b00000000000000101100011101101001;
assign LUT_3[32348] = 32'b00000000000000100000111000011110;
assign LUT_3[32349] = 32'b00000000000000100111100011111011;
assign LUT_3[32350] = 32'b00000000000000100011000000000010;
assign LUT_3[32351] = 32'b00000000000000101001101011011111;
assign LUT_3[32352] = 32'b00000000000000011100001100111111;
assign LUT_3[32353] = 32'b00000000000000100010111000011100;
assign LUT_3[32354] = 32'b00000000000000011110010100100011;
assign LUT_3[32355] = 32'b00000000000000100101000000000000;
assign LUT_3[32356] = 32'b00000000000000011001011010110101;
assign LUT_3[32357] = 32'b00000000000000100000000110010010;
assign LUT_3[32358] = 32'b00000000000000011011100010011001;
assign LUT_3[32359] = 32'b00000000000000100010001101110110;
assign LUT_3[32360] = 32'b00000000000000100001100110000101;
assign LUT_3[32361] = 32'b00000000000000101000010001100010;
assign LUT_3[32362] = 32'b00000000000000100011101101101001;
assign LUT_3[32363] = 32'b00000000000000101010011001000110;
assign LUT_3[32364] = 32'b00000000000000011110110011111011;
assign LUT_3[32365] = 32'b00000000000000100101011111011000;
assign LUT_3[32366] = 32'b00000000000000100000111011011111;
assign LUT_3[32367] = 32'b00000000000000100111100110111100;
assign LUT_3[32368] = 32'b00000000000000011111100000000010;
assign LUT_3[32369] = 32'b00000000000000100110001011011111;
assign LUT_3[32370] = 32'b00000000000000100001100111100110;
assign LUT_3[32371] = 32'b00000000000000101000010011000011;
assign LUT_3[32372] = 32'b00000000000000011100101101111000;
assign LUT_3[32373] = 32'b00000000000000100011011001010101;
assign LUT_3[32374] = 32'b00000000000000011110110101011100;
assign LUT_3[32375] = 32'b00000000000000100101100000111001;
assign LUT_3[32376] = 32'b00000000000000100100111001001000;
assign LUT_3[32377] = 32'b00000000000000101011100100100101;
assign LUT_3[32378] = 32'b00000000000000100111000000101100;
assign LUT_3[32379] = 32'b00000000000000101101101100001001;
assign LUT_3[32380] = 32'b00000000000000100010000110111110;
assign LUT_3[32381] = 32'b00000000000000101000110010011011;
assign LUT_3[32382] = 32'b00000000000000100100001110100010;
assign LUT_3[32383] = 32'b00000000000000101010111001111111;
assign LUT_3[32384] = 32'b00000000000000011101010000110010;
assign LUT_3[32385] = 32'b00000000000000100011111100001111;
assign LUT_3[32386] = 32'b00000000000000011111011000010110;
assign LUT_3[32387] = 32'b00000000000000100110000011110011;
assign LUT_3[32388] = 32'b00000000000000011010011110101000;
assign LUT_3[32389] = 32'b00000000000000100001001010000101;
assign LUT_3[32390] = 32'b00000000000000011100100110001100;
assign LUT_3[32391] = 32'b00000000000000100011010001101001;
assign LUT_3[32392] = 32'b00000000000000100010101001111000;
assign LUT_3[32393] = 32'b00000000000000101001010101010101;
assign LUT_3[32394] = 32'b00000000000000100100110001011100;
assign LUT_3[32395] = 32'b00000000000000101011011100111001;
assign LUT_3[32396] = 32'b00000000000000011111110111101110;
assign LUT_3[32397] = 32'b00000000000000100110100011001011;
assign LUT_3[32398] = 32'b00000000000000100001111111010010;
assign LUT_3[32399] = 32'b00000000000000101000101010101111;
assign LUT_3[32400] = 32'b00000000000000100000100011110101;
assign LUT_3[32401] = 32'b00000000000000100111001111010010;
assign LUT_3[32402] = 32'b00000000000000100010101011011001;
assign LUT_3[32403] = 32'b00000000000000101001010110110110;
assign LUT_3[32404] = 32'b00000000000000011101110001101011;
assign LUT_3[32405] = 32'b00000000000000100100011101001000;
assign LUT_3[32406] = 32'b00000000000000011111111001001111;
assign LUT_3[32407] = 32'b00000000000000100110100100101100;
assign LUT_3[32408] = 32'b00000000000000100101111100111011;
assign LUT_3[32409] = 32'b00000000000000101100101000011000;
assign LUT_3[32410] = 32'b00000000000000101000000100011111;
assign LUT_3[32411] = 32'b00000000000000101110101111111100;
assign LUT_3[32412] = 32'b00000000000000100011001010110001;
assign LUT_3[32413] = 32'b00000000000000101001110110001110;
assign LUT_3[32414] = 32'b00000000000000100101010010010101;
assign LUT_3[32415] = 32'b00000000000000101011111101110010;
assign LUT_3[32416] = 32'b00000000000000011110011111010010;
assign LUT_3[32417] = 32'b00000000000000100101001010101111;
assign LUT_3[32418] = 32'b00000000000000100000100110110110;
assign LUT_3[32419] = 32'b00000000000000100111010010010011;
assign LUT_3[32420] = 32'b00000000000000011011101101001000;
assign LUT_3[32421] = 32'b00000000000000100010011000100101;
assign LUT_3[32422] = 32'b00000000000000011101110100101100;
assign LUT_3[32423] = 32'b00000000000000100100100000001001;
assign LUT_3[32424] = 32'b00000000000000100011111000011000;
assign LUT_3[32425] = 32'b00000000000000101010100011110101;
assign LUT_3[32426] = 32'b00000000000000100101111111111100;
assign LUT_3[32427] = 32'b00000000000000101100101011011001;
assign LUT_3[32428] = 32'b00000000000000100001000110001110;
assign LUT_3[32429] = 32'b00000000000000100111110001101011;
assign LUT_3[32430] = 32'b00000000000000100011001101110010;
assign LUT_3[32431] = 32'b00000000000000101001111001001111;
assign LUT_3[32432] = 32'b00000000000000100001110010010101;
assign LUT_3[32433] = 32'b00000000000000101000011101110010;
assign LUT_3[32434] = 32'b00000000000000100011111001111001;
assign LUT_3[32435] = 32'b00000000000000101010100101010110;
assign LUT_3[32436] = 32'b00000000000000011111000000001011;
assign LUT_3[32437] = 32'b00000000000000100101101011101000;
assign LUT_3[32438] = 32'b00000000000000100001000111101111;
assign LUT_3[32439] = 32'b00000000000000100111110011001100;
assign LUT_3[32440] = 32'b00000000000000100111001011011011;
assign LUT_3[32441] = 32'b00000000000000101101110110111000;
assign LUT_3[32442] = 32'b00000000000000101001010010111111;
assign LUT_3[32443] = 32'b00000000000000101111111110011100;
assign LUT_3[32444] = 32'b00000000000000100100011001010001;
assign LUT_3[32445] = 32'b00000000000000101011000100101110;
assign LUT_3[32446] = 32'b00000000000000100110100000110101;
assign LUT_3[32447] = 32'b00000000000000101101001100010010;
assign LUT_3[32448] = 32'b00000000000000011101001001011101;
assign LUT_3[32449] = 32'b00000000000000100011110100111010;
assign LUT_3[32450] = 32'b00000000000000011111010001000001;
assign LUT_3[32451] = 32'b00000000000000100101111100011110;
assign LUT_3[32452] = 32'b00000000000000011010010111010011;
assign LUT_3[32453] = 32'b00000000000000100001000010110000;
assign LUT_3[32454] = 32'b00000000000000011100011110110111;
assign LUT_3[32455] = 32'b00000000000000100011001010010100;
assign LUT_3[32456] = 32'b00000000000000100010100010100011;
assign LUT_3[32457] = 32'b00000000000000101001001110000000;
assign LUT_3[32458] = 32'b00000000000000100100101010000111;
assign LUT_3[32459] = 32'b00000000000000101011010101100100;
assign LUT_3[32460] = 32'b00000000000000011111110000011001;
assign LUT_3[32461] = 32'b00000000000000100110011011110110;
assign LUT_3[32462] = 32'b00000000000000100001110111111101;
assign LUT_3[32463] = 32'b00000000000000101000100011011010;
assign LUT_3[32464] = 32'b00000000000000100000011100100000;
assign LUT_3[32465] = 32'b00000000000000100111000111111101;
assign LUT_3[32466] = 32'b00000000000000100010100100000100;
assign LUT_3[32467] = 32'b00000000000000101001001111100001;
assign LUT_3[32468] = 32'b00000000000000011101101010010110;
assign LUT_3[32469] = 32'b00000000000000100100010101110011;
assign LUT_3[32470] = 32'b00000000000000011111110001111010;
assign LUT_3[32471] = 32'b00000000000000100110011101010111;
assign LUT_3[32472] = 32'b00000000000000100101110101100110;
assign LUT_3[32473] = 32'b00000000000000101100100001000011;
assign LUT_3[32474] = 32'b00000000000000100111111101001010;
assign LUT_3[32475] = 32'b00000000000000101110101000100111;
assign LUT_3[32476] = 32'b00000000000000100011000011011100;
assign LUT_3[32477] = 32'b00000000000000101001101110111001;
assign LUT_3[32478] = 32'b00000000000000100101001011000000;
assign LUT_3[32479] = 32'b00000000000000101011110110011101;
assign LUT_3[32480] = 32'b00000000000000011110010111111101;
assign LUT_3[32481] = 32'b00000000000000100101000011011010;
assign LUT_3[32482] = 32'b00000000000000100000011111100001;
assign LUT_3[32483] = 32'b00000000000000100111001010111110;
assign LUT_3[32484] = 32'b00000000000000011011100101110011;
assign LUT_3[32485] = 32'b00000000000000100010010001010000;
assign LUT_3[32486] = 32'b00000000000000011101101101010111;
assign LUT_3[32487] = 32'b00000000000000100100011000110100;
assign LUT_3[32488] = 32'b00000000000000100011110001000011;
assign LUT_3[32489] = 32'b00000000000000101010011100100000;
assign LUT_3[32490] = 32'b00000000000000100101111000100111;
assign LUT_3[32491] = 32'b00000000000000101100100100000100;
assign LUT_3[32492] = 32'b00000000000000100000111110111001;
assign LUT_3[32493] = 32'b00000000000000100111101010010110;
assign LUT_3[32494] = 32'b00000000000000100011000110011101;
assign LUT_3[32495] = 32'b00000000000000101001110001111010;
assign LUT_3[32496] = 32'b00000000000000100001101011000000;
assign LUT_3[32497] = 32'b00000000000000101000010110011101;
assign LUT_3[32498] = 32'b00000000000000100011110010100100;
assign LUT_3[32499] = 32'b00000000000000101010011110000001;
assign LUT_3[32500] = 32'b00000000000000011110111000110110;
assign LUT_3[32501] = 32'b00000000000000100101100100010011;
assign LUT_3[32502] = 32'b00000000000000100001000000011010;
assign LUT_3[32503] = 32'b00000000000000100111101011110111;
assign LUT_3[32504] = 32'b00000000000000100111000100000110;
assign LUT_3[32505] = 32'b00000000000000101101101111100011;
assign LUT_3[32506] = 32'b00000000000000101001001011101010;
assign LUT_3[32507] = 32'b00000000000000101111110111000111;
assign LUT_3[32508] = 32'b00000000000000100100010001111100;
assign LUT_3[32509] = 32'b00000000000000101010111101011001;
assign LUT_3[32510] = 32'b00000000000000100110011001100000;
assign LUT_3[32511] = 32'b00000000000000101101000100111101;
assign LUT_3[32512] = 32'b00000000000000010111010101010101;
assign LUT_3[32513] = 32'b00000000000000011110000000110010;
assign LUT_3[32514] = 32'b00000000000000011001011100111001;
assign LUT_3[32515] = 32'b00000000000000100000001000010110;
assign LUT_3[32516] = 32'b00000000000000010100100011001011;
assign LUT_3[32517] = 32'b00000000000000011011001110101000;
assign LUT_3[32518] = 32'b00000000000000010110101010101111;
assign LUT_3[32519] = 32'b00000000000000011101010110001100;
assign LUT_3[32520] = 32'b00000000000000011100101110011011;
assign LUT_3[32521] = 32'b00000000000000100011011001111000;
assign LUT_3[32522] = 32'b00000000000000011110110101111111;
assign LUT_3[32523] = 32'b00000000000000100101100001011100;
assign LUT_3[32524] = 32'b00000000000000011001111100010001;
assign LUT_3[32525] = 32'b00000000000000100000100111101110;
assign LUT_3[32526] = 32'b00000000000000011100000011110101;
assign LUT_3[32527] = 32'b00000000000000100010101111010010;
assign LUT_3[32528] = 32'b00000000000000011010101000011000;
assign LUT_3[32529] = 32'b00000000000000100001010011110101;
assign LUT_3[32530] = 32'b00000000000000011100101111111100;
assign LUT_3[32531] = 32'b00000000000000100011011011011001;
assign LUT_3[32532] = 32'b00000000000000010111110110001110;
assign LUT_3[32533] = 32'b00000000000000011110100001101011;
assign LUT_3[32534] = 32'b00000000000000011001111101110010;
assign LUT_3[32535] = 32'b00000000000000100000101001001111;
assign LUT_3[32536] = 32'b00000000000000100000000001011110;
assign LUT_3[32537] = 32'b00000000000000100110101100111011;
assign LUT_3[32538] = 32'b00000000000000100010001001000010;
assign LUT_3[32539] = 32'b00000000000000101000110100011111;
assign LUT_3[32540] = 32'b00000000000000011101001111010100;
assign LUT_3[32541] = 32'b00000000000000100011111010110001;
assign LUT_3[32542] = 32'b00000000000000011111010110111000;
assign LUT_3[32543] = 32'b00000000000000100110000010010101;
assign LUT_3[32544] = 32'b00000000000000011000100011110101;
assign LUT_3[32545] = 32'b00000000000000011111001111010010;
assign LUT_3[32546] = 32'b00000000000000011010101011011001;
assign LUT_3[32547] = 32'b00000000000000100001010110110110;
assign LUT_3[32548] = 32'b00000000000000010101110001101011;
assign LUT_3[32549] = 32'b00000000000000011100011101001000;
assign LUT_3[32550] = 32'b00000000000000010111111001001111;
assign LUT_3[32551] = 32'b00000000000000011110100100101100;
assign LUT_3[32552] = 32'b00000000000000011101111100111011;
assign LUT_3[32553] = 32'b00000000000000100100101000011000;
assign LUT_3[32554] = 32'b00000000000000100000000100011111;
assign LUT_3[32555] = 32'b00000000000000100110101111111100;
assign LUT_3[32556] = 32'b00000000000000011011001010110001;
assign LUT_3[32557] = 32'b00000000000000100001110110001110;
assign LUT_3[32558] = 32'b00000000000000011101010010010101;
assign LUT_3[32559] = 32'b00000000000000100011111101110010;
assign LUT_3[32560] = 32'b00000000000000011011110110111000;
assign LUT_3[32561] = 32'b00000000000000100010100010010101;
assign LUT_3[32562] = 32'b00000000000000011101111110011100;
assign LUT_3[32563] = 32'b00000000000000100100101001111001;
assign LUT_3[32564] = 32'b00000000000000011001000100101110;
assign LUT_3[32565] = 32'b00000000000000011111110000001011;
assign LUT_3[32566] = 32'b00000000000000011011001100010010;
assign LUT_3[32567] = 32'b00000000000000100001110111101111;
assign LUT_3[32568] = 32'b00000000000000100001001111111110;
assign LUT_3[32569] = 32'b00000000000000100111111011011011;
assign LUT_3[32570] = 32'b00000000000000100011010111100010;
assign LUT_3[32571] = 32'b00000000000000101010000010111111;
assign LUT_3[32572] = 32'b00000000000000011110011101110100;
assign LUT_3[32573] = 32'b00000000000000100101001001010001;
assign LUT_3[32574] = 32'b00000000000000100000100101011000;
assign LUT_3[32575] = 32'b00000000000000100111010000110101;
assign LUT_3[32576] = 32'b00000000000000010111001110000000;
assign LUT_3[32577] = 32'b00000000000000011101111001011101;
assign LUT_3[32578] = 32'b00000000000000011001010101100100;
assign LUT_3[32579] = 32'b00000000000000100000000001000001;
assign LUT_3[32580] = 32'b00000000000000010100011011110110;
assign LUT_3[32581] = 32'b00000000000000011011000111010011;
assign LUT_3[32582] = 32'b00000000000000010110100011011010;
assign LUT_3[32583] = 32'b00000000000000011101001110110111;
assign LUT_3[32584] = 32'b00000000000000011100100111000110;
assign LUT_3[32585] = 32'b00000000000000100011010010100011;
assign LUT_3[32586] = 32'b00000000000000011110101110101010;
assign LUT_3[32587] = 32'b00000000000000100101011010000111;
assign LUT_3[32588] = 32'b00000000000000011001110100111100;
assign LUT_3[32589] = 32'b00000000000000100000100000011001;
assign LUT_3[32590] = 32'b00000000000000011011111100100000;
assign LUT_3[32591] = 32'b00000000000000100010100111111101;
assign LUT_3[32592] = 32'b00000000000000011010100001000011;
assign LUT_3[32593] = 32'b00000000000000100001001100100000;
assign LUT_3[32594] = 32'b00000000000000011100101000100111;
assign LUT_3[32595] = 32'b00000000000000100011010100000100;
assign LUT_3[32596] = 32'b00000000000000010111101110111001;
assign LUT_3[32597] = 32'b00000000000000011110011010010110;
assign LUT_3[32598] = 32'b00000000000000011001110110011101;
assign LUT_3[32599] = 32'b00000000000000100000100001111010;
assign LUT_3[32600] = 32'b00000000000000011111111010001001;
assign LUT_3[32601] = 32'b00000000000000100110100101100110;
assign LUT_3[32602] = 32'b00000000000000100010000001101101;
assign LUT_3[32603] = 32'b00000000000000101000101101001010;
assign LUT_3[32604] = 32'b00000000000000011101000111111111;
assign LUT_3[32605] = 32'b00000000000000100011110011011100;
assign LUT_3[32606] = 32'b00000000000000011111001111100011;
assign LUT_3[32607] = 32'b00000000000000100101111011000000;
assign LUT_3[32608] = 32'b00000000000000011000011100100000;
assign LUT_3[32609] = 32'b00000000000000011111000111111101;
assign LUT_3[32610] = 32'b00000000000000011010100100000100;
assign LUT_3[32611] = 32'b00000000000000100001001111100001;
assign LUT_3[32612] = 32'b00000000000000010101101010010110;
assign LUT_3[32613] = 32'b00000000000000011100010101110011;
assign LUT_3[32614] = 32'b00000000000000010111110001111010;
assign LUT_3[32615] = 32'b00000000000000011110011101010111;
assign LUT_3[32616] = 32'b00000000000000011101110101100110;
assign LUT_3[32617] = 32'b00000000000000100100100001000011;
assign LUT_3[32618] = 32'b00000000000000011111111101001010;
assign LUT_3[32619] = 32'b00000000000000100110101000100111;
assign LUT_3[32620] = 32'b00000000000000011011000011011100;
assign LUT_3[32621] = 32'b00000000000000100001101110111001;
assign LUT_3[32622] = 32'b00000000000000011101001011000000;
assign LUT_3[32623] = 32'b00000000000000100011110110011101;
assign LUT_3[32624] = 32'b00000000000000011011101111100011;
assign LUT_3[32625] = 32'b00000000000000100010011011000000;
assign LUT_3[32626] = 32'b00000000000000011101110111000111;
assign LUT_3[32627] = 32'b00000000000000100100100010100100;
assign LUT_3[32628] = 32'b00000000000000011000111101011001;
assign LUT_3[32629] = 32'b00000000000000011111101000110110;
assign LUT_3[32630] = 32'b00000000000000011011000100111101;
assign LUT_3[32631] = 32'b00000000000000100001110000011010;
assign LUT_3[32632] = 32'b00000000000000100001001000101001;
assign LUT_3[32633] = 32'b00000000000000100111110100000110;
assign LUT_3[32634] = 32'b00000000000000100011010000001101;
assign LUT_3[32635] = 32'b00000000000000101001111011101010;
assign LUT_3[32636] = 32'b00000000000000011110010110011111;
assign LUT_3[32637] = 32'b00000000000000100101000001111100;
assign LUT_3[32638] = 32'b00000000000000100000011110000011;
assign LUT_3[32639] = 32'b00000000000000100111001001100000;
assign LUT_3[32640] = 32'b00000000000000011001100000010011;
assign LUT_3[32641] = 32'b00000000000000100000001011110000;
assign LUT_3[32642] = 32'b00000000000000011011100111110111;
assign LUT_3[32643] = 32'b00000000000000100010010011010100;
assign LUT_3[32644] = 32'b00000000000000010110101110001001;
assign LUT_3[32645] = 32'b00000000000000011101011001100110;
assign LUT_3[32646] = 32'b00000000000000011000110101101101;
assign LUT_3[32647] = 32'b00000000000000011111100001001010;
assign LUT_3[32648] = 32'b00000000000000011110111001011001;
assign LUT_3[32649] = 32'b00000000000000100101100100110110;
assign LUT_3[32650] = 32'b00000000000000100001000000111101;
assign LUT_3[32651] = 32'b00000000000000100111101100011010;
assign LUT_3[32652] = 32'b00000000000000011100000111001111;
assign LUT_3[32653] = 32'b00000000000000100010110010101100;
assign LUT_3[32654] = 32'b00000000000000011110001110110011;
assign LUT_3[32655] = 32'b00000000000000100100111010010000;
assign LUT_3[32656] = 32'b00000000000000011100110011010110;
assign LUT_3[32657] = 32'b00000000000000100011011110110011;
assign LUT_3[32658] = 32'b00000000000000011110111010111010;
assign LUT_3[32659] = 32'b00000000000000100101100110010111;
assign LUT_3[32660] = 32'b00000000000000011010000001001100;
assign LUT_3[32661] = 32'b00000000000000100000101100101001;
assign LUT_3[32662] = 32'b00000000000000011100001000110000;
assign LUT_3[32663] = 32'b00000000000000100010110100001101;
assign LUT_3[32664] = 32'b00000000000000100010001100011100;
assign LUT_3[32665] = 32'b00000000000000101000110111111001;
assign LUT_3[32666] = 32'b00000000000000100100010100000000;
assign LUT_3[32667] = 32'b00000000000000101010111111011101;
assign LUT_3[32668] = 32'b00000000000000011111011010010010;
assign LUT_3[32669] = 32'b00000000000000100110000101101111;
assign LUT_3[32670] = 32'b00000000000000100001100001110110;
assign LUT_3[32671] = 32'b00000000000000101000001101010011;
assign LUT_3[32672] = 32'b00000000000000011010101110110011;
assign LUT_3[32673] = 32'b00000000000000100001011010010000;
assign LUT_3[32674] = 32'b00000000000000011100110110010111;
assign LUT_3[32675] = 32'b00000000000000100011100001110100;
assign LUT_3[32676] = 32'b00000000000000010111111100101001;
assign LUT_3[32677] = 32'b00000000000000011110101000000110;
assign LUT_3[32678] = 32'b00000000000000011010000100001101;
assign LUT_3[32679] = 32'b00000000000000100000101111101010;
assign LUT_3[32680] = 32'b00000000000000100000000111111001;
assign LUT_3[32681] = 32'b00000000000000100110110011010110;
assign LUT_3[32682] = 32'b00000000000000100010001111011101;
assign LUT_3[32683] = 32'b00000000000000101000111010111010;
assign LUT_3[32684] = 32'b00000000000000011101010101101111;
assign LUT_3[32685] = 32'b00000000000000100100000001001100;
assign LUT_3[32686] = 32'b00000000000000011111011101010011;
assign LUT_3[32687] = 32'b00000000000000100110001000110000;
assign LUT_3[32688] = 32'b00000000000000011110000001110110;
assign LUT_3[32689] = 32'b00000000000000100100101101010011;
assign LUT_3[32690] = 32'b00000000000000100000001001011010;
assign LUT_3[32691] = 32'b00000000000000100110110100110111;
assign LUT_3[32692] = 32'b00000000000000011011001111101100;
assign LUT_3[32693] = 32'b00000000000000100001111011001001;
assign LUT_3[32694] = 32'b00000000000000011101010111010000;
assign LUT_3[32695] = 32'b00000000000000100100000010101101;
assign LUT_3[32696] = 32'b00000000000000100011011010111100;
assign LUT_3[32697] = 32'b00000000000000101010000110011001;
assign LUT_3[32698] = 32'b00000000000000100101100010100000;
assign LUT_3[32699] = 32'b00000000000000101100001101111101;
assign LUT_3[32700] = 32'b00000000000000100000101000110010;
assign LUT_3[32701] = 32'b00000000000000100111010100001111;
assign LUT_3[32702] = 32'b00000000000000100010110000010110;
assign LUT_3[32703] = 32'b00000000000000101001011011110011;
assign LUT_3[32704] = 32'b00000000000000011001011000111110;
assign LUT_3[32705] = 32'b00000000000000100000000100011011;
assign LUT_3[32706] = 32'b00000000000000011011100000100010;
assign LUT_3[32707] = 32'b00000000000000100010001011111111;
assign LUT_3[32708] = 32'b00000000000000010110100110110100;
assign LUT_3[32709] = 32'b00000000000000011101010010010001;
assign LUT_3[32710] = 32'b00000000000000011000101110011000;
assign LUT_3[32711] = 32'b00000000000000011111011001110101;
assign LUT_3[32712] = 32'b00000000000000011110110010000100;
assign LUT_3[32713] = 32'b00000000000000100101011101100001;
assign LUT_3[32714] = 32'b00000000000000100000111001101000;
assign LUT_3[32715] = 32'b00000000000000100111100101000101;
assign LUT_3[32716] = 32'b00000000000000011011111111111010;
assign LUT_3[32717] = 32'b00000000000000100010101011010111;
assign LUT_3[32718] = 32'b00000000000000011110000111011110;
assign LUT_3[32719] = 32'b00000000000000100100110010111011;
assign LUT_3[32720] = 32'b00000000000000011100101100000001;
assign LUT_3[32721] = 32'b00000000000000100011010111011110;
assign LUT_3[32722] = 32'b00000000000000011110110011100101;
assign LUT_3[32723] = 32'b00000000000000100101011111000010;
assign LUT_3[32724] = 32'b00000000000000011001111001110111;
assign LUT_3[32725] = 32'b00000000000000100000100101010100;
assign LUT_3[32726] = 32'b00000000000000011100000001011011;
assign LUT_3[32727] = 32'b00000000000000100010101100111000;
assign LUT_3[32728] = 32'b00000000000000100010000101000111;
assign LUT_3[32729] = 32'b00000000000000101000110000100100;
assign LUT_3[32730] = 32'b00000000000000100100001100101011;
assign LUT_3[32731] = 32'b00000000000000101010111000001000;
assign LUT_3[32732] = 32'b00000000000000011111010010111101;
assign LUT_3[32733] = 32'b00000000000000100101111110011010;
assign LUT_3[32734] = 32'b00000000000000100001011010100001;
assign LUT_3[32735] = 32'b00000000000000101000000101111110;
assign LUT_3[32736] = 32'b00000000000000011010100111011110;
assign LUT_3[32737] = 32'b00000000000000100001010010111011;
assign LUT_3[32738] = 32'b00000000000000011100101111000010;
assign LUT_3[32739] = 32'b00000000000000100011011010011111;
assign LUT_3[32740] = 32'b00000000000000010111110101010100;
assign LUT_3[32741] = 32'b00000000000000011110100000110001;
assign LUT_3[32742] = 32'b00000000000000011001111100111000;
assign LUT_3[32743] = 32'b00000000000000100000101000010101;
assign LUT_3[32744] = 32'b00000000000000100000000000100100;
assign LUT_3[32745] = 32'b00000000000000100110101100000001;
assign LUT_3[32746] = 32'b00000000000000100010001000001000;
assign LUT_3[32747] = 32'b00000000000000101000110011100101;
assign LUT_3[32748] = 32'b00000000000000011101001110011010;
assign LUT_3[32749] = 32'b00000000000000100011111001110111;
assign LUT_3[32750] = 32'b00000000000000011111010101111110;
assign LUT_3[32751] = 32'b00000000000000100110000001011011;
assign LUT_3[32752] = 32'b00000000000000011101111010100001;
assign LUT_3[32753] = 32'b00000000000000100100100101111110;
assign LUT_3[32754] = 32'b00000000000000100000000010000101;
assign LUT_3[32755] = 32'b00000000000000100110101101100010;
assign LUT_3[32756] = 32'b00000000000000011011001000010111;
assign LUT_3[32757] = 32'b00000000000000100001110011110100;
assign LUT_3[32758] = 32'b00000000000000011101001111111011;
assign LUT_3[32759] = 32'b00000000000000100011111011011000;
assign LUT_3[32760] = 32'b00000000000000100011010011100111;
assign LUT_3[32761] = 32'b00000000000000101001111111000100;
assign LUT_3[32762] = 32'b00000000000000100101011011001011;
assign LUT_3[32763] = 32'b00000000000000101100000110101000;
assign LUT_3[32764] = 32'b00000000000000100000100001011101;
assign LUT_3[32765] = 32'b00000000000000100111001100111010;
assign LUT_3[32766] = 32'b00000000000000100010101001000001;
assign LUT_3[32767] = 32'b00000000000000101001010100011110;
assign LUT_3[32768] = 32'b11111111111111111000100001011110;
assign LUT_3[32769] = 32'b11111111111111111111001100111011;
assign LUT_3[32770] = 32'b11111111111111111010101001000010;
assign LUT_3[32771] = 32'b00000000000000000001010100011111;
assign LUT_3[32772] = 32'b11111111111111110101101111010100;
assign LUT_3[32773] = 32'b11111111111111111100011010110001;
assign LUT_3[32774] = 32'b11111111111111110111110110111000;
assign LUT_3[32775] = 32'b11111111111111111110100010010101;
assign LUT_3[32776] = 32'b11111111111111111101111010100100;
assign LUT_3[32777] = 32'b00000000000000000100100110000001;
assign LUT_3[32778] = 32'b00000000000000000000000010001000;
assign LUT_3[32779] = 32'b00000000000000000110101101100101;
assign LUT_3[32780] = 32'b11111111111111111011001000011010;
assign LUT_3[32781] = 32'b00000000000000000001110011110111;
assign LUT_3[32782] = 32'b11111111111111111101001111111110;
assign LUT_3[32783] = 32'b00000000000000000011111011011011;
assign LUT_3[32784] = 32'b11111111111111111011110100100001;
assign LUT_3[32785] = 32'b00000000000000000010011111111110;
assign LUT_3[32786] = 32'b11111111111111111101111100000101;
assign LUT_3[32787] = 32'b00000000000000000100100111100010;
assign LUT_3[32788] = 32'b11111111111111111001000010010111;
assign LUT_3[32789] = 32'b11111111111111111111101101110100;
assign LUT_3[32790] = 32'b11111111111111111011001001111011;
assign LUT_3[32791] = 32'b00000000000000000001110101011000;
assign LUT_3[32792] = 32'b00000000000000000001001101100111;
assign LUT_3[32793] = 32'b00000000000000000111111001000100;
assign LUT_3[32794] = 32'b00000000000000000011010101001011;
assign LUT_3[32795] = 32'b00000000000000001010000000101000;
assign LUT_3[32796] = 32'b11111111111111111110011011011101;
assign LUT_3[32797] = 32'b00000000000000000101000110111010;
assign LUT_3[32798] = 32'b00000000000000000000100011000001;
assign LUT_3[32799] = 32'b00000000000000000111001110011110;
assign LUT_3[32800] = 32'b11111111111111111001101111111110;
assign LUT_3[32801] = 32'b00000000000000000000011011011011;
assign LUT_3[32802] = 32'b11111111111111111011110111100010;
assign LUT_3[32803] = 32'b00000000000000000010100010111111;
assign LUT_3[32804] = 32'b11111111111111110110111101110100;
assign LUT_3[32805] = 32'b11111111111111111101101001010001;
assign LUT_3[32806] = 32'b11111111111111111001000101011000;
assign LUT_3[32807] = 32'b11111111111111111111110000110101;
assign LUT_3[32808] = 32'b11111111111111111111001001000100;
assign LUT_3[32809] = 32'b00000000000000000101110100100001;
assign LUT_3[32810] = 32'b00000000000000000001010000101000;
assign LUT_3[32811] = 32'b00000000000000000111111100000101;
assign LUT_3[32812] = 32'b11111111111111111100010110111010;
assign LUT_3[32813] = 32'b00000000000000000011000010010111;
assign LUT_3[32814] = 32'b11111111111111111110011110011110;
assign LUT_3[32815] = 32'b00000000000000000101001001111011;
assign LUT_3[32816] = 32'b11111111111111111101000011000001;
assign LUT_3[32817] = 32'b00000000000000000011101110011110;
assign LUT_3[32818] = 32'b11111111111111111111001010100101;
assign LUT_3[32819] = 32'b00000000000000000101110110000010;
assign LUT_3[32820] = 32'b11111111111111111010010000110111;
assign LUT_3[32821] = 32'b00000000000000000000111100010100;
assign LUT_3[32822] = 32'b11111111111111111100011000011011;
assign LUT_3[32823] = 32'b00000000000000000011000011111000;
assign LUT_3[32824] = 32'b00000000000000000010011100000111;
assign LUT_3[32825] = 32'b00000000000000001001000111100100;
assign LUT_3[32826] = 32'b00000000000000000100100011101011;
assign LUT_3[32827] = 32'b00000000000000001011001111001000;
assign LUT_3[32828] = 32'b11111111111111111111101001111101;
assign LUT_3[32829] = 32'b00000000000000000110010101011010;
assign LUT_3[32830] = 32'b00000000000000000001110001100001;
assign LUT_3[32831] = 32'b00000000000000001000011100111110;
assign LUT_3[32832] = 32'b11111111111111111000011010001001;
assign LUT_3[32833] = 32'b11111111111111111111000101100110;
assign LUT_3[32834] = 32'b11111111111111111010100001101101;
assign LUT_3[32835] = 32'b00000000000000000001001101001010;
assign LUT_3[32836] = 32'b11111111111111110101100111111111;
assign LUT_3[32837] = 32'b11111111111111111100010011011100;
assign LUT_3[32838] = 32'b11111111111111110111101111100011;
assign LUT_3[32839] = 32'b11111111111111111110011011000000;
assign LUT_3[32840] = 32'b11111111111111111101110011001111;
assign LUT_3[32841] = 32'b00000000000000000100011110101100;
assign LUT_3[32842] = 32'b11111111111111111111111010110011;
assign LUT_3[32843] = 32'b00000000000000000110100110010000;
assign LUT_3[32844] = 32'b11111111111111111011000001000101;
assign LUT_3[32845] = 32'b00000000000000000001101100100010;
assign LUT_3[32846] = 32'b11111111111111111101001000101001;
assign LUT_3[32847] = 32'b00000000000000000011110100000110;
assign LUT_3[32848] = 32'b11111111111111111011101101001100;
assign LUT_3[32849] = 32'b00000000000000000010011000101001;
assign LUT_3[32850] = 32'b11111111111111111101110100110000;
assign LUT_3[32851] = 32'b00000000000000000100100000001101;
assign LUT_3[32852] = 32'b11111111111111111000111011000010;
assign LUT_3[32853] = 32'b11111111111111111111100110011111;
assign LUT_3[32854] = 32'b11111111111111111011000010100110;
assign LUT_3[32855] = 32'b00000000000000000001101110000011;
assign LUT_3[32856] = 32'b00000000000000000001000110010010;
assign LUT_3[32857] = 32'b00000000000000000111110001101111;
assign LUT_3[32858] = 32'b00000000000000000011001101110110;
assign LUT_3[32859] = 32'b00000000000000001001111001010011;
assign LUT_3[32860] = 32'b11111111111111111110010100001000;
assign LUT_3[32861] = 32'b00000000000000000100111111100101;
assign LUT_3[32862] = 32'b00000000000000000000011011101100;
assign LUT_3[32863] = 32'b00000000000000000111000111001001;
assign LUT_3[32864] = 32'b11111111111111111001101000101001;
assign LUT_3[32865] = 32'b00000000000000000000010100000110;
assign LUT_3[32866] = 32'b11111111111111111011110000001101;
assign LUT_3[32867] = 32'b00000000000000000010011011101010;
assign LUT_3[32868] = 32'b11111111111111110110110110011111;
assign LUT_3[32869] = 32'b11111111111111111101100001111100;
assign LUT_3[32870] = 32'b11111111111111111000111110000011;
assign LUT_3[32871] = 32'b11111111111111111111101001100000;
assign LUT_3[32872] = 32'b11111111111111111111000001101111;
assign LUT_3[32873] = 32'b00000000000000000101101101001100;
assign LUT_3[32874] = 32'b00000000000000000001001001010011;
assign LUT_3[32875] = 32'b00000000000000000111110100110000;
assign LUT_3[32876] = 32'b11111111111111111100001111100101;
assign LUT_3[32877] = 32'b00000000000000000010111011000010;
assign LUT_3[32878] = 32'b11111111111111111110010111001001;
assign LUT_3[32879] = 32'b00000000000000000101000010100110;
assign LUT_3[32880] = 32'b11111111111111111100111011101100;
assign LUT_3[32881] = 32'b00000000000000000011100111001001;
assign LUT_3[32882] = 32'b11111111111111111111000011010000;
assign LUT_3[32883] = 32'b00000000000000000101101110101101;
assign LUT_3[32884] = 32'b11111111111111111010001001100010;
assign LUT_3[32885] = 32'b00000000000000000000110100111111;
assign LUT_3[32886] = 32'b11111111111111111100010001000110;
assign LUT_3[32887] = 32'b00000000000000000010111100100011;
assign LUT_3[32888] = 32'b00000000000000000010010100110010;
assign LUT_3[32889] = 32'b00000000000000001001000000001111;
assign LUT_3[32890] = 32'b00000000000000000100011100010110;
assign LUT_3[32891] = 32'b00000000000000001011000111110011;
assign LUT_3[32892] = 32'b11111111111111111111100010101000;
assign LUT_3[32893] = 32'b00000000000000000110001110000101;
assign LUT_3[32894] = 32'b00000000000000000001101010001100;
assign LUT_3[32895] = 32'b00000000000000001000010101101001;
assign LUT_3[32896] = 32'b11111111111111111010101100011100;
assign LUT_3[32897] = 32'b00000000000000000001010111111001;
assign LUT_3[32898] = 32'b11111111111111111100110100000000;
assign LUT_3[32899] = 32'b00000000000000000011011111011101;
assign LUT_3[32900] = 32'b11111111111111110111111010010010;
assign LUT_3[32901] = 32'b11111111111111111110100101101111;
assign LUT_3[32902] = 32'b11111111111111111010000001110110;
assign LUT_3[32903] = 32'b00000000000000000000101101010011;
assign LUT_3[32904] = 32'b00000000000000000000000101100010;
assign LUT_3[32905] = 32'b00000000000000000110110000111111;
assign LUT_3[32906] = 32'b00000000000000000010001101000110;
assign LUT_3[32907] = 32'b00000000000000001000111000100011;
assign LUT_3[32908] = 32'b11111111111111111101010011011000;
assign LUT_3[32909] = 32'b00000000000000000011111110110101;
assign LUT_3[32910] = 32'b11111111111111111111011010111100;
assign LUT_3[32911] = 32'b00000000000000000110000110011001;
assign LUT_3[32912] = 32'b11111111111111111101111111011111;
assign LUT_3[32913] = 32'b00000000000000000100101010111100;
assign LUT_3[32914] = 32'b00000000000000000000000111000011;
assign LUT_3[32915] = 32'b00000000000000000110110010100000;
assign LUT_3[32916] = 32'b11111111111111111011001101010101;
assign LUT_3[32917] = 32'b00000000000000000001111000110010;
assign LUT_3[32918] = 32'b11111111111111111101010100111001;
assign LUT_3[32919] = 32'b00000000000000000100000000010110;
assign LUT_3[32920] = 32'b00000000000000000011011000100101;
assign LUT_3[32921] = 32'b00000000000000001010000100000010;
assign LUT_3[32922] = 32'b00000000000000000101100000001001;
assign LUT_3[32923] = 32'b00000000000000001100001011100110;
assign LUT_3[32924] = 32'b00000000000000000000100110011011;
assign LUT_3[32925] = 32'b00000000000000000111010001111000;
assign LUT_3[32926] = 32'b00000000000000000010101101111111;
assign LUT_3[32927] = 32'b00000000000000001001011001011100;
assign LUT_3[32928] = 32'b11111111111111111011111010111100;
assign LUT_3[32929] = 32'b00000000000000000010100110011001;
assign LUT_3[32930] = 32'b11111111111111111110000010100000;
assign LUT_3[32931] = 32'b00000000000000000100101101111101;
assign LUT_3[32932] = 32'b11111111111111111001001000110010;
assign LUT_3[32933] = 32'b11111111111111111111110100001111;
assign LUT_3[32934] = 32'b11111111111111111011010000010110;
assign LUT_3[32935] = 32'b00000000000000000001111011110011;
assign LUT_3[32936] = 32'b00000000000000000001010100000010;
assign LUT_3[32937] = 32'b00000000000000000111111111011111;
assign LUT_3[32938] = 32'b00000000000000000011011011100110;
assign LUT_3[32939] = 32'b00000000000000001010000111000011;
assign LUT_3[32940] = 32'b11111111111111111110100001111000;
assign LUT_3[32941] = 32'b00000000000000000101001101010101;
assign LUT_3[32942] = 32'b00000000000000000000101001011100;
assign LUT_3[32943] = 32'b00000000000000000111010100111001;
assign LUT_3[32944] = 32'b11111111111111111111001101111111;
assign LUT_3[32945] = 32'b00000000000000000101111001011100;
assign LUT_3[32946] = 32'b00000000000000000001010101100011;
assign LUT_3[32947] = 32'b00000000000000001000000001000000;
assign LUT_3[32948] = 32'b11111111111111111100011011110101;
assign LUT_3[32949] = 32'b00000000000000000011000111010010;
assign LUT_3[32950] = 32'b11111111111111111110100011011001;
assign LUT_3[32951] = 32'b00000000000000000101001110110110;
assign LUT_3[32952] = 32'b00000000000000000100100111000101;
assign LUT_3[32953] = 32'b00000000000000001011010010100010;
assign LUT_3[32954] = 32'b00000000000000000110101110101001;
assign LUT_3[32955] = 32'b00000000000000001101011010000110;
assign LUT_3[32956] = 32'b00000000000000000001110100111011;
assign LUT_3[32957] = 32'b00000000000000001000100000011000;
assign LUT_3[32958] = 32'b00000000000000000011111100011111;
assign LUT_3[32959] = 32'b00000000000000001010100111111100;
assign LUT_3[32960] = 32'b11111111111111111010100101000111;
assign LUT_3[32961] = 32'b00000000000000000001010000100100;
assign LUT_3[32962] = 32'b11111111111111111100101100101011;
assign LUT_3[32963] = 32'b00000000000000000011011000001000;
assign LUT_3[32964] = 32'b11111111111111110111110010111101;
assign LUT_3[32965] = 32'b11111111111111111110011110011010;
assign LUT_3[32966] = 32'b11111111111111111001111010100001;
assign LUT_3[32967] = 32'b00000000000000000000100101111110;
assign LUT_3[32968] = 32'b11111111111111111111111110001101;
assign LUT_3[32969] = 32'b00000000000000000110101001101010;
assign LUT_3[32970] = 32'b00000000000000000010000101110001;
assign LUT_3[32971] = 32'b00000000000000001000110001001110;
assign LUT_3[32972] = 32'b11111111111111111101001100000011;
assign LUT_3[32973] = 32'b00000000000000000011110111100000;
assign LUT_3[32974] = 32'b11111111111111111111010011100111;
assign LUT_3[32975] = 32'b00000000000000000101111111000100;
assign LUT_3[32976] = 32'b11111111111111111101111000001010;
assign LUT_3[32977] = 32'b00000000000000000100100011100111;
assign LUT_3[32978] = 32'b11111111111111111111111111101110;
assign LUT_3[32979] = 32'b00000000000000000110101011001011;
assign LUT_3[32980] = 32'b11111111111111111011000110000000;
assign LUT_3[32981] = 32'b00000000000000000001110001011101;
assign LUT_3[32982] = 32'b11111111111111111101001101100100;
assign LUT_3[32983] = 32'b00000000000000000011111001000001;
assign LUT_3[32984] = 32'b00000000000000000011010001010000;
assign LUT_3[32985] = 32'b00000000000000001001111100101101;
assign LUT_3[32986] = 32'b00000000000000000101011000110100;
assign LUT_3[32987] = 32'b00000000000000001100000100010001;
assign LUT_3[32988] = 32'b00000000000000000000011111000110;
assign LUT_3[32989] = 32'b00000000000000000111001010100011;
assign LUT_3[32990] = 32'b00000000000000000010100110101010;
assign LUT_3[32991] = 32'b00000000000000001001010010000111;
assign LUT_3[32992] = 32'b11111111111111111011110011100111;
assign LUT_3[32993] = 32'b00000000000000000010011111000100;
assign LUT_3[32994] = 32'b11111111111111111101111011001011;
assign LUT_3[32995] = 32'b00000000000000000100100110101000;
assign LUT_3[32996] = 32'b11111111111111111001000001011101;
assign LUT_3[32997] = 32'b11111111111111111111101100111010;
assign LUT_3[32998] = 32'b11111111111111111011001001000001;
assign LUT_3[32999] = 32'b00000000000000000001110100011110;
assign LUT_3[33000] = 32'b00000000000000000001001100101101;
assign LUT_3[33001] = 32'b00000000000000000111111000001010;
assign LUT_3[33002] = 32'b00000000000000000011010100010001;
assign LUT_3[33003] = 32'b00000000000000001001111111101110;
assign LUT_3[33004] = 32'b11111111111111111110011010100011;
assign LUT_3[33005] = 32'b00000000000000000101000110000000;
assign LUT_3[33006] = 32'b00000000000000000000100010000111;
assign LUT_3[33007] = 32'b00000000000000000111001101100100;
assign LUT_3[33008] = 32'b11111111111111111111000110101010;
assign LUT_3[33009] = 32'b00000000000000000101110010000111;
assign LUT_3[33010] = 32'b00000000000000000001001110001110;
assign LUT_3[33011] = 32'b00000000000000000111111001101011;
assign LUT_3[33012] = 32'b11111111111111111100010100100000;
assign LUT_3[33013] = 32'b00000000000000000010111111111101;
assign LUT_3[33014] = 32'b11111111111111111110011100000100;
assign LUT_3[33015] = 32'b00000000000000000101000111100001;
assign LUT_3[33016] = 32'b00000000000000000100011111110000;
assign LUT_3[33017] = 32'b00000000000000001011001011001101;
assign LUT_3[33018] = 32'b00000000000000000110100111010100;
assign LUT_3[33019] = 32'b00000000000000001101010010110001;
assign LUT_3[33020] = 32'b00000000000000000001101101100110;
assign LUT_3[33021] = 32'b00000000000000001000011001000011;
assign LUT_3[33022] = 32'b00000000000000000011110101001010;
assign LUT_3[33023] = 32'b00000000000000001010100000100111;
assign LUT_3[33024] = 32'b11111111111111110100110000111111;
assign LUT_3[33025] = 32'b11111111111111111011011100011100;
assign LUT_3[33026] = 32'b11111111111111110110111000100011;
assign LUT_3[33027] = 32'b11111111111111111101100100000000;
assign LUT_3[33028] = 32'b11111111111111110001111110110101;
assign LUT_3[33029] = 32'b11111111111111111000101010010010;
assign LUT_3[33030] = 32'b11111111111111110100000110011001;
assign LUT_3[33031] = 32'b11111111111111111010110001110110;
assign LUT_3[33032] = 32'b11111111111111111010001010000101;
assign LUT_3[33033] = 32'b00000000000000000000110101100010;
assign LUT_3[33034] = 32'b11111111111111111100010001101001;
assign LUT_3[33035] = 32'b00000000000000000010111101000110;
assign LUT_3[33036] = 32'b11111111111111110111010111111011;
assign LUT_3[33037] = 32'b11111111111111111110000011011000;
assign LUT_3[33038] = 32'b11111111111111111001011111011111;
assign LUT_3[33039] = 32'b00000000000000000000001010111100;
assign LUT_3[33040] = 32'b11111111111111111000000100000010;
assign LUT_3[33041] = 32'b11111111111111111110101111011111;
assign LUT_3[33042] = 32'b11111111111111111010001011100110;
assign LUT_3[33043] = 32'b00000000000000000000110111000011;
assign LUT_3[33044] = 32'b11111111111111110101010001111000;
assign LUT_3[33045] = 32'b11111111111111111011111101010101;
assign LUT_3[33046] = 32'b11111111111111110111011001011100;
assign LUT_3[33047] = 32'b11111111111111111110000100111001;
assign LUT_3[33048] = 32'b11111111111111111101011101001000;
assign LUT_3[33049] = 32'b00000000000000000100001000100101;
assign LUT_3[33050] = 32'b11111111111111111111100100101100;
assign LUT_3[33051] = 32'b00000000000000000110010000001001;
assign LUT_3[33052] = 32'b11111111111111111010101010111110;
assign LUT_3[33053] = 32'b00000000000000000001010110011011;
assign LUT_3[33054] = 32'b11111111111111111100110010100010;
assign LUT_3[33055] = 32'b00000000000000000011011101111111;
assign LUT_3[33056] = 32'b11111111111111110101111111011111;
assign LUT_3[33057] = 32'b11111111111111111100101010111100;
assign LUT_3[33058] = 32'b11111111111111111000000111000011;
assign LUT_3[33059] = 32'b11111111111111111110110010100000;
assign LUT_3[33060] = 32'b11111111111111110011001101010101;
assign LUT_3[33061] = 32'b11111111111111111001111000110010;
assign LUT_3[33062] = 32'b11111111111111110101010100111001;
assign LUT_3[33063] = 32'b11111111111111111100000000010110;
assign LUT_3[33064] = 32'b11111111111111111011011000100101;
assign LUT_3[33065] = 32'b00000000000000000010000100000010;
assign LUT_3[33066] = 32'b11111111111111111101100000001001;
assign LUT_3[33067] = 32'b00000000000000000100001011100110;
assign LUT_3[33068] = 32'b11111111111111111000100110011011;
assign LUT_3[33069] = 32'b11111111111111111111010001111000;
assign LUT_3[33070] = 32'b11111111111111111010101101111111;
assign LUT_3[33071] = 32'b00000000000000000001011001011100;
assign LUT_3[33072] = 32'b11111111111111111001010010100010;
assign LUT_3[33073] = 32'b11111111111111111111111101111111;
assign LUT_3[33074] = 32'b11111111111111111011011010000110;
assign LUT_3[33075] = 32'b00000000000000000010000101100011;
assign LUT_3[33076] = 32'b11111111111111110110100000011000;
assign LUT_3[33077] = 32'b11111111111111111101001011110101;
assign LUT_3[33078] = 32'b11111111111111111000100111111100;
assign LUT_3[33079] = 32'b11111111111111111111010011011001;
assign LUT_3[33080] = 32'b11111111111111111110101011101000;
assign LUT_3[33081] = 32'b00000000000000000101010111000101;
assign LUT_3[33082] = 32'b00000000000000000000110011001100;
assign LUT_3[33083] = 32'b00000000000000000111011110101001;
assign LUT_3[33084] = 32'b11111111111111111011111001011110;
assign LUT_3[33085] = 32'b00000000000000000010100100111011;
assign LUT_3[33086] = 32'b11111111111111111110000001000010;
assign LUT_3[33087] = 32'b00000000000000000100101100011111;
assign LUT_3[33088] = 32'b11111111111111110100101001101010;
assign LUT_3[33089] = 32'b11111111111111111011010101000111;
assign LUT_3[33090] = 32'b11111111111111110110110001001110;
assign LUT_3[33091] = 32'b11111111111111111101011100101011;
assign LUT_3[33092] = 32'b11111111111111110001110111100000;
assign LUT_3[33093] = 32'b11111111111111111000100010111101;
assign LUT_3[33094] = 32'b11111111111111110011111111000100;
assign LUT_3[33095] = 32'b11111111111111111010101010100001;
assign LUT_3[33096] = 32'b11111111111111111010000010110000;
assign LUT_3[33097] = 32'b00000000000000000000101110001101;
assign LUT_3[33098] = 32'b11111111111111111100001010010100;
assign LUT_3[33099] = 32'b00000000000000000010110101110001;
assign LUT_3[33100] = 32'b11111111111111110111010000100110;
assign LUT_3[33101] = 32'b11111111111111111101111100000011;
assign LUT_3[33102] = 32'b11111111111111111001011000001010;
assign LUT_3[33103] = 32'b00000000000000000000000011100111;
assign LUT_3[33104] = 32'b11111111111111110111111100101101;
assign LUT_3[33105] = 32'b11111111111111111110101000001010;
assign LUT_3[33106] = 32'b11111111111111111010000100010001;
assign LUT_3[33107] = 32'b00000000000000000000101111101110;
assign LUT_3[33108] = 32'b11111111111111110101001010100011;
assign LUT_3[33109] = 32'b11111111111111111011110110000000;
assign LUT_3[33110] = 32'b11111111111111110111010010000111;
assign LUT_3[33111] = 32'b11111111111111111101111101100100;
assign LUT_3[33112] = 32'b11111111111111111101010101110011;
assign LUT_3[33113] = 32'b00000000000000000100000001010000;
assign LUT_3[33114] = 32'b11111111111111111111011101010111;
assign LUT_3[33115] = 32'b00000000000000000110001000110100;
assign LUT_3[33116] = 32'b11111111111111111010100011101001;
assign LUT_3[33117] = 32'b00000000000000000001001111000110;
assign LUT_3[33118] = 32'b11111111111111111100101011001101;
assign LUT_3[33119] = 32'b00000000000000000011010110101010;
assign LUT_3[33120] = 32'b11111111111111110101111000001010;
assign LUT_3[33121] = 32'b11111111111111111100100011100111;
assign LUT_3[33122] = 32'b11111111111111110111111111101110;
assign LUT_3[33123] = 32'b11111111111111111110101011001011;
assign LUT_3[33124] = 32'b11111111111111110011000110000000;
assign LUT_3[33125] = 32'b11111111111111111001110001011101;
assign LUT_3[33126] = 32'b11111111111111110101001101100100;
assign LUT_3[33127] = 32'b11111111111111111011111001000001;
assign LUT_3[33128] = 32'b11111111111111111011010001010000;
assign LUT_3[33129] = 32'b00000000000000000001111100101101;
assign LUT_3[33130] = 32'b11111111111111111101011000110100;
assign LUT_3[33131] = 32'b00000000000000000100000100010001;
assign LUT_3[33132] = 32'b11111111111111111000011111000110;
assign LUT_3[33133] = 32'b11111111111111111111001010100011;
assign LUT_3[33134] = 32'b11111111111111111010100110101010;
assign LUT_3[33135] = 32'b00000000000000000001010010000111;
assign LUT_3[33136] = 32'b11111111111111111001001011001101;
assign LUT_3[33137] = 32'b11111111111111111111110110101010;
assign LUT_3[33138] = 32'b11111111111111111011010010110001;
assign LUT_3[33139] = 32'b00000000000000000001111110001110;
assign LUT_3[33140] = 32'b11111111111111110110011001000011;
assign LUT_3[33141] = 32'b11111111111111111101000100100000;
assign LUT_3[33142] = 32'b11111111111111111000100000100111;
assign LUT_3[33143] = 32'b11111111111111111111001100000100;
assign LUT_3[33144] = 32'b11111111111111111110100100010011;
assign LUT_3[33145] = 32'b00000000000000000101001111110000;
assign LUT_3[33146] = 32'b00000000000000000000101011110111;
assign LUT_3[33147] = 32'b00000000000000000111010111010100;
assign LUT_3[33148] = 32'b11111111111111111011110010001001;
assign LUT_3[33149] = 32'b00000000000000000010011101100110;
assign LUT_3[33150] = 32'b11111111111111111101111001101101;
assign LUT_3[33151] = 32'b00000000000000000100100101001010;
assign LUT_3[33152] = 32'b11111111111111110110111011111101;
assign LUT_3[33153] = 32'b11111111111111111101100111011010;
assign LUT_3[33154] = 32'b11111111111111111001000011100001;
assign LUT_3[33155] = 32'b11111111111111111111101110111110;
assign LUT_3[33156] = 32'b11111111111111110100001001110011;
assign LUT_3[33157] = 32'b11111111111111111010110101010000;
assign LUT_3[33158] = 32'b11111111111111110110010001010111;
assign LUT_3[33159] = 32'b11111111111111111100111100110100;
assign LUT_3[33160] = 32'b11111111111111111100010101000011;
assign LUT_3[33161] = 32'b00000000000000000011000000100000;
assign LUT_3[33162] = 32'b11111111111111111110011100100111;
assign LUT_3[33163] = 32'b00000000000000000101001000000100;
assign LUT_3[33164] = 32'b11111111111111111001100010111001;
assign LUT_3[33165] = 32'b00000000000000000000001110010110;
assign LUT_3[33166] = 32'b11111111111111111011101010011101;
assign LUT_3[33167] = 32'b00000000000000000010010101111010;
assign LUT_3[33168] = 32'b11111111111111111010001111000000;
assign LUT_3[33169] = 32'b00000000000000000000111010011101;
assign LUT_3[33170] = 32'b11111111111111111100010110100100;
assign LUT_3[33171] = 32'b00000000000000000011000010000001;
assign LUT_3[33172] = 32'b11111111111111110111011100110110;
assign LUT_3[33173] = 32'b11111111111111111110001000010011;
assign LUT_3[33174] = 32'b11111111111111111001100100011010;
assign LUT_3[33175] = 32'b00000000000000000000001111110111;
assign LUT_3[33176] = 32'b11111111111111111111101000000110;
assign LUT_3[33177] = 32'b00000000000000000110010011100011;
assign LUT_3[33178] = 32'b00000000000000000001101111101010;
assign LUT_3[33179] = 32'b00000000000000001000011011000111;
assign LUT_3[33180] = 32'b11111111111111111100110101111100;
assign LUT_3[33181] = 32'b00000000000000000011100001011001;
assign LUT_3[33182] = 32'b11111111111111111110111101100000;
assign LUT_3[33183] = 32'b00000000000000000101101000111101;
assign LUT_3[33184] = 32'b11111111111111111000001010011101;
assign LUT_3[33185] = 32'b11111111111111111110110101111010;
assign LUT_3[33186] = 32'b11111111111111111010010010000001;
assign LUT_3[33187] = 32'b00000000000000000000111101011110;
assign LUT_3[33188] = 32'b11111111111111110101011000010011;
assign LUT_3[33189] = 32'b11111111111111111100000011110000;
assign LUT_3[33190] = 32'b11111111111111110111011111110111;
assign LUT_3[33191] = 32'b11111111111111111110001011010100;
assign LUT_3[33192] = 32'b11111111111111111101100011100011;
assign LUT_3[33193] = 32'b00000000000000000100001111000000;
assign LUT_3[33194] = 32'b11111111111111111111101011000111;
assign LUT_3[33195] = 32'b00000000000000000110010110100100;
assign LUT_3[33196] = 32'b11111111111111111010110001011001;
assign LUT_3[33197] = 32'b00000000000000000001011100110110;
assign LUT_3[33198] = 32'b11111111111111111100111000111101;
assign LUT_3[33199] = 32'b00000000000000000011100100011010;
assign LUT_3[33200] = 32'b11111111111111111011011101100000;
assign LUT_3[33201] = 32'b00000000000000000010001000111101;
assign LUT_3[33202] = 32'b11111111111111111101100101000100;
assign LUT_3[33203] = 32'b00000000000000000100010000100001;
assign LUT_3[33204] = 32'b11111111111111111000101011010110;
assign LUT_3[33205] = 32'b11111111111111111111010110110011;
assign LUT_3[33206] = 32'b11111111111111111010110010111010;
assign LUT_3[33207] = 32'b00000000000000000001011110010111;
assign LUT_3[33208] = 32'b00000000000000000000110110100110;
assign LUT_3[33209] = 32'b00000000000000000111100010000011;
assign LUT_3[33210] = 32'b00000000000000000010111110001010;
assign LUT_3[33211] = 32'b00000000000000001001101001100111;
assign LUT_3[33212] = 32'b11111111111111111110000100011100;
assign LUT_3[33213] = 32'b00000000000000000100101111111001;
assign LUT_3[33214] = 32'b00000000000000000000001100000000;
assign LUT_3[33215] = 32'b00000000000000000110110111011101;
assign LUT_3[33216] = 32'b11111111111111110110110100101000;
assign LUT_3[33217] = 32'b11111111111111111101100000000101;
assign LUT_3[33218] = 32'b11111111111111111000111100001100;
assign LUT_3[33219] = 32'b11111111111111111111100111101001;
assign LUT_3[33220] = 32'b11111111111111110100000010011110;
assign LUT_3[33221] = 32'b11111111111111111010101101111011;
assign LUT_3[33222] = 32'b11111111111111110110001010000010;
assign LUT_3[33223] = 32'b11111111111111111100110101011111;
assign LUT_3[33224] = 32'b11111111111111111100001101101110;
assign LUT_3[33225] = 32'b00000000000000000010111001001011;
assign LUT_3[33226] = 32'b11111111111111111110010101010010;
assign LUT_3[33227] = 32'b00000000000000000101000000101111;
assign LUT_3[33228] = 32'b11111111111111111001011011100100;
assign LUT_3[33229] = 32'b00000000000000000000000111000001;
assign LUT_3[33230] = 32'b11111111111111111011100011001000;
assign LUT_3[33231] = 32'b00000000000000000010001110100101;
assign LUT_3[33232] = 32'b11111111111111111010000111101011;
assign LUT_3[33233] = 32'b00000000000000000000110011001000;
assign LUT_3[33234] = 32'b11111111111111111100001111001111;
assign LUT_3[33235] = 32'b00000000000000000010111010101100;
assign LUT_3[33236] = 32'b11111111111111110111010101100001;
assign LUT_3[33237] = 32'b11111111111111111110000000111110;
assign LUT_3[33238] = 32'b11111111111111111001011101000101;
assign LUT_3[33239] = 32'b00000000000000000000001000100010;
assign LUT_3[33240] = 32'b11111111111111111111100000110001;
assign LUT_3[33241] = 32'b00000000000000000110001100001110;
assign LUT_3[33242] = 32'b00000000000000000001101000010101;
assign LUT_3[33243] = 32'b00000000000000001000010011110010;
assign LUT_3[33244] = 32'b11111111111111111100101110100111;
assign LUT_3[33245] = 32'b00000000000000000011011010000100;
assign LUT_3[33246] = 32'b11111111111111111110110110001011;
assign LUT_3[33247] = 32'b00000000000000000101100001101000;
assign LUT_3[33248] = 32'b11111111111111111000000011001000;
assign LUT_3[33249] = 32'b11111111111111111110101110100101;
assign LUT_3[33250] = 32'b11111111111111111010001010101100;
assign LUT_3[33251] = 32'b00000000000000000000110110001001;
assign LUT_3[33252] = 32'b11111111111111110101010000111110;
assign LUT_3[33253] = 32'b11111111111111111011111100011011;
assign LUT_3[33254] = 32'b11111111111111110111011000100010;
assign LUT_3[33255] = 32'b11111111111111111110000011111111;
assign LUT_3[33256] = 32'b11111111111111111101011100001110;
assign LUT_3[33257] = 32'b00000000000000000100000111101011;
assign LUT_3[33258] = 32'b11111111111111111111100011110010;
assign LUT_3[33259] = 32'b00000000000000000110001111001111;
assign LUT_3[33260] = 32'b11111111111111111010101010000100;
assign LUT_3[33261] = 32'b00000000000000000001010101100001;
assign LUT_3[33262] = 32'b11111111111111111100110001101000;
assign LUT_3[33263] = 32'b00000000000000000011011101000101;
assign LUT_3[33264] = 32'b11111111111111111011010110001011;
assign LUT_3[33265] = 32'b00000000000000000010000001101000;
assign LUT_3[33266] = 32'b11111111111111111101011101101111;
assign LUT_3[33267] = 32'b00000000000000000100001001001100;
assign LUT_3[33268] = 32'b11111111111111111000100100000001;
assign LUT_3[33269] = 32'b11111111111111111111001111011110;
assign LUT_3[33270] = 32'b11111111111111111010101011100101;
assign LUT_3[33271] = 32'b00000000000000000001010111000010;
assign LUT_3[33272] = 32'b00000000000000000000101111010001;
assign LUT_3[33273] = 32'b00000000000000000111011010101110;
assign LUT_3[33274] = 32'b00000000000000000010110110110101;
assign LUT_3[33275] = 32'b00000000000000001001100010010010;
assign LUT_3[33276] = 32'b11111111111111111101111101000111;
assign LUT_3[33277] = 32'b00000000000000000100101000100100;
assign LUT_3[33278] = 32'b00000000000000000000000100101011;
assign LUT_3[33279] = 32'b00000000000000000110110000001000;
assign LUT_3[33280] = 32'b11111111111111111011110110101010;
assign LUT_3[33281] = 32'b00000000000000000010100010000111;
assign LUT_3[33282] = 32'b11111111111111111101111110001110;
assign LUT_3[33283] = 32'b00000000000000000100101001101011;
assign LUT_3[33284] = 32'b11111111111111111001000100100000;
assign LUT_3[33285] = 32'b11111111111111111111101111111101;
assign LUT_3[33286] = 32'b11111111111111111011001100000100;
assign LUT_3[33287] = 32'b00000000000000000001110111100001;
assign LUT_3[33288] = 32'b00000000000000000001001111110000;
assign LUT_3[33289] = 32'b00000000000000000111111011001101;
assign LUT_3[33290] = 32'b00000000000000000011010111010100;
assign LUT_3[33291] = 32'b00000000000000001010000010110001;
assign LUT_3[33292] = 32'b11111111111111111110011101100110;
assign LUT_3[33293] = 32'b00000000000000000101001001000011;
assign LUT_3[33294] = 32'b00000000000000000000100101001010;
assign LUT_3[33295] = 32'b00000000000000000111010000100111;
assign LUT_3[33296] = 32'b11111111111111111111001001101101;
assign LUT_3[33297] = 32'b00000000000000000101110101001010;
assign LUT_3[33298] = 32'b00000000000000000001010001010001;
assign LUT_3[33299] = 32'b00000000000000000111111100101110;
assign LUT_3[33300] = 32'b11111111111111111100010111100011;
assign LUT_3[33301] = 32'b00000000000000000011000011000000;
assign LUT_3[33302] = 32'b11111111111111111110011111000111;
assign LUT_3[33303] = 32'b00000000000000000101001010100100;
assign LUT_3[33304] = 32'b00000000000000000100100010110011;
assign LUT_3[33305] = 32'b00000000000000001011001110010000;
assign LUT_3[33306] = 32'b00000000000000000110101010010111;
assign LUT_3[33307] = 32'b00000000000000001101010101110100;
assign LUT_3[33308] = 32'b00000000000000000001110000101001;
assign LUT_3[33309] = 32'b00000000000000001000011100000110;
assign LUT_3[33310] = 32'b00000000000000000011111000001101;
assign LUT_3[33311] = 32'b00000000000000001010100011101010;
assign LUT_3[33312] = 32'b11111111111111111101000101001010;
assign LUT_3[33313] = 32'b00000000000000000011110000100111;
assign LUT_3[33314] = 32'b11111111111111111111001100101110;
assign LUT_3[33315] = 32'b00000000000000000101111000001011;
assign LUT_3[33316] = 32'b11111111111111111010010011000000;
assign LUT_3[33317] = 32'b00000000000000000000111110011101;
assign LUT_3[33318] = 32'b11111111111111111100011010100100;
assign LUT_3[33319] = 32'b00000000000000000011000110000001;
assign LUT_3[33320] = 32'b00000000000000000010011110010000;
assign LUT_3[33321] = 32'b00000000000000001001001001101101;
assign LUT_3[33322] = 32'b00000000000000000100100101110100;
assign LUT_3[33323] = 32'b00000000000000001011010001010001;
assign LUT_3[33324] = 32'b11111111111111111111101100000110;
assign LUT_3[33325] = 32'b00000000000000000110010111100011;
assign LUT_3[33326] = 32'b00000000000000000001110011101010;
assign LUT_3[33327] = 32'b00000000000000001000011111000111;
assign LUT_3[33328] = 32'b00000000000000000000011000001101;
assign LUT_3[33329] = 32'b00000000000000000111000011101010;
assign LUT_3[33330] = 32'b00000000000000000010011111110001;
assign LUT_3[33331] = 32'b00000000000000001001001011001110;
assign LUT_3[33332] = 32'b11111111111111111101100110000011;
assign LUT_3[33333] = 32'b00000000000000000100010001100000;
assign LUT_3[33334] = 32'b11111111111111111111101101100111;
assign LUT_3[33335] = 32'b00000000000000000110011001000100;
assign LUT_3[33336] = 32'b00000000000000000101110001010011;
assign LUT_3[33337] = 32'b00000000000000001100011100110000;
assign LUT_3[33338] = 32'b00000000000000000111111000110111;
assign LUT_3[33339] = 32'b00000000000000001110100100010100;
assign LUT_3[33340] = 32'b00000000000000000010111111001001;
assign LUT_3[33341] = 32'b00000000000000001001101010100110;
assign LUT_3[33342] = 32'b00000000000000000101000110101101;
assign LUT_3[33343] = 32'b00000000000000001011110010001010;
assign LUT_3[33344] = 32'b11111111111111111011101111010101;
assign LUT_3[33345] = 32'b00000000000000000010011010110010;
assign LUT_3[33346] = 32'b11111111111111111101110110111001;
assign LUT_3[33347] = 32'b00000000000000000100100010010110;
assign LUT_3[33348] = 32'b11111111111111111000111101001011;
assign LUT_3[33349] = 32'b11111111111111111111101000101000;
assign LUT_3[33350] = 32'b11111111111111111011000100101111;
assign LUT_3[33351] = 32'b00000000000000000001110000001100;
assign LUT_3[33352] = 32'b00000000000000000001001000011011;
assign LUT_3[33353] = 32'b00000000000000000111110011111000;
assign LUT_3[33354] = 32'b00000000000000000011001111111111;
assign LUT_3[33355] = 32'b00000000000000001001111011011100;
assign LUT_3[33356] = 32'b11111111111111111110010110010001;
assign LUT_3[33357] = 32'b00000000000000000101000001101110;
assign LUT_3[33358] = 32'b00000000000000000000011101110101;
assign LUT_3[33359] = 32'b00000000000000000111001001010010;
assign LUT_3[33360] = 32'b11111111111111111111000010011000;
assign LUT_3[33361] = 32'b00000000000000000101101101110101;
assign LUT_3[33362] = 32'b00000000000000000001001001111100;
assign LUT_3[33363] = 32'b00000000000000000111110101011001;
assign LUT_3[33364] = 32'b11111111111111111100010000001110;
assign LUT_3[33365] = 32'b00000000000000000010111011101011;
assign LUT_3[33366] = 32'b11111111111111111110010111110010;
assign LUT_3[33367] = 32'b00000000000000000101000011001111;
assign LUT_3[33368] = 32'b00000000000000000100011011011110;
assign LUT_3[33369] = 32'b00000000000000001011000110111011;
assign LUT_3[33370] = 32'b00000000000000000110100011000010;
assign LUT_3[33371] = 32'b00000000000000001101001110011111;
assign LUT_3[33372] = 32'b00000000000000000001101001010100;
assign LUT_3[33373] = 32'b00000000000000001000010100110001;
assign LUT_3[33374] = 32'b00000000000000000011110000111000;
assign LUT_3[33375] = 32'b00000000000000001010011100010101;
assign LUT_3[33376] = 32'b11111111111111111100111101110101;
assign LUT_3[33377] = 32'b00000000000000000011101001010010;
assign LUT_3[33378] = 32'b11111111111111111111000101011001;
assign LUT_3[33379] = 32'b00000000000000000101110000110110;
assign LUT_3[33380] = 32'b11111111111111111010001011101011;
assign LUT_3[33381] = 32'b00000000000000000000110111001000;
assign LUT_3[33382] = 32'b11111111111111111100010011001111;
assign LUT_3[33383] = 32'b00000000000000000010111110101100;
assign LUT_3[33384] = 32'b00000000000000000010010110111011;
assign LUT_3[33385] = 32'b00000000000000001001000010011000;
assign LUT_3[33386] = 32'b00000000000000000100011110011111;
assign LUT_3[33387] = 32'b00000000000000001011001001111100;
assign LUT_3[33388] = 32'b11111111111111111111100100110001;
assign LUT_3[33389] = 32'b00000000000000000110010000001110;
assign LUT_3[33390] = 32'b00000000000000000001101100010101;
assign LUT_3[33391] = 32'b00000000000000001000010111110010;
assign LUT_3[33392] = 32'b00000000000000000000010000111000;
assign LUT_3[33393] = 32'b00000000000000000110111100010101;
assign LUT_3[33394] = 32'b00000000000000000010011000011100;
assign LUT_3[33395] = 32'b00000000000000001001000011111001;
assign LUT_3[33396] = 32'b11111111111111111101011110101110;
assign LUT_3[33397] = 32'b00000000000000000100001010001011;
assign LUT_3[33398] = 32'b11111111111111111111100110010010;
assign LUT_3[33399] = 32'b00000000000000000110010001101111;
assign LUT_3[33400] = 32'b00000000000000000101101001111110;
assign LUT_3[33401] = 32'b00000000000000001100010101011011;
assign LUT_3[33402] = 32'b00000000000000000111110001100010;
assign LUT_3[33403] = 32'b00000000000000001110011100111111;
assign LUT_3[33404] = 32'b00000000000000000010110111110100;
assign LUT_3[33405] = 32'b00000000000000001001100011010001;
assign LUT_3[33406] = 32'b00000000000000000100111111011000;
assign LUT_3[33407] = 32'b00000000000000001011101010110101;
assign LUT_3[33408] = 32'b11111111111111111110000001101000;
assign LUT_3[33409] = 32'b00000000000000000100101101000101;
assign LUT_3[33410] = 32'b00000000000000000000001001001100;
assign LUT_3[33411] = 32'b00000000000000000110110100101001;
assign LUT_3[33412] = 32'b11111111111111111011001111011110;
assign LUT_3[33413] = 32'b00000000000000000001111010111011;
assign LUT_3[33414] = 32'b11111111111111111101010111000010;
assign LUT_3[33415] = 32'b00000000000000000100000010011111;
assign LUT_3[33416] = 32'b00000000000000000011011010101110;
assign LUT_3[33417] = 32'b00000000000000001010000110001011;
assign LUT_3[33418] = 32'b00000000000000000101100010010010;
assign LUT_3[33419] = 32'b00000000000000001100001101101111;
assign LUT_3[33420] = 32'b00000000000000000000101000100100;
assign LUT_3[33421] = 32'b00000000000000000111010100000001;
assign LUT_3[33422] = 32'b00000000000000000010110000001000;
assign LUT_3[33423] = 32'b00000000000000001001011011100101;
assign LUT_3[33424] = 32'b00000000000000000001010100101011;
assign LUT_3[33425] = 32'b00000000000000001000000000001000;
assign LUT_3[33426] = 32'b00000000000000000011011100001111;
assign LUT_3[33427] = 32'b00000000000000001010000111101100;
assign LUT_3[33428] = 32'b11111111111111111110100010100001;
assign LUT_3[33429] = 32'b00000000000000000101001101111110;
assign LUT_3[33430] = 32'b00000000000000000000101010000101;
assign LUT_3[33431] = 32'b00000000000000000111010101100010;
assign LUT_3[33432] = 32'b00000000000000000110101101110001;
assign LUT_3[33433] = 32'b00000000000000001101011001001110;
assign LUT_3[33434] = 32'b00000000000000001000110101010101;
assign LUT_3[33435] = 32'b00000000000000001111100000110010;
assign LUT_3[33436] = 32'b00000000000000000011111011100111;
assign LUT_3[33437] = 32'b00000000000000001010100111000100;
assign LUT_3[33438] = 32'b00000000000000000110000011001011;
assign LUT_3[33439] = 32'b00000000000000001100101110101000;
assign LUT_3[33440] = 32'b11111111111111111111010000001000;
assign LUT_3[33441] = 32'b00000000000000000101111011100101;
assign LUT_3[33442] = 32'b00000000000000000001010111101100;
assign LUT_3[33443] = 32'b00000000000000001000000011001001;
assign LUT_3[33444] = 32'b11111111111111111100011101111110;
assign LUT_3[33445] = 32'b00000000000000000011001001011011;
assign LUT_3[33446] = 32'b11111111111111111110100101100010;
assign LUT_3[33447] = 32'b00000000000000000101010000111111;
assign LUT_3[33448] = 32'b00000000000000000100101001001110;
assign LUT_3[33449] = 32'b00000000000000001011010100101011;
assign LUT_3[33450] = 32'b00000000000000000110110000110010;
assign LUT_3[33451] = 32'b00000000000000001101011100001111;
assign LUT_3[33452] = 32'b00000000000000000001110111000100;
assign LUT_3[33453] = 32'b00000000000000001000100010100001;
assign LUT_3[33454] = 32'b00000000000000000011111110101000;
assign LUT_3[33455] = 32'b00000000000000001010101010000101;
assign LUT_3[33456] = 32'b00000000000000000010100011001011;
assign LUT_3[33457] = 32'b00000000000000001001001110101000;
assign LUT_3[33458] = 32'b00000000000000000100101010101111;
assign LUT_3[33459] = 32'b00000000000000001011010110001100;
assign LUT_3[33460] = 32'b11111111111111111111110001000001;
assign LUT_3[33461] = 32'b00000000000000000110011100011110;
assign LUT_3[33462] = 32'b00000000000000000001111000100101;
assign LUT_3[33463] = 32'b00000000000000001000100100000010;
assign LUT_3[33464] = 32'b00000000000000000111111100010001;
assign LUT_3[33465] = 32'b00000000000000001110100111101110;
assign LUT_3[33466] = 32'b00000000000000001010000011110101;
assign LUT_3[33467] = 32'b00000000000000010000101111010010;
assign LUT_3[33468] = 32'b00000000000000000101001010000111;
assign LUT_3[33469] = 32'b00000000000000001011110101100100;
assign LUT_3[33470] = 32'b00000000000000000111010001101011;
assign LUT_3[33471] = 32'b00000000000000001101111101001000;
assign LUT_3[33472] = 32'b11111111111111111101111010010011;
assign LUT_3[33473] = 32'b00000000000000000100100101110000;
assign LUT_3[33474] = 32'b00000000000000000000000001110111;
assign LUT_3[33475] = 32'b00000000000000000110101101010100;
assign LUT_3[33476] = 32'b11111111111111111011001000001001;
assign LUT_3[33477] = 32'b00000000000000000001110011100110;
assign LUT_3[33478] = 32'b11111111111111111101001111101101;
assign LUT_3[33479] = 32'b00000000000000000011111011001010;
assign LUT_3[33480] = 32'b00000000000000000011010011011001;
assign LUT_3[33481] = 32'b00000000000000001001111110110110;
assign LUT_3[33482] = 32'b00000000000000000101011010111101;
assign LUT_3[33483] = 32'b00000000000000001100000110011010;
assign LUT_3[33484] = 32'b00000000000000000000100001001111;
assign LUT_3[33485] = 32'b00000000000000000111001100101100;
assign LUT_3[33486] = 32'b00000000000000000010101000110011;
assign LUT_3[33487] = 32'b00000000000000001001010100010000;
assign LUT_3[33488] = 32'b00000000000000000001001101010110;
assign LUT_3[33489] = 32'b00000000000000000111111000110011;
assign LUT_3[33490] = 32'b00000000000000000011010100111010;
assign LUT_3[33491] = 32'b00000000000000001010000000010111;
assign LUT_3[33492] = 32'b11111111111111111110011011001100;
assign LUT_3[33493] = 32'b00000000000000000101000110101001;
assign LUT_3[33494] = 32'b00000000000000000000100010110000;
assign LUT_3[33495] = 32'b00000000000000000111001110001101;
assign LUT_3[33496] = 32'b00000000000000000110100110011100;
assign LUT_3[33497] = 32'b00000000000000001101010001111001;
assign LUT_3[33498] = 32'b00000000000000001000101110000000;
assign LUT_3[33499] = 32'b00000000000000001111011001011101;
assign LUT_3[33500] = 32'b00000000000000000011110100010010;
assign LUT_3[33501] = 32'b00000000000000001010011111101111;
assign LUT_3[33502] = 32'b00000000000000000101111011110110;
assign LUT_3[33503] = 32'b00000000000000001100100111010011;
assign LUT_3[33504] = 32'b11111111111111111111001000110011;
assign LUT_3[33505] = 32'b00000000000000000101110100010000;
assign LUT_3[33506] = 32'b00000000000000000001010000010111;
assign LUT_3[33507] = 32'b00000000000000000111111011110100;
assign LUT_3[33508] = 32'b11111111111111111100010110101001;
assign LUT_3[33509] = 32'b00000000000000000011000010000110;
assign LUT_3[33510] = 32'b11111111111111111110011110001101;
assign LUT_3[33511] = 32'b00000000000000000101001001101010;
assign LUT_3[33512] = 32'b00000000000000000100100001111001;
assign LUT_3[33513] = 32'b00000000000000001011001101010110;
assign LUT_3[33514] = 32'b00000000000000000110101001011101;
assign LUT_3[33515] = 32'b00000000000000001101010100111010;
assign LUT_3[33516] = 32'b00000000000000000001101111101111;
assign LUT_3[33517] = 32'b00000000000000001000011011001100;
assign LUT_3[33518] = 32'b00000000000000000011110111010011;
assign LUT_3[33519] = 32'b00000000000000001010100010110000;
assign LUT_3[33520] = 32'b00000000000000000010011011110110;
assign LUT_3[33521] = 32'b00000000000000001001000111010011;
assign LUT_3[33522] = 32'b00000000000000000100100011011010;
assign LUT_3[33523] = 32'b00000000000000001011001110110111;
assign LUT_3[33524] = 32'b11111111111111111111101001101100;
assign LUT_3[33525] = 32'b00000000000000000110010101001001;
assign LUT_3[33526] = 32'b00000000000000000001110001010000;
assign LUT_3[33527] = 32'b00000000000000001000011100101101;
assign LUT_3[33528] = 32'b00000000000000000111110100111100;
assign LUT_3[33529] = 32'b00000000000000001110100000011001;
assign LUT_3[33530] = 32'b00000000000000001001111100100000;
assign LUT_3[33531] = 32'b00000000000000010000100111111101;
assign LUT_3[33532] = 32'b00000000000000000101000010110010;
assign LUT_3[33533] = 32'b00000000000000001011101110001111;
assign LUT_3[33534] = 32'b00000000000000000111001010010110;
assign LUT_3[33535] = 32'b00000000000000001101110101110011;
assign LUT_3[33536] = 32'b11111111111111111000000110001011;
assign LUT_3[33537] = 32'b11111111111111111110110001101000;
assign LUT_3[33538] = 32'b11111111111111111010001101101111;
assign LUT_3[33539] = 32'b00000000000000000000111001001100;
assign LUT_3[33540] = 32'b11111111111111110101010100000001;
assign LUT_3[33541] = 32'b11111111111111111011111111011110;
assign LUT_3[33542] = 32'b11111111111111110111011011100101;
assign LUT_3[33543] = 32'b11111111111111111110000111000010;
assign LUT_3[33544] = 32'b11111111111111111101011111010001;
assign LUT_3[33545] = 32'b00000000000000000100001010101110;
assign LUT_3[33546] = 32'b11111111111111111111100110110101;
assign LUT_3[33547] = 32'b00000000000000000110010010010010;
assign LUT_3[33548] = 32'b11111111111111111010101101000111;
assign LUT_3[33549] = 32'b00000000000000000001011000100100;
assign LUT_3[33550] = 32'b11111111111111111100110100101011;
assign LUT_3[33551] = 32'b00000000000000000011100000001000;
assign LUT_3[33552] = 32'b11111111111111111011011001001110;
assign LUT_3[33553] = 32'b00000000000000000010000100101011;
assign LUT_3[33554] = 32'b11111111111111111101100000110010;
assign LUT_3[33555] = 32'b00000000000000000100001100001111;
assign LUT_3[33556] = 32'b11111111111111111000100111000100;
assign LUT_3[33557] = 32'b11111111111111111111010010100001;
assign LUT_3[33558] = 32'b11111111111111111010101110101000;
assign LUT_3[33559] = 32'b00000000000000000001011010000101;
assign LUT_3[33560] = 32'b00000000000000000000110010010100;
assign LUT_3[33561] = 32'b00000000000000000111011101110001;
assign LUT_3[33562] = 32'b00000000000000000010111001111000;
assign LUT_3[33563] = 32'b00000000000000001001100101010101;
assign LUT_3[33564] = 32'b11111111111111111110000000001010;
assign LUT_3[33565] = 32'b00000000000000000100101011100111;
assign LUT_3[33566] = 32'b00000000000000000000000111101110;
assign LUT_3[33567] = 32'b00000000000000000110110011001011;
assign LUT_3[33568] = 32'b11111111111111111001010100101011;
assign LUT_3[33569] = 32'b00000000000000000000000000001000;
assign LUT_3[33570] = 32'b11111111111111111011011100001111;
assign LUT_3[33571] = 32'b00000000000000000010000111101100;
assign LUT_3[33572] = 32'b11111111111111110110100010100001;
assign LUT_3[33573] = 32'b11111111111111111101001101111110;
assign LUT_3[33574] = 32'b11111111111111111000101010000101;
assign LUT_3[33575] = 32'b11111111111111111111010101100010;
assign LUT_3[33576] = 32'b11111111111111111110101101110001;
assign LUT_3[33577] = 32'b00000000000000000101011001001110;
assign LUT_3[33578] = 32'b00000000000000000000110101010101;
assign LUT_3[33579] = 32'b00000000000000000111100000110010;
assign LUT_3[33580] = 32'b11111111111111111011111011100111;
assign LUT_3[33581] = 32'b00000000000000000010100111000100;
assign LUT_3[33582] = 32'b11111111111111111110000011001011;
assign LUT_3[33583] = 32'b00000000000000000100101110101000;
assign LUT_3[33584] = 32'b11111111111111111100100111101110;
assign LUT_3[33585] = 32'b00000000000000000011010011001011;
assign LUT_3[33586] = 32'b11111111111111111110101111010010;
assign LUT_3[33587] = 32'b00000000000000000101011010101111;
assign LUT_3[33588] = 32'b11111111111111111001110101100100;
assign LUT_3[33589] = 32'b00000000000000000000100001000001;
assign LUT_3[33590] = 32'b11111111111111111011111101001000;
assign LUT_3[33591] = 32'b00000000000000000010101000100101;
assign LUT_3[33592] = 32'b00000000000000000010000000110100;
assign LUT_3[33593] = 32'b00000000000000001000101100010001;
assign LUT_3[33594] = 32'b00000000000000000100001000011000;
assign LUT_3[33595] = 32'b00000000000000001010110011110101;
assign LUT_3[33596] = 32'b11111111111111111111001110101010;
assign LUT_3[33597] = 32'b00000000000000000101111010000111;
assign LUT_3[33598] = 32'b00000000000000000001010110001110;
assign LUT_3[33599] = 32'b00000000000000001000000001101011;
assign LUT_3[33600] = 32'b11111111111111110111111110110110;
assign LUT_3[33601] = 32'b11111111111111111110101010010011;
assign LUT_3[33602] = 32'b11111111111111111010000110011010;
assign LUT_3[33603] = 32'b00000000000000000000110001110111;
assign LUT_3[33604] = 32'b11111111111111110101001100101100;
assign LUT_3[33605] = 32'b11111111111111111011111000001001;
assign LUT_3[33606] = 32'b11111111111111110111010100010000;
assign LUT_3[33607] = 32'b11111111111111111101111111101101;
assign LUT_3[33608] = 32'b11111111111111111101010111111100;
assign LUT_3[33609] = 32'b00000000000000000100000011011001;
assign LUT_3[33610] = 32'b11111111111111111111011111100000;
assign LUT_3[33611] = 32'b00000000000000000110001010111101;
assign LUT_3[33612] = 32'b11111111111111111010100101110010;
assign LUT_3[33613] = 32'b00000000000000000001010001001111;
assign LUT_3[33614] = 32'b11111111111111111100101101010110;
assign LUT_3[33615] = 32'b00000000000000000011011000110011;
assign LUT_3[33616] = 32'b11111111111111111011010001111001;
assign LUT_3[33617] = 32'b00000000000000000001111101010110;
assign LUT_3[33618] = 32'b11111111111111111101011001011101;
assign LUT_3[33619] = 32'b00000000000000000100000100111010;
assign LUT_3[33620] = 32'b11111111111111111000011111101111;
assign LUT_3[33621] = 32'b11111111111111111111001011001100;
assign LUT_3[33622] = 32'b11111111111111111010100111010011;
assign LUT_3[33623] = 32'b00000000000000000001010010110000;
assign LUT_3[33624] = 32'b00000000000000000000101010111111;
assign LUT_3[33625] = 32'b00000000000000000111010110011100;
assign LUT_3[33626] = 32'b00000000000000000010110010100011;
assign LUT_3[33627] = 32'b00000000000000001001011110000000;
assign LUT_3[33628] = 32'b11111111111111111101111000110101;
assign LUT_3[33629] = 32'b00000000000000000100100100010010;
assign LUT_3[33630] = 32'b00000000000000000000000000011001;
assign LUT_3[33631] = 32'b00000000000000000110101011110110;
assign LUT_3[33632] = 32'b11111111111111111001001101010110;
assign LUT_3[33633] = 32'b11111111111111111111111000110011;
assign LUT_3[33634] = 32'b11111111111111111011010100111010;
assign LUT_3[33635] = 32'b00000000000000000010000000010111;
assign LUT_3[33636] = 32'b11111111111111110110011011001100;
assign LUT_3[33637] = 32'b11111111111111111101000110101001;
assign LUT_3[33638] = 32'b11111111111111111000100010110000;
assign LUT_3[33639] = 32'b11111111111111111111001110001101;
assign LUT_3[33640] = 32'b11111111111111111110100110011100;
assign LUT_3[33641] = 32'b00000000000000000101010001111001;
assign LUT_3[33642] = 32'b00000000000000000000101110000000;
assign LUT_3[33643] = 32'b00000000000000000111011001011101;
assign LUT_3[33644] = 32'b11111111111111111011110100010010;
assign LUT_3[33645] = 32'b00000000000000000010011111101111;
assign LUT_3[33646] = 32'b11111111111111111101111011110110;
assign LUT_3[33647] = 32'b00000000000000000100100111010011;
assign LUT_3[33648] = 32'b11111111111111111100100000011001;
assign LUT_3[33649] = 32'b00000000000000000011001011110110;
assign LUT_3[33650] = 32'b11111111111111111110100111111101;
assign LUT_3[33651] = 32'b00000000000000000101010011011010;
assign LUT_3[33652] = 32'b11111111111111111001101110001111;
assign LUT_3[33653] = 32'b00000000000000000000011001101100;
assign LUT_3[33654] = 32'b11111111111111111011110101110011;
assign LUT_3[33655] = 32'b00000000000000000010100001010000;
assign LUT_3[33656] = 32'b00000000000000000001111001011111;
assign LUT_3[33657] = 32'b00000000000000001000100100111100;
assign LUT_3[33658] = 32'b00000000000000000100000001000011;
assign LUT_3[33659] = 32'b00000000000000001010101100100000;
assign LUT_3[33660] = 32'b11111111111111111111000111010101;
assign LUT_3[33661] = 32'b00000000000000000101110010110010;
assign LUT_3[33662] = 32'b00000000000000000001001110111001;
assign LUT_3[33663] = 32'b00000000000000000111111010010110;
assign LUT_3[33664] = 32'b11111111111111111010010001001001;
assign LUT_3[33665] = 32'b00000000000000000000111100100110;
assign LUT_3[33666] = 32'b11111111111111111100011000101101;
assign LUT_3[33667] = 32'b00000000000000000011000100001010;
assign LUT_3[33668] = 32'b11111111111111110111011110111111;
assign LUT_3[33669] = 32'b11111111111111111110001010011100;
assign LUT_3[33670] = 32'b11111111111111111001100110100011;
assign LUT_3[33671] = 32'b00000000000000000000010010000000;
assign LUT_3[33672] = 32'b11111111111111111111101010001111;
assign LUT_3[33673] = 32'b00000000000000000110010101101100;
assign LUT_3[33674] = 32'b00000000000000000001110001110011;
assign LUT_3[33675] = 32'b00000000000000001000011101010000;
assign LUT_3[33676] = 32'b11111111111111111100111000000101;
assign LUT_3[33677] = 32'b00000000000000000011100011100010;
assign LUT_3[33678] = 32'b11111111111111111110111111101001;
assign LUT_3[33679] = 32'b00000000000000000101101011000110;
assign LUT_3[33680] = 32'b11111111111111111101100100001100;
assign LUT_3[33681] = 32'b00000000000000000100001111101001;
assign LUT_3[33682] = 32'b11111111111111111111101011110000;
assign LUT_3[33683] = 32'b00000000000000000110010111001101;
assign LUT_3[33684] = 32'b11111111111111111010110010000010;
assign LUT_3[33685] = 32'b00000000000000000001011101011111;
assign LUT_3[33686] = 32'b11111111111111111100111001100110;
assign LUT_3[33687] = 32'b00000000000000000011100101000011;
assign LUT_3[33688] = 32'b00000000000000000010111101010010;
assign LUT_3[33689] = 32'b00000000000000001001101000101111;
assign LUT_3[33690] = 32'b00000000000000000101000100110110;
assign LUT_3[33691] = 32'b00000000000000001011110000010011;
assign LUT_3[33692] = 32'b00000000000000000000001011001000;
assign LUT_3[33693] = 32'b00000000000000000110110110100101;
assign LUT_3[33694] = 32'b00000000000000000010010010101100;
assign LUT_3[33695] = 32'b00000000000000001000111110001001;
assign LUT_3[33696] = 32'b11111111111111111011011111101001;
assign LUT_3[33697] = 32'b00000000000000000010001011000110;
assign LUT_3[33698] = 32'b11111111111111111101100111001101;
assign LUT_3[33699] = 32'b00000000000000000100010010101010;
assign LUT_3[33700] = 32'b11111111111111111000101101011111;
assign LUT_3[33701] = 32'b11111111111111111111011000111100;
assign LUT_3[33702] = 32'b11111111111111111010110101000011;
assign LUT_3[33703] = 32'b00000000000000000001100000100000;
assign LUT_3[33704] = 32'b00000000000000000000111000101111;
assign LUT_3[33705] = 32'b00000000000000000111100100001100;
assign LUT_3[33706] = 32'b00000000000000000011000000010011;
assign LUT_3[33707] = 32'b00000000000000001001101011110000;
assign LUT_3[33708] = 32'b11111111111111111110000110100101;
assign LUT_3[33709] = 32'b00000000000000000100110010000010;
assign LUT_3[33710] = 32'b00000000000000000000001110001001;
assign LUT_3[33711] = 32'b00000000000000000110111001100110;
assign LUT_3[33712] = 32'b11111111111111111110110010101100;
assign LUT_3[33713] = 32'b00000000000000000101011110001001;
assign LUT_3[33714] = 32'b00000000000000000000111010010000;
assign LUT_3[33715] = 32'b00000000000000000111100101101101;
assign LUT_3[33716] = 32'b11111111111111111100000000100010;
assign LUT_3[33717] = 32'b00000000000000000010101011111111;
assign LUT_3[33718] = 32'b11111111111111111110001000000110;
assign LUT_3[33719] = 32'b00000000000000000100110011100011;
assign LUT_3[33720] = 32'b00000000000000000100001011110010;
assign LUT_3[33721] = 32'b00000000000000001010110111001111;
assign LUT_3[33722] = 32'b00000000000000000110010011010110;
assign LUT_3[33723] = 32'b00000000000000001100111110110011;
assign LUT_3[33724] = 32'b00000000000000000001011001101000;
assign LUT_3[33725] = 32'b00000000000000001000000101000101;
assign LUT_3[33726] = 32'b00000000000000000011100001001100;
assign LUT_3[33727] = 32'b00000000000000001010001100101001;
assign LUT_3[33728] = 32'b11111111111111111010001001110100;
assign LUT_3[33729] = 32'b00000000000000000000110101010001;
assign LUT_3[33730] = 32'b11111111111111111100010001011000;
assign LUT_3[33731] = 32'b00000000000000000010111100110101;
assign LUT_3[33732] = 32'b11111111111111110111010111101010;
assign LUT_3[33733] = 32'b11111111111111111110000011000111;
assign LUT_3[33734] = 32'b11111111111111111001011111001110;
assign LUT_3[33735] = 32'b00000000000000000000001010101011;
assign LUT_3[33736] = 32'b11111111111111111111100010111010;
assign LUT_3[33737] = 32'b00000000000000000110001110010111;
assign LUT_3[33738] = 32'b00000000000000000001101010011110;
assign LUT_3[33739] = 32'b00000000000000001000010101111011;
assign LUT_3[33740] = 32'b11111111111111111100110000110000;
assign LUT_3[33741] = 32'b00000000000000000011011100001101;
assign LUT_3[33742] = 32'b11111111111111111110111000010100;
assign LUT_3[33743] = 32'b00000000000000000101100011110001;
assign LUT_3[33744] = 32'b11111111111111111101011100110111;
assign LUT_3[33745] = 32'b00000000000000000100001000010100;
assign LUT_3[33746] = 32'b11111111111111111111100100011011;
assign LUT_3[33747] = 32'b00000000000000000110001111111000;
assign LUT_3[33748] = 32'b11111111111111111010101010101101;
assign LUT_3[33749] = 32'b00000000000000000001010110001010;
assign LUT_3[33750] = 32'b11111111111111111100110010010001;
assign LUT_3[33751] = 32'b00000000000000000011011101101110;
assign LUT_3[33752] = 32'b00000000000000000010110101111101;
assign LUT_3[33753] = 32'b00000000000000001001100001011010;
assign LUT_3[33754] = 32'b00000000000000000100111101100001;
assign LUT_3[33755] = 32'b00000000000000001011101000111110;
assign LUT_3[33756] = 32'b00000000000000000000000011110011;
assign LUT_3[33757] = 32'b00000000000000000110101111010000;
assign LUT_3[33758] = 32'b00000000000000000010001011010111;
assign LUT_3[33759] = 32'b00000000000000001000110110110100;
assign LUT_3[33760] = 32'b11111111111111111011011000010100;
assign LUT_3[33761] = 32'b00000000000000000010000011110001;
assign LUT_3[33762] = 32'b11111111111111111101011111111000;
assign LUT_3[33763] = 32'b00000000000000000100001011010101;
assign LUT_3[33764] = 32'b11111111111111111000100110001010;
assign LUT_3[33765] = 32'b11111111111111111111010001100111;
assign LUT_3[33766] = 32'b11111111111111111010101101101110;
assign LUT_3[33767] = 32'b00000000000000000001011001001011;
assign LUT_3[33768] = 32'b00000000000000000000110001011010;
assign LUT_3[33769] = 32'b00000000000000000111011100110111;
assign LUT_3[33770] = 32'b00000000000000000010111000111110;
assign LUT_3[33771] = 32'b00000000000000001001100100011011;
assign LUT_3[33772] = 32'b11111111111111111101111111010000;
assign LUT_3[33773] = 32'b00000000000000000100101010101101;
assign LUT_3[33774] = 32'b00000000000000000000000110110100;
assign LUT_3[33775] = 32'b00000000000000000110110010010001;
assign LUT_3[33776] = 32'b11111111111111111110101011010111;
assign LUT_3[33777] = 32'b00000000000000000101010110110100;
assign LUT_3[33778] = 32'b00000000000000000000110010111011;
assign LUT_3[33779] = 32'b00000000000000000111011110011000;
assign LUT_3[33780] = 32'b11111111111111111011111001001101;
assign LUT_3[33781] = 32'b00000000000000000010100100101010;
assign LUT_3[33782] = 32'b11111111111111111110000000110001;
assign LUT_3[33783] = 32'b00000000000000000100101100001110;
assign LUT_3[33784] = 32'b00000000000000000100000100011101;
assign LUT_3[33785] = 32'b00000000000000001010101111111010;
assign LUT_3[33786] = 32'b00000000000000000110001100000001;
assign LUT_3[33787] = 32'b00000000000000001100110111011110;
assign LUT_3[33788] = 32'b00000000000000000001010010010011;
assign LUT_3[33789] = 32'b00000000000000000111111101110000;
assign LUT_3[33790] = 32'b00000000000000000011011001110111;
assign LUT_3[33791] = 32'b00000000000000001010000101010100;
assign LUT_3[33792] = 32'b11111111111111111111000110011011;
assign LUT_3[33793] = 32'b00000000000000000101110001111000;
assign LUT_3[33794] = 32'b00000000000000000001001101111111;
assign LUT_3[33795] = 32'b00000000000000000111111001011100;
assign LUT_3[33796] = 32'b11111111111111111100010100010001;
assign LUT_3[33797] = 32'b00000000000000000010111111101110;
assign LUT_3[33798] = 32'b11111111111111111110011011110101;
assign LUT_3[33799] = 32'b00000000000000000101000111010010;
assign LUT_3[33800] = 32'b00000000000000000100011111100001;
assign LUT_3[33801] = 32'b00000000000000001011001010111110;
assign LUT_3[33802] = 32'b00000000000000000110100111000101;
assign LUT_3[33803] = 32'b00000000000000001101010010100010;
assign LUT_3[33804] = 32'b00000000000000000001101101010111;
assign LUT_3[33805] = 32'b00000000000000001000011000110100;
assign LUT_3[33806] = 32'b00000000000000000011110100111011;
assign LUT_3[33807] = 32'b00000000000000001010100000011000;
assign LUT_3[33808] = 32'b00000000000000000010011001011110;
assign LUT_3[33809] = 32'b00000000000000001001000100111011;
assign LUT_3[33810] = 32'b00000000000000000100100001000010;
assign LUT_3[33811] = 32'b00000000000000001011001100011111;
assign LUT_3[33812] = 32'b11111111111111111111100111010100;
assign LUT_3[33813] = 32'b00000000000000000110010010110001;
assign LUT_3[33814] = 32'b00000000000000000001101110111000;
assign LUT_3[33815] = 32'b00000000000000001000011010010101;
assign LUT_3[33816] = 32'b00000000000000000111110010100100;
assign LUT_3[33817] = 32'b00000000000000001110011110000001;
assign LUT_3[33818] = 32'b00000000000000001001111010001000;
assign LUT_3[33819] = 32'b00000000000000010000100101100101;
assign LUT_3[33820] = 32'b00000000000000000101000000011010;
assign LUT_3[33821] = 32'b00000000000000001011101011110111;
assign LUT_3[33822] = 32'b00000000000000000111000111111110;
assign LUT_3[33823] = 32'b00000000000000001101110011011011;
assign LUT_3[33824] = 32'b00000000000000000000010100111011;
assign LUT_3[33825] = 32'b00000000000000000111000000011000;
assign LUT_3[33826] = 32'b00000000000000000010011100011111;
assign LUT_3[33827] = 32'b00000000000000001001000111111100;
assign LUT_3[33828] = 32'b11111111111111111101100010110001;
assign LUT_3[33829] = 32'b00000000000000000100001110001110;
assign LUT_3[33830] = 32'b11111111111111111111101010010101;
assign LUT_3[33831] = 32'b00000000000000000110010101110010;
assign LUT_3[33832] = 32'b00000000000000000101101110000001;
assign LUT_3[33833] = 32'b00000000000000001100011001011110;
assign LUT_3[33834] = 32'b00000000000000000111110101100101;
assign LUT_3[33835] = 32'b00000000000000001110100001000010;
assign LUT_3[33836] = 32'b00000000000000000010111011110111;
assign LUT_3[33837] = 32'b00000000000000001001100111010100;
assign LUT_3[33838] = 32'b00000000000000000101000011011011;
assign LUT_3[33839] = 32'b00000000000000001011101110111000;
assign LUT_3[33840] = 32'b00000000000000000011100111111110;
assign LUT_3[33841] = 32'b00000000000000001010010011011011;
assign LUT_3[33842] = 32'b00000000000000000101101111100010;
assign LUT_3[33843] = 32'b00000000000000001100011010111111;
assign LUT_3[33844] = 32'b00000000000000000000110101110100;
assign LUT_3[33845] = 32'b00000000000000000111100001010001;
assign LUT_3[33846] = 32'b00000000000000000010111101011000;
assign LUT_3[33847] = 32'b00000000000000001001101000110101;
assign LUT_3[33848] = 32'b00000000000000001001000001000100;
assign LUT_3[33849] = 32'b00000000000000001111101100100001;
assign LUT_3[33850] = 32'b00000000000000001011001000101000;
assign LUT_3[33851] = 32'b00000000000000010001110100000101;
assign LUT_3[33852] = 32'b00000000000000000110001110111010;
assign LUT_3[33853] = 32'b00000000000000001100111010010111;
assign LUT_3[33854] = 32'b00000000000000001000010110011110;
assign LUT_3[33855] = 32'b00000000000000001111000001111011;
assign LUT_3[33856] = 32'b11111111111111111110111111000110;
assign LUT_3[33857] = 32'b00000000000000000101101010100011;
assign LUT_3[33858] = 32'b00000000000000000001000110101010;
assign LUT_3[33859] = 32'b00000000000000000111110010000111;
assign LUT_3[33860] = 32'b11111111111111111100001100111100;
assign LUT_3[33861] = 32'b00000000000000000010111000011001;
assign LUT_3[33862] = 32'b11111111111111111110010100100000;
assign LUT_3[33863] = 32'b00000000000000000100111111111101;
assign LUT_3[33864] = 32'b00000000000000000100011000001100;
assign LUT_3[33865] = 32'b00000000000000001011000011101001;
assign LUT_3[33866] = 32'b00000000000000000110011111110000;
assign LUT_3[33867] = 32'b00000000000000001101001011001101;
assign LUT_3[33868] = 32'b00000000000000000001100110000010;
assign LUT_3[33869] = 32'b00000000000000001000010001011111;
assign LUT_3[33870] = 32'b00000000000000000011101101100110;
assign LUT_3[33871] = 32'b00000000000000001010011001000011;
assign LUT_3[33872] = 32'b00000000000000000010010010001001;
assign LUT_3[33873] = 32'b00000000000000001000111101100110;
assign LUT_3[33874] = 32'b00000000000000000100011001101101;
assign LUT_3[33875] = 32'b00000000000000001011000101001010;
assign LUT_3[33876] = 32'b11111111111111111111011111111111;
assign LUT_3[33877] = 32'b00000000000000000110001011011100;
assign LUT_3[33878] = 32'b00000000000000000001100111100011;
assign LUT_3[33879] = 32'b00000000000000001000010011000000;
assign LUT_3[33880] = 32'b00000000000000000111101011001111;
assign LUT_3[33881] = 32'b00000000000000001110010110101100;
assign LUT_3[33882] = 32'b00000000000000001001110010110011;
assign LUT_3[33883] = 32'b00000000000000010000011110010000;
assign LUT_3[33884] = 32'b00000000000000000100111001000101;
assign LUT_3[33885] = 32'b00000000000000001011100100100010;
assign LUT_3[33886] = 32'b00000000000000000111000000101001;
assign LUT_3[33887] = 32'b00000000000000001101101100000110;
assign LUT_3[33888] = 32'b00000000000000000000001101100110;
assign LUT_3[33889] = 32'b00000000000000000110111001000011;
assign LUT_3[33890] = 32'b00000000000000000010010101001010;
assign LUT_3[33891] = 32'b00000000000000001001000000100111;
assign LUT_3[33892] = 32'b11111111111111111101011011011100;
assign LUT_3[33893] = 32'b00000000000000000100000110111001;
assign LUT_3[33894] = 32'b11111111111111111111100011000000;
assign LUT_3[33895] = 32'b00000000000000000110001110011101;
assign LUT_3[33896] = 32'b00000000000000000101100110101100;
assign LUT_3[33897] = 32'b00000000000000001100010010001001;
assign LUT_3[33898] = 32'b00000000000000000111101110010000;
assign LUT_3[33899] = 32'b00000000000000001110011001101101;
assign LUT_3[33900] = 32'b00000000000000000010110100100010;
assign LUT_3[33901] = 32'b00000000000000001001011111111111;
assign LUT_3[33902] = 32'b00000000000000000100111100000110;
assign LUT_3[33903] = 32'b00000000000000001011100111100011;
assign LUT_3[33904] = 32'b00000000000000000011100000101001;
assign LUT_3[33905] = 32'b00000000000000001010001100000110;
assign LUT_3[33906] = 32'b00000000000000000101101000001101;
assign LUT_3[33907] = 32'b00000000000000001100010011101010;
assign LUT_3[33908] = 32'b00000000000000000000101110011111;
assign LUT_3[33909] = 32'b00000000000000000111011001111100;
assign LUT_3[33910] = 32'b00000000000000000010110110000011;
assign LUT_3[33911] = 32'b00000000000000001001100001100000;
assign LUT_3[33912] = 32'b00000000000000001000111001101111;
assign LUT_3[33913] = 32'b00000000000000001111100101001100;
assign LUT_3[33914] = 32'b00000000000000001011000001010011;
assign LUT_3[33915] = 32'b00000000000000010001101100110000;
assign LUT_3[33916] = 32'b00000000000000000110000111100101;
assign LUT_3[33917] = 32'b00000000000000001100110011000010;
assign LUT_3[33918] = 32'b00000000000000001000001111001001;
assign LUT_3[33919] = 32'b00000000000000001110111010100110;
assign LUT_3[33920] = 32'b00000000000000000001010001011001;
assign LUT_3[33921] = 32'b00000000000000000111111100110110;
assign LUT_3[33922] = 32'b00000000000000000011011000111101;
assign LUT_3[33923] = 32'b00000000000000001010000100011010;
assign LUT_3[33924] = 32'b11111111111111111110011111001111;
assign LUT_3[33925] = 32'b00000000000000000101001010101100;
assign LUT_3[33926] = 32'b00000000000000000000100110110011;
assign LUT_3[33927] = 32'b00000000000000000111010010010000;
assign LUT_3[33928] = 32'b00000000000000000110101010011111;
assign LUT_3[33929] = 32'b00000000000000001101010101111100;
assign LUT_3[33930] = 32'b00000000000000001000110010000011;
assign LUT_3[33931] = 32'b00000000000000001111011101100000;
assign LUT_3[33932] = 32'b00000000000000000011111000010101;
assign LUT_3[33933] = 32'b00000000000000001010100011110010;
assign LUT_3[33934] = 32'b00000000000000000101111111111001;
assign LUT_3[33935] = 32'b00000000000000001100101011010110;
assign LUT_3[33936] = 32'b00000000000000000100100100011100;
assign LUT_3[33937] = 32'b00000000000000001011001111111001;
assign LUT_3[33938] = 32'b00000000000000000110101100000000;
assign LUT_3[33939] = 32'b00000000000000001101010111011101;
assign LUT_3[33940] = 32'b00000000000000000001110010010010;
assign LUT_3[33941] = 32'b00000000000000001000011101101111;
assign LUT_3[33942] = 32'b00000000000000000011111001110110;
assign LUT_3[33943] = 32'b00000000000000001010100101010011;
assign LUT_3[33944] = 32'b00000000000000001001111101100010;
assign LUT_3[33945] = 32'b00000000000000010000101000111111;
assign LUT_3[33946] = 32'b00000000000000001100000101000110;
assign LUT_3[33947] = 32'b00000000000000010010110000100011;
assign LUT_3[33948] = 32'b00000000000000000111001011011000;
assign LUT_3[33949] = 32'b00000000000000001101110110110101;
assign LUT_3[33950] = 32'b00000000000000001001010010111100;
assign LUT_3[33951] = 32'b00000000000000001111111110011001;
assign LUT_3[33952] = 32'b00000000000000000010011111111001;
assign LUT_3[33953] = 32'b00000000000000001001001011010110;
assign LUT_3[33954] = 32'b00000000000000000100100111011101;
assign LUT_3[33955] = 32'b00000000000000001011010010111010;
assign LUT_3[33956] = 32'b11111111111111111111101101101111;
assign LUT_3[33957] = 32'b00000000000000000110011001001100;
assign LUT_3[33958] = 32'b00000000000000000001110101010011;
assign LUT_3[33959] = 32'b00000000000000001000100000110000;
assign LUT_3[33960] = 32'b00000000000000000111111000111111;
assign LUT_3[33961] = 32'b00000000000000001110100100011100;
assign LUT_3[33962] = 32'b00000000000000001010000000100011;
assign LUT_3[33963] = 32'b00000000000000010000101100000000;
assign LUT_3[33964] = 32'b00000000000000000101000110110101;
assign LUT_3[33965] = 32'b00000000000000001011110010010010;
assign LUT_3[33966] = 32'b00000000000000000111001110011001;
assign LUT_3[33967] = 32'b00000000000000001101111001110110;
assign LUT_3[33968] = 32'b00000000000000000101110010111100;
assign LUT_3[33969] = 32'b00000000000000001100011110011001;
assign LUT_3[33970] = 32'b00000000000000000111111010100000;
assign LUT_3[33971] = 32'b00000000000000001110100101111101;
assign LUT_3[33972] = 32'b00000000000000000011000000110010;
assign LUT_3[33973] = 32'b00000000000000001001101100001111;
assign LUT_3[33974] = 32'b00000000000000000101001000010110;
assign LUT_3[33975] = 32'b00000000000000001011110011110011;
assign LUT_3[33976] = 32'b00000000000000001011001100000010;
assign LUT_3[33977] = 32'b00000000000000010001110111011111;
assign LUT_3[33978] = 32'b00000000000000001101010011100110;
assign LUT_3[33979] = 32'b00000000000000010011111111000011;
assign LUT_3[33980] = 32'b00000000000000001000011001111000;
assign LUT_3[33981] = 32'b00000000000000001111000101010101;
assign LUT_3[33982] = 32'b00000000000000001010100001011100;
assign LUT_3[33983] = 32'b00000000000000010001001100111001;
assign LUT_3[33984] = 32'b00000000000000000001001010000100;
assign LUT_3[33985] = 32'b00000000000000000111110101100001;
assign LUT_3[33986] = 32'b00000000000000000011010001101000;
assign LUT_3[33987] = 32'b00000000000000001001111101000101;
assign LUT_3[33988] = 32'b11111111111111111110010111111010;
assign LUT_3[33989] = 32'b00000000000000000101000011010111;
assign LUT_3[33990] = 32'b00000000000000000000011111011110;
assign LUT_3[33991] = 32'b00000000000000000111001010111011;
assign LUT_3[33992] = 32'b00000000000000000110100011001010;
assign LUT_3[33993] = 32'b00000000000000001101001110100111;
assign LUT_3[33994] = 32'b00000000000000001000101010101110;
assign LUT_3[33995] = 32'b00000000000000001111010110001011;
assign LUT_3[33996] = 32'b00000000000000000011110001000000;
assign LUT_3[33997] = 32'b00000000000000001010011100011101;
assign LUT_3[33998] = 32'b00000000000000000101111000100100;
assign LUT_3[33999] = 32'b00000000000000001100100100000001;
assign LUT_3[34000] = 32'b00000000000000000100011101000111;
assign LUT_3[34001] = 32'b00000000000000001011001000100100;
assign LUT_3[34002] = 32'b00000000000000000110100100101011;
assign LUT_3[34003] = 32'b00000000000000001101010000001000;
assign LUT_3[34004] = 32'b00000000000000000001101010111101;
assign LUT_3[34005] = 32'b00000000000000001000010110011010;
assign LUT_3[34006] = 32'b00000000000000000011110010100001;
assign LUT_3[34007] = 32'b00000000000000001010011101111110;
assign LUT_3[34008] = 32'b00000000000000001001110110001101;
assign LUT_3[34009] = 32'b00000000000000010000100001101010;
assign LUT_3[34010] = 32'b00000000000000001011111101110001;
assign LUT_3[34011] = 32'b00000000000000010010101001001110;
assign LUT_3[34012] = 32'b00000000000000000111000100000011;
assign LUT_3[34013] = 32'b00000000000000001101101111100000;
assign LUT_3[34014] = 32'b00000000000000001001001011100111;
assign LUT_3[34015] = 32'b00000000000000001111110111000100;
assign LUT_3[34016] = 32'b00000000000000000010011000100100;
assign LUT_3[34017] = 32'b00000000000000001001000100000001;
assign LUT_3[34018] = 32'b00000000000000000100100000001000;
assign LUT_3[34019] = 32'b00000000000000001011001011100101;
assign LUT_3[34020] = 32'b11111111111111111111100110011010;
assign LUT_3[34021] = 32'b00000000000000000110010001110111;
assign LUT_3[34022] = 32'b00000000000000000001101101111110;
assign LUT_3[34023] = 32'b00000000000000001000011001011011;
assign LUT_3[34024] = 32'b00000000000000000111110001101010;
assign LUT_3[34025] = 32'b00000000000000001110011101000111;
assign LUT_3[34026] = 32'b00000000000000001001111001001110;
assign LUT_3[34027] = 32'b00000000000000010000100100101011;
assign LUT_3[34028] = 32'b00000000000000000100111111100000;
assign LUT_3[34029] = 32'b00000000000000001011101010111101;
assign LUT_3[34030] = 32'b00000000000000000111000111000100;
assign LUT_3[34031] = 32'b00000000000000001101110010100001;
assign LUT_3[34032] = 32'b00000000000000000101101011100111;
assign LUT_3[34033] = 32'b00000000000000001100010111000100;
assign LUT_3[34034] = 32'b00000000000000000111110011001011;
assign LUT_3[34035] = 32'b00000000000000001110011110101000;
assign LUT_3[34036] = 32'b00000000000000000010111001011101;
assign LUT_3[34037] = 32'b00000000000000001001100100111010;
assign LUT_3[34038] = 32'b00000000000000000101000001000001;
assign LUT_3[34039] = 32'b00000000000000001011101100011110;
assign LUT_3[34040] = 32'b00000000000000001011000100101101;
assign LUT_3[34041] = 32'b00000000000000010001110000001010;
assign LUT_3[34042] = 32'b00000000000000001101001100010001;
assign LUT_3[34043] = 32'b00000000000000010011110111101110;
assign LUT_3[34044] = 32'b00000000000000001000010010100011;
assign LUT_3[34045] = 32'b00000000000000001110111110000000;
assign LUT_3[34046] = 32'b00000000000000001010011010000111;
assign LUT_3[34047] = 32'b00000000000000010001000101100100;
assign LUT_3[34048] = 32'b11111111111111111011010101111100;
assign LUT_3[34049] = 32'b00000000000000000010000001011001;
assign LUT_3[34050] = 32'b11111111111111111101011101100000;
assign LUT_3[34051] = 32'b00000000000000000100001000111101;
assign LUT_3[34052] = 32'b11111111111111111000100011110010;
assign LUT_3[34053] = 32'b11111111111111111111001111001111;
assign LUT_3[34054] = 32'b11111111111111111010101011010110;
assign LUT_3[34055] = 32'b00000000000000000001010110110011;
assign LUT_3[34056] = 32'b00000000000000000000101111000010;
assign LUT_3[34057] = 32'b00000000000000000111011010011111;
assign LUT_3[34058] = 32'b00000000000000000010110110100110;
assign LUT_3[34059] = 32'b00000000000000001001100010000011;
assign LUT_3[34060] = 32'b11111111111111111101111100111000;
assign LUT_3[34061] = 32'b00000000000000000100101000010101;
assign LUT_3[34062] = 32'b00000000000000000000000100011100;
assign LUT_3[34063] = 32'b00000000000000000110101111111001;
assign LUT_3[34064] = 32'b11111111111111111110101000111111;
assign LUT_3[34065] = 32'b00000000000000000101010100011100;
assign LUT_3[34066] = 32'b00000000000000000000110000100011;
assign LUT_3[34067] = 32'b00000000000000000111011100000000;
assign LUT_3[34068] = 32'b11111111111111111011110110110101;
assign LUT_3[34069] = 32'b00000000000000000010100010010010;
assign LUT_3[34070] = 32'b11111111111111111101111110011001;
assign LUT_3[34071] = 32'b00000000000000000100101001110110;
assign LUT_3[34072] = 32'b00000000000000000100000010000101;
assign LUT_3[34073] = 32'b00000000000000001010101101100010;
assign LUT_3[34074] = 32'b00000000000000000110001001101001;
assign LUT_3[34075] = 32'b00000000000000001100110101000110;
assign LUT_3[34076] = 32'b00000000000000000001001111111011;
assign LUT_3[34077] = 32'b00000000000000000111111011011000;
assign LUT_3[34078] = 32'b00000000000000000011010111011111;
assign LUT_3[34079] = 32'b00000000000000001010000010111100;
assign LUT_3[34080] = 32'b11111111111111111100100100011100;
assign LUT_3[34081] = 32'b00000000000000000011001111111001;
assign LUT_3[34082] = 32'b11111111111111111110101100000000;
assign LUT_3[34083] = 32'b00000000000000000101010111011101;
assign LUT_3[34084] = 32'b11111111111111111001110010010010;
assign LUT_3[34085] = 32'b00000000000000000000011101101111;
assign LUT_3[34086] = 32'b11111111111111111011111001110110;
assign LUT_3[34087] = 32'b00000000000000000010100101010011;
assign LUT_3[34088] = 32'b00000000000000000001111101100010;
assign LUT_3[34089] = 32'b00000000000000001000101000111111;
assign LUT_3[34090] = 32'b00000000000000000100000101000110;
assign LUT_3[34091] = 32'b00000000000000001010110000100011;
assign LUT_3[34092] = 32'b11111111111111111111001011011000;
assign LUT_3[34093] = 32'b00000000000000000101110110110101;
assign LUT_3[34094] = 32'b00000000000000000001010010111100;
assign LUT_3[34095] = 32'b00000000000000000111111110011001;
assign LUT_3[34096] = 32'b11111111111111111111110111011111;
assign LUT_3[34097] = 32'b00000000000000000110100010111100;
assign LUT_3[34098] = 32'b00000000000000000001111111000011;
assign LUT_3[34099] = 32'b00000000000000001000101010100000;
assign LUT_3[34100] = 32'b11111111111111111101000101010101;
assign LUT_3[34101] = 32'b00000000000000000011110000110010;
assign LUT_3[34102] = 32'b11111111111111111111001100111001;
assign LUT_3[34103] = 32'b00000000000000000101111000010110;
assign LUT_3[34104] = 32'b00000000000000000101010000100101;
assign LUT_3[34105] = 32'b00000000000000001011111100000010;
assign LUT_3[34106] = 32'b00000000000000000111011000001001;
assign LUT_3[34107] = 32'b00000000000000001110000011100110;
assign LUT_3[34108] = 32'b00000000000000000010011110011011;
assign LUT_3[34109] = 32'b00000000000000001001001001111000;
assign LUT_3[34110] = 32'b00000000000000000100100101111111;
assign LUT_3[34111] = 32'b00000000000000001011010001011100;
assign LUT_3[34112] = 32'b11111111111111111011001110100111;
assign LUT_3[34113] = 32'b00000000000000000001111010000100;
assign LUT_3[34114] = 32'b11111111111111111101010110001011;
assign LUT_3[34115] = 32'b00000000000000000100000001101000;
assign LUT_3[34116] = 32'b11111111111111111000011100011101;
assign LUT_3[34117] = 32'b11111111111111111111000111111010;
assign LUT_3[34118] = 32'b11111111111111111010100100000001;
assign LUT_3[34119] = 32'b00000000000000000001001111011110;
assign LUT_3[34120] = 32'b00000000000000000000100111101101;
assign LUT_3[34121] = 32'b00000000000000000111010011001010;
assign LUT_3[34122] = 32'b00000000000000000010101111010001;
assign LUT_3[34123] = 32'b00000000000000001001011010101110;
assign LUT_3[34124] = 32'b11111111111111111101110101100011;
assign LUT_3[34125] = 32'b00000000000000000100100001000000;
assign LUT_3[34126] = 32'b11111111111111111111111101000111;
assign LUT_3[34127] = 32'b00000000000000000110101000100100;
assign LUT_3[34128] = 32'b11111111111111111110100001101010;
assign LUT_3[34129] = 32'b00000000000000000101001101000111;
assign LUT_3[34130] = 32'b00000000000000000000101001001110;
assign LUT_3[34131] = 32'b00000000000000000111010100101011;
assign LUT_3[34132] = 32'b11111111111111111011101111100000;
assign LUT_3[34133] = 32'b00000000000000000010011010111101;
assign LUT_3[34134] = 32'b11111111111111111101110111000100;
assign LUT_3[34135] = 32'b00000000000000000100100010100001;
assign LUT_3[34136] = 32'b00000000000000000011111010110000;
assign LUT_3[34137] = 32'b00000000000000001010100110001101;
assign LUT_3[34138] = 32'b00000000000000000110000010010100;
assign LUT_3[34139] = 32'b00000000000000001100101101110001;
assign LUT_3[34140] = 32'b00000000000000000001001000100110;
assign LUT_3[34141] = 32'b00000000000000000111110100000011;
assign LUT_3[34142] = 32'b00000000000000000011010000001010;
assign LUT_3[34143] = 32'b00000000000000001001111011100111;
assign LUT_3[34144] = 32'b11111111111111111100011101000111;
assign LUT_3[34145] = 32'b00000000000000000011001000100100;
assign LUT_3[34146] = 32'b11111111111111111110100100101011;
assign LUT_3[34147] = 32'b00000000000000000101010000001000;
assign LUT_3[34148] = 32'b11111111111111111001101010111101;
assign LUT_3[34149] = 32'b00000000000000000000010110011010;
assign LUT_3[34150] = 32'b11111111111111111011110010100001;
assign LUT_3[34151] = 32'b00000000000000000010011101111110;
assign LUT_3[34152] = 32'b00000000000000000001110110001101;
assign LUT_3[34153] = 32'b00000000000000001000100001101010;
assign LUT_3[34154] = 32'b00000000000000000011111101110001;
assign LUT_3[34155] = 32'b00000000000000001010101001001110;
assign LUT_3[34156] = 32'b11111111111111111111000100000011;
assign LUT_3[34157] = 32'b00000000000000000101101111100000;
assign LUT_3[34158] = 32'b00000000000000000001001011100111;
assign LUT_3[34159] = 32'b00000000000000000111110111000100;
assign LUT_3[34160] = 32'b11111111111111111111110000001010;
assign LUT_3[34161] = 32'b00000000000000000110011011100111;
assign LUT_3[34162] = 32'b00000000000000000001110111101110;
assign LUT_3[34163] = 32'b00000000000000001000100011001011;
assign LUT_3[34164] = 32'b11111111111111111100111110000000;
assign LUT_3[34165] = 32'b00000000000000000011101001011101;
assign LUT_3[34166] = 32'b11111111111111111111000101100100;
assign LUT_3[34167] = 32'b00000000000000000101110001000001;
assign LUT_3[34168] = 32'b00000000000000000101001001010000;
assign LUT_3[34169] = 32'b00000000000000001011110100101101;
assign LUT_3[34170] = 32'b00000000000000000111010000110100;
assign LUT_3[34171] = 32'b00000000000000001101111100010001;
assign LUT_3[34172] = 32'b00000000000000000010010111000110;
assign LUT_3[34173] = 32'b00000000000000001001000010100011;
assign LUT_3[34174] = 32'b00000000000000000100011110101010;
assign LUT_3[34175] = 32'b00000000000000001011001010000111;
assign LUT_3[34176] = 32'b11111111111111111101100000111010;
assign LUT_3[34177] = 32'b00000000000000000100001100010111;
assign LUT_3[34178] = 32'b11111111111111111111101000011110;
assign LUT_3[34179] = 32'b00000000000000000110010011111011;
assign LUT_3[34180] = 32'b11111111111111111010101110110000;
assign LUT_3[34181] = 32'b00000000000000000001011010001101;
assign LUT_3[34182] = 32'b11111111111111111100110110010100;
assign LUT_3[34183] = 32'b00000000000000000011100001110001;
assign LUT_3[34184] = 32'b00000000000000000010111010000000;
assign LUT_3[34185] = 32'b00000000000000001001100101011101;
assign LUT_3[34186] = 32'b00000000000000000101000001100100;
assign LUT_3[34187] = 32'b00000000000000001011101101000001;
assign LUT_3[34188] = 32'b00000000000000000000000111110110;
assign LUT_3[34189] = 32'b00000000000000000110110011010011;
assign LUT_3[34190] = 32'b00000000000000000010001111011010;
assign LUT_3[34191] = 32'b00000000000000001000111010110111;
assign LUT_3[34192] = 32'b00000000000000000000110011111101;
assign LUT_3[34193] = 32'b00000000000000000111011111011010;
assign LUT_3[34194] = 32'b00000000000000000010111011100001;
assign LUT_3[34195] = 32'b00000000000000001001100110111110;
assign LUT_3[34196] = 32'b11111111111111111110000001110011;
assign LUT_3[34197] = 32'b00000000000000000100101101010000;
assign LUT_3[34198] = 32'b00000000000000000000001001010111;
assign LUT_3[34199] = 32'b00000000000000000110110100110100;
assign LUT_3[34200] = 32'b00000000000000000110001101000011;
assign LUT_3[34201] = 32'b00000000000000001100111000100000;
assign LUT_3[34202] = 32'b00000000000000001000010100100111;
assign LUT_3[34203] = 32'b00000000000000001111000000000100;
assign LUT_3[34204] = 32'b00000000000000000011011010111001;
assign LUT_3[34205] = 32'b00000000000000001010000110010110;
assign LUT_3[34206] = 32'b00000000000000000101100010011101;
assign LUT_3[34207] = 32'b00000000000000001100001101111010;
assign LUT_3[34208] = 32'b11111111111111111110101111011010;
assign LUT_3[34209] = 32'b00000000000000000101011010110111;
assign LUT_3[34210] = 32'b00000000000000000000110110111110;
assign LUT_3[34211] = 32'b00000000000000000111100010011011;
assign LUT_3[34212] = 32'b11111111111111111011111101010000;
assign LUT_3[34213] = 32'b00000000000000000010101000101101;
assign LUT_3[34214] = 32'b11111111111111111110000100110100;
assign LUT_3[34215] = 32'b00000000000000000100110000010001;
assign LUT_3[34216] = 32'b00000000000000000100001000100000;
assign LUT_3[34217] = 32'b00000000000000001010110011111101;
assign LUT_3[34218] = 32'b00000000000000000110010000000100;
assign LUT_3[34219] = 32'b00000000000000001100111011100001;
assign LUT_3[34220] = 32'b00000000000000000001010110010110;
assign LUT_3[34221] = 32'b00000000000000001000000001110011;
assign LUT_3[34222] = 32'b00000000000000000011011101111010;
assign LUT_3[34223] = 32'b00000000000000001010001001010111;
assign LUT_3[34224] = 32'b00000000000000000010000010011101;
assign LUT_3[34225] = 32'b00000000000000001000101101111010;
assign LUT_3[34226] = 32'b00000000000000000100001010000001;
assign LUT_3[34227] = 32'b00000000000000001010110101011110;
assign LUT_3[34228] = 32'b11111111111111111111010000010011;
assign LUT_3[34229] = 32'b00000000000000000101111011110000;
assign LUT_3[34230] = 32'b00000000000000000001010111110111;
assign LUT_3[34231] = 32'b00000000000000001000000011010100;
assign LUT_3[34232] = 32'b00000000000000000111011011100011;
assign LUT_3[34233] = 32'b00000000000000001110000111000000;
assign LUT_3[34234] = 32'b00000000000000001001100011000111;
assign LUT_3[34235] = 32'b00000000000000010000001110100100;
assign LUT_3[34236] = 32'b00000000000000000100101001011001;
assign LUT_3[34237] = 32'b00000000000000001011010100110110;
assign LUT_3[34238] = 32'b00000000000000000110110000111101;
assign LUT_3[34239] = 32'b00000000000000001101011100011010;
assign LUT_3[34240] = 32'b11111111111111111101011001100101;
assign LUT_3[34241] = 32'b00000000000000000100000101000010;
assign LUT_3[34242] = 32'b11111111111111111111100001001001;
assign LUT_3[34243] = 32'b00000000000000000110001100100110;
assign LUT_3[34244] = 32'b11111111111111111010100111011011;
assign LUT_3[34245] = 32'b00000000000000000001010010111000;
assign LUT_3[34246] = 32'b11111111111111111100101110111111;
assign LUT_3[34247] = 32'b00000000000000000011011010011100;
assign LUT_3[34248] = 32'b00000000000000000010110010101011;
assign LUT_3[34249] = 32'b00000000000000001001011110001000;
assign LUT_3[34250] = 32'b00000000000000000100111010001111;
assign LUT_3[34251] = 32'b00000000000000001011100101101100;
assign LUT_3[34252] = 32'b00000000000000000000000000100001;
assign LUT_3[34253] = 32'b00000000000000000110101011111110;
assign LUT_3[34254] = 32'b00000000000000000010001000000101;
assign LUT_3[34255] = 32'b00000000000000001000110011100010;
assign LUT_3[34256] = 32'b00000000000000000000101100101000;
assign LUT_3[34257] = 32'b00000000000000000111011000000101;
assign LUT_3[34258] = 32'b00000000000000000010110100001100;
assign LUT_3[34259] = 32'b00000000000000001001011111101001;
assign LUT_3[34260] = 32'b11111111111111111101111010011110;
assign LUT_3[34261] = 32'b00000000000000000100100101111011;
assign LUT_3[34262] = 32'b00000000000000000000000010000010;
assign LUT_3[34263] = 32'b00000000000000000110101101011111;
assign LUT_3[34264] = 32'b00000000000000000110000101101110;
assign LUT_3[34265] = 32'b00000000000000001100110001001011;
assign LUT_3[34266] = 32'b00000000000000001000001101010010;
assign LUT_3[34267] = 32'b00000000000000001110111000101111;
assign LUT_3[34268] = 32'b00000000000000000011010011100100;
assign LUT_3[34269] = 32'b00000000000000001001111111000001;
assign LUT_3[34270] = 32'b00000000000000000101011011001000;
assign LUT_3[34271] = 32'b00000000000000001100000110100101;
assign LUT_3[34272] = 32'b11111111111111111110101000000101;
assign LUT_3[34273] = 32'b00000000000000000101010011100010;
assign LUT_3[34274] = 32'b00000000000000000000101111101001;
assign LUT_3[34275] = 32'b00000000000000000111011011000110;
assign LUT_3[34276] = 32'b11111111111111111011110101111011;
assign LUT_3[34277] = 32'b00000000000000000010100001011000;
assign LUT_3[34278] = 32'b11111111111111111101111101011111;
assign LUT_3[34279] = 32'b00000000000000000100101000111100;
assign LUT_3[34280] = 32'b00000000000000000100000001001011;
assign LUT_3[34281] = 32'b00000000000000001010101100101000;
assign LUT_3[34282] = 32'b00000000000000000110001000101111;
assign LUT_3[34283] = 32'b00000000000000001100110100001100;
assign LUT_3[34284] = 32'b00000000000000000001001111000001;
assign LUT_3[34285] = 32'b00000000000000000111111010011110;
assign LUT_3[34286] = 32'b00000000000000000011010110100101;
assign LUT_3[34287] = 32'b00000000000000001010000010000010;
assign LUT_3[34288] = 32'b00000000000000000001111011001000;
assign LUT_3[34289] = 32'b00000000000000001000100110100101;
assign LUT_3[34290] = 32'b00000000000000000100000010101100;
assign LUT_3[34291] = 32'b00000000000000001010101110001001;
assign LUT_3[34292] = 32'b11111111111111111111001000111110;
assign LUT_3[34293] = 32'b00000000000000000101110100011011;
assign LUT_3[34294] = 32'b00000000000000000001010000100010;
assign LUT_3[34295] = 32'b00000000000000000111111011111111;
assign LUT_3[34296] = 32'b00000000000000000111010100001110;
assign LUT_3[34297] = 32'b00000000000000001101111111101011;
assign LUT_3[34298] = 32'b00000000000000001001011011110010;
assign LUT_3[34299] = 32'b00000000000000010000000111001111;
assign LUT_3[34300] = 32'b00000000000000000100100010000100;
assign LUT_3[34301] = 32'b00000000000000001011001101100001;
assign LUT_3[34302] = 32'b00000000000000000110101001101000;
assign LUT_3[34303] = 32'b00000000000000001101010101000101;
assign LUT_3[34304] = 32'b00000000000000000010011011100111;
assign LUT_3[34305] = 32'b00000000000000001001000111000100;
assign LUT_3[34306] = 32'b00000000000000000100100011001011;
assign LUT_3[34307] = 32'b00000000000000001011001110101000;
assign LUT_3[34308] = 32'b11111111111111111111101001011101;
assign LUT_3[34309] = 32'b00000000000000000110010100111010;
assign LUT_3[34310] = 32'b00000000000000000001110001000001;
assign LUT_3[34311] = 32'b00000000000000001000011100011110;
assign LUT_3[34312] = 32'b00000000000000000111110100101101;
assign LUT_3[34313] = 32'b00000000000000001110100000001010;
assign LUT_3[34314] = 32'b00000000000000001001111100010001;
assign LUT_3[34315] = 32'b00000000000000010000100111101110;
assign LUT_3[34316] = 32'b00000000000000000101000010100011;
assign LUT_3[34317] = 32'b00000000000000001011101110000000;
assign LUT_3[34318] = 32'b00000000000000000111001010000111;
assign LUT_3[34319] = 32'b00000000000000001101110101100100;
assign LUT_3[34320] = 32'b00000000000000000101101110101010;
assign LUT_3[34321] = 32'b00000000000000001100011010000111;
assign LUT_3[34322] = 32'b00000000000000000111110110001110;
assign LUT_3[34323] = 32'b00000000000000001110100001101011;
assign LUT_3[34324] = 32'b00000000000000000010111100100000;
assign LUT_3[34325] = 32'b00000000000000001001100111111101;
assign LUT_3[34326] = 32'b00000000000000000101000100000100;
assign LUT_3[34327] = 32'b00000000000000001011101111100001;
assign LUT_3[34328] = 32'b00000000000000001011000111110000;
assign LUT_3[34329] = 32'b00000000000000010001110011001101;
assign LUT_3[34330] = 32'b00000000000000001101001111010100;
assign LUT_3[34331] = 32'b00000000000000010011111010110001;
assign LUT_3[34332] = 32'b00000000000000001000010101100110;
assign LUT_3[34333] = 32'b00000000000000001111000001000011;
assign LUT_3[34334] = 32'b00000000000000001010011101001010;
assign LUT_3[34335] = 32'b00000000000000010001001000100111;
assign LUT_3[34336] = 32'b00000000000000000011101010000111;
assign LUT_3[34337] = 32'b00000000000000001010010101100100;
assign LUT_3[34338] = 32'b00000000000000000101110001101011;
assign LUT_3[34339] = 32'b00000000000000001100011101001000;
assign LUT_3[34340] = 32'b00000000000000000000110111111101;
assign LUT_3[34341] = 32'b00000000000000000111100011011010;
assign LUT_3[34342] = 32'b00000000000000000010111111100001;
assign LUT_3[34343] = 32'b00000000000000001001101010111110;
assign LUT_3[34344] = 32'b00000000000000001001000011001101;
assign LUT_3[34345] = 32'b00000000000000001111101110101010;
assign LUT_3[34346] = 32'b00000000000000001011001010110001;
assign LUT_3[34347] = 32'b00000000000000010001110110001110;
assign LUT_3[34348] = 32'b00000000000000000110010001000011;
assign LUT_3[34349] = 32'b00000000000000001100111100100000;
assign LUT_3[34350] = 32'b00000000000000001000011000100111;
assign LUT_3[34351] = 32'b00000000000000001111000100000100;
assign LUT_3[34352] = 32'b00000000000000000110111101001010;
assign LUT_3[34353] = 32'b00000000000000001101101000100111;
assign LUT_3[34354] = 32'b00000000000000001001000100101110;
assign LUT_3[34355] = 32'b00000000000000001111110000001011;
assign LUT_3[34356] = 32'b00000000000000000100001011000000;
assign LUT_3[34357] = 32'b00000000000000001010110110011101;
assign LUT_3[34358] = 32'b00000000000000000110010010100100;
assign LUT_3[34359] = 32'b00000000000000001100111110000001;
assign LUT_3[34360] = 32'b00000000000000001100010110010000;
assign LUT_3[34361] = 32'b00000000000000010011000001101101;
assign LUT_3[34362] = 32'b00000000000000001110011101110100;
assign LUT_3[34363] = 32'b00000000000000010101001001010001;
assign LUT_3[34364] = 32'b00000000000000001001100100000110;
assign LUT_3[34365] = 32'b00000000000000010000001111100011;
assign LUT_3[34366] = 32'b00000000000000001011101011101010;
assign LUT_3[34367] = 32'b00000000000000010010010111000111;
assign LUT_3[34368] = 32'b00000000000000000010010100010010;
assign LUT_3[34369] = 32'b00000000000000001000111111101111;
assign LUT_3[34370] = 32'b00000000000000000100011011110110;
assign LUT_3[34371] = 32'b00000000000000001011000111010011;
assign LUT_3[34372] = 32'b11111111111111111111100010001000;
assign LUT_3[34373] = 32'b00000000000000000110001101100101;
assign LUT_3[34374] = 32'b00000000000000000001101001101100;
assign LUT_3[34375] = 32'b00000000000000001000010101001001;
assign LUT_3[34376] = 32'b00000000000000000111101101011000;
assign LUT_3[34377] = 32'b00000000000000001110011000110101;
assign LUT_3[34378] = 32'b00000000000000001001110100111100;
assign LUT_3[34379] = 32'b00000000000000010000100000011001;
assign LUT_3[34380] = 32'b00000000000000000100111011001110;
assign LUT_3[34381] = 32'b00000000000000001011100110101011;
assign LUT_3[34382] = 32'b00000000000000000111000010110010;
assign LUT_3[34383] = 32'b00000000000000001101101110001111;
assign LUT_3[34384] = 32'b00000000000000000101100111010101;
assign LUT_3[34385] = 32'b00000000000000001100010010110010;
assign LUT_3[34386] = 32'b00000000000000000111101110111001;
assign LUT_3[34387] = 32'b00000000000000001110011010010110;
assign LUT_3[34388] = 32'b00000000000000000010110101001011;
assign LUT_3[34389] = 32'b00000000000000001001100000101000;
assign LUT_3[34390] = 32'b00000000000000000100111100101111;
assign LUT_3[34391] = 32'b00000000000000001011101000001100;
assign LUT_3[34392] = 32'b00000000000000001011000000011011;
assign LUT_3[34393] = 32'b00000000000000010001101011111000;
assign LUT_3[34394] = 32'b00000000000000001101000111111111;
assign LUT_3[34395] = 32'b00000000000000010011110011011100;
assign LUT_3[34396] = 32'b00000000000000001000001110010001;
assign LUT_3[34397] = 32'b00000000000000001110111001101110;
assign LUT_3[34398] = 32'b00000000000000001010010101110101;
assign LUT_3[34399] = 32'b00000000000000010001000001010010;
assign LUT_3[34400] = 32'b00000000000000000011100010110010;
assign LUT_3[34401] = 32'b00000000000000001010001110001111;
assign LUT_3[34402] = 32'b00000000000000000101101010010110;
assign LUT_3[34403] = 32'b00000000000000001100010101110011;
assign LUT_3[34404] = 32'b00000000000000000000110000101000;
assign LUT_3[34405] = 32'b00000000000000000111011100000101;
assign LUT_3[34406] = 32'b00000000000000000010111000001100;
assign LUT_3[34407] = 32'b00000000000000001001100011101001;
assign LUT_3[34408] = 32'b00000000000000001000111011111000;
assign LUT_3[34409] = 32'b00000000000000001111100111010101;
assign LUT_3[34410] = 32'b00000000000000001011000011011100;
assign LUT_3[34411] = 32'b00000000000000010001101110111001;
assign LUT_3[34412] = 32'b00000000000000000110001001101110;
assign LUT_3[34413] = 32'b00000000000000001100110101001011;
assign LUT_3[34414] = 32'b00000000000000001000010001010010;
assign LUT_3[34415] = 32'b00000000000000001110111100101111;
assign LUT_3[34416] = 32'b00000000000000000110110101110101;
assign LUT_3[34417] = 32'b00000000000000001101100001010010;
assign LUT_3[34418] = 32'b00000000000000001000111101011001;
assign LUT_3[34419] = 32'b00000000000000001111101000110110;
assign LUT_3[34420] = 32'b00000000000000000100000011101011;
assign LUT_3[34421] = 32'b00000000000000001010101111001000;
assign LUT_3[34422] = 32'b00000000000000000110001011001111;
assign LUT_3[34423] = 32'b00000000000000001100110110101100;
assign LUT_3[34424] = 32'b00000000000000001100001110111011;
assign LUT_3[34425] = 32'b00000000000000010010111010011000;
assign LUT_3[34426] = 32'b00000000000000001110010110011111;
assign LUT_3[34427] = 32'b00000000000000010101000001111100;
assign LUT_3[34428] = 32'b00000000000000001001011100110001;
assign LUT_3[34429] = 32'b00000000000000010000001000001110;
assign LUT_3[34430] = 32'b00000000000000001011100100010101;
assign LUT_3[34431] = 32'b00000000000000010010001111110010;
assign LUT_3[34432] = 32'b00000000000000000100100110100101;
assign LUT_3[34433] = 32'b00000000000000001011010010000010;
assign LUT_3[34434] = 32'b00000000000000000110101110001001;
assign LUT_3[34435] = 32'b00000000000000001101011001100110;
assign LUT_3[34436] = 32'b00000000000000000001110100011011;
assign LUT_3[34437] = 32'b00000000000000001000011111111000;
assign LUT_3[34438] = 32'b00000000000000000011111011111111;
assign LUT_3[34439] = 32'b00000000000000001010100111011100;
assign LUT_3[34440] = 32'b00000000000000001001111111101011;
assign LUT_3[34441] = 32'b00000000000000010000101011001000;
assign LUT_3[34442] = 32'b00000000000000001100000111001111;
assign LUT_3[34443] = 32'b00000000000000010010110010101100;
assign LUT_3[34444] = 32'b00000000000000000111001101100001;
assign LUT_3[34445] = 32'b00000000000000001101111000111110;
assign LUT_3[34446] = 32'b00000000000000001001010101000101;
assign LUT_3[34447] = 32'b00000000000000010000000000100010;
assign LUT_3[34448] = 32'b00000000000000000111111001101000;
assign LUT_3[34449] = 32'b00000000000000001110100101000101;
assign LUT_3[34450] = 32'b00000000000000001010000001001100;
assign LUT_3[34451] = 32'b00000000000000010000101100101001;
assign LUT_3[34452] = 32'b00000000000000000101000111011110;
assign LUT_3[34453] = 32'b00000000000000001011110010111011;
assign LUT_3[34454] = 32'b00000000000000000111001111000010;
assign LUT_3[34455] = 32'b00000000000000001101111010011111;
assign LUT_3[34456] = 32'b00000000000000001101010010101110;
assign LUT_3[34457] = 32'b00000000000000010011111110001011;
assign LUT_3[34458] = 32'b00000000000000001111011010010010;
assign LUT_3[34459] = 32'b00000000000000010110000101101111;
assign LUT_3[34460] = 32'b00000000000000001010100000100100;
assign LUT_3[34461] = 32'b00000000000000010001001100000001;
assign LUT_3[34462] = 32'b00000000000000001100101000001000;
assign LUT_3[34463] = 32'b00000000000000010011010011100101;
assign LUT_3[34464] = 32'b00000000000000000101110101000101;
assign LUT_3[34465] = 32'b00000000000000001100100000100010;
assign LUT_3[34466] = 32'b00000000000000000111111100101001;
assign LUT_3[34467] = 32'b00000000000000001110101000000110;
assign LUT_3[34468] = 32'b00000000000000000011000010111011;
assign LUT_3[34469] = 32'b00000000000000001001101110011000;
assign LUT_3[34470] = 32'b00000000000000000101001010011111;
assign LUT_3[34471] = 32'b00000000000000001011110101111100;
assign LUT_3[34472] = 32'b00000000000000001011001110001011;
assign LUT_3[34473] = 32'b00000000000000010001111001101000;
assign LUT_3[34474] = 32'b00000000000000001101010101101111;
assign LUT_3[34475] = 32'b00000000000000010100000001001100;
assign LUT_3[34476] = 32'b00000000000000001000011100000001;
assign LUT_3[34477] = 32'b00000000000000001111000111011110;
assign LUT_3[34478] = 32'b00000000000000001010100011100101;
assign LUT_3[34479] = 32'b00000000000000010001001111000010;
assign LUT_3[34480] = 32'b00000000000000001001001000001000;
assign LUT_3[34481] = 32'b00000000000000001111110011100101;
assign LUT_3[34482] = 32'b00000000000000001011001111101100;
assign LUT_3[34483] = 32'b00000000000000010001111011001001;
assign LUT_3[34484] = 32'b00000000000000000110010101111110;
assign LUT_3[34485] = 32'b00000000000000001101000001011011;
assign LUT_3[34486] = 32'b00000000000000001000011101100010;
assign LUT_3[34487] = 32'b00000000000000001111001000111111;
assign LUT_3[34488] = 32'b00000000000000001110100001001110;
assign LUT_3[34489] = 32'b00000000000000010101001100101011;
assign LUT_3[34490] = 32'b00000000000000010000101000110010;
assign LUT_3[34491] = 32'b00000000000000010111010100001111;
assign LUT_3[34492] = 32'b00000000000000001011101111000100;
assign LUT_3[34493] = 32'b00000000000000010010011010100001;
assign LUT_3[34494] = 32'b00000000000000001101110110101000;
assign LUT_3[34495] = 32'b00000000000000010100100010000101;
assign LUT_3[34496] = 32'b00000000000000000100011111010000;
assign LUT_3[34497] = 32'b00000000000000001011001010101101;
assign LUT_3[34498] = 32'b00000000000000000110100110110100;
assign LUT_3[34499] = 32'b00000000000000001101010010010001;
assign LUT_3[34500] = 32'b00000000000000000001101101000110;
assign LUT_3[34501] = 32'b00000000000000001000011000100011;
assign LUT_3[34502] = 32'b00000000000000000011110100101010;
assign LUT_3[34503] = 32'b00000000000000001010100000000111;
assign LUT_3[34504] = 32'b00000000000000001001111000010110;
assign LUT_3[34505] = 32'b00000000000000010000100011110011;
assign LUT_3[34506] = 32'b00000000000000001011111111111010;
assign LUT_3[34507] = 32'b00000000000000010010101011010111;
assign LUT_3[34508] = 32'b00000000000000000111000110001100;
assign LUT_3[34509] = 32'b00000000000000001101110001101001;
assign LUT_3[34510] = 32'b00000000000000001001001101110000;
assign LUT_3[34511] = 32'b00000000000000001111111001001101;
assign LUT_3[34512] = 32'b00000000000000000111110010010011;
assign LUT_3[34513] = 32'b00000000000000001110011101110000;
assign LUT_3[34514] = 32'b00000000000000001001111001110111;
assign LUT_3[34515] = 32'b00000000000000010000100101010100;
assign LUT_3[34516] = 32'b00000000000000000101000000001001;
assign LUT_3[34517] = 32'b00000000000000001011101011100110;
assign LUT_3[34518] = 32'b00000000000000000111000111101101;
assign LUT_3[34519] = 32'b00000000000000001101110011001010;
assign LUT_3[34520] = 32'b00000000000000001101001011011001;
assign LUT_3[34521] = 32'b00000000000000010011110110110110;
assign LUT_3[34522] = 32'b00000000000000001111010010111101;
assign LUT_3[34523] = 32'b00000000000000010101111110011010;
assign LUT_3[34524] = 32'b00000000000000001010011001001111;
assign LUT_3[34525] = 32'b00000000000000010001000100101100;
assign LUT_3[34526] = 32'b00000000000000001100100000110011;
assign LUT_3[34527] = 32'b00000000000000010011001100010000;
assign LUT_3[34528] = 32'b00000000000000000101101101110000;
assign LUT_3[34529] = 32'b00000000000000001100011001001101;
assign LUT_3[34530] = 32'b00000000000000000111110101010100;
assign LUT_3[34531] = 32'b00000000000000001110100000110001;
assign LUT_3[34532] = 32'b00000000000000000010111011100110;
assign LUT_3[34533] = 32'b00000000000000001001100111000011;
assign LUT_3[34534] = 32'b00000000000000000101000011001010;
assign LUT_3[34535] = 32'b00000000000000001011101110100111;
assign LUT_3[34536] = 32'b00000000000000001011000110110110;
assign LUT_3[34537] = 32'b00000000000000010001110010010011;
assign LUT_3[34538] = 32'b00000000000000001101001110011010;
assign LUT_3[34539] = 32'b00000000000000010011111001110111;
assign LUT_3[34540] = 32'b00000000000000001000010100101100;
assign LUT_3[34541] = 32'b00000000000000001111000000001001;
assign LUT_3[34542] = 32'b00000000000000001010011100010000;
assign LUT_3[34543] = 32'b00000000000000010001000111101101;
assign LUT_3[34544] = 32'b00000000000000001001000000110011;
assign LUT_3[34545] = 32'b00000000000000001111101100010000;
assign LUT_3[34546] = 32'b00000000000000001011001000010111;
assign LUT_3[34547] = 32'b00000000000000010001110011110100;
assign LUT_3[34548] = 32'b00000000000000000110001110101001;
assign LUT_3[34549] = 32'b00000000000000001100111010000110;
assign LUT_3[34550] = 32'b00000000000000001000010110001101;
assign LUT_3[34551] = 32'b00000000000000001111000001101010;
assign LUT_3[34552] = 32'b00000000000000001110011001111001;
assign LUT_3[34553] = 32'b00000000000000010101000101010110;
assign LUT_3[34554] = 32'b00000000000000010000100001011101;
assign LUT_3[34555] = 32'b00000000000000010111001100111010;
assign LUT_3[34556] = 32'b00000000000000001011100111101111;
assign LUT_3[34557] = 32'b00000000000000010010010011001100;
assign LUT_3[34558] = 32'b00000000000000001101101111010011;
assign LUT_3[34559] = 32'b00000000000000010100011010110000;
assign LUT_3[34560] = 32'b11111111111111111110101011001000;
assign LUT_3[34561] = 32'b00000000000000000101010110100101;
assign LUT_3[34562] = 32'b00000000000000000000110010101100;
assign LUT_3[34563] = 32'b00000000000000000111011110001001;
assign LUT_3[34564] = 32'b11111111111111111011111000111110;
assign LUT_3[34565] = 32'b00000000000000000010100100011011;
assign LUT_3[34566] = 32'b11111111111111111110000000100010;
assign LUT_3[34567] = 32'b00000000000000000100101011111111;
assign LUT_3[34568] = 32'b00000000000000000100000100001110;
assign LUT_3[34569] = 32'b00000000000000001010101111101011;
assign LUT_3[34570] = 32'b00000000000000000110001011110010;
assign LUT_3[34571] = 32'b00000000000000001100110111001111;
assign LUT_3[34572] = 32'b00000000000000000001010010000100;
assign LUT_3[34573] = 32'b00000000000000000111111101100001;
assign LUT_3[34574] = 32'b00000000000000000011011001101000;
assign LUT_3[34575] = 32'b00000000000000001010000101000101;
assign LUT_3[34576] = 32'b00000000000000000001111110001011;
assign LUT_3[34577] = 32'b00000000000000001000101001101000;
assign LUT_3[34578] = 32'b00000000000000000100000101101111;
assign LUT_3[34579] = 32'b00000000000000001010110001001100;
assign LUT_3[34580] = 32'b11111111111111111111001100000001;
assign LUT_3[34581] = 32'b00000000000000000101110111011110;
assign LUT_3[34582] = 32'b00000000000000000001010011100101;
assign LUT_3[34583] = 32'b00000000000000000111111111000010;
assign LUT_3[34584] = 32'b00000000000000000111010111010001;
assign LUT_3[34585] = 32'b00000000000000001110000010101110;
assign LUT_3[34586] = 32'b00000000000000001001011110110101;
assign LUT_3[34587] = 32'b00000000000000010000001010010010;
assign LUT_3[34588] = 32'b00000000000000000100100101000111;
assign LUT_3[34589] = 32'b00000000000000001011010000100100;
assign LUT_3[34590] = 32'b00000000000000000110101100101011;
assign LUT_3[34591] = 32'b00000000000000001101011000001000;
assign LUT_3[34592] = 32'b11111111111111111111111001101000;
assign LUT_3[34593] = 32'b00000000000000000110100101000101;
assign LUT_3[34594] = 32'b00000000000000000010000001001100;
assign LUT_3[34595] = 32'b00000000000000001000101100101001;
assign LUT_3[34596] = 32'b11111111111111111101000111011110;
assign LUT_3[34597] = 32'b00000000000000000011110010111011;
assign LUT_3[34598] = 32'b11111111111111111111001111000010;
assign LUT_3[34599] = 32'b00000000000000000101111010011111;
assign LUT_3[34600] = 32'b00000000000000000101010010101110;
assign LUT_3[34601] = 32'b00000000000000001011111110001011;
assign LUT_3[34602] = 32'b00000000000000000111011010010010;
assign LUT_3[34603] = 32'b00000000000000001110000101101111;
assign LUT_3[34604] = 32'b00000000000000000010100000100100;
assign LUT_3[34605] = 32'b00000000000000001001001100000001;
assign LUT_3[34606] = 32'b00000000000000000100101000001000;
assign LUT_3[34607] = 32'b00000000000000001011010011100101;
assign LUT_3[34608] = 32'b00000000000000000011001100101011;
assign LUT_3[34609] = 32'b00000000000000001001111000001000;
assign LUT_3[34610] = 32'b00000000000000000101010100001111;
assign LUT_3[34611] = 32'b00000000000000001011111111101100;
assign LUT_3[34612] = 32'b00000000000000000000011010100001;
assign LUT_3[34613] = 32'b00000000000000000111000101111110;
assign LUT_3[34614] = 32'b00000000000000000010100010000101;
assign LUT_3[34615] = 32'b00000000000000001001001101100010;
assign LUT_3[34616] = 32'b00000000000000001000100101110001;
assign LUT_3[34617] = 32'b00000000000000001111010001001110;
assign LUT_3[34618] = 32'b00000000000000001010101101010101;
assign LUT_3[34619] = 32'b00000000000000010001011000110010;
assign LUT_3[34620] = 32'b00000000000000000101110011100111;
assign LUT_3[34621] = 32'b00000000000000001100011111000100;
assign LUT_3[34622] = 32'b00000000000000000111111011001011;
assign LUT_3[34623] = 32'b00000000000000001110100110101000;
assign LUT_3[34624] = 32'b11111111111111111110100011110011;
assign LUT_3[34625] = 32'b00000000000000000101001111010000;
assign LUT_3[34626] = 32'b00000000000000000000101011010111;
assign LUT_3[34627] = 32'b00000000000000000111010110110100;
assign LUT_3[34628] = 32'b11111111111111111011110001101001;
assign LUT_3[34629] = 32'b00000000000000000010011101000110;
assign LUT_3[34630] = 32'b11111111111111111101111001001101;
assign LUT_3[34631] = 32'b00000000000000000100100100101010;
assign LUT_3[34632] = 32'b00000000000000000011111100111001;
assign LUT_3[34633] = 32'b00000000000000001010101000010110;
assign LUT_3[34634] = 32'b00000000000000000110000100011101;
assign LUT_3[34635] = 32'b00000000000000001100101111111010;
assign LUT_3[34636] = 32'b00000000000000000001001010101111;
assign LUT_3[34637] = 32'b00000000000000000111110110001100;
assign LUT_3[34638] = 32'b00000000000000000011010010010011;
assign LUT_3[34639] = 32'b00000000000000001001111101110000;
assign LUT_3[34640] = 32'b00000000000000000001110110110110;
assign LUT_3[34641] = 32'b00000000000000001000100010010011;
assign LUT_3[34642] = 32'b00000000000000000011111110011010;
assign LUT_3[34643] = 32'b00000000000000001010101001110111;
assign LUT_3[34644] = 32'b11111111111111111111000100101100;
assign LUT_3[34645] = 32'b00000000000000000101110000001001;
assign LUT_3[34646] = 32'b00000000000000000001001100010000;
assign LUT_3[34647] = 32'b00000000000000000111110111101101;
assign LUT_3[34648] = 32'b00000000000000000111001111111100;
assign LUT_3[34649] = 32'b00000000000000001101111011011001;
assign LUT_3[34650] = 32'b00000000000000001001010111100000;
assign LUT_3[34651] = 32'b00000000000000010000000010111101;
assign LUT_3[34652] = 32'b00000000000000000100011101110010;
assign LUT_3[34653] = 32'b00000000000000001011001001001111;
assign LUT_3[34654] = 32'b00000000000000000110100101010110;
assign LUT_3[34655] = 32'b00000000000000001101010000110011;
assign LUT_3[34656] = 32'b11111111111111111111110010010011;
assign LUT_3[34657] = 32'b00000000000000000110011101110000;
assign LUT_3[34658] = 32'b00000000000000000001111001110111;
assign LUT_3[34659] = 32'b00000000000000001000100101010100;
assign LUT_3[34660] = 32'b11111111111111111101000000001001;
assign LUT_3[34661] = 32'b00000000000000000011101011100110;
assign LUT_3[34662] = 32'b11111111111111111111000111101101;
assign LUT_3[34663] = 32'b00000000000000000101110011001010;
assign LUT_3[34664] = 32'b00000000000000000101001011011001;
assign LUT_3[34665] = 32'b00000000000000001011110110110110;
assign LUT_3[34666] = 32'b00000000000000000111010010111101;
assign LUT_3[34667] = 32'b00000000000000001101111110011010;
assign LUT_3[34668] = 32'b00000000000000000010011001001111;
assign LUT_3[34669] = 32'b00000000000000001001000100101100;
assign LUT_3[34670] = 32'b00000000000000000100100000110011;
assign LUT_3[34671] = 32'b00000000000000001011001100010000;
assign LUT_3[34672] = 32'b00000000000000000011000101010110;
assign LUT_3[34673] = 32'b00000000000000001001110000110011;
assign LUT_3[34674] = 32'b00000000000000000101001100111010;
assign LUT_3[34675] = 32'b00000000000000001011111000010111;
assign LUT_3[34676] = 32'b00000000000000000000010011001100;
assign LUT_3[34677] = 32'b00000000000000000110111110101001;
assign LUT_3[34678] = 32'b00000000000000000010011010110000;
assign LUT_3[34679] = 32'b00000000000000001001000110001101;
assign LUT_3[34680] = 32'b00000000000000001000011110011100;
assign LUT_3[34681] = 32'b00000000000000001111001001111001;
assign LUT_3[34682] = 32'b00000000000000001010100110000000;
assign LUT_3[34683] = 32'b00000000000000010001010001011101;
assign LUT_3[34684] = 32'b00000000000000000101101100010010;
assign LUT_3[34685] = 32'b00000000000000001100010111101111;
assign LUT_3[34686] = 32'b00000000000000000111110011110110;
assign LUT_3[34687] = 32'b00000000000000001110011111010011;
assign LUT_3[34688] = 32'b00000000000000000000110110000110;
assign LUT_3[34689] = 32'b00000000000000000111100001100011;
assign LUT_3[34690] = 32'b00000000000000000010111101101010;
assign LUT_3[34691] = 32'b00000000000000001001101001000111;
assign LUT_3[34692] = 32'b11111111111111111110000011111100;
assign LUT_3[34693] = 32'b00000000000000000100101111011001;
assign LUT_3[34694] = 32'b00000000000000000000001011100000;
assign LUT_3[34695] = 32'b00000000000000000110110110111101;
assign LUT_3[34696] = 32'b00000000000000000110001111001100;
assign LUT_3[34697] = 32'b00000000000000001100111010101001;
assign LUT_3[34698] = 32'b00000000000000001000010110110000;
assign LUT_3[34699] = 32'b00000000000000001111000010001101;
assign LUT_3[34700] = 32'b00000000000000000011011101000010;
assign LUT_3[34701] = 32'b00000000000000001010001000011111;
assign LUT_3[34702] = 32'b00000000000000000101100100100110;
assign LUT_3[34703] = 32'b00000000000000001100010000000011;
assign LUT_3[34704] = 32'b00000000000000000100001001001001;
assign LUT_3[34705] = 32'b00000000000000001010110100100110;
assign LUT_3[34706] = 32'b00000000000000000110010000101101;
assign LUT_3[34707] = 32'b00000000000000001100111100001010;
assign LUT_3[34708] = 32'b00000000000000000001010110111111;
assign LUT_3[34709] = 32'b00000000000000001000000010011100;
assign LUT_3[34710] = 32'b00000000000000000011011110100011;
assign LUT_3[34711] = 32'b00000000000000001010001010000000;
assign LUT_3[34712] = 32'b00000000000000001001100010001111;
assign LUT_3[34713] = 32'b00000000000000010000001101101100;
assign LUT_3[34714] = 32'b00000000000000001011101001110011;
assign LUT_3[34715] = 32'b00000000000000010010010101010000;
assign LUT_3[34716] = 32'b00000000000000000110110000000101;
assign LUT_3[34717] = 32'b00000000000000001101011011100010;
assign LUT_3[34718] = 32'b00000000000000001000110111101001;
assign LUT_3[34719] = 32'b00000000000000001111100011000110;
assign LUT_3[34720] = 32'b00000000000000000010000100100110;
assign LUT_3[34721] = 32'b00000000000000001000110000000011;
assign LUT_3[34722] = 32'b00000000000000000100001100001010;
assign LUT_3[34723] = 32'b00000000000000001010110111100111;
assign LUT_3[34724] = 32'b11111111111111111111010010011100;
assign LUT_3[34725] = 32'b00000000000000000101111101111001;
assign LUT_3[34726] = 32'b00000000000000000001011010000000;
assign LUT_3[34727] = 32'b00000000000000001000000101011101;
assign LUT_3[34728] = 32'b00000000000000000111011101101100;
assign LUT_3[34729] = 32'b00000000000000001110001001001001;
assign LUT_3[34730] = 32'b00000000000000001001100101010000;
assign LUT_3[34731] = 32'b00000000000000010000010000101101;
assign LUT_3[34732] = 32'b00000000000000000100101011100010;
assign LUT_3[34733] = 32'b00000000000000001011010110111111;
assign LUT_3[34734] = 32'b00000000000000000110110011000110;
assign LUT_3[34735] = 32'b00000000000000001101011110100011;
assign LUT_3[34736] = 32'b00000000000000000101010111101001;
assign LUT_3[34737] = 32'b00000000000000001100000011000110;
assign LUT_3[34738] = 32'b00000000000000000111011111001101;
assign LUT_3[34739] = 32'b00000000000000001110001010101010;
assign LUT_3[34740] = 32'b00000000000000000010100101011111;
assign LUT_3[34741] = 32'b00000000000000001001010000111100;
assign LUT_3[34742] = 32'b00000000000000000100101101000011;
assign LUT_3[34743] = 32'b00000000000000001011011000100000;
assign LUT_3[34744] = 32'b00000000000000001010110000101111;
assign LUT_3[34745] = 32'b00000000000000010001011100001100;
assign LUT_3[34746] = 32'b00000000000000001100111000010011;
assign LUT_3[34747] = 32'b00000000000000010011100011110000;
assign LUT_3[34748] = 32'b00000000000000000111111110100101;
assign LUT_3[34749] = 32'b00000000000000001110101010000010;
assign LUT_3[34750] = 32'b00000000000000001010000110001001;
assign LUT_3[34751] = 32'b00000000000000010000110001100110;
assign LUT_3[34752] = 32'b00000000000000000000101110110001;
assign LUT_3[34753] = 32'b00000000000000000111011010001110;
assign LUT_3[34754] = 32'b00000000000000000010110110010101;
assign LUT_3[34755] = 32'b00000000000000001001100001110010;
assign LUT_3[34756] = 32'b11111111111111111101111100100111;
assign LUT_3[34757] = 32'b00000000000000000100101000000100;
assign LUT_3[34758] = 32'b00000000000000000000000100001011;
assign LUT_3[34759] = 32'b00000000000000000110101111101000;
assign LUT_3[34760] = 32'b00000000000000000110000111110111;
assign LUT_3[34761] = 32'b00000000000000001100110011010100;
assign LUT_3[34762] = 32'b00000000000000001000001111011011;
assign LUT_3[34763] = 32'b00000000000000001110111010111000;
assign LUT_3[34764] = 32'b00000000000000000011010101101101;
assign LUT_3[34765] = 32'b00000000000000001010000001001010;
assign LUT_3[34766] = 32'b00000000000000000101011101010001;
assign LUT_3[34767] = 32'b00000000000000001100001000101110;
assign LUT_3[34768] = 32'b00000000000000000100000001110100;
assign LUT_3[34769] = 32'b00000000000000001010101101010001;
assign LUT_3[34770] = 32'b00000000000000000110001001011000;
assign LUT_3[34771] = 32'b00000000000000001100110100110101;
assign LUT_3[34772] = 32'b00000000000000000001001111101010;
assign LUT_3[34773] = 32'b00000000000000000111111011000111;
assign LUT_3[34774] = 32'b00000000000000000011010111001110;
assign LUT_3[34775] = 32'b00000000000000001010000010101011;
assign LUT_3[34776] = 32'b00000000000000001001011010111010;
assign LUT_3[34777] = 32'b00000000000000010000000110010111;
assign LUT_3[34778] = 32'b00000000000000001011100010011110;
assign LUT_3[34779] = 32'b00000000000000010010001101111011;
assign LUT_3[34780] = 32'b00000000000000000110101000110000;
assign LUT_3[34781] = 32'b00000000000000001101010100001101;
assign LUT_3[34782] = 32'b00000000000000001000110000010100;
assign LUT_3[34783] = 32'b00000000000000001111011011110001;
assign LUT_3[34784] = 32'b00000000000000000001111101010001;
assign LUT_3[34785] = 32'b00000000000000001000101000101110;
assign LUT_3[34786] = 32'b00000000000000000100000100110101;
assign LUT_3[34787] = 32'b00000000000000001010110000010010;
assign LUT_3[34788] = 32'b11111111111111111111001011000111;
assign LUT_3[34789] = 32'b00000000000000000101110110100100;
assign LUT_3[34790] = 32'b00000000000000000001010010101011;
assign LUT_3[34791] = 32'b00000000000000000111111110001000;
assign LUT_3[34792] = 32'b00000000000000000111010110010111;
assign LUT_3[34793] = 32'b00000000000000001110000001110100;
assign LUT_3[34794] = 32'b00000000000000001001011101111011;
assign LUT_3[34795] = 32'b00000000000000010000001001011000;
assign LUT_3[34796] = 32'b00000000000000000100100100001101;
assign LUT_3[34797] = 32'b00000000000000001011001111101010;
assign LUT_3[34798] = 32'b00000000000000000110101011110001;
assign LUT_3[34799] = 32'b00000000000000001101010111001110;
assign LUT_3[34800] = 32'b00000000000000000101010000010100;
assign LUT_3[34801] = 32'b00000000000000001011111011110001;
assign LUT_3[34802] = 32'b00000000000000000111010111111000;
assign LUT_3[34803] = 32'b00000000000000001110000011010101;
assign LUT_3[34804] = 32'b00000000000000000010011110001010;
assign LUT_3[34805] = 32'b00000000000000001001001001100111;
assign LUT_3[34806] = 32'b00000000000000000100100101101110;
assign LUT_3[34807] = 32'b00000000000000001011010001001011;
assign LUT_3[34808] = 32'b00000000000000001010101001011010;
assign LUT_3[34809] = 32'b00000000000000010001010100110111;
assign LUT_3[34810] = 32'b00000000000000001100110000111110;
assign LUT_3[34811] = 32'b00000000000000010011011100011011;
assign LUT_3[34812] = 32'b00000000000000000111110111010000;
assign LUT_3[34813] = 32'b00000000000000001110100010101101;
assign LUT_3[34814] = 32'b00000000000000001001111110110100;
assign LUT_3[34815] = 32'b00000000000000010000101010010001;
assign LUT_3[34816] = 32'b11111111111111111010010111101100;
assign LUT_3[34817] = 32'b00000000000000000001000011001001;
assign LUT_3[34818] = 32'b11111111111111111100011111010000;
assign LUT_3[34819] = 32'b00000000000000000011001010101101;
assign LUT_3[34820] = 32'b11111111111111110111100101100010;
assign LUT_3[34821] = 32'b11111111111111111110010000111111;
assign LUT_3[34822] = 32'b11111111111111111001101101000110;
assign LUT_3[34823] = 32'b00000000000000000000011000100011;
assign LUT_3[34824] = 32'b11111111111111111111110000110010;
assign LUT_3[34825] = 32'b00000000000000000110011100001111;
assign LUT_3[34826] = 32'b00000000000000000001111000010110;
assign LUT_3[34827] = 32'b00000000000000001000100011110011;
assign LUT_3[34828] = 32'b11111111111111111100111110101000;
assign LUT_3[34829] = 32'b00000000000000000011101010000101;
assign LUT_3[34830] = 32'b11111111111111111111000110001100;
assign LUT_3[34831] = 32'b00000000000000000101110001101001;
assign LUT_3[34832] = 32'b11111111111111111101101010101111;
assign LUT_3[34833] = 32'b00000000000000000100010110001100;
assign LUT_3[34834] = 32'b11111111111111111111110010010011;
assign LUT_3[34835] = 32'b00000000000000000110011101110000;
assign LUT_3[34836] = 32'b11111111111111111010111000100101;
assign LUT_3[34837] = 32'b00000000000000000001100100000010;
assign LUT_3[34838] = 32'b11111111111111111101000000001001;
assign LUT_3[34839] = 32'b00000000000000000011101011100110;
assign LUT_3[34840] = 32'b00000000000000000011000011110101;
assign LUT_3[34841] = 32'b00000000000000001001101111010010;
assign LUT_3[34842] = 32'b00000000000000000101001011011001;
assign LUT_3[34843] = 32'b00000000000000001011110110110110;
assign LUT_3[34844] = 32'b00000000000000000000010001101011;
assign LUT_3[34845] = 32'b00000000000000000110111101001000;
assign LUT_3[34846] = 32'b00000000000000000010011001001111;
assign LUT_3[34847] = 32'b00000000000000001001000100101100;
assign LUT_3[34848] = 32'b11111111111111111011100110001100;
assign LUT_3[34849] = 32'b00000000000000000010010001101001;
assign LUT_3[34850] = 32'b11111111111111111101101101110000;
assign LUT_3[34851] = 32'b00000000000000000100011001001101;
assign LUT_3[34852] = 32'b11111111111111111000110100000010;
assign LUT_3[34853] = 32'b11111111111111111111011111011111;
assign LUT_3[34854] = 32'b11111111111111111010111011100110;
assign LUT_3[34855] = 32'b00000000000000000001100111000011;
assign LUT_3[34856] = 32'b00000000000000000000111111010010;
assign LUT_3[34857] = 32'b00000000000000000111101010101111;
assign LUT_3[34858] = 32'b00000000000000000011000110110110;
assign LUT_3[34859] = 32'b00000000000000001001110010010011;
assign LUT_3[34860] = 32'b11111111111111111110001101001000;
assign LUT_3[34861] = 32'b00000000000000000100111000100101;
assign LUT_3[34862] = 32'b00000000000000000000010100101100;
assign LUT_3[34863] = 32'b00000000000000000111000000001001;
assign LUT_3[34864] = 32'b11111111111111111110111001001111;
assign LUT_3[34865] = 32'b00000000000000000101100100101100;
assign LUT_3[34866] = 32'b00000000000000000001000000110011;
assign LUT_3[34867] = 32'b00000000000000000111101100010000;
assign LUT_3[34868] = 32'b11111111111111111100000111000101;
assign LUT_3[34869] = 32'b00000000000000000010110010100010;
assign LUT_3[34870] = 32'b11111111111111111110001110101001;
assign LUT_3[34871] = 32'b00000000000000000100111010000110;
assign LUT_3[34872] = 32'b00000000000000000100010010010101;
assign LUT_3[34873] = 32'b00000000000000001010111101110010;
assign LUT_3[34874] = 32'b00000000000000000110011001111001;
assign LUT_3[34875] = 32'b00000000000000001101000101010110;
assign LUT_3[34876] = 32'b00000000000000000001100000001011;
assign LUT_3[34877] = 32'b00000000000000001000001011101000;
assign LUT_3[34878] = 32'b00000000000000000011100111101111;
assign LUT_3[34879] = 32'b00000000000000001010010011001100;
assign LUT_3[34880] = 32'b11111111111111111010010000010111;
assign LUT_3[34881] = 32'b00000000000000000000111011110100;
assign LUT_3[34882] = 32'b11111111111111111100010111111011;
assign LUT_3[34883] = 32'b00000000000000000011000011011000;
assign LUT_3[34884] = 32'b11111111111111110111011110001101;
assign LUT_3[34885] = 32'b11111111111111111110001001101010;
assign LUT_3[34886] = 32'b11111111111111111001100101110001;
assign LUT_3[34887] = 32'b00000000000000000000010001001110;
assign LUT_3[34888] = 32'b11111111111111111111101001011101;
assign LUT_3[34889] = 32'b00000000000000000110010100111010;
assign LUT_3[34890] = 32'b00000000000000000001110001000001;
assign LUT_3[34891] = 32'b00000000000000001000011100011110;
assign LUT_3[34892] = 32'b11111111111111111100110111010011;
assign LUT_3[34893] = 32'b00000000000000000011100010110000;
assign LUT_3[34894] = 32'b11111111111111111110111110110111;
assign LUT_3[34895] = 32'b00000000000000000101101010010100;
assign LUT_3[34896] = 32'b11111111111111111101100011011010;
assign LUT_3[34897] = 32'b00000000000000000100001110110111;
assign LUT_3[34898] = 32'b11111111111111111111101010111110;
assign LUT_3[34899] = 32'b00000000000000000110010110011011;
assign LUT_3[34900] = 32'b11111111111111111010110001010000;
assign LUT_3[34901] = 32'b00000000000000000001011100101101;
assign LUT_3[34902] = 32'b11111111111111111100111000110100;
assign LUT_3[34903] = 32'b00000000000000000011100100010001;
assign LUT_3[34904] = 32'b00000000000000000010111100100000;
assign LUT_3[34905] = 32'b00000000000000001001100111111101;
assign LUT_3[34906] = 32'b00000000000000000101000100000100;
assign LUT_3[34907] = 32'b00000000000000001011101111100001;
assign LUT_3[34908] = 32'b00000000000000000000001010010110;
assign LUT_3[34909] = 32'b00000000000000000110110101110011;
assign LUT_3[34910] = 32'b00000000000000000010010001111010;
assign LUT_3[34911] = 32'b00000000000000001000111101010111;
assign LUT_3[34912] = 32'b11111111111111111011011110110111;
assign LUT_3[34913] = 32'b00000000000000000010001010010100;
assign LUT_3[34914] = 32'b11111111111111111101100110011011;
assign LUT_3[34915] = 32'b00000000000000000100010001111000;
assign LUT_3[34916] = 32'b11111111111111111000101100101101;
assign LUT_3[34917] = 32'b11111111111111111111011000001010;
assign LUT_3[34918] = 32'b11111111111111111010110100010001;
assign LUT_3[34919] = 32'b00000000000000000001011111101110;
assign LUT_3[34920] = 32'b00000000000000000000110111111101;
assign LUT_3[34921] = 32'b00000000000000000111100011011010;
assign LUT_3[34922] = 32'b00000000000000000010111111100001;
assign LUT_3[34923] = 32'b00000000000000001001101010111110;
assign LUT_3[34924] = 32'b11111111111111111110000101110011;
assign LUT_3[34925] = 32'b00000000000000000100110001010000;
assign LUT_3[34926] = 32'b00000000000000000000001101010111;
assign LUT_3[34927] = 32'b00000000000000000110111000110100;
assign LUT_3[34928] = 32'b11111111111111111110110001111010;
assign LUT_3[34929] = 32'b00000000000000000101011101010111;
assign LUT_3[34930] = 32'b00000000000000000000111001011110;
assign LUT_3[34931] = 32'b00000000000000000111100100111011;
assign LUT_3[34932] = 32'b11111111111111111011111111110000;
assign LUT_3[34933] = 32'b00000000000000000010101011001101;
assign LUT_3[34934] = 32'b11111111111111111110000111010100;
assign LUT_3[34935] = 32'b00000000000000000100110010110001;
assign LUT_3[34936] = 32'b00000000000000000100001011000000;
assign LUT_3[34937] = 32'b00000000000000001010110110011101;
assign LUT_3[34938] = 32'b00000000000000000110010010100100;
assign LUT_3[34939] = 32'b00000000000000001100111110000001;
assign LUT_3[34940] = 32'b00000000000000000001011000110110;
assign LUT_3[34941] = 32'b00000000000000001000000100010011;
assign LUT_3[34942] = 32'b00000000000000000011100000011010;
assign LUT_3[34943] = 32'b00000000000000001010001011110111;
assign LUT_3[34944] = 32'b11111111111111111100100010101010;
assign LUT_3[34945] = 32'b00000000000000000011001110000111;
assign LUT_3[34946] = 32'b11111111111111111110101010001110;
assign LUT_3[34947] = 32'b00000000000000000101010101101011;
assign LUT_3[34948] = 32'b11111111111111111001110000100000;
assign LUT_3[34949] = 32'b00000000000000000000011011111101;
assign LUT_3[34950] = 32'b11111111111111111011111000000100;
assign LUT_3[34951] = 32'b00000000000000000010100011100001;
assign LUT_3[34952] = 32'b00000000000000000001111011110000;
assign LUT_3[34953] = 32'b00000000000000001000100111001101;
assign LUT_3[34954] = 32'b00000000000000000100000011010100;
assign LUT_3[34955] = 32'b00000000000000001010101110110001;
assign LUT_3[34956] = 32'b11111111111111111111001001100110;
assign LUT_3[34957] = 32'b00000000000000000101110101000011;
assign LUT_3[34958] = 32'b00000000000000000001010001001010;
assign LUT_3[34959] = 32'b00000000000000000111111100100111;
assign LUT_3[34960] = 32'b11111111111111111111110101101101;
assign LUT_3[34961] = 32'b00000000000000000110100001001010;
assign LUT_3[34962] = 32'b00000000000000000001111101010001;
assign LUT_3[34963] = 32'b00000000000000001000101000101110;
assign LUT_3[34964] = 32'b11111111111111111101000011100011;
assign LUT_3[34965] = 32'b00000000000000000011101111000000;
assign LUT_3[34966] = 32'b11111111111111111111001011000111;
assign LUT_3[34967] = 32'b00000000000000000101110110100100;
assign LUT_3[34968] = 32'b00000000000000000101001110110011;
assign LUT_3[34969] = 32'b00000000000000001011111010010000;
assign LUT_3[34970] = 32'b00000000000000000111010110010111;
assign LUT_3[34971] = 32'b00000000000000001110000001110100;
assign LUT_3[34972] = 32'b00000000000000000010011100101001;
assign LUT_3[34973] = 32'b00000000000000001001001000000110;
assign LUT_3[34974] = 32'b00000000000000000100100100001101;
assign LUT_3[34975] = 32'b00000000000000001011001111101010;
assign LUT_3[34976] = 32'b11111111111111111101110001001010;
assign LUT_3[34977] = 32'b00000000000000000100011100100111;
assign LUT_3[34978] = 32'b11111111111111111111111000101110;
assign LUT_3[34979] = 32'b00000000000000000110100100001011;
assign LUT_3[34980] = 32'b11111111111111111010111111000000;
assign LUT_3[34981] = 32'b00000000000000000001101010011101;
assign LUT_3[34982] = 32'b11111111111111111101000110100100;
assign LUT_3[34983] = 32'b00000000000000000011110010000001;
assign LUT_3[34984] = 32'b00000000000000000011001010010000;
assign LUT_3[34985] = 32'b00000000000000001001110101101101;
assign LUT_3[34986] = 32'b00000000000000000101010001110100;
assign LUT_3[34987] = 32'b00000000000000001011111101010001;
assign LUT_3[34988] = 32'b00000000000000000000011000000110;
assign LUT_3[34989] = 32'b00000000000000000111000011100011;
assign LUT_3[34990] = 32'b00000000000000000010011111101010;
assign LUT_3[34991] = 32'b00000000000000001001001011000111;
assign LUT_3[34992] = 32'b00000000000000000001000100001101;
assign LUT_3[34993] = 32'b00000000000000000111101111101010;
assign LUT_3[34994] = 32'b00000000000000000011001011110001;
assign LUT_3[34995] = 32'b00000000000000001001110111001110;
assign LUT_3[34996] = 32'b11111111111111111110010010000011;
assign LUT_3[34997] = 32'b00000000000000000100111101100000;
assign LUT_3[34998] = 32'b00000000000000000000011001100111;
assign LUT_3[34999] = 32'b00000000000000000111000101000100;
assign LUT_3[35000] = 32'b00000000000000000110011101010011;
assign LUT_3[35001] = 32'b00000000000000001101001000110000;
assign LUT_3[35002] = 32'b00000000000000001000100100110111;
assign LUT_3[35003] = 32'b00000000000000001111010000010100;
assign LUT_3[35004] = 32'b00000000000000000011101011001001;
assign LUT_3[35005] = 32'b00000000000000001010010110100110;
assign LUT_3[35006] = 32'b00000000000000000101110010101101;
assign LUT_3[35007] = 32'b00000000000000001100011110001010;
assign LUT_3[35008] = 32'b11111111111111111100011011010101;
assign LUT_3[35009] = 32'b00000000000000000011000110110010;
assign LUT_3[35010] = 32'b11111111111111111110100010111001;
assign LUT_3[35011] = 32'b00000000000000000101001110010110;
assign LUT_3[35012] = 32'b11111111111111111001101001001011;
assign LUT_3[35013] = 32'b00000000000000000000010100101000;
assign LUT_3[35014] = 32'b11111111111111111011110000101111;
assign LUT_3[35015] = 32'b00000000000000000010011100001100;
assign LUT_3[35016] = 32'b00000000000000000001110100011011;
assign LUT_3[35017] = 32'b00000000000000001000011111111000;
assign LUT_3[35018] = 32'b00000000000000000011111011111111;
assign LUT_3[35019] = 32'b00000000000000001010100111011100;
assign LUT_3[35020] = 32'b11111111111111111111000010010001;
assign LUT_3[35021] = 32'b00000000000000000101101101101110;
assign LUT_3[35022] = 32'b00000000000000000001001001110101;
assign LUT_3[35023] = 32'b00000000000000000111110101010010;
assign LUT_3[35024] = 32'b11111111111111111111101110011000;
assign LUT_3[35025] = 32'b00000000000000000110011001110101;
assign LUT_3[35026] = 32'b00000000000000000001110101111100;
assign LUT_3[35027] = 32'b00000000000000001000100001011001;
assign LUT_3[35028] = 32'b11111111111111111100111100001110;
assign LUT_3[35029] = 32'b00000000000000000011100111101011;
assign LUT_3[35030] = 32'b11111111111111111111000011110010;
assign LUT_3[35031] = 32'b00000000000000000101101111001111;
assign LUT_3[35032] = 32'b00000000000000000101000111011110;
assign LUT_3[35033] = 32'b00000000000000001011110010111011;
assign LUT_3[35034] = 32'b00000000000000000111001111000010;
assign LUT_3[35035] = 32'b00000000000000001101111010011111;
assign LUT_3[35036] = 32'b00000000000000000010010101010100;
assign LUT_3[35037] = 32'b00000000000000001001000000110001;
assign LUT_3[35038] = 32'b00000000000000000100011100111000;
assign LUT_3[35039] = 32'b00000000000000001011001000010101;
assign LUT_3[35040] = 32'b11111111111111111101101001110101;
assign LUT_3[35041] = 32'b00000000000000000100010101010010;
assign LUT_3[35042] = 32'b11111111111111111111110001011001;
assign LUT_3[35043] = 32'b00000000000000000110011100110110;
assign LUT_3[35044] = 32'b11111111111111111010110111101011;
assign LUT_3[35045] = 32'b00000000000000000001100011001000;
assign LUT_3[35046] = 32'b11111111111111111100111111001111;
assign LUT_3[35047] = 32'b00000000000000000011101010101100;
assign LUT_3[35048] = 32'b00000000000000000011000010111011;
assign LUT_3[35049] = 32'b00000000000000001001101110011000;
assign LUT_3[35050] = 32'b00000000000000000101001010011111;
assign LUT_3[35051] = 32'b00000000000000001011110101111100;
assign LUT_3[35052] = 32'b00000000000000000000010000110001;
assign LUT_3[35053] = 32'b00000000000000000110111100001110;
assign LUT_3[35054] = 32'b00000000000000000010011000010101;
assign LUT_3[35055] = 32'b00000000000000001001000011110010;
assign LUT_3[35056] = 32'b00000000000000000000111100111000;
assign LUT_3[35057] = 32'b00000000000000000111101000010101;
assign LUT_3[35058] = 32'b00000000000000000011000100011100;
assign LUT_3[35059] = 32'b00000000000000001001101111111001;
assign LUT_3[35060] = 32'b11111111111111111110001010101110;
assign LUT_3[35061] = 32'b00000000000000000100110110001011;
assign LUT_3[35062] = 32'b00000000000000000000010010010010;
assign LUT_3[35063] = 32'b00000000000000000110111101101111;
assign LUT_3[35064] = 32'b00000000000000000110010101111110;
assign LUT_3[35065] = 32'b00000000000000001101000001011011;
assign LUT_3[35066] = 32'b00000000000000001000011101100010;
assign LUT_3[35067] = 32'b00000000000000001111001000111111;
assign LUT_3[35068] = 32'b00000000000000000011100011110100;
assign LUT_3[35069] = 32'b00000000000000001010001111010001;
assign LUT_3[35070] = 32'b00000000000000000101101011011000;
assign LUT_3[35071] = 32'b00000000000000001100010110110101;
assign LUT_3[35072] = 32'b11111111111111110110100111001101;
assign LUT_3[35073] = 32'b11111111111111111101010010101010;
assign LUT_3[35074] = 32'b11111111111111111000101110110001;
assign LUT_3[35075] = 32'b11111111111111111111011010001110;
assign LUT_3[35076] = 32'b11111111111111110011110101000011;
assign LUT_3[35077] = 32'b11111111111111111010100000100000;
assign LUT_3[35078] = 32'b11111111111111110101111100100111;
assign LUT_3[35079] = 32'b11111111111111111100101000000100;
assign LUT_3[35080] = 32'b11111111111111111100000000010011;
assign LUT_3[35081] = 32'b00000000000000000010101011110000;
assign LUT_3[35082] = 32'b11111111111111111110000111110111;
assign LUT_3[35083] = 32'b00000000000000000100110011010100;
assign LUT_3[35084] = 32'b11111111111111111001001110001001;
assign LUT_3[35085] = 32'b11111111111111111111111001100110;
assign LUT_3[35086] = 32'b11111111111111111011010101101101;
assign LUT_3[35087] = 32'b00000000000000000010000001001010;
assign LUT_3[35088] = 32'b11111111111111111001111010010000;
assign LUT_3[35089] = 32'b00000000000000000000100101101101;
assign LUT_3[35090] = 32'b11111111111111111100000001110100;
assign LUT_3[35091] = 32'b00000000000000000010101101010001;
assign LUT_3[35092] = 32'b11111111111111110111001000000110;
assign LUT_3[35093] = 32'b11111111111111111101110011100011;
assign LUT_3[35094] = 32'b11111111111111111001001111101010;
assign LUT_3[35095] = 32'b11111111111111111111111011000111;
assign LUT_3[35096] = 32'b11111111111111111111010011010110;
assign LUT_3[35097] = 32'b00000000000000000101111110110011;
assign LUT_3[35098] = 32'b00000000000000000001011010111010;
assign LUT_3[35099] = 32'b00000000000000001000000110010111;
assign LUT_3[35100] = 32'b11111111111111111100100001001100;
assign LUT_3[35101] = 32'b00000000000000000011001100101001;
assign LUT_3[35102] = 32'b11111111111111111110101000110000;
assign LUT_3[35103] = 32'b00000000000000000101010100001101;
assign LUT_3[35104] = 32'b11111111111111110111110101101101;
assign LUT_3[35105] = 32'b11111111111111111110100001001010;
assign LUT_3[35106] = 32'b11111111111111111001111101010001;
assign LUT_3[35107] = 32'b00000000000000000000101000101110;
assign LUT_3[35108] = 32'b11111111111111110101000011100011;
assign LUT_3[35109] = 32'b11111111111111111011101111000000;
assign LUT_3[35110] = 32'b11111111111111110111001011000111;
assign LUT_3[35111] = 32'b11111111111111111101110110100100;
assign LUT_3[35112] = 32'b11111111111111111101001110110011;
assign LUT_3[35113] = 32'b00000000000000000011111010010000;
assign LUT_3[35114] = 32'b11111111111111111111010110010111;
assign LUT_3[35115] = 32'b00000000000000000110000001110100;
assign LUT_3[35116] = 32'b11111111111111111010011100101001;
assign LUT_3[35117] = 32'b00000000000000000001001000000110;
assign LUT_3[35118] = 32'b11111111111111111100100100001101;
assign LUT_3[35119] = 32'b00000000000000000011001111101010;
assign LUT_3[35120] = 32'b11111111111111111011001000110000;
assign LUT_3[35121] = 32'b00000000000000000001110100001101;
assign LUT_3[35122] = 32'b11111111111111111101010000010100;
assign LUT_3[35123] = 32'b00000000000000000011111011110001;
assign LUT_3[35124] = 32'b11111111111111111000010110100110;
assign LUT_3[35125] = 32'b11111111111111111111000010000011;
assign LUT_3[35126] = 32'b11111111111111111010011110001010;
assign LUT_3[35127] = 32'b00000000000000000001001001100111;
assign LUT_3[35128] = 32'b00000000000000000000100001110110;
assign LUT_3[35129] = 32'b00000000000000000111001101010011;
assign LUT_3[35130] = 32'b00000000000000000010101001011010;
assign LUT_3[35131] = 32'b00000000000000001001010100110111;
assign LUT_3[35132] = 32'b11111111111111111101101111101100;
assign LUT_3[35133] = 32'b00000000000000000100011011001001;
assign LUT_3[35134] = 32'b11111111111111111111110111010000;
assign LUT_3[35135] = 32'b00000000000000000110100010101101;
assign LUT_3[35136] = 32'b11111111111111110110011111111000;
assign LUT_3[35137] = 32'b11111111111111111101001011010101;
assign LUT_3[35138] = 32'b11111111111111111000100111011100;
assign LUT_3[35139] = 32'b11111111111111111111010010111001;
assign LUT_3[35140] = 32'b11111111111111110011101101101110;
assign LUT_3[35141] = 32'b11111111111111111010011001001011;
assign LUT_3[35142] = 32'b11111111111111110101110101010010;
assign LUT_3[35143] = 32'b11111111111111111100100000101111;
assign LUT_3[35144] = 32'b11111111111111111011111000111110;
assign LUT_3[35145] = 32'b00000000000000000010100100011011;
assign LUT_3[35146] = 32'b11111111111111111110000000100010;
assign LUT_3[35147] = 32'b00000000000000000100101011111111;
assign LUT_3[35148] = 32'b11111111111111111001000110110100;
assign LUT_3[35149] = 32'b11111111111111111111110010010001;
assign LUT_3[35150] = 32'b11111111111111111011001110011000;
assign LUT_3[35151] = 32'b00000000000000000001111001110101;
assign LUT_3[35152] = 32'b11111111111111111001110010111011;
assign LUT_3[35153] = 32'b00000000000000000000011110011000;
assign LUT_3[35154] = 32'b11111111111111111011111010011111;
assign LUT_3[35155] = 32'b00000000000000000010100101111100;
assign LUT_3[35156] = 32'b11111111111111110111000000110001;
assign LUT_3[35157] = 32'b11111111111111111101101100001110;
assign LUT_3[35158] = 32'b11111111111111111001001000010101;
assign LUT_3[35159] = 32'b11111111111111111111110011110010;
assign LUT_3[35160] = 32'b11111111111111111111001100000001;
assign LUT_3[35161] = 32'b00000000000000000101110111011110;
assign LUT_3[35162] = 32'b00000000000000000001010011100101;
assign LUT_3[35163] = 32'b00000000000000000111111111000010;
assign LUT_3[35164] = 32'b11111111111111111100011001110111;
assign LUT_3[35165] = 32'b00000000000000000011000101010100;
assign LUT_3[35166] = 32'b11111111111111111110100001011011;
assign LUT_3[35167] = 32'b00000000000000000101001100111000;
assign LUT_3[35168] = 32'b11111111111111110111101110011000;
assign LUT_3[35169] = 32'b11111111111111111110011001110101;
assign LUT_3[35170] = 32'b11111111111111111001110101111100;
assign LUT_3[35171] = 32'b00000000000000000000100001011001;
assign LUT_3[35172] = 32'b11111111111111110100111100001110;
assign LUT_3[35173] = 32'b11111111111111111011100111101011;
assign LUT_3[35174] = 32'b11111111111111110111000011110010;
assign LUT_3[35175] = 32'b11111111111111111101101111001111;
assign LUT_3[35176] = 32'b11111111111111111101000111011110;
assign LUT_3[35177] = 32'b00000000000000000011110010111011;
assign LUT_3[35178] = 32'b11111111111111111111001111000010;
assign LUT_3[35179] = 32'b00000000000000000101111010011111;
assign LUT_3[35180] = 32'b11111111111111111010010101010100;
assign LUT_3[35181] = 32'b00000000000000000001000000110001;
assign LUT_3[35182] = 32'b11111111111111111100011100111000;
assign LUT_3[35183] = 32'b00000000000000000011001000010101;
assign LUT_3[35184] = 32'b11111111111111111011000001011011;
assign LUT_3[35185] = 32'b00000000000000000001101100111000;
assign LUT_3[35186] = 32'b11111111111111111101001000111111;
assign LUT_3[35187] = 32'b00000000000000000011110100011100;
assign LUT_3[35188] = 32'b11111111111111111000001111010001;
assign LUT_3[35189] = 32'b11111111111111111110111010101110;
assign LUT_3[35190] = 32'b11111111111111111010010110110101;
assign LUT_3[35191] = 32'b00000000000000000001000010010010;
assign LUT_3[35192] = 32'b00000000000000000000011010100001;
assign LUT_3[35193] = 32'b00000000000000000111000101111110;
assign LUT_3[35194] = 32'b00000000000000000010100010000101;
assign LUT_3[35195] = 32'b00000000000000001001001101100010;
assign LUT_3[35196] = 32'b11111111111111111101101000010111;
assign LUT_3[35197] = 32'b00000000000000000100010011110100;
assign LUT_3[35198] = 32'b11111111111111111111101111111011;
assign LUT_3[35199] = 32'b00000000000000000110011011011000;
assign LUT_3[35200] = 32'b11111111111111111000110010001011;
assign LUT_3[35201] = 32'b11111111111111111111011101101000;
assign LUT_3[35202] = 32'b11111111111111111010111001101111;
assign LUT_3[35203] = 32'b00000000000000000001100101001100;
assign LUT_3[35204] = 32'b11111111111111110110000000000001;
assign LUT_3[35205] = 32'b11111111111111111100101011011110;
assign LUT_3[35206] = 32'b11111111111111111000000111100101;
assign LUT_3[35207] = 32'b11111111111111111110110011000010;
assign LUT_3[35208] = 32'b11111111111111111110001011010001;
assign LUT_3[35209] = 32'b00000000000000000100110110101110;
assign LUT_3[35210] = 32'b00000000000000000000010010110101;
assign LUT_3[35211] = 32'b00000000000000000110111110010010;
assign LUT_3[35212] = 32'b11111111111111111011011001000111;
assign LUT_3[35213] = 32'b00000000000000000010000100100100;
assign LUT_3[35214] = 32'b11111111111111111101100000101011;
assign LUT_3[35215] = 32'b00000000000000000100001100001000;
assign LUT_3[35216] = 32'b11111111111111111100000101001110;
assign LUT_3[35217] = 32'b00000000000000000010110000101011;
assign LUT_3[35218] = 32'b11111111111111111110001100110010;
assign LUT_3[35219] = 32'b00000000000000000100111000001111;
assign LUT_3[35220] = 32'b11111111111111111001010011000100;
assign LUT_3[35221] = 32'b11111111111111111111111110100001;
assign LUT_3[35222] = 32'b11111111111111111011011010101000;
assign LUT_3[35223] = 32'b00000000000000000010000110000101;
assign LUT_3[35224] = 32'b00000000000000000001011110010100;
assign LUT_3[35225] = 32'b00000000000000001000001001110001;
assign LUT_3[35226] = 32'b00000000000000000011100101111000;
assign LUT_3[35227] = 32'b00000000000000001010010001010101;
assign LUT_3[35228] = 32'b11111111111111111110101100001010;
assign LUT_3[35229] = 32'b00000000000000000101010111100111;
assign LUT_3[35230] = 32'b00000000000000000000110011101110;
assign LUT_3[35231] = 32'b00000000000000000111011111001011;
assign LUT_3[35232] = 32'b11111111111111111010000000101011;
assign LUT_3[35233] = 32'b00000000000000000000101100001000;
assign LUT_3[35234] = 32'b11111111111111111100001000001111;
assign LUT_3[35235] = 32'b00000000000000000010110011101100;
assign LUT_3[35236] = 32'b11111111111111110111001110100001;
assign LUT_3[35237] = 32'b11111111111111111101111001111110;
assign LUT_3[35238] = 32'b11111111111111111001010110000101;
assign LUT_3[35239] = 32'b00000000000000000000000001100010;
assign LUT_3[35240] = 32'b11111111111111111111011001110001;
assign LUT_3[35241] = 32'b00000000000000000110000101001110;
assign LUT_3[35242] = 32'b00000000000000000001100001010101;
assign LUT_3[35243] = 32'b00000000000000001000001100110010;
assign LUT_3[35244] = 32'b11111111111111111100100111100111;
assign LUT_3[35245] = 32'b00000000000000000011010011000100;
assign LUT_3[35246] = 32'b11111111111111111110101111001011;
assign LUT_3[35247] = 32'b00000000000000000101011010101000;
assign LUT_3[35248] = 32'b11111111111111111101010011101110;
assign LUT_3[35249] = 32'b00000000000000000011111111001011;
assign LUT_3[35250] = 32'b11111111111111111111011011010010;
assign LUT_3[35251] = 32'b00000000000000000110000110101111;
assign LUT_3[35252] = 32'b11111111111111111010100001100100;
assign LUT_3[35253] = 32'b00000000000000000001001101000001;
assign LUT_3[35254] = 32'b11111111111111111100101001001000;
assign LUT_3[35255] = 32'b00000000000000000011010100100101;
assign LUT_3[35256] = 32'b00000000000000000010101100110100;
assign LUT_3[35257] = 32'b00000000000000001001011000010001;
assign LUT_3[35258] = 32'b00000000000000000100110100011000;
assign LUT_3[35259] = 32'b00000000000000001011011111110101;
assign LUT_3[35260] = 32'b11111111111111111111111010101010;
assign LUT_3[35261] = 32'b00000000000000000110100110000111;
assign LUT_3[35262] = 32'b00000000000000000010000010001110;
assign LUT_3[35263] = 32'b00000000000000001000101101101011;
assign LUT_3[35264] = 32'b11111111111111111000101010110110;
assign LUT_3[35265] = 32'b11111111111111111111010110010011;
assign LUT_3[35266] = 32'b11111111111111111010110010011010;
assign LUT_3[35267] = 32'b00000000000000000001011101110111;
assign LUT_3[35268] = 32'b11111111111111110101111000101100;
assign LUT_3[35269] = 32'b11111111111111111100100100001001;
assign LUT_3[35270] = 32'b11111111111111111000000000010000;
assign LUT_3[35271] = 32'b11111111111111111110101011101101;
assign LUT_3[35272] = 32'b11111111111111111110000011111100;
assign LUT_3[35273] = 32'b00000000000000000100101111011001;
assign LUT_3[35274] = 32'b00000000000000000000001011100000;
assign LUT_3[35275] = 32'b00000000000000000110110110111101;
assign LUT_3[35276] = 32'b11111111111111111011010001110010;
assign LUT_3[35277] = 32'b00000000000000000001111101001111;
assign LUT_3[35278] = 32'b11111111111111111101011001010110;
assign LUT_3[35279] = 32'b00000000000000000100000100110011;
assign LUT_3[35280] = 32'b11111111111111111011111101111001;
assign LUT_3[35281] = 32'b00000000000000000010101001010110;
assign LUT_3[35282] = 32'b11111111111111111110000101011101;
assign LUT_3[35283] = 32'b00000000000000000100110000111010;
assign LUT_3[35284] = 32'b11111111111111111001001011101111;
assign LUT_3[35285] = 32'b11111111111111111111110111001100;
assign LUT_3[35286] = 32'b11111111111111111011010011010011;
assign LUT_3[35287] = 32'b00000000000000000001111110110000;
assign LUT_3[35288] = 32'b00000000000000000001010110111111;
assign LUT_3[35289] = 32'b00000000000000001000000010011100;
assign LUT_3[35290] = 32'b00000000000000000011011110100011;
assign LUT_3[35291] = 32'b00000000000000001010001010000000;
assign LUT_3[35292] = 32'b11111111111111111110100100110101;
assign LUT_3[35293] = 32'b00000000000000000101010000010010;
assign LUT_3[35294] = 32'b00000000000000000000101100011001;
assign LUT_3[35295] = 32'b00000000000000000111010111110110;
assign LUT_3[35296] = 32'b11111111111111111001111001010110;
assign LUT_3[35297] = 32'b00000000000000000000100100110011;
assign LUT_3[35298] = 32'b11111111111111111100000000111010;
assign LUT_3[35299] = 32'b00000000000000000010101100010111;
assign LUT_3[35300] = 32'b11111111111111110111000111001100;
assign LUT_3[35301] = 32'b11111111111111111101110010101001;
assign LUT_3[35302] = 32'b11111111111111111001001110110000;
assign LUT_3[35303] = 32'b11111111111111111111111010001101;
assign LUT_3[35304] = 32'b11111111111111111111010010011100;
assign LUT_3[35305] = 32'b00000000000000000101111101111001;
assign LUT_3[35306] = 32'b00000000000000000001011010000000;
assign LUT_3[35307] = 32'b00000000000000001000000101011101;
assign LUT_3[35308] = 32'b11111111111111111100100000010010;
assign LUT_3[35309] = 32'b00000000000000000011001011101111;
assign LUT_3[35310] = 32'b11111111111111111110100111110110;
assign LUT_3[35311] = 32'b00000000000000000101010011010011;
assign LUT_3[35312] = 32'b11111111111111111101001100011001;
assign LUT_3[35313] = 32'b00000000000000000011110111110110;
assign LUT_3[35314] = 32'b11111111111111111111010011111101;
assign LUT_3[35315] = 32'b00000000000000000101111111011010;
assign LUT_3[35316] = 32'b11111111111111111010011010001111;
assign LUT_3[35317] = 32'b00000000000000000001000101101100;
assign LUT_3[35318] = 32'b11111111111111111100100001110011;
assign LUT_3[35319] = 32'b00000000000000000011001101010000;
assign LUT_3[35320] = 32'b00000000000000000010100101011111;
assign LUT_3[35321] = 32'b00000000000000001001010000111100;
assign LUT_3[35322] = 32'b00000000000000000100101101000011;
assign LUT_3[35323] = 32'b00000000000000001011011000100000;
assign LUT_3[35324] = 32'b11111111111111111111110011010101;
assign LUT_3[35325] = 32'b00000000000000000110011110110010;
assign LUT_3[35326] = 32'b00000000000000000001111010111001;
assign LUT_3[35327] = 32'b00000000000000001000100110010110;
assign LUT_3[35328] = 32'b11111111111111111101101100111000;
assign LUT_3[35329] = 32'b00000000000000000100011000010101;
assign LUT_3[35330] = 32'b11111111111111111111110100011100;
assign LUT_3[35331] = 32'b00000000000000000110011111111001;
assign LUT_3[35332] = 32'b11111111111111111010111010101110;
assign LUT_3[35333] = 32'b00000000000000000001100110001011;
assign LUT_3[35334] = 32'b11111111111111111101000010010010;
assign LUT_3[35335] = 32'b00000000000000000011101101101111;
assign LUT_3[35336] = 32'b00000000000000000011000101111110;
assign LUT_3[35337] = 32'b00000000000000001001110001011011;
assign LUT_3[35338] = 32'b00000000000000000101001101100010;
assign LUT_3[35339] = 32'b00000000000000001011111000111111;
assign LUT_3[35340] = 32'b00000000000000000000010011110100;
assign LUT_3[35341] = 32'b00000000000000000110111111010001;
assign LUT_3[35342] = 32'b00000000000000000010011011011000;
assign LUT_3[35343] = 32'b00000000000000001001000110110101;
assign LUT_3[35344] = 32'b00000000000000000000111111111011;
assign LUT_3[35345] = 32'b00000000000000000111101011011000;
assign LUT_3[35346] = 32'b00000000000000000011000111011111;
assign LUT_3[35347] = 32'b00000000000000001001110010111100;
assign LUT_3[35348] = 32'b11111111111111111110001101110001;
assign LUT_3[35349] = 32'b00000000000000000100111001001110;
assign LUT_3[35350] = 32'b00000000000000000000010101010101;
assign LUT_3[35351] = 32'b00000000000000000111000000110010;
assign LUT_3[35352] = 32'b00000000000000000110011001000001;
assign LUT_3[35353] = 32'b00000000000000001101000100011110;
assign LUT_3[35354] = 32'b00000000000000001000100000100101;
assign LUT_3[35355] = 32'b00000000000000001111001100000010;
assign LUT_3[35356] = 32'b00000000000000000011100110110111;
assign LUT_3[35357] = 32'b00000000000000001010010010010100;
assign LUT_3[35358] = 32'b00000000000000000101101110011011;
assign LUT_3[35359] = 32'b00000000000000001100011001111000;
assign LUT_3[35360] = 32'b11111111111111111110111011011000;
assign LUT_3[35361] = 32'b00000000000000000101100110110101;
assign LUT_3[35362] = 32'b00000000000000000001000010111100;
assign LUT_3[35363] = 32'b00000000000000000111101110011001;
assign LUT_3[35364] = 32'b11111111111111111100001001001110;
assign LUT_3[35365] = 32'b00000000000000000010110100101011;
assign LUT_3[35366] = 32'b11111111111111111110010000110010;
assign LUT_3[35367] = 32'b00000000000000000100111100001111;
assign LUT_3[35368] = 32'b00000000000000000100010100011110;
assign LUT_3[35369] = 32'b00000000000000001010111111111011;
assign LUT_3[35370] = 32'b00000000000000000110011100000010;
assign LUT_3[35371] = 32'b00000000000000001101000111011111;
assign LUT_3[35372] = 32'b00000000000000000001100010010100;
assign LUT_3[35373] = 32'b00000000000000001000001101110001;
assign LUT_3[35374] = 32'b00000000000000000011101001111000;
assign LUT_3[35375] = 32'b00000000000000001010010101010101;
assign LUT_3[35376] = 32'b00000000000000000010001110011011;
assign LUT_3[35377] = 32'b00000000000000001000111001111000;
assign LUT_3[35378] = 32'b00000000000000000100010101111111;
assign LUT_3[35379] = 32'b00000000000000001011000001011100;
assign LUT_3[35380] = 32'b11111111111111111111011100010001;
assign LUT_3[35381] = 32'b00000000000000000110000111101110;
assign LUT_3[35382] = 32'b00000000000000000001100011110101;
assign LUT_3[35383] = 32'b00000000000000001000001111010010;
assign LUT_3[35384] = 32'b00000000000000000111100111100001;
assign LUT_3[35385] = 32'b00000000000000001110010010111110;
assign LUT_3[35386] = 32'b00000000000000001001101111000101;
assign LUT_3[35387] = 32'b00000000000000010000011010100010;
assign LUT_3[35388] = 32'b00000000000000000100110101010111;
assign LUT_3[35389] = 32'b00000000000000001011100000110100;
assign LUT_3[35390] = 32'b00000000000000000110111100111011;
assign LUT_3[35391] = 32'b00000000000000001101101000011000;
assign LUT_3[35392] = 32'b11111111111111111101100101100011;
assign LUT_3[35393] = 32'b00000000000000000100010001000000;
assign LUT_3[35394] = 32'b11111111111111111111101101000111;
assign LUT_3[35395] = 32'b00000000000000000110011000100100;
assign LUT_3[35396] = 32'b11111111111111111010110011011001;
assign LUT_3[35397] = 32'b00000000000000000001011110110110;
assign LUT_3[35398] = 32'b11111111111111111100111010111101;
assign LUT_3[35399] = 32'b00000000000000000011100110011010;
assign LUT_3[35400] = 32'b00000000000000000010111110101001;
assign LUT_3[35401] = 32'b00000000000000001001101010000110;
assign LUT_3[35402] = 32'b00000000000000000101000110001101;
assign LUT_3[35403] = 32'b00000000000000001011110001101010;
assign LUT_3[35404] = 32'b00000000000000000000001100011111;
assign LUT_3[35405] = 32'b00000000000000000110110111111100;
assign LUT_3[35406] = 32'b00000000000000000010010100000011;
assign LUT_3[35407] = 32'b00000000000000001000111111100000;
assign LUT_3[35408] = 32'b00000000000000000000111000100110;
assign LUT_3[35409] = 32'b00000000000000000111100100000011;
assign LUT_3[35410] = 32'b00000000000000000011000000001010;
assign LUT_3[35411] = 32'b00000000000000001001101011100111;
assign LUT_3[35412] = 32'b11111111111111111110000110011100;
assign LUT_3[35413] = 32'b00000000000000000100110001111001;
assign LUT_3[35414] = 32'b00000000000000000000001110000000;
assign LUT_3[35415] = 32'b00000000000000000110111001011101;
assign LUT_3[35416] = 32'b00000000000000000110010001101100;
assign LUT_3[35417] = 32'b00000000000000001100111101001001;
assign LUT_3[35418] = 32'b00000000000000001000011001010000;
assign LUT_3[35419] = 32'b00000000000000001111000100101101;
assign LUT_3[35420] = 32'b00000000000000000011011111100010;
assign LUT_3[35421] = 32'b00000000000000001010001010111111;
assign LUT_3[35422] = 32'b00000000000000000101100111000110;
assign LUT_3[35423] = 32'b00000000000000001100010010100011;
assign LUT_3[35424] = 32'b11111111111111111110110100000011;
assign LUT_3[35425] = 32'b00000000000000000101011111100000;
assign LUT_3[35426] = 32'b00000000000000000000111011100111;
assign LUT_3[35427] = 32'b00000000000000000111100111000100;
assign LUT_3[35428] = 32'b11111111111111111100000001111001;
assign LUT_3[35429] = 32'b00000000000000000010101101010110;
assign LUT_3[35430] = 32'b11111111111111111110001001011101;
assign LUT_3[35431] = 32'b00000000000000000100110100111010;
assign LUT_3[35432] = 32'b00000000000000000100001101001001;
assign LUT_3[35433] = 32'b00000000000000001010111000100110;
assign LUT_3[35434] = 32'b00000000000000000110010100101101;
assign LUT_3[35435] = 32'b00000000000000001101000000001010;
assign LUT_3[35436] = 32'b00000000000000000001011010111111;
assign LUT_3[35437] = 32'b00000000000000001000000110011100;
assign LUT_3[35438] = 32'b00000000000000000011100010100011;
assign LUT_3[35439] = 32'b00000000000000001010001110000000;
assign LUT_3[35440] = 32'b00000000000000000010000111000110;
assign LUT_3[35441] = 32'b00000000000000001000110010100011;
assign LUT_3[35442] = 32'b00000000000000000100001110101010;
assign LUT_3[35443] = 32'b00000000000000001010111010000111;
assign LUT_3[35444] = 32'b11111111111111111111010100111100;
assign LUT_3[35445] = 32'b00000000000000000110000000011001;
assign LUT_3[35446] = 32'b00000000000000000001011100100000;
assign LUT_3[35447] = 32'b00000000000000001000000111111101;
assign LUT_3[35448] = 32'b00000000000000000111100000001100;
assign LUT_3[35449] = 32'b00000000000000001110001011101001;
assign LUT_3[35450] = 32'b00000000000000001001100111110000;
assign LUT_3[35451] = 32'b00000000000000010000010011001101;
assign LUT_3[35452] = 32'b00000000000000000100101110000010;
assign LUT_3[35453] = 32'b00000000000000001011011001011111;
assign LUT_3[35454] = 32'b00000000000000000110110101100110;
assign LUT_3[35455] = 32'b00000000000000001101100001000011;
assign LUT_3[35456] = 32'b11111111111111111111110111110110;
assign LUT_3[35457] = 32'b00000000000000000110100011010011;
assign LUT_3[35458] = 32'b00000000000000000001111111011010;
assign LUT_3[35459] = 32'b00000000000000001000101010110111;
assign LUT_3[35460] = 32'b11111111111111111101000101101100;
assign LUT_3[35461] = 32'b00000000000000000011110001001001;
assign LUT_3[35462] = 32'b11111111111111111111001101010000;
assign LUT_3[35463] = 32'b00000000000000000101111000101101;
assign LUT_3[35464] = 32'b00000000000000000101010000111100;
assign LUT_3[35465] = 32'b00000000000000001011111100011001;
assign LUT_3[35466] = 32'b00000000000000000111011000100000;
assign LUT_3[35467] = 32'b00000000000000001110000011111101;
assign LUT_3[35468] = 32'b00000000000000000010011110110010;
assign LUT_3[35469] = 32'b00000000000000001001001010001111;
assign LUT_3[35470] = 32'b00000000000000000100100110010110;
assign LUT_3[35471] = 32'b00000000000000001011010001110011;
assign LUT_3[35472] = 32'b00000000000000000011001010111001;
assign LUT_3[35473] = 32'b00000000000000001001110110010110;
assign LUT_3[35474] = 32'b00000000000000000101010010011101;
assign LUT_3[35475] = 32'b00000000000000001011111101111010;
assign LUT_3[35476] = 32'b00000000000000000000011000101111;
assign LUT_3[35477] = 32'b00000000000000000111000100001100;
assign LUT_3[35478] = 32'b00000000000000000010100000010011;
assign LUT_3[35479] = 32'b00000000000000001001001011110000;
assign LUT_3[35480] = 32'b00000000000000001000100011111111;
assign LUT_3[35481] = 32'b00000000000000001111001111011100;
assign LUT_3[35482] = 32'b00000000000000001010101011100011;
assign LUT_3[35483] = 32'b00000000000000010001010111000000;
assign LUT_3[35484] = 32'b00000000000000000101110001110101;
assign LUT_3[35485] = 32'b00000000000000001100011101010010;
assign LUT_3[35486] = 32'b00000000000000000111111001011001;
assign LUT_3[35487] = 32'b00000000000000001110100100110110;
assign LUT_3[35488] = 32'b00000000000000000001000110010110;
assign LUT_3[35489] = 32'b00000000000000000111110001110011;
assign LUT_3[35490] = 32'b00000000000000000011001101111010;
assign LUT_3[35491] = 32'b00000000000000001001111001010111;
assign LUT_3[35492] = 32'b11111111111111111110010100001100;
assign LUT_3[35493] = 32'b00000000000000000100111111101001;
assign LUT_3[35494] = 32'b00000000000000000000011011110000;
assign LUT_3[35495] = 32'b00000000000000000111000111001101;
assign LUT_3[35496] = 32'b00000000000000000110011111011100;
assign LUT_3[35497] = 32'b00000000000000001101001010111001;
assign LUT_3[35498] = 32'b00000000000000001000100111000000;
assign LUT_3[35499] = 32'b00000000000000001111010010011101;
assign LUT_3[35500] = 32'b00000000000000000011101101010010;
assign LUT_3[35501] = 32'b00000000000000001010011000101111;
assign LUT_3[35502] = 32'b00000000000000000101110100110110;
assign LUT_3[35503] = 32'b00000000000000001100100000010011;
assign LUT_3[35504] = 32'b00000000000000000100011001011001;
assign LUT_3[35505] = 32'b00000000000000001011000100110110;
assign LUT_3[35506] = 32'b00000000000000000110100000111101;
assign LUT_3[35507] = 32'b00000000000000001101001100011010;
assign LUT_3[35508] = 32'b00000000000000000001100111001111;
assign LUT_3[35509] = 32'b00000000000000001000010010101100;
assign LUT_3[35510] = 32'b00000000000000000011101110110011;
assign LUT_3[35511] = 32'b00000000000000001010011010010000;
assign LUT_3[35512] = 32'b00000000000000001001110010011111;
assign LUT_3[35513] = 32'b00000000000000010000011101111100;
assign LUT_3[35514] = 32'b00000000000000001011111010000011;
assign LUT_3[35515] = 32'b00000000000000010010100101100000;
assign LUT_3[35516] = 32'b00000000000000000111000000010101;
assign LUT_3[35517] = 32'b00000000000000001101101011110010;
assign LUT_3[35518] = 32'b00000000000000001001000111111001;
assign LUT_3[35519] = 32'b00000000000000001111110011010110;
assign LUT_3[35520] = 32'b11111111111111111111110000100001;
assign LUT_3[35521] = 32'b00000000000000000110011011111110;
assign LUT_3[35522] = 32'b00000000000000000001111000000101;
assign LUT_3[35523] = 32'b00000000000000001000100011100010;
assign LUT_3[35524] = 32'b11111111111111111100111110010111;
assign LUT_3[35525] = 32'b00000000000000000011101001110100;
assign LUT_3[35526] = 32'b11111111111111111111000101111011;
assign LUT_3[35527] = 32'b00000000000000000101110001011000;
assign LUT_3[35528] = 32'b00000000000000000101001001100111;
assign LUT_3[35529] = 32'b00000000000000001011110101000100;
assign LUT_3[35530] = 32'b00000000000000000111010001001011;
assign LUT_3[35531] = 32'b00000000000000001101111100101000;
assign LUT_3[35532] = 32'b00000000000000000010010111011101;
assign LUT_3[35533] = 32'b00000000000000001001000010111010;
assign LUT_3[35534] = 32'b00000000000000000100011111000001;
assign LUT_3[35535] = 32'b00000000000000001011001010011110;
assign LUT_3[35536] = 32'b00000000000000000011000011100100;
assign LUT_3[35537] = 32'b00000000000000001001101111000001;
assign LUT_3[35538] = 32'b00000000000000000101001011001000;
assign LUT_3[35539] = 32'b00000000000000001011110110100101;
assign LUT_3[35540] = 32'b00000000000000000000010001011010;
assign LUT_3[35541] = 32'b00000000000000000110111100110111;
assign LUT_3[35542] = 32'b00000000000000000010011000111110;
assign LUT_3[35543] = 32'b00000000000000001001000100011011;
assign LUT_3[35544] = 32'b00000000000000001000011100101010;
assign LUT_3[35545] = 32'b00000000000000001111001000000111;
assign LUT_3[35546] = 32'b00000000000000001010100100001110;
assign LUT_3[35547] = 32'b00000000000000010001001111101011;
assign LUT_3[35548] = 32'b00000000000000000101101010100000;
assign LUT_3[35549] = 32'b00000000000000001100010101111101;
assign LUT_3[35550] = 32'b00000000000000000111110010000100;
assign LUT_3[35551] = 32'b00000000000000001110011101100001;
assign LUT_3[35552] = 32'b00000000000000000000111111000001;
assign LUT_3[35553] = 32'b00000000000000000111101010011110;
assign LUT_3[35554] = 32'b00000000000000000011000110100101;
assign LUT_3[35555] = 32'b00000000000000001001110010000010;
assign LUT_3[35556] = 32'b11111111111111111110001100110111;
assign LUT_3[35557] = 32'b00000000000000000100111000010100;
assign LUT_3[35558] = 32'b00000000000000000000010100011011;
assign LUT_3[35559] = 32'b00000000000000000110111111111000;
assign LUT_3[35560] = 32'b00000000000000000110011000000111;
assign LUT_3[35561] = 32'b00000000000000001101000011100100;
assign LUT_3[35562] = 32'b00000000000000001000011111101011;
assign LUT_3[35563] = 32'b00000000000000001111001011001000;
assign LUT_3[35564] = 32'b00000000000000000011100101111101;
assign LUT_3[35565] = 32'b00000000000000001010010001011010;
assign LUT_3[35566] = 32'b00000000000000000101101101100001;
assign LUT_3[35567] = 32'b00000000000000001100011000111110;
assign LUT_3[35568] = 32'b00000000000000000100010010000100;
assign LUT_3[35569] = 32'b00000000000000001010111101100001;
assign LUT_3[35570] = 32'b00000000000000000110011001101000;
assign LUT_3[35571] = 32'b00000000000000001101000101000101;
assign LUT_3[35572] = 32'b00000000000000000001011111111010;
assign LUT_3[35573] = 32'b00000000000000001000001011010111;
assign LUT_3[35574] = 32'b00000000000000000011100111011110;
assign LUT_3[35575] = 32'b00000000000000001010010010111011;
assign LUT_3[35576] = 32'b00000000000000001001101011001010;
assign LUT_3[35577] = 32'b00000000000000010000010110100111;
assign LUT_3[35578] = 32'b00000000000000001011110010101110;
assign LUT_3[35579] = 32'b00000000000000010010011110001011;
assign LUT_3[35580] = 32'b00000000000000000110111001000000;
assign LUT_3[35581] = 32'b00000000000000001101100100011101;
assign LUT_3[35582] = 32'b00000000000000001001000000100100;
assign LUT_3[35583] = 32'b00000000000000001111101100000001;
assign LUT_3[35584] = 32'b11111111111111111001111100011001;
assign LUT_3[35585] = 32'b00000000000000000000100111110110;
assign LUT_3[35586] = 32'b11111111111111111100000011111101;
assign LUT_3[35587] = 32'b00000000000000000010101111011010;
assign LUT_3[35588] = 32'b11111111111111110111001010001111;
assign LUT_3[35589] = 32'b11111111111111111101110101101100;
assign LUT_3[35590] = 32'b11111111111111111001010001110011;
assign LUT_3[35591] = 32'b11111111111111111111111101010000;
assign LUT_3[35592] = 32'b11111111111111111111010101011111;
assign LUT_3[35593] = 32'b00000000000000000110000000111100;
assign LUT_3[35594] = 32'b00000000000000000001011101000011;
assign LUT_3[35595] = 32'b00000000000000001000001000100000;
assign LUT_3[35596] = 32'b11111111111111111100100011010101;
assign LUT_3[35597] = 32'b00000000000000000011001110110010;
assign LUT_3[35598] = 32'b11111111111111111110101010111001;
assign LUT_3[35599] = 32'b00000000000000000101010110010110;
assign LUT_3[35600] = 32'b11111111111111111101001111011100;
assign LUT_3[35601] = 32'b00000000000000000011111010111001;
assign LUT_3[35602] = 32'b11111111111111111111010111000000;
assign LUT_3[35603] = 32'b00000000000000000110000010011101;
assign LUT_3[35604] = 32'b11111111111111111010011101010010;
assign LUT_3[35605] = 32'b00000000000000000001001000101111;
assign LUT_3[35606] = 32'b11111111111111111100100100110110;
assign LUT_3[35607] = 32'b00000000000000000011010000010011;
assign LUT_3[35608] = 32'b00000000000000000010101000100010;
assign LUT_3[35609] = 32'b00000000000000001001010011111111;
assign LUT_3[35610] = 32'b00000000000000000100110000000110;
assign LUT_3[35611] = 32'b00000000000000001011011011100011;
assign LUT_3[35612] = 32'b11111111111111111111110110011000;
assign LUT_3[35613] = 32'b00000000000000000110100001110101;
assign LUT_3[35614] = 32'b00000000000000000001111101111100;
assign LUT_3[35615] = 32'b00000000000000001000101001011001;
assign LUT_3[35616] = 32'b11111111111111111011001010111001;
assign LUT_3[35617] = 32'b00000000000000000001110110010110;
assign LUT_3[35618] = 32'b11111111111111111101010010011101;
assign LUT_3[35619] = 32'b00000000000000000011111101111010;
assign LUT_3[35620] = 32'b11111111111111111000011000101111;
assign LUT_3[35621] = 32'b11111111111111111111000100001100;
assign LUT_3[35622] = 32'b11111111111111111010100000010011;
assign LUT_3[35623] = 32'b00000000000000000001001011110000;
assign LUT_3[35624] = 32'b00000000000000000000100011111111;
assign LUT_3[35625] = 32'b00000000000000000111001111011100;
assign LUT_3[35626] = 32'b00000000000000000010101011100011;
assign LUT_3[35627] = 32'b00000000000000001001010111000000;
assign LUT_3[35628] = 32'b11111111111111111101110001110101;
assign LUT_3[35629] = 32'b00000000000000000100011101010010;
assign LUT_3[35630] = 32'b11111111111111111111111001011001;
assign LUT_3[35631] = 32'b00000000000000000110100100110110;
assign LUT_3[35632] = 32'b11111111111111111110011101111100;
assign LUT_3[35633] = 32'b00000000000000000101001001011001;
assign LUT_3[35634] = 32'b00000000000000000000100101100000;
assign LUT_3[35635] = 32'b00000000000000000111010000111101;
assign LUT_3[35636] = 32'b11111111111111111011101011110010;
assign LUT_3[35637] = 32'b00000000000000000010010111001111;
assign LUT_3[35638] = 32'b11111111111111111101110011010110;
assign LUT_3[35639] = 32'b00000000000000000100011110110011;
assign LUT_3[35640] = 32'b00000000000000000011110111000010;
assign LUT_3[35641] = 32'b00000000000000001010100010011111;
assign LUT_3[35642] = 32'b00000000000000000101111110100110;
assign LUT_3[35643] = 32'b00000000000000001100101010000011;
assign LUT_3[35644] = 32'b00000000000000000001000100111000;
assign LUT_3[35645] = 32'b00000000000000000111110000010101;
assign LUT_3[35646] = 32'b00000000000000000011001100011100;
assign LUT_3[35647] = 32'b00000000000000001001110111111001;
assign LUT_3[35648] = 32'b11111111111111111001110101000100;
assign LUT_3[35649] = 32'b00000000000000000000100000100001;
assign LUT_3[35650] = 32'b11111111111111111011111100101000;
assign LUT_3[35651] = 32'b00000000000000000010101000000101;
assign LUT_3[35652] = 32'b11111111111111110111000010111010;
assign LUT_3[35653] = 32'b11111111111111111101101110010111;
assign LUT_3[35654] = 32'b11111111111111111001001010011110;
assign LUT_3[35655] = 32'b11111111111111111111110101111011;
assign LUT_3[35656] = 32'b11111111111111111111001110001010;
assign LUT_3[35657] = 32'b00000000000000000101111001100111;
assign LUT_3[35658] = 32'b00000000000000000001010101101110;
assign LUT_3[35659] = 32'b00000000000000001000000001001011;
assign LUT_3[35660] = 32'b11111111111111111100011100000000;
assign LUT_3[35661] = 32'b00000000000000000011000111011101;
assign LUT_3[35662] = 32'b11111111111111111110100011100100;
assign LUT_3[35663] = 32'b00000000000000000101001111000001;
assign LUT_3[35664] = 32'b11111111111111111101001000000111;
assign LUT_3[35665] = 32'b00000000000000000011110011100100;
assign LUT_3[35666] = 32'b11111111111111111111001111101011;
assign LUT_3[35667] = 32'b00000000000000000101111011001000;
assign LUT_3[35668] = 32'b11111111111111111010010101111101;
assign LUT_3[35669] = 32'b00000000000000000001000001011010;
assign LUT_3[35670] = 32'b11111111111111111100011101100001;
assign LUT_3[35671] = 32'b00000000000000000011001000111110;
assign LUT_3[35672] = 32'b00000000000000000010100001001101;
assign LUT_3[35673] = 32'b00000000000000001001001100101010;
assign LUT_3[35674] = 32'b00000000000000000100101000110001;
assign LUT_3[35675] = 32'b00000000000000001011010100001110;
assign LUT_3[35676] = 32'b11111111111111111111101111000011;
assign LUT_3[35677] = 32'b00000000000000000110011010100000;
assign LUT_3[35678] = 32'b00000000000000000001110110100111;
assign LUT_3[35679] = 32'b00000000000000001000100010000100;
assign LUT_3[35680] = 32'b11111111111111111011000011100100;
assign LUT_3[35681] = 32'b00000000000000000001101111000001;
assign LUT_3[35682] = 32'b11111111111111111101001011001000;
assign LUT_3[35683] = 32'b00000000000000000011110110100101;
assign LUT_3[35684] = 32'b11111111111111111000010001011010;
assign LUT_3[35685] = 32'b11111111111111111110111100110111;
assign LUT_3[35686] = 32'b11111111111111111010011000111110;
assign LUT_3[35687] = 32'b00000000000000000001000100011011;
assign LUT_3[35688] = 32'b00000000000000000000011100101010;
assign LUT_3[35689] = 32'b00000000000000000111001000000111;
assign LUT_3[35690] = 32'b00000000000000000010100100001110;
assign LUT_3[35691] = 32'b00000000000000001001001111101011;
assign LUT_3[35692] = 32'b11111111111111111101101010100000;
assign LUT_3[35693] = 32'b00000000000000000100010101111101;
assign LUT_3[35694] = 32'b11111111111111111111110010000100;
assign LUT_3[35695] = 32'b00000000000000000110011101100001;
assign LUT_3[35696] = 32'b11111111111111111110010110100111;
assign LUT_3[35697] = 32'b00000000000000000101000010000100;
assign LUT_3[35698] = 32'b00000000000000000000011110001011;
assign LUT_3[35699] = 32'b00000000000000000111001001101000;
assign LUT_3[35700] = 32'b11111111111111111011100100011101;
assign LUT_3[35701] = 32'b00000000000000000010001111111010;
assign LUT_3[35702] = 32'b11111111111111111101101100000001;
assign LUT_3[35703] = 32'b00000000000000000100010111011110;
assign LUT_3[35704] = 32'b00000000000000000011101111101101;
assign LUT_3[35705] = 32'b00000000000000001010011011001010;
assign LUT_3[35706] = 32'b00000000000000000101110111010001;
assign LUT_3[35707] = 32'b00000000000000001100100010101110;
assign LUT_3[35708] = 32'b00000000000000000000111101100011;
assign LUT_3[35709] = 32'b00000000000000000111101001000000;
assign LUT_3[35710] = 32'b00000000000000000011000101000111;
assign LUT_3[35711] = 32'b00000000000000001001110000100100;
assign LUT_3[35712] = 32'b11111111111111111100000111010111;
assign LUT_3[35713] = 32'b00000000000000000010110010110100;
assign LUT_3[35714] = 32'b11111111111111111110001110111011;
assign LUT_3[35715] = 32'b00000000000000000100111010011000;
assign LUT_3[35716] = 32'b11111111111111111001010101001101;
assign LUT_3[35717] = 32'b00000000000000000000000000101010;
assign LUT_3[35718] = 32'b11111111111111111011011100110001;
assign LUT_3[35719] = 32'b00000000000000000010001000001110;
assign LUT_3[35720] = 32'b00000000000000000001100000011101;
assign LUT_3[35721] = 32'b00000000000000001000001011111010;
assign LUT_3[35722] = 32'b00000000000000000011101000000001;
assign LUT_3[35723] = 32'b00000000000000001010010011011110;
assign LUT_3[35724] = 32'b11111111111111111110101110010011;
assign LUT_3[35725] = 32'b00000000000000000101011001110000;
assign LUT_3[35726] = 32'b00000000000000000000110101110111;
assign LUT_3[35727] = 32'b00000000000000000111100001010100;
assign LUT_3[35728] = 32'b11111111111111111111011010011010;
assign LUT_3[35729] = 32'b00000000000000000110000101110111;
assign LUT_3[35730] = 32'b00000000000000000001100001111110;
assign LUT_3[35731] = 32'b00000000000000001000001101011011;
assign LUT_3[35732] = 32'b11111111111111111100101000010000;
assign LUT_3[35733] = 32'b00000000000000000011010011101101;
assign LUT_3[35734] = 32'b11111111111111111110101111110100;
assign LUT_3[35735] = 32'b00000000000000000101011011010001;
assign LUT_3[35736] = 32'b00000000000000000100110011100000;
assign LUT_3[35737] = 32'b00000000000000001011011110111101;
assign LUT_3[35738] = 32'b00000000000000000110111011000100;
assign LUT_3[35739] = 32'b00000000000000001101100110100001;
assign LUT_3[35740] = 32'b00000000000000000010000001010110;
assign LUT_3[35741] = 32'b00000000000000001000101100110011;
assign LUT_3[35742] = 32'b00000000000000000100001000111010;
assign LUT_3[35743] = 32'b00000000000000001010110100010111;
assign LUT_3[35744] = 32'b11111111111111111101010101110111;
assign LUT_3[35745] = 32'b00000000000000000100000001010100;
assign LUT_3[35746] = 32'b11111111111111111111011101011011;
assign LUT_3[35747] = 32'b00000000000000000110001000111000;
assign LUT_3[35748] = 32'b11111111111111111010100011101101;
assign LUT_3[35749] = 32'b00000000000000000001001111001010;
assign LUT_3[35750] = 32'b11111111111111111100101011010001;
assign LUT_3[35751] = 32'b00000000000000000011010110101110;
assign LUT_3[35752] = 32'b00000000000000000010101110111101;
assign LUT_3[35753] = 32'b00000000000000001001011010011010;
assign LUT_3[35754] = 32'b00000000000000000100110110100001;
assign LUT_3[35755] = 32'b00000000000000001011100001111110;
assign LUT_3[35756] = 32'b11111111111111111111111100110011;
assign LUT_3[35757] = 32'b00000000000000000110101000010000;
assign LUT_3[35758] = 32'b00000000000000000010000100010111;
assign LUT_3[35759] = 32'b00000000000000001000101111110100;
assign LUT_3[35760] = 32'b00000000000000000000101000111010;
assign LUT_3[35761] = 32'b00000000000000000111010100010111;
assign LUT_3[35762] = 32'b00000000000000000010110000011110;
assign LUT_3[35763] = 32'b00000000000000001001011011111011;
assign LUT_3[35764] = 32'b11111111111111111101110110110000;
assign LUT_3[35765] = 32'b00000000000000000100100010001101;
assign LUT_3[35766] = 32'b11111111111111111111111110010100;
assign LUT_3[35767] = 32'b00000000000000000110101001110001;
assign LUT_3[35768] = 32'b00000000000000000110000010000000;
assign LUT_3[35769] = 32'b00000000000000001100101101011101;
assign LUT_3[35770] = 32'b00000000000000001000001001100100;
assign LUT_3[35771] = 32'b00000000000000001110110101000001;
assign LUT_3[35772] = 32'b00000000000000000011001111110110;
assign LUT_3[35773] = 32'b00000000000000001001111011010011;
assign LUT_3[35774] = 32'b00000000000000000101010111011010;
assign LUT_3[35775] = 32'b00000000000000001100000010110111;
assign LUT_3[35776] = 32'b11111111111111111100000000000010;
assign LUT_3[35777] = 32'b00000000000000000010101011011111;
assign LUT_3[35778] = 32'b11111111111111111110000111100110;
assign LUT_3[35779] = 32'b00000000000000000100110011000011;
assign LUT_3[35780] = 32'b11111111111111111001001101111000;
assign LUT_3[35781] = 32'b11111111111111111111111001010101;
assign LUT_3[35782] = 32'b11111111111111111011010101011100;
assign LUT_3[35783] = 32'b00000000000000000010000000111001;
assign LUT_3[35784] = 32'b00000000000000000001011001001000;
assign LUT_3[35785] = 32'b00000000000000001000000100100101;
assign LUT_3[35786] = 32'b00000000000000000011100000101100;
assign LUT_3[35787] = 32'b00000000000000001010001100001001;
assign LUT_3[35788] = 32'b11111111111111111110100110111110;
assign LUT_3[35789] = 32'b00000000000000000101010010011011;
assign LUT_3[35790] = 32'b00000000000000000000101110100010;
assign LUT_3[35791] = 32'b00000000000000000111011001111111;
assign LUT_3[35792] = 32'b11111111111111111111010011000101;
assign LUT_3[35793] = 32'b00000000000000000101111110100010;
assign LUT_3[35794] = 32'b00000000000000000001011010101001;
assign LUT_3[35795] = 32'b00000000000000001000000110000110;
assign LUT_3[35796] = 32'b11111111111111111100100000111011;
assign LUT_3[35797] = 32'b00000000000000000011001100011000;
assign LUT_3[35798] = 32'b11111111111111111110101000011111;
assign LUT_3[35799] = 32'b00000000000000000101010011111100;
assign LUT_3[35800] = 32'b00000000000000000100101100001011;
assign LUT_3[35801] = 32'b00000000000000001011010111101000;
assign LUT_3[35802] = 32'b00000000000000000110110011101111;
assign LUT_3[35803] = 32'b00000000000000001101011111001100;
assign LUT_3[35804] = 32'b00000000000000000001111010000001;
assign LUT_3[35805] = 32'b00000000000000001000100101011110;
assign LUT_3[35806] = 32'b00000000000000000100000001100101;
assign LUT_3[35807] = 32'b00000000000000001010101101000010;
assign LUT_3[35808] = 32'b11111111111111111101001110100010;
assign LUT_3[35809] = 32'b00000000000000000011111001111111;
assign LUT_3[35810] = 32'b11111111111111111111010110000110;
assign LUT_3[35811] = 32'b00000000000000000110000001100011;
assign LUT_3[35812] = 32'b11111111111111111010011100011000;
assign LUT_3[35813] = 32'b00000000000000000001000111110101;
assign LUT_3[35814] = 32'b11111111111111111100100011111100;
assign LUT_3[35815] = 32'b00000000000000000011001111011001;
assign LUT_3[35816] = 32'b00000000000000000010100111101000;
assign LUT_3[35817] = 32'b00000000000000001001010011000101;
assign LUT_3[35818] = 32'b00000000000000000100101111001100;
assign LUT_3[35819] = 32'b00000000000000001011011010101001;
assign LUT_3[35820] = 32'b11111111111111111111110101011110;
assign LUT_3[35821] = 32'b00000000000000000110100000111011;
assign LUT_3[35822] = 32'b00000000000000000001111101000010;
assign LUT_3[35823] = 32'b00000000000000001000101000011111;
assign LUT_3[35824] = 32'b00000000000000000000100001100101;
assign LUT_3[35825] = 32'b00000000000000000111001101000010;
assign LUT_3[35826] = 32'b00000000000000000010101001001001;
assign LUT_3[35827] = 32'b00000000000000001001010100100110;
assign LUT_3[35828] = 32'b11111111111111111101101111011011;
assign LUT_3[35829] = 32'b00000000000000000100011010111000;
assign LUT_3[35830] = 32'b11111111111111111111110110111111;
assign LUT_3[35831] = 32'b00000000000000000110100010011100;
assign LUT_3[35832] = 32'b00000000000000000101111010101011;
assign LUT_3[35833] = 32'b00000000000000001100100110001000;
assign LUT_3[35834] = 32'b00000000000000001000000010001111;
assign LUT_3[35835] = 32'b00000000000000001110101101101100;
assign LUT_3[35836] = 32'b00000000000000000011001000100001;
assign LUT_3[35837] = 32'b00000000000000001001110011111110;
assign LUT_3[35838] = 32'b00000000000000000101010000000101;
assign LUT_3[35839] = 32'b00000000000000001011111011100010;
assign LUT_3[35840] = 32'b00000000000000000000111100101001;
assign LUT_3[35841] = 32'b00000000000000000111101000000110;
assign LUT_3[35842] = 32'b00000000000000000011000100001101;
assign LUT_3[35843] = 32'b00000000000000001001101111101010;
assign LUT_3[35844] = 32'b11111111111111111110001010011111;
assign LUT_3[35845] = 32'b00000000000000000100110101111100;
assign LUT_3[35846] = 32'b00000000000000000000010010000011;
assign LUT_3[35847] = 32'b00000000000000000110111101100000;
assign LUT_3[35848] = 32'b00000000000000000110010101101111;
assign LUT_3[35849] = 32'b00000000000000001101000001001100;
assign LUT_3[35850] = 32'b00000000000000001000011101010011;
assign LUT_3[35851] = 32'b00000000000000001111001000110000;
assign LUT_3[35852] = 32'b00000000000000000011100011100101;
assign LUT_3[35853] = 32'b00000000000000001010001111000010;
assign LUT_3[35854] = 32'b00000000000000000101101011001001;
assign LUT_3[35855] = 32'b00000000000000001100010110100110;
assign LUT_3[35856] = 32'b00000000000000000100001111101100;
assign LUT_3[35857] = 32'b00000000000000001010111011001001;
assign LUT_3[35858] = 32'b00000000000000000110010111010000;
assign LUT_3[35859] = 32'b00000000000000001101000010101101;
assign LUT_3[35860] = 32'b00000000000000000001011101100010;
assign LUT_3[35861] = 32'b00000000000000001000001000111111;
assign LUT_3[35862] = 32'b00000000000000000011100101000110;
assign LUT_3[35863] = 32'b00000000000000001010010000100011;
assign LUT_3[35864] = 32'b00000000000000001001101000110010;
assign LUT_3[35865] = 32'b00000000000000010000010100001111;
assign LUT_3[35866] = 32'b00000000000000001011110000010110;
assign LUT_3[35867] = 32'b00000000000000010010011011110011;
assign LUT_3[35868] = 32'b00000000000000000110110110101000;
assign LUT_3[35869] = 32'b00000000000000001101100010000101;
assign LUT_3[35870] = 32'b00000000000000001000111110001100;
assign LUT_3[35871] = 32'b00000000000000001111101001101001;
assign LUT_3[35872] = 32'b00000000000000000010001011001001;
assign LUT_3[35873] = 32'b00000000000000001000110110100110;
assign LUT_3[35874] = 32'b00000000000000000100010010101101;
assign LUT_3[35875] = 32'b00000000000000001010111110001010;
assign LUT_3[35876] = 32'b11111111111111111111011000111111;
assign LUT_3[35877] = 32'b00000000000000000110000100011100;
assign LUT_3[35878] = 32'b00000000000000000001100000100011;
assign LUT_3[35879] = 32'b00000000000000001000001100000000;
assign LUT_3[35880] = 32'b00000000000000000111100100001111;
assign LUT_3[35881] = 32'b00000000000000001110001111101100;
assign LUT_3[35882] = 32'b00000000000000001001101011110011;
assign LUT_3[35883] = 32'b00000000000000010000010111010000;
assign LUT_3[35884] = 32'b00000000000000000100110010000101;
assign LUT_3[35885] = 32'b00000000000000001011011101100010;
assign LUT_3[35886] = 32'b00000000000000000110111001101001;
assign LUT_3[35887] = 32'b00000000000000001101100101000110;
assign LUT_3[35888] = 32'b00000000000000000101011110001100;
assign LUT_3[35889] = 32'b00000000000000001100001001101001;
assign LUT_3[35890] = 32'b00000000000000000111100101110000;
assign LUT_3[35891] = 32'b00000000000000001110010001001101;
assign LUT_3[35892] = 32'b00000000000000000010101100000010;
assign LUT_3[35893] = 32'b00000000000000001001010111011111;
assign LUT_3[35894] = 32'b00000000000000000100110011100110;
assign LUT_3[35895] = 32'b00000000000000001011011111000011;
assign LUT_3[35896] = 32'b00000000000000001010110111010010;
assign LUT_3[35897] = 32'b00000000000000010001100010101111;
assign LUT_3[35898] = 32'b00000000000000001100111110110110;
assign LUT_3[35899] = 32'b00000000000000010011101010010011;
assign LUT_3[35900] = 32'b00000000000000001000000101001000;
assign LUT_3[35901] = 32'b00000000000000001110110000100101;
assign LUT_3[35902] = 32'b00000000000000001010001100101100;
assign LUT_3[35903] = 32'b00000000000000010000111000001001;
assign LUT_3[35904] = 32'b00000000000000000000110101010100;
assign LUT_3[35905] = 32'b00000000000000000111100000110001;
assign LUT_3[35906] = 32'b00000000000000000010111100111000;
assign LUT_3[35907] = 32'b00000000000000001001101000010101;
assign LUT_3[35908] = 32'b11111111111111111110000011001010;
assign LUT_3[35909] = 32'b00000000000000000100101110100111;
assign LUT_3[35910] = 32'b00000000000000000000001010101110;
assign LUT_3[35911] = 32'b00000000000000000110110110001011;
assign LUT_3[35912] = 32'b00000000000000000110001110011010;
assign LUT_3[35913] = 32'b00000000000000001100111001110111;
assign LUT_3[35914] = 32'b00000000000000001000010101111110;
assign LUT_3[35915] = 32'b00000000000000001111000001011011;
assign LUT_3[35916] = 32'b00000000000000000011011100010000;
assign LUT_3[35917] = 32'b00000000000000001010000111101101;
assign LUT_3[35918] = 32'b00000000000000000101100011110100;
assign LUT_3[35919] = 32'b00000000000000001100001111010001;
assign LUT_3[35920] = 32'b00000000000000000100001000010111;
assign LUT_3[35921] = 32'b00000000000000001010110011110100;
assign LUT_3[35922] = 32'b00000000000000000110001111111011;
assign LUT_3[35923] = 32'b00000000000000001100111011011000;
assign LUT_3[35924] = 32'b00000000000000000001010110001101;
assign LUT_3[35925] = 32'b00000000000000001000000001101010;
assign LUT_3[35926] = 32'b00000000000000000011011101110001;
assign LUT_3[35927] = 32'b00000000000000001010001001001110;
assign LUT_3[35928] = 32'b00000000000000001001100001011101;
assign LUT_3[35929] = 32'b00000000000000010000001100111010;
assign LUT_3[35930] = 32'b00000000000000001011101001000001;
assign LUT_3[35931] = 32'b00000000000000010010010100011110;
assign LUT_3[35932] = 32'b00000000000000000110101111010011;
assign LUT_3[35933] = 32'b00000000000000001101011010110000;
assign LUT_3[35934] = 32'b00000000000000001000110110110111;
assign LUT_3[35935] = 32'b00000000000000001111100010010100;
assign LUT_3[35936] = 32'b00000000000000000010000011110100;
assign LUT_3[35937] = 32'b00000000000000001000101111010001;
assign LUT_3[35938] = 32'b00000000000000000100001011011000;
assign LUT_3[35939] = 32'b00000000000000001010110110110101;
assign LUT_3[35940] = 32'b11111111111111111111010001101010;
assign LUT_3[35941] = 32'b00000000000000000101111101000111;
assign LUT_3[35942] = 32'b00000000000000000001011001001110;
assign LUT_3[35943] = 32'b00000000000000001000000100101011;
assign LUT_3[35944] = 32'b00000000000000000111011100111010;
assign LUT_3[35945] = 32'b00000000000000001110001000010111;
assign LUT_3[35946] = 32'b00000000000000001001100100011110;
assign LUT_3[35947] = 32'b00000000000000010000001111111011;
assign LUT_3[35948] = 32'b00000000000000000100101010110000;
assign LUT_3[35949] = 32'b00000000000000001011010110001101;
assign LUT_3[35950] = 32'b00000000000000000110110010010100;
assign LUT_3[35951] = 32'b00000000000000001101011101110001;
assign LUT_3[35952] = 32'b00000000000000000101010110110111;
assign LUT_3[35953] = 32'b00000000000000001100000010010100;
assign LUT_3[35954] = 32'b00000000000000000111011110011011;
assign LUT_3[35955] = 32'b00000000000000001110001001111000;
assign LUT_3[35956] = 32'b00000000000000000010100100101101;
assign LUT_3[35957] = 32'b00000000000000001001010000001010;
assign LUT_3[35958] = 32'b00000000000000000100101100010001;
assign LUT_3[35959] = 32'b00000000000000001011010111101110;
assign LUT_3[35960] = 32'b00000000000000001010101111111101;
assign LUT_3[35961] = 32'b00000000000000010001011011011010;
assign LUT_3[35962] = 32'b00000000000000001100110111100001;
assign LUT_3[35963] = 32'b00000000000000010011100010111110;
assign LUT_3[35964] = 32'b00000000000000000111111101110011;
assign LUT_3[35965] = 32'b00000000000000001110101001010000;
assign LUT_3[35966] = 32'b00000000000000001010000101010111;
assign LUT_3[35967] = 32'b00000000000000010000110000110100;
assign LUT_3[35968] = 32'b00000000000000000011000111100111;
assign LUT_3[35969] = 32'b00000000000000001001110011000100;
assign LUT_3[35970] = 32'b00000000000000000101001111001011;
assign LUT_3[35971] = 32'b00000000000000001011111010101000;
assign LUT_3[35972] = 32'b00000000000000000000010101011101;
assign LUT_3[35973] = 32'b00000000000000000111000000111010;
assign LUT_3[35974] = 32'b00000000000000000010011101000001;
assign LUT_3[35975] = 32'b00000000000000001001001000011110;
assign LUT_3[35976] = 32'b00000000000000001000100000101101;
assign LUT_3[35977] = 32'b00000000000000001111001100001010;
assign LUT_3[35978] = 32'b00000000000000001010101000010001;
assign LUT_3[35979] = 32'b00000000000000010001010011101110;
assign LUT_3[35980] = 32'b00000000000000000101101110100011;
assign LUT_3[35981] = 32'b00000000000000001100011010000000;
assign LUT_3[35982] = 32'b00000000000000000111110110000111;
assign LUT_3[35983] = 32'b00000000000000001110100001100100;
assign LUT_3[35984] = 32'b00000000000000000110011010101010;
assign LUT_3[35985] = 32'b00000000000000001101000110000111;
assign LUT_3[35986] = 32'b00000000000000001000100010001110;
assign LUT_3[35987] = 32'b00000000000000001111001101101011;
assign LUT_3[35988] = 32'b00000000000000000011101000100000;
assign LUT_3[35989] = 32'b00000000000000001010010011111101;
assign LUT_3[35990] = 32'b00000000000000000101110000000100;
assign LUT_3[35991] = 32'b00000000000000001100011011100001;
assign LUT_3[35992] = 32'b00000000000000001011110011110000;
assign LUT_3[35993] = 32'b00000000000000010010011111001101;
assign LUT_3[35994] = 32'b00000000000000001101111011010100;
assign LUT_3[35995] = 32'b00000000000000010100100110110001;
assign LUT_3[35996] = 32'b00000000000000001001000001100110;
assign LUT_3[35997] = 32'b00000000000000001111101101000011;
assign LUT_3[35998] = 32'b00000000000000001011001001001010;
assign LUT_3[35999] = 32'b00000000000000010001110100100111;
assign LUT_3[36000] = 32'b00000000000000000100010110000111;
assign LUT_3[36001] = 32'b00000000000000001011000001100100;
assign LUT_3[36002] = 32'b00000000000000000110011101101011;
assign LUT_3[36003] = 32'b00000000000000001101001001001000;
assign LUT_3[36004] = 32'b00000000000000000001100011111101;
assign LUT_3[36005] = 32'b00000000000000001000001111011010;
assign LUT_3[36006] = 32'b00000000000000000011101011100001;
assign LUT_3[36007] = 32'b00000000000000001010010110111110;
assign LUT_3[36008] = 32'b00000000000000001001101111001101;
assign LUT_3[36009] = 32'b00000000000000010000011010101010;
assign LUT_3[36010] = 32'b00000000000000001011110110110001;
assign LUT_3[36011] = 32'b00000000000000010010100010001110;
assign LUT_3[36012] = 32'b00000000000000000110111101000011;
assign LUT_3[36013] = 32'b00000000000000001101101000100000;
assign LUT_3[36014] = 32'b00000000000000001001000100100111;
assign LUT_3[36015] = 32'b00000000000000001111110000000100;
assign LUT_3[36016] = 32'b00000000000000000111101001001010;
assign LUT_3[36017] = 32'b00000000000000001110010100100111;
assign LUT_3[36018] = 32'b00000000000000001001110000101110;
assign LUT_3[36019] = 32'b00000000000000010000011100001011;
assign LUT_3[36020] = 32'b00000000000000000100110111000000;
assign LUT_3[36021] = 32'b00000000000000001011100010011101;
assign LUT_3[36022] = 32'b00000000000000000110111110100100;
assign LUT_3[36023] = 32'b00000000000000001101101010000001;
assign LUT_3[36024] = 32'b00000000000000001101000010010000;
assign LUT_3[36025] = 32'b00000000000000010011101101101101;
assign LUT_3[36026] = 32'b00000000000000001111001001110100;
assign LUT_3[36027] = 32'b00000000000000010101110101010001;
assign LUT_3[36028] = 32'b00000000000000001010010000000110;
assign LUT_3[36029] = 32'b00000000000000010000111011100011;
assign LUT_3[36030] = 32'b00000000000000001100010111101010;
assign LUT_3[36031] = 32'b00000000000000010011000011000111;
assign LUT_3[36032] = 32'b00000000000000000011000000010010;
assign LUT_3[36033] = 32'b00000000000000001001101011101111;
assign LUT_3[36034] = 32'b00000000000000000101000111110110;
assign LUT_3[36035] = 32'b00000000000000001011110011010011;
assign LUT_3[36036] = 32'b00000000000000000000001110001000;
assign LUT_3[36037] = 32'b00000000000000000110111001100101;
assign LUT_3[36038] = 32'b00000000000000000010010101101100;
assign LUT_3[36039] = 32'b00000000000000001001000001001001;
assign LUT_3[36040] = 32'b00000000000000001000011001011000;
assign LUT_3[36041] = 32'b00000000000000001111000100110101;
assign LUT_3[36042] = 32'b00000000000000001010100000111100;
assign LUT_3[36043] = 32'b00000000000000010001001100011001;
assign LUT_3[36044] = 32'b00000000000000000101100111001110;
assign LUT_3[36045] = 32'b00000000000000001100010010101011;
assign LUT_3[36046] = 32'b00000000000000000111101110110010;
assign LUT_3[36047] = 32'b00000000000000001110011010001111;
assign LUT_3[36048] = 32'b00000000000000000110010011010101;
assign LUT_3[36049] = 32'b00000000000000001100111110110010;
assign LUT_3[36050] = 32'b00000000000000001000011010111001;
assign LUT_3[36051] = 32'b00000000000000001111000110010110;
assign LUT_3[36052] = 32'b00000000000000000011100001001011;
assign LUT_3[36053] = 32'b00000000000000001010001100101000;
assign LUT_3[36054] = 32'b00000000000000000101101000101111;
assign LUT_3[36055] = 32'b00000000000000001100010100001100;
assign LUT_3[36056] = 32'b00000000000000001011101100011011;
assign LUT_3[36057] = 32'b00000000000000010010010111111000;
assign LUT_3[36058] = 32'b00000000000000001101110011111111;
assign LUT_3[36059] = 32'b00000000000000010100011111011100;
assign LUT_3[36060] = 32'b00000000000000001000111010010001;
assign LUT_3[36061] = 32'b00000000000000001111100101101110;
assign LUT_3[36062] = 32'b00000000000000001011000001110101;
assign LUT_3[36063] = 32'b00000000000000010001101101010010;
assign LUT_3[36064] = 32'b00000000000000000100001110110010;
assign LUT_3[36065] = 32'b00000000000000001010111010001111;
assign LUT_3[36066] = 32'b00000000000000000110010110010110;
assign LUT_3[36067] = 32'b00000000000000001101000001110011;
assign LUT_3[36068] = 32'b00000000000000000001011100101000;
assign LUT_3[36069] = 32'b00000000000000001000001000000101;
assign LUT_3[36070] = 32'b00000000000000000011100100001100;
assign LUT_3[36071] = 32'b00000000000000001010001111101001;
assign LUT_3[36072] = 32'b00000000000000001001100111111000;
assign LUT_3[36073] = 32'b00000000000000010000010011010101;
assign LUT_3[36074] = 32'b00000000000000001011101111011100;
assign LUT_3[36075] = 32'b00000000000000010010011010111001;
assign LUT_3[36076] = 32'b00000000000000000110110101101110;
assign LUT_3[36077] = 32'b00000000000000001101100001001011;
assign LUT_3[36078] = 32'b00000000000000001000111101010010;
assign LUT_3[36079] = 32'b00000000000000001111101000101111;
assign LUT_3[36080] = 32'b00000000000000000111100001110101;
assign LUT_3[36081] = 32'b00000000000000001110001101010010;
assign LUT_3[36082] = 32'b00000000000000001001101001011001;
assign LUT_3[36083] = 32'b00000000000000010000010100110110;
assign LUT_3[36084] = 32'b00000000000000000100101111101011;
assign LUT_3[36085] = 32'b00000000000000001011011011001000;
assign LUT_3[36086] = 32'b00000000000000000110110111001111;
assign LUT_3[36087] = 32'b00000000000000001101100010101100;
assign LUT_3[36088] = 32'b00000000000000001100111010111011;
assign LUT_3[36089] = 32'b00000000000000010011100110011000;
assign LUT_3[36090] = 32'b00000000000000001111000010011111;
assign LUT_3[36091] = 32'b00000000000000010101101101111100;
assign LUT_3[36092] = 32'b00000000000000001010001000110001;
assign LUT_3[36093] = 32'b00000000000000010000110100001110;
assign LUT_3[36094] = 32'b00000000000000001100010000010101;
assign LUT_3[36095] = 32'b00000000000000010010111011110010;
assign LUT_3[36096] = 32'b11111111111111111101001100001010;
assign LUT_3[36097] = 32'b00000000000000000011110111100111;
assign LUT_3[36098] = 32'b11111111111111111111010011101110;
assign LUT_3[36099] = 32'b00000000000000000101111111001011;
assign LUT_3[36100] = 32'b11111111111111111010011010000000;
assign LUT_3[36101] = 32'b00000000000000000001000101011101;
assign LUT_3[36102] = 32'b11111111111111111100100001100100;
assign LUT_3[36103] = 32'b00000000000000000011001101000001;
assign LUT_3[36104] = 32'b00000000000000000010100101010000;
assign LUT_3[36105] = 32'b00000000000000001001010000101101;
assign LUT_3[36106] = 32'b00000000000000000100101100110100;
assign LUT_3[36107] = 32'b00000000000000001011011000010001;
assign LUT_3[36108] = 32'b11111111111111111111110011000110;
assign LUT_3[36109] = 32'b00000000000000000110011110100011;
assign LUT_3[36110] = 32'b00000000000000000001111010101010;
assign LUT_3[36111] = 32'b00000000000000001000100110000111;
assign LUT_3[36112] = 32'b00000000000000000000011111001101;
assign LUT_3[36113] = 32'b00000000000000000111001010101010;
assign LUT_3[36114] = 32'b00000000000000000010100110110001;
assign LUT_3[36115] = 32'b00000000000000001001010010001110;
assign LUT_3[36116] = 32'b11111111111111111101101101000011;
assign LUT_3[36117] = 32'b00000000000000000100011000100000;
assign LUT_3[36118] = 32'b11111111111111111111110100100111;
assign LUT_3[36119] = 32'b00000000000000000110100000000100;
assign LUT_3[36120] = 32'b00000000000000000101111000010011;
assign LUT_3[36121] = 32'b00000000000000001100100011110000;
assign LUT_3[36122] = 32'b00000000000000000111111111110111;
assign LUT_3[36123] = 32'b00000000000000001110101011010100;
assign LUT_3[36124] = 32'b00000000000000000011000110001001;
assign LUT_3[36125] = 32'b00000000000000001001110001100110;
assign LUT_3[36126] = 32'b00000000000000000101001101101101;
assign LUT_3[36127] = 32'b00000000000000001011111001001010;
assign LUT_3[36128] = 32'b11111111111111111110011010101010;
assign LUT_3[36129] = 32'b00000000000000000101000110000111;
assign LUT_3[36130] = 32'b00000000000000000000100010001110;
assign LUT_3[36131] = 32'b00000000000000000111001101101011;
assign LUT_3[36132] = 32'b11111111111111111011101000100000;
assign LUT_3[36133] = 32'b00000000000000000010010011111101;
assign LUT_3[36134] = 32'b11111111111111111101110000000100;
assign LUT_3[36135] = 32'b00000000000000000100011011100001;
assign LUT_3[36136] = 32'b00000000000000000011110011110000;
assign LUT_3[36137] = 32'b00000000000000001010011111001101;
assign LUT_3[36138] = 32'b00000000000000000101111011010100;
assign LUT_3[36139] = 32'b00000000000000001100100110110001;
assign LUT_3[36140] = 32'b00000000000000000001000001100110;
assign LUT_3[36141] = 32'b00000000000000000111101101000011;
assign LUT_3[36142] = 32'b00000000000000000011001001001010;
assign LUT_3[36143] = 32'b00000000000000001001110100100111;
assign LUT_3[36144] = 32'b00000000000000000001101101101101;
assign LUT_3[36145] = 32'b00000000000000001000011001001010;
assign LUT_3[36146] = 32'b00000000000000000011110101010001;
assign LUT_3[36147] = 32'b00000000000000001010100000101110;
assign LUT_3[36148] = 32'b11111111111111111110111011100011;
assign LUT_3[36149] = 32'b00000000000000000101100111000000;
assign LUT_3[36150] = 32'b00000000000000000001000011000111;
assign LUT_3[36151] = 32'b00000000000000000111101110100100;
assign LUT_3[36152] = 32'b00000000000000000111000110110011;
assign LUT_3[36153] = 32'b00000000000000001101110010010000;
assign LUT_3[36154] = 32'b00000000000000001001001110010111;
assign LUT_3[36155] = 32'b00000000000000001111111001110100;
assign LUT_3[36156] = 32'b00000000000000000100010100101001;
assign LUT_3[36157] = 32'b00000000000000001011000000000110;
assign LUT_3[36158] = 32'b00000000000000000110011100001101;
assign LUT_3[36159] = 32'b00000000000000001101000111101010;
assign LUT_3[36160] = 32'b11111111111111111101000100110101;
assign LUT_3[36161] = 32'b00000000000000000011110000010010;
assign LUT_3[36162] = 32'b11111111111111111111001100011001;
assign LUT_3[36163] = 32'b00000000000000000101110111110110;
assign LUT_3[36164] = 32'b11111111111111111010010010101011;
assign LUT_3[36165] = 32'b00000000000000000000111110001000;
assign LUT_3[36166] = 32'b11111111111111111100011010001111;
assign LUT_3[36167] = 32'b00000000000000000011000101101100;
assign LUT_3[36168] = 32'b00000000000000000010011101111011;
assign LUT_3[36169] = 32'b00000000000000001001001001011000;
assign LUT_3[36170] = 32'b00000000000000000100100101011111;
assign LUT_3[36171] = 32'b00000000000000001011010000111100;
assign LUT_3[36172] = 32'b11111111111111111111101011110001;
assign LUT_3[36173] = 32'b00000000000000000110010111001110;
assign LUT_3[36174] = 32'b00000000000000000001110011010101;
assign LUT_3[36175] = 32'b00000000000000001000011110110010;
assign LUT_3[36176] = 32'b00000000000000000000010111111000;
assign LUT_3[36177] = 32'b00000000000000000111000011010101;
assign LUT_3[36178] = 32'b00000000000000000010011111011100;
assign LUT_3[36179] = 32'b00000000000000001001001010111001;
assign LUT_3[36180] = 32'b11111111111111111101100101101110;
assign LUT_3[36181] = 32'b00000000000000000100010001001011;
assign LUT_3[36182] = 32'b11111111111111111111101101010010;
assign LUT_3[36183] = 32'b00000000000000000110011000101111;
assign LUT_3[36184] = 32'b00000000000000000101110000111110;
assign LUT_3[36185] = 32'b00000000000000001100011100011011;
assign LUT_3[36186] = 32'b00000000000000000111111000100010;
assign LUT_3[36187] = 32'b00000000000000001110100011111111;
assign LUT_3[36188] = 32'b00000000000000000010111110110100;
assign LUT_3[36189] = 32'b00000000000000001001101010010001;
assign LUT_3[36190] = 32'b00000000000000000101000110011000;
assign LUT_3[36191] = 32'b00000000000000001011110001110101;
assign LUT_3[36192] = 32'b11111111111111111110010011010101;
assign LUT_3[36193] = 32'b00000000000000000100111110110010;
assign LUT_3[36194] = 32'b00000000000000000000011010111001;
assign LUT_3[36195] = 32'b00000000000000000111000110010110;
assign LUT_3[36196] = 32'b11111111111111111011100001001011;
assign LUT_3[36197] = 32'b00000000000000000010001100101000;
assign LUT_3[36198] = 32'b11111111111111111101101000101111;
assign LUT_3[36199] = 32'b00000000000000000100010100001100;
assign LUT_3[36200] = 32'b00000000000000000011101100011011;
assign LUT_3[36201] = 32'b00000000000000001010010111111000;
assign LUT_3[36202] = 32'b00000000000000000101110011111111;
assign LUT_3[36203] = 32'b00000000000000001100011111011100;
assign LUT_3[36204] = 32'b00000000000000000000111010010001;
assign LUT_3[36205] = 32'b00000000000000000111100101101110;
assign LUT_3[36206] = 32'b00000000000000000011000001110101;
assign LUT_3[36207] = 32'b00000000000000001001101101010010;
assign LUT_3[36208] = 32'b00000000000000000001100110011000;
assign LUT_3[36209] = 32'b00000000000000001000010001110101;
assign LUT_3[36210] = 32'b00000000000000000011101101111100;
assign LUT_3[36211] = 32'b00000000000000001010011001011001;
assign LUT_3[36212] = 32'b11111111111111111110110100001110;
assign LUT_3[36213] = 32'b00000000000000000101011111101011;
assign LUT_3[36214] = 32'b00000000000000000000111011110010;
assign LUT_3[36215] = 32'b00000000000000000111100111001111;
assign LUT_3[36216] = 32'b00000000000000000110111111011110;
assign LUT_3[36217] = 32'b00000000000000001101101010111011;
assign LUT_3[36218] = 32'b00000000000000001001000111000010;
assign LUT_3[36219] = 32'b00000000000000001111110010011111;
assign LUT_3[36220] = 32'b00000000000000000100001101010100;
assign LUT_3[36221] = 32'b00000000000000001010111000110001;
assign LUT_3[36222] = 32'b00000000000000000110010100111000;
assign LUT_3[36223] = 32'b00000000000000001101000000010101;
assign LUT_3[36224] = 32'b11111111111111111111010111001000;
assign LUT_3[36225] = 32'b00000000000000000110000010100101;
assign LUT_3[36226] = 32'b00000000000000000001011110101100;
assign LUT_3[36227] = 32'b00000000000000001000001010001001;
assign LUT_3[36228] = 32'b11111111111111111100100100111110;
assign LUT_3[36229] = 32'b00000000000000000011010000011011;
assign LUT_3[36230] = 32'b11111111111111111110101100100010;
assign LUT_3[36231] = 32'b00000000000000000101010111111111;
assign LUT_3[36232] = 32'b00000000000000000100110000001110;
assign LUT_3[36233] = 32'b00000000000000001011011011101011;
assign LUT_3[36234] = 32'b00000000000000000110110111110010;
assign LUT_3[36235] = 32'b00000000000000001101100011001111;
assign LUT_3[36236] = 32'b00000000000000000001111110000100;
assign LUT_3[36237] = 32'b00000000000000001000101001100001;
assign LUT_3[36238] = 32'b00000000000000000100000101101000;
assign LUT_3[36239] = 32'b00000000000000001010110001000101;
assign LUT_3[36240] = 32'b00000000000000000010101010001011;
assign LUT_3[36241] = 32'b00000000000000001001010101101000;
assign LUT_3[36242] = 32'b00000000000000000100110001101111;
assign LUT_3[36243] = 32'b00000000000000001011011101001100;
assign LUT_3[36244] = 32'b11111111111111111111111000000001;
assign LUT_3[36245] = 32'b00000000000000000110100011011110;
assign LUT_3[36246] = 32'b00000000000000000001111111100101;
assign LUT_3[36247] = 32'b00000000000000001000101011000010;
assign LUT_3[36248] = 32'b00000000000000001000000011010001;
assign LUT_3[36249] = 32'b00000000000000001110101110101110;
assign LUT_3[36250] = 32'b00000000000000001010001010110101;
assign LUT_3[36251] = 32'b00000000000000010000110110010010;
assign LUT_3[36252] = 32'b00000000000000000101010001000111;
assign LUT_3[36253] = 32'b00000000000000001011111100100100;
assign LUT_3[36254] = 32'b00000000000000000111011000101011;
assign LUT_3[36255] = 32'b00000000000000001110000100001000;
assign LUT_3[36256] = 32'b00000000000000000000100101101000;
assign LUT_3[36257] = 32'b00000000000000000111010001000101;
assign LUT_3[36258] = 32'b00000000000000000010101101001100;
assign LUT_3[36259] = 32'b00000000000000001001011000101001;
assign LUT_3[36260] = 32'b11111111111111111101110011011110;
assign LUT_3[36261] = 32'b00000000000000000100011110111011;
assign LUT_3[36262] = 32'b11111111111111111111111011000010;
assign LUT_3[36263] = 32'b00000000000000000110100110011111;
assign LUT_3[36264] = 32'b00000000000000000101111110101110;
assign LUT_3[36265] = 32'b00000000000000001100101010001011;
assign LUT_3[36266] = 32'b00000000000000001000000110010010;
assign LUT_3[36267] = 32'b00000000000000001110110001101111;
assign LUT_3[36268] = 32'b00000000000000000011001100100100;
assign LUT_3[36269] = 32'b00000000000000001001111000000001;
assign LUT_3[36270] = 32'b00000000000000000101010100001000;
assign LUT_3[36271] = 32'b00000000000000001011111111100101;
assign LUT_3[36272] = 32'b00000000000000000011111000101011;
assign LUT_3[36273] = 32'b00000000000000001010100100001000;
assign LUT_3[36274] = 32'b00000000000000000110000000001111;
assign LUT_3[36275] = 32'b00000000000000001100101011101100;
assign LUT_3[36276] = 32'b00000000000000000001000110100001;
assign LUT_3[36277] = 32'b00000000000000000111110001111110;
assign LUT_3[36278] = 32'b00000000000000000011001110000101;
assign LUT_3[36279] = 32'b00000000000000001001111001100010;
assign LUT_3[36280] = 32'b00000000000000001001010001110001;
assign LUT_3[36281] = 32'b00000000000000001111111101001110;
assign LUT_3[36282] = 32'b00000000000000001011011001010101;
assign LUT_3[36283] = 32'b00000000000000010010000100110010;
assign LUT_3[36284] = 32'b00000000000000000110011111100111;
assign LUT_3[36285] = 32'b00000000000000001101001011000100;
assign LUT_3[36286] = 32'b00000000000000001000100111001011;
assign LUT_3[36287] = 32'b00000000000000001111010010101000;
assign LUT_3[36288] = 32'b11111111111111111111001111110011;
assign LUT_3[36289] = 32'b00000000000000000101111011010000;
assign LUT_3[36290] = 32'b00000000000000000001010111010111;
assign LUT_3[36291] = 32'b00000000000000001000000010110100;
assign LUT_3[36292] = 32'b11111111111111111100011101101001;
assign LUT_3[36293] = 32'b00000000000000000011001001000110;
assign LUT_3[36294] = 32'b11111111111111111110100101001101;
assign LUT_3[36295] = 32'b00000000000000000101010000101010;
assign LUT_3[36296] = 32'b00000000000000000100101000111001;
assign LUT_3[36297] = 32'b00000000000000001011010100010110;
assign LUT_3[36298] = 32'b00000000000000000110110000011101;
assign LUT_3[36299] = 32'b00000000000000001101011011111010;
assign LUT_3[36300] = 32'b00000000000000000001110110101111;
assign LUT_3[36301] = 32'b00000000000000001000100010001100;
assign LUT_3[36302] = 32'b00000000000000000011111110010011;
assign LUT_3[36303] = 32'b00000000000000001010101001110000;
assign LUT_3[36304] = 32'b00000000000000000010100010110110;
assign LUT_3[36305] = 32'b00000000000000001001001110010011;
assign LUT_3[36306] = 32'b00000000000000000100101010011010;
assign LUT_3[36307] = 32'b00000000000000001011010101110111;
assign LUT_3[36308] = 32'b11111111111111111111110000101100;
assign LUT_3[36309] = 32'b00000000000000000110011100001001;
assign LUT_3[36310] = 32'b00000000000000000001111000010000;
assign LUT_3[36311] = 32'b00000000000000001000100011101101;
assign LUT_3[36312] = 32'b00000000000000000111111011111100;
assign LUT_3[36313] = 32'b00000000000000001110100111011001;
assign LUT_3[36314] = 32'b00000000000000001010000011100000;
assign LUT_3[36315] = 32'b00000000000000010000101110111101;
assign LUT_3[36316] = 32'b00000000000000000101001001110010;
assign LUT_3[36317] = 32'b00000000000000001011110101001111;
assign LUT_3[36318] = 32'b00000000000000000111010001010110;
assign LUT_3[36319] = 32'b00000000000000001101111100110011;
assign LUT_3[36320] = 32'b00000000000000000000011110010011;
assign LUT_3[36321] = 32'b00000000000000000111001001110000;
assign LUT_3[36322] = 32'b00000000000000000010100101110111;
assign LUT_3[36323] = 32'b00000000000000001001010001010100;
assign LUT_3[36324] = 32'b11111111111111111101101100001001;
assign LUT_3[36325] = 32'b00000000000000000100010111100110;
assign LUT_3[36326] = 32'b11111111111111111111110011101101;
assign LUT_3[36327] = 32'b00000000000000000110011111001010;
assign LUT_3[36328] = 32'b00000000000000000101110111011001;
assign LUT_3[36329] = 32'b00000000000000001100100010110110;
assign LUT_3[36330] = 32'b00000000000000000111111110111101;
assign LUT_3[36331] = 32'b00000000000000001110101010011010;
assign LUT_3[36332] = 32'b00000000000000000011000101001111;
assign LUT_3[36333] = 32'b00000000000000001001110000101100;
assign LUT_3[36334] = 32'b00000000000000000101001100110011;
assign LUT_3[36335] = 32'b00000000000000001011111000010000;
assign LUT_3[36336] = 32'b00000000000000000011110001010110;
assign LUT_3[36337] = 32'b00000000000000001010011100110011;
assign LUT_3[36338] = 32'b00000000000000000101111000111010;
assign LUT_3[36339] = 32'b00000000000000001100100100010111;
assign LUT_3[36340] = 32'b00000000000000000000111111001100;
assign LUT_3[36341] = 32'b00000000000000000111101010101001;
assign LUT_3[36342] = 32'b00000000000000000011000110110000;
assign LUT_3[36343] = 32'b00000000000000001001110010001101;
assign LUT_3[36344] = 32'b00000000000000001001001010011100;
assign LUT_3[36345] = 32'b00000000000000001111110101111001;
assign LUT_3[36346] = 32'b00000000000000001011010010000000;
assign LUT_3[36347] = 32'b00000000000000010001111101011101;
assign LUT_3[36348] = 32'b00000000000000000110011000010010;
assign LUT_3[36349] = 32'b00000000000000001101000011101111;
assign LUT_3[36350] = 32'b00000000000000001000011111110110;
assign LUT_3[36351] = 32'b00000000000000001111001011010011;
assign LUT_3[36352] = 32'b00000000000000000100010001110101;
assign LUT_3[36353] = 32'b00000000000000001010111101010010;
assign LUT_3[36354] = 32'b00000000000000000110011001011001;
assign LUT_3[36355] = 32'b00000000000000001101000100110110;
assign LUT_3[36356] = 32'b00000000000000000001011111101011;
assign LUT_3[36357] = 32'b00000000000000001000001011001000;
assign LUT_3[36358] = 32'b00000000000000000011100111001111;
assign LUT_3[36359] = 32'b00000000000000001010010010101100;
assign LUT_3[36360] = 32'b00000000000000001001101010111011;
assign LUT_3[36361] = 32'b00000000000000010000010110011000;
assign LUT_3[36362] = 32'b00000000000000001011110010011111;
assign LUT_3[36363] = 32'b00000000000000010010011101111100;
assign LUT_3[36364] = 32'b00000000000000000110111000110001;
assign LUT_3[36365] = 32'b00000000000000001101100100001110;
assign LUT_3[36366] = 32'b00000000000000001001000000010101;
assign LUT_3[36367] = 32'b00000000000000001111101011110010;
assign LUT_3[36368] = 32'b00000000000000000111100100111000;
assign LUT_3[36369] = 32'b00000000000000001110010000010101;
assign LUT_3[36370] = 32'b00000000000000001001101100011100;
assign LUT_3[36371] = 32'b00000000000000010000010111111001;
assign LUT_3[36372] = 32'b00000000000000000100110010101110;
assign LUT_3[36373] = 32'b00000000000000001011011110001011;
assign LUT_3[36374] = 32'b00000000000000000110111010010010;
assign LUT_3[36375] = 32'b00000000000000001101100101101111;
assign LUT_3[36376] = 32'b00000000000000001100111101111110;
assign LUT_3[36377] = 32'b00000000000000010011101001011011;
assign LUT_3[36378] = 32'b00000000000000001111000101100010;
assign LUT_3[36379] = 32'b00000000000000010101110000111111;
assign LUT_3[36380] = 32'b00000000000000001010001011110100;
assign LUT_3[36381] = 32'b00000000000000010000110111010001;
assign LUT_3[36382] = 32'b00000000000000001100010011011000;
assign LUT_3[36383] = 32'b00000000000000010010111110110101;
assign LUT_3[36384] = 32'b00000000000000000101100000010101;
assign LUT_3[36385] = 32'b00000000000000001100001011110010;
assign LUT_3[36386] = 32'b00000000000000000111100111111001;
assign LUT_3[36387] = 32'b00000000000000001110010011010110;
assign LUT_3[36388] = 32'b00000000000000000010101110001011;
assign LUT_3[36389] = 32'b00000000000000001001011001101000;
assign LUT_3[36390] = 32'b00000000000000000100110101101111;
assign LUT_3[36391] = 32'b00000000000000001011100001001100;
assign LUT_3[36392] = 32'b00000000000000001010111001011011;
assign LUT_3[36393] = 32'b00000000000000010001100100111000;
assign LUT_3[36394] = 32'b00000000000000001101000000111111;
assign LUT_3[36395] = 32'b00000000000000010011101100011100;
assign LUT_3[36396] = 32'b00000000000000001000000111010001;
assign LUT_3[36397] = 32'b00000000000000001110110010101110;
assign LUT_3[36398] = 32'b00000000000000001010001110110101;
assign LUT_3[36399] = 32'b00000000000000010000111010010010;
assign LUT_3[36400] = 32'b00000000000000001000110011011000;
assign LUT_3[36401] = 32'b00000000000000001111011110110101;
assign LUT_3[36402] = 32'b00000000000000001010111010111100;
assign LUT_3[36403] = 32'b00000000000000010001100110011001;
assign LUT_3[36404] = 32'b00000000000000000110000001001110;
assign LUT_3[36405] = 32'b00000000000000001100101100101011;
assign LUT_3[36406] = 32'b00000000000000001000001000110010;
assign LUT_3[36407] = 32'b00000000000000001110110100001111;
assign LUT_3[36408] = 32'b00000000000000001110001100011110;
assign LUT_3[36409] = 32'b00000000000000010100110111111011;
assign LUT_3[36410] = 32'b00000000000000010000010100000010;
assign LUT_3[36411] = 32'b00000000000000010110111111011111;
assign LUT_3[36412] = 32'b00000000000000001011011010010100;
assign LUT_3[36413] = 32'b00000000000000010010000101110001;
assign LUT_3[36414] = 32'b00000000000000001101100001111000;
assign LUT_3[36415] = 32'b00000000000000010100001101010101;
assign LUT_3[36416] = 32'b00000000000000000100001010100000;
assign LUT_3[36417] = 32'b00000000000000001010110101111101;
assign LUT_3[36418] = 32'b00000000000000000110010010000100;
assign LUT_3[36419] = 32'b00000000000000001100111101100001;
assign LUT_3[36420] = 32'b00000000000000000001011000010110;
assign LUT_3[36421] = 32'b00000000000000001000000011110011;
assign LUT_3[36422] = 32'b00000000000000000011011111111010;
assign LUT_3[36423] = 32'b00000000000000001010001011010111;
assign LUT_3[36424] = 32'b00000000000000001001100011100110;
assign LUT_3[36425] = 32'b00000000000000010000001111000011;
assign LUT_3[36426] = 32'b00000000000000001011101011001010;
assign LUT_3[36427] = 32'b00000000000000010010010110100111;
assign LUT_3[36428] = 32'b00000000000000000110110001011100;
assign LUT_3[36429] = 32'b00000000000000001101011100111001;
assign LUT_3[36430] = 32'b00000000000000001000111001000000;
assign LUT_3[36431] = 32'b00000000000000001111100100011101;
assign LUT_3[36432] = 32'b00000000000000000111011101100011;
assign LUT_3[36433] = 32'b00000000000000001110001001000000;
assign LUT_3[36434] = 32'b00000000000000001001100101000111;
assign LUT_3[36435] = 32'b00000000000000010000010000100100;
assign LUT_3[36436] = 32'b00000000000000000100101011011001;
assign LUT_3[36437] = 32'b00000000000000001011010110110110;
assign LUT_3[36438] = 32'b00000000000000000110110010111101;
assign LUT_3[36439] = 32'b00000000000000001101011110011010;
assign LUT_3[36440] = 32'b00000000000000001100110110101001;
assign LUT_3[36441] = 32'b00000000000000010011100010000110;
assign LUT_3[36442] = 32'b00000000000000001110111110001101;
assign LUT_3[36443] = 32'b00000000000000010101101001101010;
assign LUT_3[36444] = 32'b00000000000000001010000100011111;
assign LUT_3[36445] = 32'b00000000000000010000101111111100;
assign LUT_3[36446] = 32'b00000000000000001100001100000011;
assign LUT_3[36447] = 32'b00000000000000010010110111100000;
assign LUT_3[36448] = 32'b00000000000000000101011001000000;
assign LUT_3[36449] = 32'b00000000000000001100000100011101;
assign LUT_3[36450] = 32'b00000000000000000111100000100100;
assign LUT_3[36451] = 32'b00000000000000001110001100000001;
assign LUT_3[36452] = 32'b00000000000000000010100110110110;
assign LUT_3[36453] = 32'b00000000000000001001010010010011;
assign LUT_3[36454] = 32'b00000000000000000100101110011010;
assign LUT_3[36455] = 32'b00000000000000001011011001110111;
assign LUT_3[36456] = 32'b00000000000000001010110010000110;
assign LUT_3[36457] = 32'b00000000000000010001011101100011;
assign LUT_3[36458] = 32'b00000000000000001100111001101010;
assign LUT_3[36459] = 32'b00000000000000010011100101000111;
assign LUT_3[36460] = 32'b00000000000000000111111111111100;
assign LUT_3[36461] = 32'b00000000000000001110101011011001;
assign LUT_3[36462] = 32'b00000000000000001010000111100000;
assign LUT_3[36463] = 32'b00000000000000010000110010111101;
assign LUT_3[36464] = 32'b00000000000000001000101100000011;
assign LUT_3[36465] = 32'b00000000000000001111010111100000;
assign LUT_3[36466] = 32'b00000000000000001010110011100111;
assign LUT_3[36467] = 32'b00000000000000010001011111000100;
assign LUT_3[36468] = 32'b00000000000000000101111001111001;
assign LUT_3[36469] = 32'b00000000000000001100100101010110;
assign LUT_3[36470] = 32'b00000000000000001000000001011101;
assign LUT_3[36471] = 32'b00000000000000001110101100111010;
assign LUT_3[36472] = 32'b00000000000000001110000101001001;
assign LUT_3[36473] = 32'b00000000000000010100110000100110;
assign LUT_3[36474] = 32'b00000000000000010000001100101101;
assign LUT_3[36475] = 32'b00000000000000010110111000001010;
assign LUT_3[36476] = 32'b00000000000000001011010010111111;
assign LUT_3[36477] = 32'b00000000000000010001111110011100;
assign LUT_3[36478] = 32'b00000000000000001101011010100011;
assign LUT_3[36479] = 32'b00000000000000010100000110000000;
assign LUT_3[36480] = 32'b00000000000000000110011100110011;
assign LUT_3[36481] = 32'b00000000000000001101001000010000;
assign LUT_3[36482] = 32'b00000000000000001000100100010111;
assign LUT_3[36483] = 32'b00000000000000001111001111110100;
assign LUT_3[36484] = 32'b00000000000000000011101010101001;
assign LUT_3[36485] = 32'b00000000000000001010010110000110;
assign LUT_3[36486] = 32'b00000000000000000101110010001101;
assign LUT_3[36487] = 32'b00000000000000001100011101101010;
assign LUT_3[36488] = 32'b00000000000000001011110101111001;
assign LUT_3[36489] = 32'b00000000000000010010100001010110;
assign LUT_3[36490] = 32'b00000000000000001101111101011101;
assign LUT_3[36491] = 32'b00000000000000010100101000111010;
assign LUT_3[36492] = 32'b00000000000000001001000011101111;
assign LUT_3[36493] = 32'b00000000000000001111101111001100;
assign LUT_3[36494] = 32'b00000000000000001011001011010011;
assign LUT_3[36495] = 32'b00000000000000010001110110110000;
assign LUT_3[36496] = 32'b00000000000000001001101111110110;
assign LUT_3[36497] = 32'b00000000000000010000011011010011;
assign LUT_3[36498] = 32'b00000000000000001011110111011010;
assign LUT_3[36499] = 32'b00000000000000010010100010110111;
assign LUT_3[36500] = 32'b00000000000000000110111101101100;
assign LUT_3[36501] = 32'b00000000000000001101101001001001;
assign LUT_3[36502] = 32'b00000000000000001001000101010000;
assign LUT_3[36503] = 32'b00000000000000001111110000101101;
assign LUT_3[36504] = 32'b00000000000000001111001000111100;
assign LUT_3[36505] = 32'b00000000000000010101110100011001;
assign LUT_3[36506] = 32'b00000000000000010001010000100000;
assign LUT_3[36507] = 32'b00000000000000010111111011111101;
assign LUT_3[36508] = 32'b00000000000000001100010110110010;
assign LUT_3[36509] = 32'b00000000000000010011000010001111;
assign LUT_3[36510] = 32'b00000000000000001110011110010110;
assign LUT_3[36511] = 32'b00000000000000010101001001110011;
assign LUT_3[36512] = 32'b00000000000000000111101011010011;
assign LUT_3[36513] = 32'b00000000000000001110010110110000;
assign LUT_3[36514] = 32'b00000000000000001001110010110111;
assign LUT_3[36515] = 32'b00000000000000010000011110010100;
assign LUT_3[36516] = 32'b00000000000000000100111001001001;
assign LUT_3[36517] = 32'b00000000000000001011100100100110;
assign LUT_3[36518] = 32'b00000000000000000111000000101101;
assign LUT_3[36519] = 32'b00000000000000001101101100001010;
assign LUT_3[36520] = 32'b00000000000000001101000100011001;
assign LUT_3[36521] = 32'b00000000000000010011101111110110;
assign LUT_3[36522] = 32'b00000000000000001111001011111101;
assign LUT_3[36523] = 32'b00000000000000010101110111011010;
assign LUT_3[36524] = 32'b00000000000000001010010010001111;
assign LUT_3[36525] = 32'b00000000000000010000111101101100;
assign LUT_3[36526] = 32'b00000000000000001100011001110011;
assign LUT_3[36527] = 32'b00000000000000010011000101010000;
assign LUT_3[36528] = 32'b00000000000000001010111110010110;
assign LUT_3[36529] = 32'b00000000000000010001101001110011;
assign LUT_3[36530] = 32'b00000000000000001101000101111010;
assign LUT_3[36531] = 32'b00000000000000010011110001010111;
assign LUT_3[36532] = 32'b00000000000000001000001100001100;
assign LUT_3[36533] = 32'b00000000000000001110110111101001;
assign LUT_3[36534] = 32'b00000000000000001010010011110000;
assign LUT_3[36535] = 32'b00000000000000010000111111001101;
assign LUT_3[36536] = 32'b00000000000000010000010111011100;
assign LUT_3[36537] = 32'b00000000000000010111000010111001;
assign LUT_3[36538] = 32'b00000000000000010010011111000000;
assign LUT_3[36539] = 32'b00000000000000011001001010011101;
assign LUT_3[36540] = 32'b00000000000000001101100101010010;
assign LUT_3[36541] = 32'b00000000000000010100010000101111;
assign LUT_3[36542] = 32'b00000000000000001111101100110110;
assign LUT_3[36543] = 32'b00000000000000010110011000010011;
assign LUT_3[36544] = 32'b00000000000000000110010101011110;
assign LUT_3[36545] = 32'b00000000000000001101000000111011;
assign LUT_3[36546] = 32'b00000000000000001000011101000010;
assign LUT_3[36547] = 32'b00000000000000001111001000011111;
assign LUT_3[36548] = 32'b00000000000000000011100011010100;
assign LUT_3[36549] = 32'b00000000000000001010001110110001;
assign LUT_3[36550] = 32'b00000000000000000101101010111000;
assign LUT_3[36551] = 32'b00000000000000001100010110010101;
assign LUT_3[36552] = 32'b00000000000000001011101110100100;
assign LUT_3[36553] = 32'b00000000000000010010011010000001;
assign LUT_3[36554] = 32'b00000000000000001101110110001000;
assign LUT_3[36555] = 32'b00000000000000010100100001100101;
assign LUT_3[36556] = 32'b00000000000000001000111100011010;
assign LUT_3[36557] = 32'b00000000000000001111100111110111;
assign LUT_3[36558] = 32'b00000000000000001011000011111110;
assign LUT_3[36559] = 32'b00000000000000010001101111011011;
assign LUT_3[36560] = 32'b00000000000000001001101000100001;
assign LUT_3[36561] = 32'b00000000000000010000010011111110;
assign LUT_3[36562] = 32'b00000000000000001011110000000101;
assign LUT_3[36563] = 32'b00000000000000010010011011100010;
assign LUT_3[36564] = 32'b00000000000000000110110110010111;
assign LUT_3[36565] = 32'b00000000000000001101100001110100;
assign LUT_3[36566] = 32'b00000000000000001000111101111011;
assign LUT_3[36567] = 32'b00000000000000001111101001011000;
assign LUT_3[36568] = 32'b00000000000000001111000001100111;
assign LUT_3[36569] = 32'b00000000000000010101101101000100;
assign LUT_3[36570] = 32'b00000000000000010001001001001011;
assign LUT_3[36571] = 32'b00000000000000010111110100101000;
assign LUT_3[36572] = 32'b00000000000000001100001111011101;
assign LUT_3[36573] = 32'b00000000000000010010111010111010;
assign LUT_3[36574] = 32'b00000000000000001110010111000001;
assign LUT_3[36575] = 32'b00000000000000010101000010011110;
assign LUT_3[36576] = 32'b00000000000000000111100011111110;
assign LUT_3[36577] = 32'b00000000000000001110001111011011;
assign LUT_3[36578] = 32'b00000000000000001001101011100010;
assign LUT_3[36579] = 32'b00000000000000010000010110111111;
assign LUT_3[36580] = 32'b00000000000000000100110001110100;
assign LUT_3[36581] = 32'b00000000000000001011011101010001;
assign LUT_3[36582] = 32'b00000000000000000110111001011000;
assign LUT_3[36583] = 32'b00000000000000001101100100110101;
assign LUT_3[36584] = 32'b00000000000000001100111101000100;
assign LUT_3[36585] = 32'b00000000000000010011101000100001;
assign LUT_3[36586] = 32'b00000000000000001111000100101000;
assign LUT_3[36587] = 32'b00000000000000010101110000000101;
assign LUT_3[36588] = 32'b00000000000000001010001010111010;
assign LUT_3[36589] = 32'b00000000000000010000110110010111;
assign LUT_3[36590] = 32'b00000000000000001100010010011110;
assign LUT_3[36591] = 32'b00000000000000010010111101111011;
assign LUT_3[36592] = 32'b00000000000000001010110111000001;
assign LUT_3[36593] = 32'b00000000000000010001100010011110;
assign LUT_3[36594] = 32'b00000000000000001100111110100101;
assign LUT_3[36595] = 32'b00000000000000010011101010000010;
assign LUT_3[36596] = 32'b00000000000000001000000100110111;
assign LUT_3[36597] = 32'b00000000000000001110110000010100;
assign LUT_3[36598] = 32'b00000000000000001010001100011011;
assign LUT_3[36599] = 32'b00000000000000010000110111111000;
assign LUT_3[36600] = 32'b00000000000000010000010000000111;
assign LUT_3[36601] = 32'b00000000000000010110111011100100;
assign LUT_3[36602] = 32'b00000000000000010010010111101011;
assign LUT_3[36603] = 32'b00000000000000011001000011001000;
assign LUT_3[36604] = 32'b00000000000000001101011101111101;
assign LUT_3[36605] = 32'b00000000000000010100001001011010;
assign LUT_3[36606] = 32'b00000000000000001111100101100001;
assign LUT_3[36607] = 32'b00000000000000010110010000111110;
assign LUT_3[36608] = 32'b00000000000000000000100001010110;
assign LUT_3[36609] = 32'b00000000000000000111001100110011;
assign LUT_3[36610] = 32'b00000000000000000010101000111010;
assign LUT_3[36611] = 32'b00000000000000001001010100010111;
assign LUT_3[36612] = 32'b11111111111111111101101111001100;
assign LUT_3[36613] = 32'b00000000000000000100011010101001;
assign LUT_3[36614] = 32'b11111111111111111111110110110000;
assign LUT_3[36615] = 32'b00000000000000000110100010001101;
assign LUT_3[36616] = 32'b00000000000000000101111010011100;
assign LUT_3[36617] = 32'b00000000000000001100100101111001;
assign LUT_3[36618] = 32'b00000000000000001000000010000000;
assign LUT_3[36619] = 32'b00000000000000001110101101011101;
assign LUT_3[36620] = 32'b00000000000000000011001000010010;
assign LUT_3[36621] = 32'b00000000000000001001110011101111;
assign LUT_3[36622] = 32'b00000000000000000101001111110110;
assign LUT_3[36623] = 32'b00000000000000001011111011010011;
assign LUT_3[36624] = 32'b00000000000000000011110100011001;
assign LUT_3[36625] = 32'b00000000000000001010011111110110;
assign LUT_3[36626] = 32'b00000000000000000101111011111101;
assign LUT_3[36627] = 32'b00000000000000001100100111011010;
assign LUT_3[36628] = 32'b00000000000000000001000010001111;
assign LUT_3[36629] = 32'b00000000000000000111101101101100;
assign LUT_3[36630] = 32'b00000000000000000011001001110011;
assign LUT_3[36631] = 32'b00000000000000001001110101010000;
assign LUT_3[36632] = 32'b00000000000000001001001101011111;
assign LUT_3[36633] = 32'b00000000000000001111111000111100;
assign LUT_3[36634] = 32'b00000000000000001011010101000011;
assign LUT_3[36635] = 32'b00000000000000010010000000100000;
assign LUT_3[36636] = 32'b00000000000000000110011011010101;
assign LUT_3[36637] = 32'b00000000000000001101000110110010;
assign LUT_3[36638] = 32'b00000000000000001000100010111001;
assign LUT_3[36639] = 32'b00000000000000001111001110010110;
assign LUT_3[36640] = 32'b00000000000000000001101111110110;
assign LUT_3[36641] = 32'b00000000000000001000011011010011;
assign LUT_3[36642] = 32'b00000000000000000011110111011010;
assign LUT_3[36643] = 32'b00000000000000001010100010110111;
assign LUT_3[36644] = 32'b11111111111111111110111101101100;
assign LUT_3[36645] = 32'b00000000000000000101101001001001;
assign LUT_3[36646] = 32'b00000000000000000001000101010000;
assign LUT_3[36647] = 32'b00000000000000000111110000101101;
assign LUT_3[36648] = 32'b00000000000000000111001000111100;
assign LUT_3[36649] = 32'b00000000000000001101110100011001;
assign LUT_3[36650] = 32'b00000000000000001001010000100000;
assign LUT_3[36651] = 32'b00000000000000001111111011111101;
assign LUT_3[36652] = 32'b00000000000000000100010110110010;
assign LUT_3[36653] = 32'b00000000000000001011000010001111;
assign LUT_3[36654] = 32'b00000000000000000110011110010110;
assign LUT_3[36655] = 32'b00000000000000001101001001110011;
assign LUT_3[36656] = 32'b00000000000000000101000010111001;
assign LUT_3[36657] = 32'b00000000000000001011101110010110;
assign LUT_3[36658] = 32'b00000000000000000111001010011101;
assign LUT_3[36659] = 32'b00000000000000001101110101111010;
assign LUT_3[36660] = 32'b00000000000000000010010000101111;
assign LUT_3[36661] = 32'b00000000000000001000111100001100;
assign LUT_3[36662] = 32'b00000000000000000100011000010011;
assign LUT_3[36663] = 32'b00000000000000001011000011110000;
assign LUT_3[36664] = 32'b00000000000000001010011011111111;
assign LUT_3[36665] = 32'b00000000000000010001000111011100;
assign LUT_3[36666] = 32'b00000000000000001100100011100011;
assign LUT_3[36667] = 32'b00000000000000010011001111000000;
assign LUT_3[36668] = 32'b00000000000000000111101001110101;
assign LUT_3[36669] = 32'b00000000000000001110010101010010;
assign LUT_3[36670] = 32'b00000000000000001001110001011001;
assign LUT_3[36671] = 32'b00000000000000010000011100110110;
assign LUT_3[36672] = 32'b00000000000000000000011010000001;
assign LUT_3[36673] = 32'b00000000000000000111000101011110;
assign LUT_3[36674] = 32'b00000000000000000010100001100101;
assign LUT_3[36675] = 32'b00000000000000001001001101000010;
assign LUT_3[36676] = 32'b11111111111111111101100111110111;
assign LUT_3[36677] = 32'b00000000000000000100010011010100;
assign LUT_3[36678] = 32'b11111111111111111111101111011011;
assign LUT_3[36679] = 32'b00000000000000000110011010111000;
assign LUT_3[36680] = 32'b00000000000000000101110011000111;
assign LUT_3[36681] = 32'b00000000000000001100011110100100;
assign LUT_3[36682] = 32'b00000000000000000111111010101011;
assign LUT_3[36683] = 32'b00000000000000001110100110001000;
assign LUT_3[36684] = 32'b00000000000000000011000000111101;
assign LUT_3[36685] = 32'b00000000000000001001101100011010;
assign LUT_3[36686] = 32'b00000000000000000101001000100001;
assign LUT_3[36687] = 32'b00000000000000001011110011111110;
assign LUT_3[36688] = 32'b00000000000000000011101101000100;
assign LUT_3[36689] = 32'b00000000000000001010011000100001;
assign LUT_3[36690] = 32'b00000000000000000101110100101000;
assign LUT_3[36691] = 32'b00000000000000001100100000000101;
assign LUT_3[36692] = 32'b00000000000000000000111010111010;
assign LUT_3[36693] = 32'b00000000000000000111100110010111;
assign LUT_3[36694] = 32'b00000000000000000011000010011110;
assign LUT_3[36695] = 32'b00000000000000001001101101111011;
assign LUT_3[36696] = 32'b00000000000000001001000110001010;
assign LUT_3[36697] = 32'b00000000000000001111110001100111;
assign LUT_3[36698] = 32'b00000000000000001011001101101110;
assign LUT_3[36699] = 32'b00000000000000010001111001001011;
assign LUT_3[36700] = 32'b00000000000000000110010100000000;
assign LUT_3[36701] = 32'b00000000000000001100111111011101;
assign LUT_3[36702] = 32'b00000000000000001000011011100100;
assign LUT_3[36703] = 32'b00000000000000001111000111000001;
assign LUT_3[36704] = 32'b00000000000000000001101000100001;
assign LUT_3[36705] = 32'b00000000000000001000010011111110;
assign LUT_3[36706] = 32'b00000000000000000011110000000101;
assign LUT_3[36707] = 32'b00000000000000001010011011100010;
assign LUT_3[36708] = 32'b11111111111111111110110110010111;
assign LUT_3[36709] = 32'b00000000000000000101100001110100;
assign LUT_3[36710] = 32'b00000000000000000000111101111011;
assign LUT_3[36711] = 32'b00000000000000000111101001011000;
assign LUT_3[36712] = 32'b00000000000000000111000001100111;
assign LUT_3[36713] = 32'b00000000000000001101101101000100;
assign LUT_3[36714] = 32'b00000000000000001001001001001011;
assign LUT_3[36715] = 32'b00000000000000001111110100101000;
assign LUT_3[36716] = 32'b00000000000000000100001111011101;
assign LUT_3[36717] = 32'b00000000000000001010111010111010;
assign LUT_3[36718] = 32'b00000000000000000110010111000001;
assign LUT_3[36719] = 32'b00000000000000001101000010011110;
assign LUT_3[36720] = 32'b00000000000000000100111011100100;
assign LUT_3[36721] = 32'b00000000000000001011100111000001;
assign LUT_3[36722] = 32'b00000000000000000111000011001000;
assign LUT_3[36723] = 32'b00000000000000001101101110100101;
assign LUT_3[36724] = 32'b00000000000000000010001001011010;
assign LUT_3[36725] = 32'b00000000000000001000110100110111;
assign LUT_3[36726] = 32'b00000000000000000100010000111110;
assign LUT_3[36727] = 32'b00000000000000001010111100011011;
assign LUT_3[36728] = 32'b00000000000000001010010100101010;
assign LUT_3[36729] = 32'b00000000000000010001000000000111;
assign LUT_3[36730] = 32'b00000000000000001100011100001110;
assign LUT_3[36731] = 32'b00000000000000010011000111101011;
assign LUT_3[36732] = 32'b00000000000000000111100010100000;
assign LUT_3[36733] = 32'b00000000000000001110001101111101;
assign LUT_3[36734] = 32'b00000000000000001001101010000100;
assign LUT_3[36735] = 32'b00000000000000010000010101100001;
assign LUT_3[36736] = 32'b00000000000000000010101100010100;
assign LUT_3[36737] = 32'b00000000000000001001010111110001;
assign LUT_3[36738] = 32'b00000000000000000100110011111000;
assign LUT_3[36739] = 32'b00000000000000001011011111010101;
assign LUT_3[36740] = 32'b11111111111111111111111010001010;
assign LUT_3[36741] = 32'b00000000000000000110100101100111;
assign LUT_3[36742] = 32'b00000000000000000010000001101110;
assign LUT_3[36743] = 32'b00000000000000001000101101001011;
assign LUT_3[36744] = 32'b00000000000000001000000101011010;
assign LUT_3[36745] = 32'b00000000000000001110110000110111;
assign LUT_3[36746] = 32'b00000000000000001010001100111110;
assign LUT_3[36747] = 32'b00000000000000010000111000011011;
assign LUT_3[36748] = 32'b00000000000000000101010011010000;
assign LUT_3[36749] = 32'b00000000000000001011111110101101;
assign LUT_3[36750] = 32'b00000000000000000111011010110100;
assign LUT_3[36751] = 32'b00000000000000001110000110010001;
assign LUT_3[36752] = 32'b00000000000000000101111111010111;
assign LUT_3[36753] = 32'b00000000000000001100101010110100;
assign LUT_3[36754] = 32'b00000000000000001000000110111011;
assign LUT_3[36755] = 32'b00000000000000001110110010011000;
assign LUT_3[36756] = 32'b00000000000000000011001101001101;
assign LUT_3[36757] = 32'b00000000000000001001111000101010;
assign LUT_3[36758] = 32'b00000000000000000101010100110001;
assign LUT_3[36759] = 32'b00000000000000001100000000001110;
assign LUT_3[36760] = 32'b00000000000000001011011000011101;
assign LUT_3[36761] = 32'b00000000000000010010000011111010;
assign LUT_3[36762] = 32'b00000000000000001101100000000001;
assign LUT_3[36763] = 32'b00000000000000010100001011011110;
assign LUT_3[36764] = 32'b00000000000000001000100110010011;
assign LUT_3[36765] = 32'b00000000000000001111010001110000;
assign LUT_3[36766] = 32'b00000000000000001010101101110111;
assign LUT_3[36767] = 32'b00000000000000010001011001010100;
assign LUT_3[36768] = 32'b00000000000000000011111010110100;
assign LUT_3[36769] = 32'b00000000000000001010100110010001;
assign LUT_3[36770] = 32'b00000000000000000110000010011000;
assign LUT_3[36771] = 32'b00000000000000001100101101110101;
assign LUT_3[36772] = 32'b00000000000000000001001000101010;
assign LUT_3[36773] = 32'b00000000000000000111110100000111;
assign LUT_3[36774] = 32'b00000000000000000011010000001110;
assign LUT_3[36775] = 32'b00000000000000001001111011101011;
assign LUT_3[36776] = 32'b00000000000000001001010011111010;
assign LUT_3[36777] = 32'b00000000000000001111111111010111;
assign LUT_3[36778] = 32'b00000000000000001011011011011110;
assign LUT_3[36779] = 32'b00000000000000010010000110111011;
assign LUT_3[36780] = 32'b00000000000000000110100001110000;
assign LUT_3[36781] = 32'b00000000000000001101001101001101;
assign LUT_3[36782] = 32'b00000000000000001000101001010100;
assign LUT_3[36783] = 32'b00000000000000001111010100110001;
assign LUT_3[36784] = 32'b00000000000000000111001101110111;
assign LUT_3[36785] = 32'b00000000000000001101111001010100;
assign LUT_3[36786] = 32'b00000000000000001001010101011011;
assign LUT_3[36787] = 32'b00000000000000010000000000111000;
assign LUT_3[36788] = 32'b00000000000000000100011011101101;
assign LUT_3[36789] = 32'b00000000000000001011000111001010;
assign LUT_3[36790] = 32'b00000000000000000110100011010001;
assign LUT_3[36791] = 32'b00000000000000001101001110101110;
assign LUT_3[36792] = 32'b00000000000000001100100110111101;
assign LUT_3[36793] = 32'b00000000000000010011010010011010;
assign LUT_3[36794] = 32'b00000000000000001110101110100001;
assign LUT_3[36795] = 32'b00000000000000010101011001111110;
assign LUT_3[36796] = 32'b00000000000000001001110100110011;
assign LUT_3[36797] = 32'b00000000000000010000100000010000;
assign LUT_3[36798] = 32'b00000000000000001011111100010111;
assign LUT_3[36799] = 32'b00000000000000010010100111110100;
assign LUT_3[36800] = 32'b00000000000000000010100100111111;
assign LUT_3[36801] = 32'b00000000000000001001010000011100;
assign LUT_3[36802] = 32'b00000000000000000100101100100011;
assign LUT_3[36803] = 32'b00000000000000001011011000000000;
assign LUT_3[36804] = 32'b11111111111111111111110010110101;
assign LUT_3[36805] = 32'b00000000000000000110011110010010;
assign LUT_3[36806] = 32'b00000000000000000001111010011001;
assign LUT_3[36807] = 32'b00000000000000001000100101110110;
assign LUT_3[36808] = 32'b00000000000000000111111110000101;
assign LUT_3[36809] = 32'b00000000000000001110101001100010;
assign LUT_3[36810] = 32'b00000000000000001010000101101001;
assign LUT_3[36811] = 32'b00000000000000010000110001000110;
assign LUT_3[36812] = 32'b00000000000000000101001011111011;
assign LUT_3[36813] = 32'b00000000000000001011110111011000;
assign LUT_3[36814] = 32'b00000000000000000111010011011111;
assign LUT_3[36815] = 32'b00000000000000001101111110111100;
assign LUT_3[36816] = 32'b00000000000000000101111000000010;
assign LUT_3[36817] = 32'b00000000000000001100100011011111;
assign LUT_3[36818] = 32'b00000000000000000111111111100110;
assign LUT_3[36819] = 32'b00000000000000001110101011000011;
assign LUT_3[36820] = 32'b00000000000000000011000101111000;
assign LUT_3[36821] = 32'b00000000000000001001110001010101;
assign LUT_3[36822] = 32'b00000000000000000101001101011100;
assign LUT_3[36823] = 32'b00000000000000001011111000111001;
assign LUT_3[36824] = 32'b00000000000000001011010001001000;
assign LUT_3[36825] = 32'b00000000000000010001111100100101;
assign LUT_3[36826] = 32'b00000000000000001101011000101100;
assign LUT_3[36827] = 32'b00000000000000010100000100001001;
assign LUT_3[36828] = 32'b00000000000000001000011110111110;
assign LUT_3[36829] = 32'b00000000000000001111001010011011;
assign LUT_3[36830] = 32'b00000000000000001010100110100010;
assign LUT_3[36831] = 32'b00000000000000010001010001111111;
assign LUT_3[36832] = 32'b00000000000000000011110011011111;
assign LUT_3[36833] = 32'b00000000000000001010011110111100;
assign LUT_3[36834] = 32'b00000000000000000101111011000011;
assign LUT_3[36835] = 32'b00000000000000001100100110100000;
assign LUT_3[36836] = 32'b00000000000000000001000001010101;
assign LUT_3[36837] = 32'b00000000000000000111101100110010;
assign LUT_3[36838] = 32'b00000000000000000011001000111001;
assign LUT_3[36839] = 32'b00000000000000001001110100010110;
assign LUT_3[36840] = 32'b00000000000000001001001100100101;
assign LUT_3[36841] = 32'b00000000000000001111111000000010;
assign LUT_3[36842] = 32'b00000000000000001011010100001001;
assign LUT_3[36843] = 32'b00000000000000010001111111100110;
assign LUT_3[36844] = 32'b00000000000000000110011010011011;
assign LUT_3[36845] = 32'b00000000000000001101000101111000;
assign LUT_3[36846] = 32'b00000000000000001000100001111111;
assign LUT_3[36847] = 32'b00000000000000001111001101011100;
assign LUT_3[36848] = 32'b00000000000000000111000110100010;
assign LUT_3[36849] = 32'b00000000000000001101110001111111;
assign LUT_3[36850] = 32'b00000000000000001001001110000110;
assign LUT_3[36851] = 32'b00000000000000001111111001100011;
assign LUT_3[36852] = 32'b00000000000000000100010100011000;
assign LUT_3[36853] = 32'b00000000000000001010111111110101;
assign LUT_3[36854] = 32'b00000000000000000110011011111100;
assign LUT_3[36855] = 32'b00000000000000001101000111011001;
assign LUT_3[36856] = 32'b00000000000000001100011111101000;
assign LUT_3[36857] = 32'b00000000000000010011001011000101;
assign LUT_3[36858] = 32'b00000000000000001110100111001100;
assign LUT_3[36859] = 32'b00000000000000010101010010101001;
assign LUT_3[36860] = 32'b00000000000000001001101101011110;
assign LUT_3[36861] = 32'b00000000000000010000011000111011;
assign LUT_3[36862] = 32'b00000000000000001011110101000010;
assign LUT_3[36863] = 32'b00000000000000010010100000011111;
assign LUT_3[36864] = 32'b11111111111111111100110010111001;
assign LUT_3[36865] = 32'b00000000000000000011011110010110;
assign LUT_3[36866] = 32'b11111111111111111110111010011101;
assign LUT_3[36867] = 32'b00000000000000000101100101111010;
assign LUT_3[36868] = 32'b11111111111111111010000000101111;
assign LUT_3[36869] = 32'b00000000000000000000101100001100;
assign LUT_3[36870] = 32'b11111111111111111100001000010011;
assign LUT_3[36871] = 32'b00000000000000000010110011110000;
assign LUT_3[36872] = 32'b00000000000000000010001011111111;
assign LUT_3[36873] = 32'b00000000000000001000110111011100;
assign LUT_3[36874] = 32'b00000000000000000100010011100011;
assign LUT_3[36875] = 32'b00000000000000001010111111000000;
assign LUT_3[36876] = 32'b11111111111111111111011001110101;
assign LUT_3[36877] = 32'b00000000000000000110000101010010;
assign LUT_3[36878] = 32'b00000000000000000001100001011001;
assign LUT_3[36879] = 32'b00000000000000001000001100110110;
assign LUT_3[36880] = 32'b00000000000000000000000101111100;
assign LUT_3[36881] = 32'b00000000000000000110110001011001;
assign LUT_3[36882] = 32'b00000000000000000010001101100000;
assign LUT_3[36883] = 32'b00000000000000001000111000111101;
assign LUT_3[36884] = 32'b11111111111111111101010011110010;
assign LUT_3[36885] = 32'b00000000000000000011111111001111;
assign LUT_3[36886] = 32'b11111111111111111111011011010110;
assign LUT_3[36887] = 32'b00000000000000000110000110110011;
assign LUT_3[36888] = 32'b00000000000000000101011111000010;
assign LUT_3[36889] = 32'b00000000000000001100001010011111;
assign LUT_3[36890] = 32'b00000000000000000111100110100110;
assign LUT_3[36891] = 32'b00000000000000001110010010000011;
assign LUT_3[36892] = 32'b00000000000000000010101100111000;
assign LUT_3[36893] = 32'b00000000000000001001011000010101;
assign LUT_3[36894] = 32'b00000000000000000100110100011100;
assign LUT_3[36895] = 32'b00000000000000001011011111111001;
assign LUT_3[36896] = 32'b11111111111111111110000001011001;
assign LUT_3[36897] = 32'b00000000000000000100101100110110;
assign LUT_3[36898] = 32'b00000000000000000000001000111101;
assign LUT_3[36899] = 32'b00000000000000000110110100011010;
assign LUT_3[36900] = 32'b11111111111111111011001111001111;
assign LUT_3[36901] = 32'b00000000000000000001111010101100;
assign LUT_3[36902] = 32'b11111111111111111101010110110011;
assign LUT_3[36903] = 32'b00000000000000000100000010010000;
assign LUT_3[36904] = 32'b00000000000000000011011010011111;
assign LUT_3[36905] = 32'b00000000000000001010000101111100;
assign LUT_3[36906] = 32'b00000000000000000101100010000011;
assign LUT_3[36907] = 32'b00000000000000001100001101100000;
assign LUT_3[36908] = 32'b00000000000000000000101000010101;
assign LUT_3[36909] = 32'b00000000000000000111010011110010;
assign LUT_3[36910] = 32'b00000000000000000010101111111001;
assign LUT_3[36911] = 32'b00000000000000001001011011010110;
assign LUT_3[36912] = 32'b00000000000000000001010100011100;
assign LUT_3[36913] = 32'b00000000000000000111111111111001;
assign LUT_3[36914] = 32'b00000000000000000011011100000000;
assign LUT_3[36915] = 32'b00000000000000001010000111011101;
assign LUT_3[36916] = 32'b11111111111111111110100010010010;
assign LUT_3[36917] = 32'b00000000000000000101001101101111;
assign LUT_3[36918] = 32'b00000000000000000000101001110110;
assign LUT_3[36919] = 32'b00000000000000000111010101010011;
assign LUT_3[36920] = 32'b00000000000000000110101101100010;
assign LUT_3[36921] = 32'b00000000000000001101011000111111;
assign LUT_3[36922] = 32'b00000000000000001000110101000110;
assign LUT_3[36923] = 32'b00000000000000001111100000100011;
assign LUT_3[36924] = 32'b00000000000000000011111011011000;
assign LUT_3[36925] = 32'b00000000000000001010100110110101;
assign LUT_3[36926] = 32'b00000000000000000110000010111100;
assign LUT_3[36927] = 32'b00000000000000001100101110011001;
assign LUT_3[36928] = 32'b11111111111111111100101011100100;
assign LUT_3[36929] = 32'b00000000000000000011010111000001;
assign LUT_3[36930] = 32'b11111111111111111110110011001000;
assign LUT_3[36931] = 32'b00000000000000000101011110100101;
assign LUT_3[36932] = 32'b11111111111111111001111001011010;
assign LUT_3[36933] = 32'b00000000000000000000100100110111;
assign LUT_3[36934] = 32'b11111111111111111100000000111110;
assign LUT_3[36935] = 32'b00000000000000000010101100011011;
assign LUT_3[36936] = 32'b00000000000000000010000100101010;
assign LUT_3[36937] = 32'b00000000000000001000110000000111;
assign LUT_3[36938] = 32'b00000000000000000100001100001110;
assign LUT_3[36939] = 32'b00000000000000001010110111101011;
assign LUT_3[36940] = 32'b11111111111111111111010010100000;
assign LUT_3[36941] = 32'b00000000000000000101111101111101;
assign LUT_3[36942] = 32'b00000000000000000001011010000100;
assign LUT_3[36943] = 32'b00000000000000001000000101100001;
assign LUT_3[36944] = 32'b11111111111111111111111110100111;
assign LUT_3[36945] = 32'b00000000000000000110101010000100;
assign LUT_3[36946] = 32'b00000000000000000010000110001011;
assign LUT_3[36947] = 32'b00000000000000001000110001101000;
assign LUT_3[36948] = 32'b11111111111111111101001100011101;
assign LUT_3[36949] = 32'b00000000000000000011110111111010;
assign LUT_3[36950] = 32'b11111111111111111111010100000001;
assign LUT_3[36951] = 32'b00000000000000000101111111011110;
assign LUT_3[36952] = 32'b00000000000000000101010111101101;
assign LUT_3[36953] = 32'b00000000000000001100000011001010;
assign LUT_3[36954] = 32'b00000000000000000111011111010001;
assign LUT_3[36955] = 32'b00000000000000001110001010101110;
assign LUT_3[36956] = 32'b00000000000000000010100101100011;
assign LUT_3[36957] = 32'b00000000000000001001010001000000;
assign LUT_3[36958] = 32'b00000000000000000100101101000111;
assign LUT_3[36959] = 32'b00000000000000001011011000100100;
assign LUT_3[36960] = 32'b11111111111111111101111010000100;
assign LUT_3[36961] = 32'b00000000000000000100100101100001;
assign LUT_3[36962] = 32'b00000000000000000000000001101000;
assign LUT_3[36963] = 32'b00000000000000000110101101000101;
assign LUT_3[36964] = 32'b11111111111111111011000111111010;
assign LUT_3[36965] = 32'b00000000000000000001110011010111;
assign LUT_3[36966] = 32'b11111111111111111101001111011110;
assign LUT_3[36967] = 32'b00000000000000000011111010111011;
assign LUT_3[36968] = 32'b00000000000000000011010011001010;
assign LUT_3[36969] = 32'b00000000000000001001111110100111;
assign LUT_3[36970] = 32'b00000000000000000101011010101110;
assign LUT_3[36971] = 32'b00000000000000001100000110001011;
assign LUT_3[36972] = 32'b00000000000000000000100001000000;
assign LUT_3[36973] = 32'b00000000000000000111001100011101;
assign LUT_3[36974] = 32'b00000000000000000010101000100100;
assign LUT_3[36975] = 32'b00000000000000001001010100000001;
assign LUT_3[36976] = 32'b00000000000000000001001101000111;
assign LUT_3[36977] = 32'b00000000000000000111111000100100;
assign LUT_3[36978] = 32'b00000000000000000011010100101011;
assign LUT_3[36979] = 32'b00000000000000001010000000001000;
assign LUT_3[36980] = 32'b11111111111111111110011010111101;
assign LUT_3[36981] = 32'b00000000000000000101000110011010;
assign LUT_3[36982] = 32'b00000000000000000000100010100001;
assign LUT_3[36983] = 32'b00000000000000000111001101111110;
assign LUT_3[36984] = 32'b00000000000000000110100110001101;
assign LUT_3[36985] = 32'b00000000000000001101010001101010;
assign LUT_3[36986] = 32'b00000000000000001000101101110001;
assign LUT_3[36987] = 32'b00000000000000001111011001001110;
assign LUT_3[36988] = 32'b00000000000000000011110100000011;
assign LUT_3[36989] = 32'b00000000000000001010011111100000;
assign LUT_3[36990] = 32'b00000000000000000101111011100111;
assign LUT_3[36991] = 32'b00000000000000001100100111000100;
assign LUT_3[36992] = 32'b11111111111111111110111101110111;
assign LUT_3[36993] = 32'b00000000000000000101101001010100;
assign LUT_3[36994] = 32'b00000000000000000001000101011011;
assign LUT_3[36995] = 32'b00000000000000000111110000111000;
assign LUT_3[36996] = 32'b11111111111111111100001011101101;
assign LUT_3[36997] = 32'b00000000000000000010110111001010;
assign LUT_3[36998] = 32'b11111111111111111110010011010001;
assign LUT_3[36999] = 32'b00000000000000000100111110101110;
assign LUT_3[37000] = 32'b00000000000000000100010110111101;
assign LUT_3[37001] = 32'b00000000000000001011000010011010;
assign LUT_3[37002] = 32'b00000000000000000110011110100001;
assign LUT_3[37003] = 32'b00000000000000001101001001111110;
assign LUT_3[37004] = 32'b00000000000000000001100100110011;
assign LUT_3[37005] = 32'b00000000000000001000010000010000;
assign LUT_3[37006] = 32'b00000000000000000011101100010111;
assign LUT_3[37007] = 32'b00000000000000001010010111110100;
assign LUT_3[37008] = 32'b00000000000000000010010000111010;
assign LUT_3[37009] = 32'b00000000000000001000111100010111;
assign LUT_3[37010] = 32'b00000000000000000100011000011110;
assign LUT_3[37011] = 32'b00000000000000001011000011111011;
assign LUT_3[37012] = 32'b11111111111111111111011110110000;
assign LUT_3[37013] = 32'b00000000000000000110001010001101;
assign LUT_3[37014] = 32'b00000000000000000001100110010100;
assign LUT_3[37015] = 32'b00000000000000001000010001110001;
assign LUT_3[37016] = 32'b00000000000000000111101010000000;
assign LUT_3[37017] = 32'b00000000000000001110010101011101;
assign LUT_3[37018] = 32'b00000000000000001001110001100100;
assign LUT_3[37019] = 32'b00000000000000010000011101000001;
assign LUT_3[37020] = 32'b00000000000000000100110111110110;
assign LUT_3[37021] = 32'b00000000000000001011100011010011;
assign LUT_3[37022] = 32'b00000000000000000110111111011010;
assign LUT_3[37023] = 32'b00000000000000001101101010110111;
assign LUT_3[37024] = 32'b00000000000000000000001100010111;
assign LUT_3[37025] = 32'b00000000000000000110110111110100;
assign LUT_3[37026] = 32'b00000000000000000010010011111011;
assign LUT_3[37027] = 32'b00000000000000001000111111011000;
assign LUT_3[37028] = 32'b11111111111111111101011010001101;
assign LUT_3[37029] = 32'b00000000000000000100000101101010;
assign LUT_3[37030] = 32'b11111111111111111111100001110001;
assign LUT_3[37031] = 32'b00000000000000000110001101001110;
assign LUT_3[37032] = 32'b00000000000000000101100101011101;
assign LUT_3[37033] = 32'b00000000000000001100010000111010;
assign LUT_3[37034] = 32'b00000000000000000111101101000001;
assign LUT_3[37035] = 32'b00000000000000001110011000011110;
assign LUT_3[37036] = 32'b00000000000000000010110011010011;
assign LUT_3[37037] = 32'b00000000000000001001011110110000;
assign LUT_3[37038] = 32'b00000000000000000100111010110111;
assign LUT_3[37039] = 32'b00000000000000001011100110010100;
assign LUT_3[37040] = 32'b00000000000000000011011111011010;
assign LUT_3[37041] = 32'b00000000000000001010001010110111;
assign LUT_3[37042] = 32'b00000000000000000101100110111110;
assign LUT_3[37043] = 32'b00000000000000001100010010011011;
assign LUT_3[37044] = 32'b00000000000000000000101101010000;
assign LUT_3[37045] = 32'b00000000000000000111011000101101;
assign LUT_3[37046] = 32'b00000000000000000010110100110100;
assign LUT_3[37047] = 32'b00000000000000001001100000010001;
assign LUT_3[37048] = 32'b00000000000000001000111000100000;
assign LUT_3[37049] = 32'b00000000000000001111100011111101;
assign LUT_3[37050] = 32'b00000000000000001011000000000100;
assign LUT_3[37051] = 32'b00000000000000010001101011100001;
assign LUT_3[37052] = 32'b00000000000000000110000110010110;
assign LUT_3[37053] = 32'b00000000000000001100110001110011;
assign LUT_3[37054] = 32'b00000000000000001000001101111010;
assign LUT_3[37055] = 32'b00000000000000001110111001010111;
assign LUT_3[37056] = 32'b11111111111111111110110110100010;
assign LUT_3[37057] = 32'b00000000000000000101100001111111;
assign LUT_3[37058] = 32'b00000000000000000000111110000110;
assign LUT_3[37059] = 32'b00000000000000000111101001100011;
assign LUT_3[37060] = 32'b11111111111111111100000100011000;
assign LUT_3[37061] = 32'b00000000000000000010101111110101;
assign LUT_3[37062] = 32'b11111111111111111110001011111100;
assign LUT_3[37063] = 32'b00000000000000000100110111011001;
assign LUT_3[37064] = 32'b00000000000000000100001111101000;
assign LUT_3[37065] = 32'b00000000000000001010111011000101;
assign LUT_3[37066] = 32'b00000000000000000110010111001100;
assign LUT_3[37067] = 32'b00000000000000001101000010101001;
assign LUT_3[37068] = 32'b00000000000000000001011101011110;
assign LUT_3[37069] = 32'b00000000000000001000001000111011;
assign LUT_3[37070] = 32'b00000000000000000011100101000010;
assign LUT_3[37071] = 32'b00000000000000001010010000011111;
assign LUT_3[37072] = 32'b00000000000000000010001001100101;
assign LUT_3[37073] = 32'b00000000000000001000110101000010;
assign LUT_3[37074] = 32'b00000000000000000100010001001001;
assign LUT_3[37075] = 32'b00000000000000001010111100100110;
assign LUT_3[37076] = 32'b11111111111111111111010111011011;
assign LUT_3[37077] = 32'b00000000000000000110000010111000;
assign LUT_3[37078] = 32'b00000000000000000001011110111111;
assign LUT_3[37079] = 32'b00000000000000001000001010011100;
assign LUT_3[37080] = 32'b00000000000000000111100010101011;
assign LUT_3[37081] = 32'b00000000000000001110001110001000;
assign LUT_3[37082] = 32'b00000000000000001001101010001111;
assign LUT_3[37083] = 32'b00000000000000010000010101101100;
assign LUT_3[37084] = 32'b00000000000000000100110000100001;
assign LUT_3[37085] = 32'b00000000000000001011011011111110;
assign LUT_3[37086] = 32'b00000000000000000110111000000101;
assign LUT_3[37087] = 32'b00000000000000001101100011100010;
assign LUT_3[37088] = 32'b00000000000000000000000101000010;
assign LUT_3[37089] = 32'b00000000000000000110110000011111;
assign LUT_3[37090] = 32'b00000000000000000010001100100110;
assign LUT_3[37091] = 32'b00000000000000001000111000000011;
assign LUT_3[37092] = 32'b11111111111111111101010010111000;
assign LUT_3[37093] = 32'b00000000000000000011111110010101;
assign LUT_3[37094] = 32'b11111111111111111111011010011100;
assign LUT_3[37095] = 32'b00000000000000000110000101111001;
assign LUT_3[37096] = 32'b00000000000000000101011110001000;
assign LUT_3[37097] = 32'b00000000000000001100001001100101;
assign LUT_3[37098] = 32'b00000000000000000111100101101100;
assign LUT_3[37099] = 32'b00000000000000001110010001001001;
assign LUT_3[37100] = 32'b00000000000000000010101011111110;
assign LUT_3[37101] = 32'b00000000000000001001010111011011;
assign LUT_3[37102] = 32'b00000000000000000100110011100010;
assign LUT_3[37103] = 32'b00000000000000001011011110111111;
assign LUT_3[37104] = 32'b00000000000000000011011000000101;
assign LUT_3[37105] = 32'b00000000000000001010000011100010;
assign LUT_3[37106] = 32'b00000000000000000101011111101001;
assign LUT_3[37107] = 32'b00000000000000001100001011000110;
assign LUT_3[37108] = 32'b00000000000000000000100101111011;
assign LUT_3[37109] = 32'b00000000000000000111010001011000;
assign LUT_3[37110] = 32'b00000000000000000010101101011111;
assign LUT_3[37111] = 32'b00000000000000001001011000111100;
assign LUT_3[37112] = 32'b00000000000000001000110001001011;
assign LUT_3[37113] = 32'b00000000000000001111011100101000;
assign LUT_3[37114] = 32'b00000000000000001010111000101111;
assign LUT_3[37115] = 32'b00000000000000010001100100001100;
assign LUT_3[37116] = 32'b00000000000000000101111111000001;
assign LUT_3[37117] = 32'b00000000000000001100101010011110;
assign LUT_3[37118] = 32'b00000000000000001000000110100101;
assign LUT_3[37119] = 32'b00000000000000001110110010000010;
assign LUT_3[37120] = 32'b11111111111111111001000010011010;
assign LUT_3[37121] = 32'b11111111111111111111101101110111;
assign LUT_3[37122] = 32'b11111111111111111011001001111110;
assign LUT_3[37123] = 32'b00000000000000000001110101011011;
assign LUT_3[37124] = 32'b11111111111111110110010000010000;
assign LUT_3[37125] = 32'b11111111111111111100111011101101;
assign LUT_3[37126] = 32'b11111111111111111000010111110100;
assign LUT_3[37127] = 32'b11111111111111111111000011010001;
assign LUT_3[37128] = 32'b11111111111111111110011011100000;
assign LUT_3[37129] = 32'b00000000000000000101000110111101;
assign LUT_3[37130] = 32'b00000000000000000000100011000100;
assign LUT_3[37131] = 32'b00000000000000000111001110100001;
assign LUT_3[37132] = 32'b11111111111111111011101001010110;
assign LUT_3[37133] = 32'b00000000000000000010010100110011;
assign LUT_3[37134] = 32'b11111111111111111101110000111010;
assign LUT_3[37135] = 32'b00000000000000000100011100010111;
assign LUT_3[37136] = 32'b11111111111111111100010101011101;
assign LUT_3[37137] = 32'b00000000000000000011000000111010;
assign LUT_3[37138] = 32'b11111111111111111110011101000001;
assign LUT_3[37139] = 32'b00000000000000000101001000011110;
assign LUT_3[37140] = 32'b11111111111111111001100011010011;
assign LUT_3[37141] = 32'b00000000000000000000001110110000;
assign LUT_3[37142] = 32'b11111111111111111011101010110111;
assign LUT_3[37143] = 32'b00000000000000000010010110010100;
assign LUT_3[37144] = 32'b00000000000000000001101110100011;
assign LUT_3[37145] = 32'b00000000000000001000011010000000;
assign LUT_3[37146] = 32'b00000000000000000011110110000111;
assign LUT_3[37147] = 32'b00000000000000001010100001100100;
assign LUT_3[37148] = 32'b11111111111111111110111100011001;
assign LUT_3[37149] = 32'b00000000000000000101100111110110;
assign LUT_3[37150] = 32'b00000000000000000001000011111101;
assign LUT_3[37151] = 32'b00000000000000000111101111011010;
assign LUT_3[37152] = 32'b11111111111111111010010000111010;
assign LUT_3[37153] = 32'b00000000000000000000111100010111;
assign LUT_3[37154] = 32'b11111111111111111100011000011110;
assign LUT_3[37155] = 32'b00000000000000000011000011111011;
assign LUT_3[37156] = 32'b11111111111111110111011110110000;
assign LUT_3[37157] = 32'b11111111111111111110001010001101;
assign LUT_3[37158] = 32'b11111111111111111001100110010100;
assign LUT_3[37159] = 32'b00000000000000000000010001110001;
assign LUT_3[37160] = 32'b11111111111111111111101010000000;
assign LUT_3[37161] = 32'b00000000000000000110010101011101;
assign LUT_3[37162] = 32'b00000000000000000001110001100100;
assign LUT_3[37163] = 32'b00000000000000001000011101000001;
assign LUT_3[37164] = 32'b11111111111111111100110111110110;
assign LUT_3[37165] = 32'b00000000000000000011100011010011;
assign LUT_3[37166] = 32'b11111111111111111110111111011010;
assign LUT_3[37167] = 32'b00000000000000000101101010110111;
assign LUT_3[37168] = 32'b11111111111111111101100011111101;
assign LUT_3[37169] = 32'b00000000000000000100001111011010;
assign LUT_3[37170] = 32'b11111111111111111111101011100001;
assign LUT_3[37171] = 32'b00000000000000000110010110111110;
assign LUT_3[37172] = 32'b11111111111111111010110001110011;
assign LUT_3[37173] = 32'b00000000000000000001011101010000;
assign LUT_3[37174] = 32'b11111111111111111100111001010111;
assign LUT_3[37175] = 32'b00000000000000000011100100110100;
assign LUT_3[37176] = 32'b00000000000000000010111101000011;
assign LUT_3[37177] = 32'b00000000000000001001101000100000;
assign LUT_3[37178] = 32'b00000000000000000101000100100111;
assign LUT_3[37179] = 32'b00000000000000001011110000000100;
assign LUT_3[37180] = 32'b00000000000000000000001010111001;
assign LUT_3[37181] = 32'b00000000000000000110110110010110;
assign LUT_3[37182] = 32'b00000000000000000010010010011101;
assign LUT_3[37183] = 32'b00000000000000001000111101111010;
assign LUT_3[37184] = 32'b11111111111111111000111011000101;
assign LUT_3[37185] = 32'b11111111111111111111100110100010;
assign LUT_3[37186] = 32'b11111111111111111011000010101001;
assign LUT_3[37187] = 32'b00000000000000000001101110000110;
assign LUT_3[37188] = 32'b11111111111111110110001000111011;
assign LUT_3[37189] = 32'b11111111111111111100110100011000;
assign LUT_3[37190] = 32'b11111111111111111000010000011111;
assign LUT_3[37191] = 32'b11111111111111111110111011111100;
assign LUT_3[37192] = 32'b11111111111111111110010100001011;
assign LUT_3[37193] = 32'b00000000000000000100111111101000;
assign LUT_3[37194] = 32'b00000000000000000000011011101111;
assign LUT_3[37195] = 32'b00000000000000000111000111001100;
assign LUT_3[37196] = 32'b11111111111111111011100010000001;
assign LUT_3[37197] = 32'b00000000000000000010001101011110;
assign LUT_3[37198] = 32'b11111111111111111101101001100101;
assign LUT_3[37199] = 32'b00000000000000000100010101000010;
assign LUT_3[37200] = 32'b11111111111111111100001110001000;
assign LUT_3[37201] = 32'b00000000000000000010111001100101;
assign LUT_3[37202] = 32'b11111111111111111110010101101100;
assign LUT_3[37203] = 32'b00000000000000000101000001001001;
assign LUT_3[37204] = 32'b11111111111111111001011011111110;
assign LUT_3[37205] = 32'b00000000000000000000000111011011;
assign LUT_3[37206] = 32'b11111111111111111011100011100010;
assign LUT_3[37207] = 32'b00000000000000000010001110111111;
assign LUT_3[37208] = 32'b00000000000000000001100111001110;
assign LUT_3[37209] = 32'b00000000000000001000010010101011;
assign LUT_3[37210] = 32'b00000000000000000011101110110010;
assign LUT_3[37211] = 32'b00000000000000001010011010001111;
assign LUT_3[37212] = 32'b11111111111111111110110101000100;
assign LUT_3[37213] = 32'b00000000000000000101100000100001;
assign LUT_3[37214] = 32'b00000000000000000000111100101000;
assign LUT_3[37215] = 32'b00000000000000000111101000000101;
assign LUT_3[37216] = 32'b11111111111111111010001001100101;
assign LUT_3[37217] = 32'b00000000000000000000110101000010;
assign LUT_3[37218] = 32'b11111111111111111100010001001001;
assign LUT_3[37219] = 32'b00000000000000000010111100100110;
assign LUT_3[37220] = 32'b11111111111111110111010111011011;
assign LUT_3[37221] = 32'b11111111111111111110000010111000;
assign LUT_3[37222] = 32'b11111111111111111001011110111111;
assign LUT_3[37223] = 32'b00000000000000000000001010011100;
assign LUT_3[37224] = 32'b11111111111111111111100010101011;
assign LUT_3[37225] = 32'b00000000000000000110001110001000;
assign LUT_3[37226] = 32'b00000000000000000001101010001111;
assign LUT_3[37227] = 32'b00000000000000001000010101101100;
assign LUT_3[37228] = 32'b11111111111111111100110000100001;
assign LUT_3[37229] = 32'b00000000000000000011011011111110;
assign LUT_3[37230] = 32'b11111111111111111110111000000101;
assign LUT_3[37231] = 32'b00000000000000000101100011100010;
assign LUT_3[37232] = 32'b11111111111111111101011100101000;
assign LUT_3[37233] = 32'b00000000000000000100001000000101;
assign LUT_3[37234] = 32'b11111111111111111111100100001100;
assign LUT_3[37235] = 32'b00000000000000000110001111101001;
assign LUT_3[37236] = 32'b11111111111111111010101010011110;
assign LUT_3[37237] = 32'b00000000000000000001010101111011;
assign LUT_3[37238] = 32'b11111111111111111100110010000010;
assign LUT_3[37239] = 32'b00000000000000000011011101011111;
assign LUT_3[37240] = 32'b00000000000000000010110101101110;
assign LUT_3[37241] = 32'b00000000000000001001100001001011;
assign LUT_3[37242] = 32'b00000000000000000100111101010010;
assign LUT_3[37243] = 32'b00000000000000001011101000101111;
assign LUT_3[37244] = 32'b00000000000000000000000011100100;
assign LUT_3[37245] = 32'b00000000000000000110101111000001;
assign LUT_3[37246] = 32'b00000000000000000010001011001000;
assign LUT_3[37247] = 32'b00000000000000001000110110100101;
assign LUT_3[37248] = 32'b11111111111111111011001101011000;
assign LUT_3[37249] = 32'b00000000000000000001111000110101;
assign LUT_3[37250] = 32'b11111111111111111101010100111100;
assign LUT_3[37251] = 32'b00000000000000000100000000011001;
assign LUT_3[37252] = 32'b11111111111111111000011011001110;
assign LUT_3[37253] = 32'b11111111111111111111000110101011;
assign LUT_3[37254] = 32'b11111111111111111010100010110010;
assign LUT_3[37255] = 32'b00000000000000000001001110001111;
assign LUT_3[37256] = 32'b00000000000000000000100110011110;
assign LUT_3[37257] = 32'b00000000000000000111010001111011;
assign LUT_3[37258] = 32'b00000000000000000010101110000010;
assign LUT_3[37259] = 32'b00000000000000001001011001011111;
assign LUT_3[37260] = 32'b11111111111111111101110100010100;
assign LUT_3[37261] = 32'b00000000000000000100011111110001;
assign LUT_3[37262] = 32'b11111111111111111111111011111000;
assign LUT_3[37263] = 32'b00000000000000000110100111010101;
assign LUT_3[37264] = 32'b11111111111111111110100000011011;
assign LUT_3[37265] = 32'b00000000000000000101001011111000;
assign LUT_3[37266] = 32'b00000000000000000000100111111111;
assign LUT_3[37267] = 32'b00000000000000000111010011011100;
assign LUT_3[37268] = 32'b11111111111111111011101110010001;
assign LUT_3[37269] = 32'b00000000000000000010011001101110;
assign LUT_3[37270] = 32'b11111111111111111101110101110101;
assign LUT_3[37271] = 32'b00000000000000000100100001010010;
assign LUT_3[37272] = 32'b00000000000000000011111001100001;
assign LUT_3[37273] = 32'b00000000000000001010100100111110;
assign LUT_3[37274] = 32'b00000000000000000110000001000101;
assign LUT_3[37275] = 32'b00000000000000001100101100100010;
assign LUT_3[37276] = 32'b00000000000000000001000111010111;
assign LUT_3[37277] = 32'b00000000000000000111110010110100;
assign LUT_3[37278] = 32'b00000000000000000011001110111011;
assign LUT_3[37279] = 32'b00000000000000001001111010011000;
assign LUT_3[37280] = 32'b11111111111111111100011011111000;
assign LUT_3[37281] = 32'b00000000000000000011000111010101;
assign LUT_3[37282] = 32'b11111111111111111110100011011100;
assign LUT_3[37283] = 32'b00000000000000000101001110111001;
assign LUT_3[37284] = 32'b11111111111111111001101001101110;
assign LUT_3[37285] = 32'b00000000000000000000010101001011;
assign LUT_3[37286] = 32'b11111111111111111011110001010010;
assign LUT_3[37287] = 32'b00000000000000000010011100101111;
assign LUT_3[37288] = 32'b00000000000000000001110100111110;
assign LUT_3[37289] = 32'b00000000000000001000100000011011;
assign LUT_3[37290] = 32'b00000000000000000011111100100010;
assign LUT_3[37291] = 32'b00000000000000001010100111111111;
assign LUT_3[37292] = 32'b11111111111111111111000010110100;
assign LUT_3[37293] = 32'b00000000000000000101101110010001;
assign LUT_3[37294] = 32'b00000000000000000001001010011000;
assign LUT_3[37295] = 32'b00000000000000000111110101110101;
assign LUT_3[37296] = 32'b11111111111111111111101110111011;
assign LUT_3[37297] = 32'b00000000000000000110011010011000;
assign LUT_3[37298] = 32'b00000000000000000001110110011111;
assign LUT_3[37299] = 32'b00000000000000001000100001111100;
assign LUT_3[37300] = 32'b11111111111111111100111100110001;
assign LUT_3[37301] = 32'b00000000000000000011101000001110;
assign LUT_3[37302] = 32'b11111111111111111111000100010101;
assign LUT_3[37303] = 32'b00000000000000000101101111110010;
assign LUT_3[37304] = 32'b00000000000000000101001000000001;
assign LUT_3[37305] = 32'b00000000000000001011110011011110;
assign LUT_3[37306] = 32'b00000000000000000111001111100101;
assign LUT_3[37307] = 32'b00000000000000001101111011000010;
assign LUT_3[37308] = 32'b00000000000000000010010101110111;
assign LUT_3[37309] = 32'b00000000000000001001000001010100;
assign LUT_3[37310] = 32'b00000000000000000100011101011011;
assign LUT_3[37311] = 32'b00000000000000001011001000111000;
assign LUT_3[37312] = 32'b11111111111111111011000110000011;
assign LUT_3[37313] = 32'b00000000000000000001110001100000;
assign LUT_3[37314] = 32'b11111111111111111101001101100111;
assign LUT_3[37315] = 32'b00000000000000000011111001000100;
assign LUT_3[37316] = 32'b11111111111111111000010011111001;
assign LUT_3[37317] = 32'b11111111111111111110111111010110;
assign LUT_3[37318] = 32'b11111111111111111010011011011101;
assign LUT_3[37319] = 32'b00000000000000000001000110111010;
assign LUT_3[37320] = 32'b00000000000000000000011111001001;
assign LUT_3[37321] = 32'b00000000000000000111001010100110;
assign LUT_3[37322] = 32'b00000000000000000010100110101101;
assign LUT_3[37323] = 32'b00000000000000001001010010001010;
assign LUT_3[37324] = 32'b11111111111111111101101100111111;
assign LUT_3[37325] = 32'b00000000000000000100011000011100;
assign LUT_3[37326] = 32'b11111111111111111111110100100011;
assign LUT_3[37327] = 32'b00000000000000000110100000000000;
assign LUT_3[37328] = 32'b11111111111111111110011001000110;
assign LUT_3[37329] = 32'b00000000000000000101000100100011;
assign LUT_3[37330] = 32'b00000000000000000000100000101010;
assign LUT_3[37331] = 32'b00000000000000000111001100000111;
assign LUT_3[37332] = 32'b11111111111111111011100110111100;
assign LUT_3[37333] = 32'b00000000000000000010010010011001;
assign LUT_3[37334] = 32'b11111111111111111101101110100000;
assign LUT_3[37335] = 32'b00000000000000000100011001111101;
assign LUT_3[37336] = 32'b00000000000000000011110010001100;
assign LUT_3[37337] = 32'b00000000000000001010011101101001;
assign LUT_3[37338] = 32'b00000000000000000101111001110000;
assign LUT_3[37339] = 32'b00000000000000001100100101001101;
assign LUT_3[37340] = 32'b00000000000000000001000000000010;
assign LUT_3[37341] = 32'b00000000000000000111101011011111;
assign LUT_3[37342] = 32'b00000000000000000011000111100110;
assign LUT_3[37343] = 32'b00000000000000001001110011000011;
assign LUT_3[37344] = 32'b11111111111111111100010100100011;
assign LUT_3[37345] = 32'b00000000000000000011000000000000;
assign LUT_3[37346] = 32'b11111111111111111110011100000111;
assign LUT_3[37347] = 32'b00000000000000000101000111100100;
assign LUT_3[37348] = 32'b11111111111111111001100010011001;
assign LUT_3[37349] = 32'b00000000000000000000001101110110;
assign LUT_3[37350] = 32'b11111111111111111011101001111101;
assign LUT_3[37351] = 32'b00000000000000000010010101011010;
assign LUT_3[37352] = 32'b00000000000000000001101101101001;
assign LUT_3[37353] = 32'b00000000000000001000011001000110;
assign LUT_3[37354] = 32'b00000000000000000011110101001101;
assign LUT_3[37355] = 32'b00000000000000001010100000101010;
assign LUT_3[37356] = 32'b11111111111111111110111011011111;
assign LUT_3[37357] = 32'b00000000000000000101100110111100;
assign LUT_3[37358] = 32'b00000000000000000001000011000011;
assign LUT_3[37359] = 32'b00000000000000000111101110100000;
assign LUT_3[37360] = 32'b11111111111111111111100111100110;
assign LUT_3[37361] = 32'b00000000000000000110010011000011;
assign LUT_3[37362] = 32'b00000000000000000001101111001010;
assign LUT_3[37363] = 32'b00000000000000001000011010100111;
assign LUT_3[37364] = 32'b11111111111111111100110101011100;
assign LUT_3[37365] = 32'b00000000000000000011100000111001;
assign LUT_3[37366] = 32'b11111111111111111110111101000000;
assign LUT_3[37367] = 32'b00000000000000000101101000011101;
assign LUT_3[37368] = 32'b00000000000000000101000000101100;
assign LUT_3[37369] = 32'b00000000000000001011101100001001;
assign LUT_3[37370] = 32'b00000000000000000111001000010000;
assign LUT_3[37371] = 32'b00000000000000001101110011101101;
assign LUT_3[37372] = 32'b00000000000000000010001110100010;
assign LUT_3[37373] = 32'b00000000000000001000111001111111;
assign LUT_3[37374] = 32'b00000000000000000100010110000110;
assign LUT_3[37375] = 32'b00000000000000001011000001100011;
assign LUT_3[37376] = 32'b00000000000000000000001000000101;
assign LUT_3[37377] = 32'b00000000000000000110110011100010;
assign LUT_3[37378] = 32'b00000000000000000010001111101001;
assign LUT_3[37379] = 32'b00000000000000001000111011000110;
assign LUT_3[37380] = 32'b11111111111111111101010101111011;
assign LUT_3[37381] = 32'b00000000000000000100000001011000;
assign LUT_3[37382] = 32'b11111111111111111111011101011111;
assign LUT_3[37383] = 32'b00000000000000000110001000111100;
assign LUT_3[37384] = 32'b00000000000000000101100001001011;
assign LUT_3[37385] = 32'b00000000000000001100001100101000;
assign LUT_3[37386] = 32'b00000000000000000111101000101111;
assign LUT_3[37387] = 32'b00000000000000001110010100001100;
assign LUT_3[37388] = 32'b00000000000000000010101111000001;
assign LUT_3[37389] = 32'b00000000000000001001011010011110;
assign LUT_3[37390] = 32'b00000000000000000100110110100101;
assign LUT_3[37391] = 32'b00000000000000001011100010000010;
assign LUT_3[37392] = 32'b00000000000000000011011011001000;
assign LUT_3[37393] = 32'b00000000000000001010000110100101;
assign LUT_3[37394] = 32'b00000000000000000101100010101100;
assign LUT_3[37395] = 32'b00000000000000001100001110001001;
assign LUT_3[37396] = 32'b00000000000000000000101000111110;
assign LUT_3[37397] = 32'b00000000000000000111010100011011;
assign LUT_3[37398] = 32'b00000000000000000010110000100010;
assign LUT_3[37399] = 32'b00000000000000001001011011111111;
assign LUT_3[37400] = 32'b00000000000000001000110100001110;
assign LUT_3[37401] = 32'b00000000000000001111011111101011;
assign LUT_3[37402] = 32'b00000000000000001010111011110010;
assign LUT_3[37403] = 32'b00000000000000010001100111001111;
assign LUT_3[37404] = 32'b00000000000000000110000010000100;
assign LUT_3[37405] = 32'b00000000000000001100101101100001;
assign LUT_3[37406] = 32'b00000000000000001000001001101000;
assign LUT_3[37407] = 32'b00000000000000001110110101000101;
assign LUT_3[37408] = 32'b00000000000000000001010110100101;
assign LUT_3[37409] = 32'b00000000000000001000000010000010;
assign LUT_3[37410] = 32'b00000000000000000011011110001001;
assign LUT_3[37411] = 32'b00000000000000001010001001100110;
assign LUT_3[37412] = 32'b11111111111111111110100100011011;
assign LUT_3[37413] = 32'b00000000000000000101001111111000;
assign LUT_3[37414] = 32'b00000000000000000000101011111111;
assign LUT_3[37415] = 32'b00000000000000000111010111011100;
assign LUT_3[37416] = 32'b00000000000000000110101111101011;
assign LUT_3[37417] = 32'b00000000000000001101011011001000;
assign LUT_3[37418] = 32'b00000000000000001000110111001111;
assign LUT_3[37419] = 32'b00000000000000001111100010101100;
assign LUT_3[37420] = 32'b00000000000000000011111101100001;
assign LUT_3[37421] = 32'b00000000000000001010101000111110;
assign LUT_3[37422] = 32'b00000000000000000110000101000101;
assign LUT_3[37423] = 32'b00000000000000001100110000100010;
assign LUT_3[37424] = 32'b00000000000000000100101001101000;
assign LUT_3[37425] = 32'b00000000000000001011010101000101;
assign LUT_3[37426] = 32'b00000000000000000110110001001100;
assign LUT_3[37427] = 32'b00000000000000001101011100101001;
assign LUT_3[37428] = 32'b00000000000000000001110111011110;
assign LUT_3[37429] = 32'b00000000000000001000100010111011;
assign LUT_3[37430] = 32'b00000000000000000011111111000010;
assign LUT_3[37431] = 32'b00000000000000001010101010011111;
assign LUT_3[37432] = 32'b00000000000000001010000010101110;
assign LUT_3[37433] = 32'b00000000000000010000101110001011;
assign LUT_3[37434] = 32'b00000000000000001100001010010010;
assign LUT_3[37435] = 32'b00000000000000010010110101101111;
assign LUT_3[37436] = 32'b00000000000000000111010000100100;
assign LUT_3[37437] = 32'b00000000000000001101111100000001;
assign LUT_3[37438] = 32'b00000000000000001001011000001000;
assign LUT_3[37439] = 32'b00000000000000010000000011100101;
assign LUT_3[37440] = 32'b00000000000000000000000000110000;
assign LUT_3[37441] = 32'b00000000000000000110101100001101;
assign LUT_3[37442] = 32'b00000000000000000010001000010100;
assign LUT_3[37443] = 32'b00000000000000001000110011110001;
assign LUT_3[37444] = 32'b11111111111111111101001110100110;
assign LUT_3[37445] = 32'b00000000000000000011111010000011;
assign LUT_3[37446] = 32'b11111111111111111111010110001010;
assign LUT_3[37447] = 32'b00000000000000000110000001100111;
assign LUT_3[37448] = 32'b00000000000000000101011001110110;
assign LUT_3[37449] = 32'b00000000000000001100000101010011;
assign LUT_3[37450] = 32'b00000000000000000111100001011010;
assign LUT_3[37451] = 32'b00000000000000001110001100110111;
assign LUT_3[37452] = 32'b00000000000000000010100111101100;
assign LUT_3[37453] = 32'b00000000000000001001010011001001;
assign LUT_3[37454] = 32'b00000000000000000100101111010000;
assign LUT_3[37455] = 32'b00000000000000001011011010101101;
assign LUT_3[37456] = 32'b00000000000000000011010011110011;
assign LUT_3[37457] = 32'b00000000000000001001111111010000;
assign LUT_3[37458] = 32'b00000000000000000101011011010111;
assign LUT_3[37459] = 32'b00000000000000001100000110110100;
assign LUT_3[37460] = 32'b00000000000000000000100001101001;
assign LUT_3[37461] = 32'b00000000000000000111001101000110;
assign LUT_3[37462] = 32'b00000000000000000010101001001101;
assign LUT_3[37463] = 32'b00000000000000001001010100101010;
assign LUT_3[37464] = 32'b00000000000000001000101100111001;
assign LUT_3[37465] = 32'b00000000000000001111011000010110;
assign LUT_3[37466] = 32'b00000000000000001010110100011101;
assign LUT_3[37467] = 32'b00000000000000010001011111111010;
assign LUT_3[37468] = 32'b00000000000000000101111010101111;
assign LUT_3[37469] = 32'b00000000000000001100100110001100;
assign LUT_3[37470] = 32'b00000000000000001000000010010011;
assign LUT_3[37471] = 32'b00000000000000001110101101110000;
assign LUT_3[37472] = 32'b00000000000000000001001111010000;
assign LUT_3[37473] = 32'b00000000000000000111111010101101;
assign LUT_3[37474] = 32'b00000000000000000011010110110100;
assign LUT_3[37475] = 32'b00000000000000001010000010010001;
assign LUT_3[37476] = 32'b11111111111111111110011101000110;
assign LUT_3[37477] = 32'b00000000000000000101001000100011;
assign LUT_3[37478] = 32'b00000000000000000000100100101010;
assign LUT_3[37479] = 32'b00000000000000000111010000000111;
assign LUT_3[37480] = 32'b00000000000000000110101000010110;
assign LUT_3[37481] = 32'b00000000000000001101010011110011;
assign LUT_3[37482] = 32'b00000000000000001000101111111010;
assign LUT_3[37483] = 32'b00000000000000001111011011010111;
assign LUT_3[37484] = 32'b00000000000000000011110110001100;
assign LUT_3[37485] = 32'b00000000000000001010100001101001;
assign LUT_3[37486] = 32'b00000000000000000101111101110000;
assign LUT_3[37487] = 32'b00000000000000001100101001001101;
assign LUT_3[37488] = 32'b00000000000000000100100010010011;
assign LUT_3[37489] = 32'b00000000000000001011001101110000;
assign LUT_3[37490] = 32'b00000000000000000110101001110111;
assign LUT_3[37491] = 32'b00000000000000001101010101010100;
assign LUT_3[37492] = 32'b00000000000000000001110000001001;
assign LUT_3[37493] = 32'b00000000000000001000011011100110;
assign LUT_3[37494] = 32'b00000000000000000011110111101101;
assign LUT_3[37495] = 32'b00000000000000001010100011001010;
assign LUT_3[37496] = 32'b00000000000000001001111011011001;
assign LUT_3[37497] = 32'b00000000000000010000100110110110;
assign LUT_3[37498] = 32'b00000000000000001100000010111101;
assign LUT_3[37499] = 32'b00000000000000010010101110011010;
assign LUT_3[37500] = 32'b00000000000000000111001001001111;
assign LUT_3[37501] = 32'b00000000000000001101110100101100;
assign LUT_3[37502] = 32'b00000000000000001001010000110011;
assign LUT_3[37503] = 32'b00000000000000001111111100010000;
assign LUT_3[37504] = 32'b00000000000000000010010011000011;
assign LUT_3[37505] = 32'b00000000000000001000111110100000;
assign LUT_3[37506] = 32'b00000000000000000100011010100111;
assign LUT_3[37507] = 32'b00000000000000001011000110000100;
assign LUT_3[37508] = 32'b11111111111111111111100000111001;
assign LUT_3[37509] = 32'b00000000000000000110001100010110;
assign LUT_3[37510] = 32'b00000000000000000001101000011101;
assign LUT_3[37511] = 32'b00000000000000001000010011111010;
assign LUT_3[37512] = 32'b00000000000000000111101100001001;
assign LUT_3[37513] = 32'b00000000000000001110010111100110;
assign LUT_3[37514] = 32'b00000000000000001001110011101101;
assign LUT_3[37515] = 32'b00000000000000010000011111001010;
assign LUT_3[37516] = 32'b00000000000000000100111001111111;
assign LUT_3[37517] = 32'b00000000000000001011100101011100;
assign LUT_3[37518] = 32'b00000000000000000111000001100011;
assign LUT_3[37519] = 32'b00000000000000001101101101000000;
assign LUT_3[37520] = 32'b00000000000000000101100110000110;
assign LUT_3[37521] = 32'b00000000000000001100010001100011;
assign LUT_3[37522] = 32'b00000000000000000111101101101010;
assign LUT_3[37523] = 32'b00000000000000001110011001000111;
assign LUT_3[37524] = 32'b00000000000000000010110011111100;
assign LUT_3[37525] = 32'b00000000000000001001011111011001;
assign LUT_3[37526] = 32'b00000000000000000100111011100000;
assign LUT_3[37527] = 32'b00000000000000001011100110111101;
assign LUT_3[37528] = 32'b00000000000000001010111111001100;
assign LUT_3[37529] = 32'b00000000000000010001101010101001;
assign LUT_3[37530] = 32'b00000000000000001101000110110000;
assign LUT_3[37531] = 32'b00000000000000010011110010001101;
assign LUT_3[37532] = 32'b00000000000000001000001101000010;
assign LUT_3[37533] = 32'b00000000000000001110111000011111;
assign LUT_3[37534] = 32'b00000000000000001010010100100110;
assign LUT_3[37535] = 32'b00000000000000010001000000000011;
assign LUT_3[37536] = 32'b00000000000000000011100001100011;
assign LUT_3[37537] = 32'b00000000000000001010001101000000;
assign LUT_3[37538] = 32'b00000000000000000101101001000111;
assign LUT_3[37539] = 32'b00000000000000001100010100100100;
assign LUT_3[37540] = 32'b00000000000000000000101111011001;
assign LUT_3[37541] = 32'b00000000000000000111011010110110;
assign LUT_3[37542] = 32'b00000000000000000010110110111101;
assign LUT_3[37543] = 32'b00000000000000001001100010011010;
assign LUT_3[37544] = 32'b00000000000000001000111010101001;
assign LUT_3[37545] = 32'b00000000000000001111100110000110;
assign LUT_3[37546] = 32'b00000000000000001011000010001101;
assign LUT_3[37547] = 32'b00000000000000010001101101101010;
assign LUT_3[37548] = 32'b00000000000000000110001000011111;
assign LUT_3[37549] = 32'b00000000000000001100110011111100;
assign LUT_3[37550] = 32'b00000000000000001000010000000011;
assign LUT_3[37551] = 32'b00000000000000001110111011100000;
assign LUT_3[37552] = 32'b00000000000000000110110100100110;
assign LUT_3[37553] = 32'b00000000000000001101100000000011;
assign LUT_3[37554] = 32'b00000000000000001000111100001010;
assign LUT_3[37555] = 32'b00000000000000001111100111100111;
assign LUT_3[37556] = 32'b00000000000000000100000010011100;
assign LUT_3[37557] = 32'b00000000000000001010101101111001;
assign LUT_3[37558] = 32'b00000000000000000110001010000000;
assign LUT_3[37559] = 32'b00000000000000001100110101011101;
assign LUT_3[37560] = 32'b00000000000000001100001101101100;
assign LUT_3[37561] = 32'b00000000000000010010111001001001;
assign LUT_3[37562] = 32'b00000000000000001110010101010000;
assign LUT_3[37563] = 32'b00000000000000010101000000101101;
assign LUT_3[37564] = 32'b00000000000000001001011011100010;
assign LUT_3[37565] = 32'b00000000000000010000000110111111;
assign LUT_3[37566] = 32'b00000000000000001011100011000110;
assign LUT_3[37567] = 32'b00000000000000010010001110100011;
assign LUT_3[37568] = 32'b00000000000000000010001011101110;
assign LUT_3[37569] = 32'b00000000000000001000110111001011;
assign LUT_3[37570] = 32'b00000000000000000100010011010010;
assign LUT_3[37571] = 32'b00000000000000001010111110101111;
assign LUT_3[37572] = 32'b11111111111111111111011001100100;
assign LUT_3[37573] = 32'b00000000000000000110000101000001;
assign LUT_3[37574] = 32'b00000000000000000001100001001000;
assign LUT_3[37575] = 32'b00000000000000001000001100100101;
assign LUT_3[37576] = 32'b00000000000000000111100100110100;
assign LUT_3[37577] = 32'b00000000000000001110010000010001;
assign LUT_3[37578] = 32'b00000000000000001001101100011000;
assign LUT_3[37579] = 32'b00000000000000010000010111110101;
assign LUT_3[37580] = 32'b00000000000000000100110010101010;
assign LUT_3[37581] = 32'b00000000000000001011011110000111;
assign LUT_3[37582] = 32'b00000000000000000110111010001110;
assign LUT_3[37583] = 32'b00000000000000001101100101101011;
assign LUT_3[37584] = 32'b00000000000000000101011110110001;
assign LUT_3[37585] = 32'b00000000000000001100001010001110;
assign LUT_3[37586] = 32'b00000000000000000111100110010101;
assign LUT_3[37587] = 32'b00000000000000001110010001110010;
assign LUT_3[37588] = 32'b00000000000000000010101100100111;
assign LUT_3[37589] = 32'b00000000000000001001011000000100;
assign LUT_3[37590] = 32'b00000000000000000100110100001011;
assign LUT_3[37591] = 32'b00000000000000001011011111101000;
assign LUT_3[37592] = 32'b00000000000000001010110111110111;
assign LUT_3[37593] = 32'b00000000000000010001100011010100;
assign LUT_3[37594] = 32'b00000000000000001100111111011011;
assign LUT_3[37595] = 32'b00000000000000010011101010111000;
assign LUT_3[37596] = 32'b00000000000000001000000101101101;
assign LUT_3[37597] = 32'b00000000000000001110110001001010;
assign LUT_3[37598] = 32'b00000000000000001010001101010001;
assign LUT_3[37599] = 32'b00000000000000010000111000101110;
assign LUT_3[37600] = 32'b00000000000000000011011010001110;
assign LUT_3[37601] = 32'b00000000000000001010000101101011;
assign LUT_3[37602] = 32'b00000000000000000101100001110010;
assign LUT_3[37603] = 32'b00000000000000001100001101001111;
assign LUT_3[37604] = 32'b00000000000000000000101000000100;
assign LUT_3[37605] = 32'b00000000000000000111010011100001;
assign LUT_3[37606] = 32'b00000000000000000010101111101000;
assign LUT_3[37607] = 32'b00000000000000001001011011000101;
assign LUT_3[37608] = 32'b00000000000000001000110011010100;
assign LUT_3[37609] = 32'b00000000000000001111011110110001;
assign LUT_3[37610] = 32'b00000000000000001010111010111000;
assign LUT_3[37611] = 32'b00000000000000010001100110010101;
assign LUT_3[37612] = 32'b00000000000000000110000001001010;
assign LUT_3[37613] = 32'b00000000000000001100101100100111;
assign LUT_3[37614] = 32'b00000000000000001000001000101110;
assign LUT_3[37615] = 32'b00000000000000001110110100001011;
assign LUT_3[37616] = 32'b00000000000000000110101101010001;
assign LUT_3[37617] = 32'b00000000000000001101011000101110;
assign LUT_3[37618] = 32'b00000000000000001000110100110101;
assign LUT_3[37619] = 32'b00000000000000001111100000010010;
assign LUT_3[37620] = 32'b00000000000000000011111011000111;
assign LUT_3[37621] = 32'b00000000000000001010100110100100;
assign LUT_3[37622] = 32'b00000000000000000110000010101011;
assign LUT_3[37623] = 32'b00000000000000001100101110001000;
assign LUT_3[37624] = 32'b00000000000000001100000110010111;
assign LUT_3[37625] = 32'b00000000000000010010110001110100;
assign LUT_3[37626] = 32'b00000000000000001110001101111011;
assign LUT_3[37627] = 32'b00000000000000010100111001011000;
assign LUT_3[37628] = 32'b00000000000000001001010100001101;
assign LUT_3[37629] = 32'b00000000000000001111111111101010;
assign LUT_3[37630] = 32'b00000000000000001011011011110001;
assign LUT_3[37631] = 32'b00000000000000010010000111001110;
assign LUT_3[37632] = 32'b11111111111111111100010111100110;
assign LUT_3[37633] = 32'b00000000000000000011000011000011;
assign LUT_3[37634] = 32'b11111111111111111110011111001010;
assign LUT_3[37635] = 32'b00000000000000000101001010100111;
assign LUT_3[37636] = 32'b11111111111111111001100101011100;
assign LUT_3[37637] = 32'b00000000000000000000010000111001;
assign LUT_3[37638] = 32'b11111111111111111011101101000000;
assign LUT_3[37639] = 32'b00000000000000000010011000011101;
assign LUT_3[37640] = 32'b00000000000000000001110000101100;
assign LUT_3[37641] = 32'b00000000000000001000011100001001;
assign LUT_3[37642] = 32'b00000000000000000011111000010000;
assign LUT_3[37643] = 32'b00000000000000001010100011101101;
assign LUT_3[37644] = 32'b11111111111111111110111110100010;
assign LUT_3[37645] = 32'b00000000000000000101101001111111;
assign LUT_3[37646] = 32'b00000000000000000001000110000110;
assign LUT_3[37647] = 32'b00000000000000000111110001100011;
assign LUT_3[37648] = 32'b11111111111111111111101010101001;
assign LUT_3[37649] = 32'b00000000000000000110010110000110;
assign LUT_3[37650] = 32'b00000000000000000001110010001101;
assign LUT_3[37651] = 32'b00000000000000001000011101101010;
assign LUT_3[37652] = 32'b11111111111111111100111000011111;
assign LUT_3[37653] = 32'b00000000000000000011100011111100;
assign LUT_3[37654] = 32'b11111111111111111111000000000011;
assign LUT_3[37655] = 32'b00000000000000000101101011100000;
assign LUT_3[37656] = 32'b00000000000000000101000011101111;
assign LUT_3[37657] = 32'b00000000000000001011101111001100;
assign LUT_3[37658] = 32'b00000000000000000111001011010011;
assign LUT_3[37659] = 32'b00000000000000001101110110110000;
assign LUT_3[37660] = 32'b00000000000000000010010001100101;
assign LUT_3[37661] = 32'b00000000000000001000111101000010;
assign LUT_3[37662] = 32'b00000000000000000100011001001001;
assign LUT_3[37663] = 32'b00000000000000001011000100100110;
assign LUT_3[37664] = 32'b11111111111111111101100110000110;
assign LUT_3[37665] = 32'b00000000000000000100010001100011;
assign LUT_3[37666] = 32'b11111111111111111111101101101010;
assign LUT_3[37667] = 32'b00000000000000000110011001000111;
assign LUT_3[37668] = 32'b11111111111111111010110011111100;
assign LUT_3[37669] = 32'b00000000000000000001011111011001;
assign LUT_3[37670] = 32'b11111111111111111100111011100000;
assign LUT_3[37671] = 32'b00000000000000000011100110111101;
assign LUT_3[37672] = 32'b00000000000000000010111111001100;
assign LUT_3[37673] = 32'b00000000000000001001101010101001;
assign LUT_3[37674] = 32'b00000000000000000101000110110000;
assign LUT_3[37675] = 32'b00000000000000001011110010001101;
assign LUT_3[37676] = 32'b00000000000000000000001101000010;
assign LUT_3[37677] = 32'b00000000000000000110111000011111;
assign LUT_3[37678] = 32'b00000000000000000010010100100110;
assign LUT_3[37679] = 32'b00000000000000001001000000000011;
assign LUT_3[37680] = 32'b00000000000000000000111001001001;
assign LUT_3[37681] = 32'b00000000000000000111100100100110;
assign LUT_3[37682] = 32'b00000000000000000011000000101101;
assign LUT_3[37683] = 32'b00000000000000001001101100001010;
assign LUT_3[37684] = 32'b11111111111111111110000110111111;
assign LUT_3[37685] = 32'b00000000000000000100110010011100;
assign LUT_3[37686] = 32'b00000000000000000000001110100011;
assign LUT_3[37687] = 32'b00000000000000000110111010000000;
assign LUT_3[37688] = 32'b00000000000000000110010010001111;
assign LUT_3[37689] = 32'b00000000000000001100111101101100;
assign LUT_3[37690] = 32'b00000000000000001000011001110011;
assign LUT_3[37691] = 32'b00000000000000001111000101010000;
assign LUT_3[37692] = 32'b00000000000000000011100000000101;
assign LUT_3[37693] = 32'b00000000000000001010001011100010;
assign LUT_3[37694] = 32'b00000000000000000101100111101001;
assign LUT_3[37695] = 32'b00000000000000001100010011000110;
assign LUT_3[37696] = 32'b11111111111111111100010000010001;
assign LUT_3[37697] = 32'b00000000000000000010111011101110;
assign LUT_3[37698] = 32'b11111111111111111110010111110101;
assign LUT_3[37699] = 32'b00000000000000000101000011010010;
assign LUT_3[37700] = 32'b11111111111111111001011110000111;
assign LUT_3[37701] = 32'b00000000000000000000001001100100;
assign LUT_3[37702] = 32'b11111111111111111011100101101011;
assign LUT_3[37703] = 32'b00000000000000000010010001001000;
assign LUT_3[37704] = 32'b00000000000000000001101001010111;
assign LUT_3[37705] = 32'b00000000000000001000010100110100;
assign LUT_3[37706] = 32'b00000000000000000011110000111011;
assign LUT_3[37707] = 32'b00000000000000001010011100011000;
assign LUT_3[37708] = 32'b11111111111111111110110111001101;
assign LUT_3[37709] = 32'b00000000000000000101100010101010;
assign LUT_3[37710] = 32'b00000000000000000000111110110001;
assign LUT_3[37711] = 32'b00000000000000000111101010001110;
assign LUT_3[37712] = 32'b11111111111111111111100011010100;
assign LUT_3[37713] = 32'b00000000000000000110001110110001;
assign LUT_3[37714] = 32'b00000000000000000001101010111000;
assign LUT_3[37715] = 32'b00000000000000001000010110010101;
assign LUT_3[37716] = 32'b11111111111111111100110001001010;
assign LUT_3[37717] = 32'b00000000000000000011011100100111;
assign LUT_3[37718] = 32'b11111111111111111110111000101110;
assign LUT_3[37719] = 32'b00000000000000000101100100001011;
assign LUT_3[37720] = 32'b00000000000000000100111100011010;
assign LUT_3[37721] = 32'b00000000000000001011100111110111;
assign LUT_3[37722] = 32'b00000000000000000111000011111110;
assign LUT_3[37723] = 32'b00000000000000001101101111011011;
assign LUT_3[37724] = 32'b00000000000000000010001010010000;
assign LUT_3[37725] = 32'b00000000000000001000110101101101;
assign LUT_3[37726] = 32'b00000000000000000100010001110100;
assign LUT_3[37727] = 32'b00000000000000001010111101010001;
assign LUT_3[37728] = 32'b11111111111111111101011110110001;
assign LUT_3[37729] = 32'b00000000000000000100001010001110;
assign LUT_3[37730] = 32'b11111111111111111111100110010101;
assign LUT_3[37731] = 32'b00000000000000000110010001110010;
assign LUT_3[37732] = 32'b11111111111111111010101100100111;
assign LUT_3[37733] = 32'b00000000000000000001011000000100;
assign LUT_3[37734] = 32'b11111111111111111100110100001011;
assign LUT_3[37735] = 32'b00000000000000000011011111101000;
assign LUT_3[37736] = 32'b00000000000000000010110111110111;
assign LUT_3[37737] = 32'b00000000000000001001100011010100;
assign LUT_3[37738] = 32'b00000000000000000100111111011011;
assign LUT_3[37739] = 32'b00000000000000001011101010111000;
assign LUT_3[37740] = 32'b00000000000000000000000101101101;
assign LUT_3[37741] = 32'b00000000000000000110110001001010;
assign LUT_3[37742] = 32'b00000000000000000010001101010001;
assign LUT_3[37743] = 32'b00000000000000001000111000101110;
assign LUT_3[37744] = 32'b00000000000000000000110001110100;
assign LUT_3[37745] = 32'b00000000000000000111011101010001;
assign LUT_3[37746] = 32'b00000000000000000010111001011000;
assign LUT_3[37747] = 32'b00000000000000001001100100110101;
assign LUT_3[37748] = 32'b11111111111111111101111111101010;
assign LUT_3[37749] = 32'b00000000000000000100101011000111;
assign LUT_3[37750] = 32'b00000000000000000000000111001110;
assign LUT_3[37751] = 32'b00000000000000000110110010101011;
assign LUT_3[37752] = 32'b00000000000000000110001010111010;
assign LUT_3[37753] = 32'b00000000000000001100110110010111;
assign LUT_3[37754] = 32'b00000000000000001000010010011110;
assign LUT_3[37755] = 32'b00000000000000001110111101111011;
assign LUT_3[37756] = 32'b00000000000000000011011000110000;
assign LUT_3[37757] = 32'b00000000000000001010000100001101;
assign LUT_3[37758] = 32'b00000000000000000101100000010100;
assign LUT_3[37759] = 32'b00000000000000001100001011110001;
assign LUT_3[37760] = 32'b11111111111111111110100010100100;
assign LUT_3[37761] = 32'b00000000000000000101001110000001;
assign LUT_3[37762] = 32'b00000000000000000000101010001000;
assign LUT_3[37763] = 32'b00000000000000000111010101100101;
assign LUT_3[37764] = 32'b11111111111111111011110000011010;
assign LUT_3[37765] = 32'b00000000000000000010011011110111;
assign LUT_3[37766] = 32'b11111111111111111101110111111110;
assign LUT_3[37767] = 32'b00000000000000000100100011011011;
assign LUT_3[37768] = 32'b00000000000000000011111011101010;
assign LUT_3[37769] = 32'b00000000000000001010100111000111;
assign LUT_3[37770] = 32'b00000000000000000110000011001110;
assign LUT_3[37771] = 32'b00000000000000001100101110101011;
assign LUT_3[37772] = 32'b00000000000000000001001001100000;
assign LUT_3[37773] = 32'b00000000000000000111110100111101;
assign LUT_3[37774] = 32'b00000000000000000011010001000100;
assign LUT_3[37775] = 32'b00000000000000001001111100100001;
assign LUT_3[37776] = 32'b00000000000000000001110101100111;
assign LUT_3[37777] = 32'b00000000000000001000100001000100;
assign LUT_3[37778] = 32'b00000000000000000011111101001011;
assign LUT_3[37779] = 32'b00000000000000001010101000101000;
assign LUT_3[37780] = 32'b11111111111111111111000011011101;
assign LUT_3[37781] = 32'b00000000000000000101101110111010;
assign LUT_3[37782] = 32'b00000000000000000001001011000001;
assign LUT_3[37783] = 32'b00000000000000000111110110011110;
assign LUT_3[37784] = 32'b00000000000000000111001110101101;
assign LUT_3[37785] = 32'b00000000000000001101111010001010;
assign LUT_3[37786] = 32'b00000000000000001001010110010001;
assign LUT_3[37787] = 32'b00000000000000010000000001101110;
assign LUT_3[37788] = 32'b00000000000000000100011100100011;
assign LUT_3[37789] = 32'b00000000000000001011001000000000;
assign LUT_3[37790] = 32'b00000000000000000110100100000111;
assign LUT_3[37791] = 32'b00000000000000001101001111100100;
assign LUT_3[37792] = 32'b11111111111111111111110001000100;
assign LUT_3[37793] = 32'b00000000000000000110011100100001;
assign LUT_3[37794] = 32'b00000000000000000001111000101000;
assign LUT_3[37795] = 32'b00000000000000001000100100000101;
assign LUT_3[37796] = 32'b11111111111111111100111110111010;
assign LUT_3[37797] = 32'b00000000000000000011101010010111;
assign LUT_3[37798] = 32'b11111111111111111111000110011110;
assign LUT_3[37799] = 32'b00000000000000000101110001111011;
assign LUT_3[37800] = 32'b00000000000000000101001010001010;
assign LUT_3[37801] = 32'b00000000000000001011110101100111;
assign LUT_3[37802] = 32'b00000000000000000111010001101110;
assign LUT_3[37803] = 32'b00000000000000001101111101001011;
assign LUT_3[37804] = 32'b00000000000000000010011000000000;
assign LUT_3[37805] = 32'b00000000000000001001000011011101;
assign LUT_3[37806] = 32'b00000000000000000100011111100100;
assign LUT_3[37807] = 32'b00000000000000001011001011000001;
assign LUT_3[37808] = 32'b00000000000000000011000100000111;
assign LUT_3[37809] = 32'b00000000000000001001101111100100;
assign LUT_3[37810] = 32'b00000000000000000101001011101011;
assign LUT_3[37811] = 32'b00000000000000001011110111001000;
assign LUT_3[37812] = 32'b00000000000000000000010001111101;
assign LUT_3[37813] = 32'b00000000000000000110111101011010;
assign LUT_3[37814] = 32'b00000000000000000010011001100001;
assign LUT_3[37815] = 32'b00000000000000001001000100111110;
assign LUT_3[37816] = 32'b00000000000000001000011101001101;
assign LUT_3[37817] = 32'b00000000000000001111001000101010;
assign LUT_3[37818] = 32'b00000000000000001010100100110001;
assign LUT_3[37819] = 32'b00000000000000010001010000001110;
assign LUT_3[37820] = 32'b00000000000000000101101011000011;
assign LUT_3[37821] = 32'b00000000000000001100010110100000;
assign LUT_3[37822] = 32'b00000000000000000111110010100111;
assign LUT_3[37823] = 32'b00000000000000001110011110000100;
assign LUT_3[37824] = 32'b11111111111111111110011011001111;
assign LUT_3[37825] = 32'b00000000000000000101000110101100;
assign LUT_3[37826] = 32'b00000000000000000000100010110011;
assign LUT_3[37827] = 32'b00000000000000000111001110010000;
assign LUT_3[37828] = 32'b11111111111111111011101001000101;
assign LUT_3[37829] = 32'b00000000000000000010010100100010;
assign LUT_3[37830] = 32'b11111111111111111101110000101001;
assign LUT_3[37831] = 32'b00000000000000000100011100000110;
assign LUT_3[37832] = 32'b00000000000000000011110100010101;
assign LUT_3[37833] = 32'b00000000000000001010011111110010;
assign LUT_3[37834] = 32'b00000000000000000101111011111001;
assign LUT_3[37835] = 32'b00000000000000001100100111010110;
assign LUT_3[37836] = 32'b00000000000000000001000010001011;
assign LUT_3[37837] = 32'b00000000000000000111101101101000;
assign LUT_3[37838] = 32'b00000000000000000011001001101111;
assign LUT_3[37839] = 32'b00000000000000001001110101001100;
assign LUT_3[37840] = 32'b00000000000000000001101110010010;
assign LUT_3[37841] = 32'b00000000000000001000011001101111;
assign LUT_3[37842] = 32'b00000000000000000011110101110110;
assign LUT_3[37843] = 32'b00000000000000001010100001010011;
assign LUT_3[37844] = 32'b11111111111111111110111100001000;
assign LUT_3[37845] = 32'b00000000000000000101100111100101;
assign LUT_3[37846] = 32'b00000000000000000001000011101100;
assign LUT_3[37847] = 32'b00000000000000000111101111001001;
assign LUT_3[37848] = 32'b00000000000000000111000111011000;
assign LUT_3[37849] = 32'b00000000000000001101110010110101;
assign LUT_3[37850] = 32'b00000000000000001001001110111100;
assign LUT_3[37851] = 32'b00000000000000001111111010011001;
assign LUT_3[37852] = 32'b00000000000000000100010101001110;
assign LUT_3[37853] = 32'b00000000000000001011000000101011;
assign LUT_3[37854] = 32'b00000000000000000110011100110010;
assign LUT_3[37855] = 32'b00000000000000001101001000001111;
assign LUT_3[37856] = 32'b11111111111111111111101001101111;
assign LUT_3[37857] = 32'b00000000000000000110010101001100;
assign LUT_3[37858] = 32'b00000000000000000001110001010011;
assign LUT_3[37859] = 32'b00000000000000001000011100110000;
assign LUT_3[37860] = 32'b11111111111111111100110111100101;
assign LUT_3[37861] = 32'b00000000000000000011100011000010;
assign LUT_3[37862] = 32'b11111111111111111110111111001001;
assign LUT_3[37863] = 32'b00000000000000000101101010100110;
assign LUT_3[37864] = 32'b00000000000000000101000010110101;
assign LUT_3[37865] = 32'b00000000000000001011101110010010;
assign LUT_3[37866] = 32'b00000000000000000111001010011001;
assign LUT_3[37867] = 32'b00000000000000001101110101110110;
assign LUT_3[37868] = 32'b00000000000000000010010000101011;
assign LUT_3[37869] = 32'b00000000000000001000111100001000;
assign LUT_3[37870] = 32'b00000000000000000100011000001111;
assign LUT_3[37871] = 32'b00000000000000001011000011101100;
assign LUT_3[37872] = 32'b00000000000000000010111100110010;
assign LUT_3[37873] = 32'b00000000000000001001101000001111;
assign LUT_3[37874] = 32'b00000000000000000101000100010110;
assign LUT_3[37875] = 32'b00000000000000001011101111110011;
assign LUT_3[37876] = 32'b00000000000000000000001010101000;
assign LUT_3[37877] = 32'b00000000000000000110110110000101;
assign LUT_3[37878] = 32'b00000000000000000010010010001100;
assign LUT_3[37879] = 32'b00000000000000001000111101101001;
assign LUT_3[37880] = 32'b00000000000000001000010101111000;
assign LUT_3[37881] = 32'b00000000000000001111000001010101;
assign LUT_3[37882] = 32'b00000000000000001010011101011100;
assign LUT_3[37883] = 32'b00000000000000010001001000111001;
assign LUT_3[37884] = 32'b00000000000000000101100011101110;
assign LUT_3[37885] = 32'b00000000000000001100001111001011;
assign LUT_3[37886] = 32'b00000000000000000111101011010010;
assign LUT_3[37887] = 32'b00000000000000001110010110101111;
assign LUT_3[37888] = 32'b00000000000000000011010111110110;
assign LUT_3[37889] = 32'b00000000000000001010000011010011;
assign LUT_3[37890] = 32'b00000000000000000101011111011010;
assign LUT_3[37891] = 32'b00000000000000001100001010110111;
assign LUT_3[37892] = 32'b00000000000000000000100101101100;
assign LUT_3[37893] = 32'b00000000000000000111010001001001;
assign LUT_3[37894] = 32'b00000000000000000010101101010000;
assign LUT_3[37895] = 32'b00000000000000001001011000101101;
assign LUT_3[37896] = 32'b00000000000000001000110000111100;
assign LUT_3[37897] = 32'b00000000000000001111011100011001;
assign LUT_3[37898] = 32'b00000000000000001010111000100000;
assign LUT_3[37899] = 32'b00000000000000010001100011111101;
assign LUT_3[37900] = 32'b00000000000000000101111110110010;
assign LUT_3[37901] = 32'b00000000000000001100101010001111;
assign LUT_3[37902] = 32'b00000000000000001000000110010110;
assign LUT_3[37903] = 32'b00000000000000001110110001110011;
assign LUT_3[37904] = 32'b00000000000000000110101010111001;
assign LUT_3[37905] = 32'b00000000000000001101010110010110;
assign LUT_3[37906] = 32'b00000000000000001000110010011101;
assign LUT_3[37907] = 32'b00000000000000001111011101111010;
assign LUT_3[37908] = 32'b00000000000000000011111000101111;
assign LUT_3[37909] = 32'b00000000000000001010100100001100;
assign LUT_3[37910] = 32'b00000000000000000110000000010011;
assign LUT_3[37911] = 32'b00000000000000001100101011110000;
assign LUT_3[37912] = 32'b00000000000000001100000011111111;
assign LUT_3[37913] = 32'b00000000000000010010101111011100;
assign LUT_3[37914] = 32'b00000000000000001110001011100011;
assign LUT_3[37915] = 32'b00000000000000010100110111000000;
assign LUT_3[37916] = 32'b00000000000000001001010001110101;
assign LUT_3[37917] = 32'b00000000000000001111111101010010;
assign LUT_3[37918] = 32'b00000000000000001011011001011001;
assign LUT_3[37919] = 32'b00000000000000010010000100110110;
assign LUT_3[37920] = 32'b00000000000000000100100110010110;
assign LUT_3[37921] = 32'b00000000000000001011010001110011;
assign LUT_3[37922] = 32'b00000000000000000110101101111010;
assign LUT_3[37923] = 32'b00000000000000001101011001010111;
assign LUT_3[37924] = 32'b00000000000000000001110100001100;
assign LUT_3[37925] = 32'b00000000000000001000011111101001;
assign LUT_3[37926] = 32'b00000000000000000011111011110000;
assign LUT_3[37927] = 32'b00000000000000001010100111001101;
assign LUT_3[37928] = 32'b00000000000000001001111111011100;
assign LUT_3[37929] = 32'b00000000000000010000101010111001;
assign LUT_3[37930] = 32'b00000000000000001100000111000000;
assign LUT_3[37931] = 32'b00000000000000010010110010011101;
assign LUT_3[37932] = 32'b00000000000000000111001101010010;
assign LUT_3[37933] = 32'b00000000000000001101111000101111;
assign LUT_3[37934] = 32'b00000000000000001001010100110110;
assign LUT_3[37935] = 32'b00000000000000010000000000010011;
assign LUT_3[37936] = 32'b00000000000000000111111001011001;
assign LUT_3[37937] = 32'b00000000000000001110100100110110;
assign LUT_3[37938] = 32'b00000000000000001010000000111101;
assign LUT_3[37939] = 32'b00000000000000010000101100011010;
assign LUT_3[37940] = 32'b00000000000000000101000111001111;
assign LUT_3[37941] = 32'b00000000000000001011110010101100;
assign LUT_3[37942] = 32'b00000000000000000111001110110011;
assign LUT_3[37943] = 32'b00000000000000001101111010010000;
assign LUT_3[37944] = 32'b00000000000000001101010010011111;
assign LUT_3[37945] = 32'b00000000000000010011111101111100;
assign LUT_3[37946] = 32'b00000000000000001111011010000011;
assign LUT_3[37947] = 32'b00000000000000010110000101100000;
assign LUT_3[37948] = 32'b00000000000000001010100000010101;
assign LUT_3[37949] = 32'b00000000000000010001001011110010;
assign LUT_3[37950] = 32'b00000000000000001100100111111001;
assign LUT_3[37951] = 32'b00000000000000010011010011010110;
assign LUT_3[37952] = 32'b00000000000000000011010000100001;
assign LUT_3[37953] = 32'b00000000000000001001111011111110;
assign LUT_3[37954] = 32'b00000000000000000101011000000101;
assign LUT_3[37955] = 32'b00000000000000001100000011100010;
assign LUT_3[37956] = 32'b00000000000000000000011110010111;
assign LUT_3[37957] = 32'b00000000000000000111001001110100;
assign LUT_3[37958] = 32'b00000000000000000010100101111011;
assign LUT_3[37959] = 32'b00000000000000001001010001011000;
assign LUT_3[37960] = 32'b00000000000000001000101001100111;
assign LUT_3[37961] = 32'b00000000000000001111010101000100;
assign LUT_3[37962] = 32'b00000000000000001010110001001011;
assign LUT_3[37963] = 32'b00000000000000010001011100101000;
assign LUT_3[37964] = 32'b00000000000000000101110111011101;
assign LUT_3[37965] = 32'b00000000000000001100100010111010;
assign LUT_3[37966] = 32'b00000000000000000111111111000001;
assign LUT_3[37967] = 32'b00000000000000001110101010011110;
assign LUT_3[37968] = 32'b00000000000000000110100011100100;
assign LUT_3[37969] = 32'b00000000000000001101001111000001;
assign LUT_3[37970] = 32'b00000000000000001000101011001000;
assign LUT_3[37971] = 32'b00000000000000001111010110100101;
assign LUT_3[37972] = 32'b00000000000000000011110001011010;
assign LUT_3[37973] = 32'b00000000000000001010011100110111;
assign LUT_3[37974] = 32'b00000000000000000101111000111110;
assign LUT_3[37975] = 32'b00000000000000001100100100011011;
assign LUT_3[37976] = 32'b00000000000000001011111100101010;
assign LUT_3[37977] = 32'b00000000000000010010101000000111;
assign LUT_3[37978] = 32'b00000000000000001110000100001110;
assign LUT_3[37979] = 32'b00000000000000010100101111101011;
assign LUT_3[37980] = 32'b00000000000000001001001010100000;
assign LUT_3[37981] = 32'b00000000000000001111110101111101;
assign LUT_3[37982] = 32'b00000000000000001011010010000100;
assign LUT_3[37983] = 32'b00000000000000010001111101100001;
assign LUT_3[37984] = 32'b00000000000000000100011111000001;
assign LUT_3[37985] = 32'b00000000000000001011001010011110;
assign LUT_3[37986] = 32'b00000000000000000110100110100101;
assign LUT_3[37987] = 32'b00000000000000001101010010000010;
assign LUT_3[37988] = 32'b00000000000000000001101100110111;
assign LUT_3[37989] = 32'b00000000000000001000011000010100;
assign LUT_3[37990] = 32'b00000000000000000011110100011011;
assign LUT_3[37991] = 32'b00000000000000001010011111111000;
assign LUT_3[37992] = 32'b00000000000000001001111000000111;
assign LUT_3[37993] = 32'b00000000000000010000100011100100;
assign LUT_3[37994] = 32'b00000000000000001011111111101011;
assign LUT_3[37995] = 32'b00000000000000010010101011001000;
assign LUT_3[37996] = 32'b00000000000000000111000101111101;
assign LUT_3[37997] = 32'b00000000000000001101110001011010;
assign LUT_3[37998] = 32'b00000000000000001001001101100001;
assign LUT_3[37999] = 32'b00000000000000001111111000111110;
assign LUT_3[38000] = 32'b00000000000000000111110010000100;
assign LUT_3[38001] = 32'b00000000000000001110011101100001;
assign LUT_3[38002] = 32'b00000000000000001001111001101000;
assign LUT_3[38003] = 32'b00000000000000010000100101000101;
assign LUT_3[38004] = 32'b00000000000000000100111111111010;
assign LUT_3[38005] = 32'b00000000000000001011101011010111;
assign LUT_3[38006] = 32'b00000000000000000111000111011110;
assign LUT_3[38007] = 32'b00000000000000001101110010111011;
assign LUT_3[38008] = 32'b00000000000000001101001011001010;
assign LUT_3[38009] = 32'b00000000000000010011110110100111;
assign LUT_3[38010] = 32'b00000000000000001111010010101110;
assign LUT_3[38011] = 32'b00000000000000010101111110001011;
assign LUT_3[38012] = 32'b00000000000000001010011001000000;
assign LUT_3[38013] = 32'b00000000000000010001000100011101;
assign LUT_3[38014] = 32'b00000000000000001100100000100100;
assign LUT_3[38015] = 32'b00000000000000010011001100000001;
assign LUT_3[38016] = 32'b00000000000000000101100010110100;
assign LUT_3[38017] = 32'b00000000000000001100001110010001;
assign LUT_3[38018] = 32'b00000000000000000111101010011000;
assign LUT_3[38019] = 32'b00000000000000001110010101110101;
assign LUT_3[38020] = 32'b00000000000000000010110000101010;
assign LUT_3[38021] = 32'b00000000000000001001011100000111;
assign LUT_3[38022] = 32'b00000000000000000100111000001110;
assign LUT_3[38023] = 32'b00000000000000001011100011101011;
assign LUT_3[38024] = 32'b00000000000000001010111011111010;
assign LUT_3[38025] = 32'b00000000000000010001100111010111;
assign LUT_3[38026] = 32'b00000000000000001101000011011110;
assign LUT_3[38027] = 32'b00000000000000010011101110111011;
assign LUT_3[38028] = 32'b00000000000000001000001001110000;
assign LUT_3[38029] = 32'b00000000000000001110110101001101;
assign LUT_3[38030] = 32'b00000000000000001010010001010100;
assign LUT_3[38031] = 32'b00000000000000010000111100110001;
assign LUT_3[38032] = 32'b00000000000000001000110101110111;
assign LUT_3[38033] = 32'b00000000000000001111100001010100;
assign LUT_3[38034] = 32'b00000000000000001010111101011011;
assign LUT_3[38035] = 32'b00000000000000010001101000111000;
assign LUT_3[38036] = 32'b00000000000000000110000011101101;
assign LUT_3[38037] = 32'b00000000000000001100101111001010;
assign LUT_3[38038] = 32'b00000000000000001000001011010001;
assign LUT_3[38039] = 32'b00000000000000001110110110101110;
assign LUT_3[38040] = 32'b00000000000000001110001110111101;
assign LUT_3[38041] = 32'b00000000000000010100111010011010;
assign LUT_3[38042] = 32'b00000000000000010000010110100001;
assign LUT_3[38043] = 32'b00000000000000010111000001111110;
assign LUT_3[38044] = 32'b00000000000000001011011100110011;
assign LUT_3[38045] = 32'b00000000000000010010001000010000;
assign LUT_3[38046] = 32'b00000000000000001101100100010111;
assign LUT_3[38047] = 32'b00000000000000010100001111110100;
assign LUT_3[38048] = 32'b00000000000000000110110001010100;
assign LUT_3[38049] = 32'b00000000000000001101011100110001;
assign LUT_3[38050] = 32'b00000000000000001000111000111000;
assign LUT_3[38051] = 32'b00000000000000001111100100010101;
assign LUT_3[38052] = 32'b00000000000000000011111111001010;
assign LUT_3[38053] = 32'b00000000000000001010101010100111;
assign LUT_3[38054] = 32'b00000000000000000110000110101110;
assign LUT_3[38055] = 32'b00000000000000001100110010001011;
assign LUT_3[38056] = 32'b00000000000000001100001010011010;
assign LUT_3[38057] = 32'b00000000000000010010110101110111;
assign LUT_3[38058] = 32'b00000000000000001110010001111110;
assign LUT_3[38059] = 32'b00000000000000010100111101011011;
assign LUT_3[38060] = 32'b00000000000000001001011000010000;
assign LUT_3[38061] = 32'b00000000000000010000000011101101;
assign LUT_3[38062] = 32'b00000000000000001011011111110100;
assign LUT_3[38063] = 32'b00000000000000010010001011010001;
assign LUT_3[38064] = 32'b00000000000000001010000100010111;
assign LUT_3[38065] = 32'b00000000000000010000101111110100;
assign LUT_3[38066] = 32'b00000000000000001100001011111011;
assign LUT_3[38067] = 32'b00000000000000010010110111011000;
assign LUT_3[38068] = 32'b00000000000000000111010010001101;
assign LUT_3[38069] = 32'b00000000000000001101111101101010;
assign LUT_3[38070] = 32'b00000000000000001001011001110001;
assign LUT_3[38071] = 32'b00000000000000010000000101001110;
assign LUT_3[38072] = 32'b00000000000000001111011101011101;
assign LUT_3[38073] = 32'b00000000000000010110001000111010;
assign LUT_3[38074] = 32'b00000000000000010001100101000001;
assign LUT_3[38075] = 32'b00000000000000011000010000011110;
assign LUT_3[38076] = 32'b00000000000000001100101011010011;
assign LUT_3[38077] = 32'b00000000000000010011010110110000;
assign LUT_3[38078] = 32'b00000000000000001110110010110111;
assign LUT_3[38079] = 32'b00000000000000010101011110010100;
assign LUT_3[38080] = 32'b00000000000000000101011011011111;
assign LUT_3[38081] = 32'b00000000000000001100000110111100;
assign LUT_3[38082] = 32'b00000000000000000111100011000011;
assign LUT_3[38083] = 32'b00000000000000001110001110100000;
assign LUT_3[38084] = 32'b00000000000000000010101001010101;
assign LUT_3[38085] = 32'b00000000000000001001010100110010;
assign LUT_3[38086] = 32'b00000000000000000100110000111001;
assign LUT_3[38087] = 32'b00000000000000001011011100010110;
assign LUT_3[38088] = 32'b00000000000000001010110100100101;
assign LUT_3[38089] = 32'b00000000000000010001100000000010;
assign LUT_3[38090] = 32'b00000000000000001100111100001001;
assign LUT_3[38091] = 32'b00000000000000010011100111100110;
assign LUT_3[38092] = 32'b00000000000000001000000010011011;
assign LUT_3[38093] = 32'b00000000000000001110101101111000;
assign LUT_3[38094] = 32'b00000000000000001010001001111111;
assign LUT_3[38095] = 32'b00000000000000010000110101011100;
assign LUT_3[38096] = 32'b00000000000000001000101110100010;
assign LUT_3[38097] = 32'b00000000000000001111011001111111;
assign LUT_3[38098] = 32'b00000000000000001010110110000110;
assign LUT_3[38099] = 32'b00000000000000010001100001100011;
assign LUT_3[38100] = 32'b00000000000000000101111100011000;
assign LUT_3[38101] = 32'b00000000000000001100100111110101;
assign LUT_3[38102] = 32'b00000000000000001000000011111100;
assign LUT_3[38103] = 32'b00000000000000001110101111011001;
assign LUT_3[38104] = 32'b00000000000000001110000111101000;
assign LUT_3[38105] = 32'b00000000000000010100110011000101;
assign LUT_3[38106] = 32'b00000000000000010000001111001100;
assign LUT_3[38107] = 32'b00000000000000010110111010101001;
assign LUT_3[38108] = 32'b00000000000000001011010101011110;
assign LUT_3[38109] = 32'b00000000000000010010000000111011;
assign LUT_3[38110] = 32'b00000000000000001101011101000010;
assign LUT_3[38111] = 32'b00000000000000010100001000011111;
assign LUT_3[38112] = 32'b00000000000000000110101001111111;
assign LUT_3[38113] = 32'b00000000000000001101010101011100;
assign LUT_3[38114] = 32'b00000000000000001000110001100011;
assign LUT_3[38115] = 32'b00000000000000001111011101000000;
assign LUT_3[38116] = 32'b00000000000000000011110111110101;
assign LUT_3[38117] = 32'b00000000000000001010100011010010;
assign LUT_3[38118] = 32'b00000000000000000101111111011001;
assign LUT_3[38119] = 32'b00000000000000001100101010110110;
assign LUT_3[38120] = 32'b00000000000000001100000011000101;
assign LUT_3[38121] = 32'b00000000000000010010101110100010;
assign LUT_3[38122] = 32'b00000000000000001110001010101001;
assign LUT_3[38123] = 32'b00000000000000010100110110000110;
assign LUT_3[38124] = 32'b00000000000000001001010000111011;
assign LUT_3[38125] = 32'b00000000000000001111111100011000;
assign LUT_3[38126] = 32'b00000000000000001011011000011111;
assign LUT_3[38127] = 32'b00000000000000010010000011111100;
assign LUT_3[38128] = 32'b00000000000000001001111101000010;
assign LUT_3[38129] = 32'b00000000000000010000101000011111;
assign LUT_3[38130] = 32'b00000000000000001100000100100110;
assign LUT_3[38131] = 32'b00000000000000010010110000000011;
assign LUT_3[38132] = 32'b00000000000000000111001010111000;
assign LUT_3[38133] = 32'b00000000000000001101110110010101;
assign LUT_3[38134] = 32'b00000000000000001001010010011100;
assign LUT_3[38135] = 32'b00000000000000001111111101111001;
assign LUT_3[38136] = 32'b00000000000000001111010110001000;
assign LUT_3[38137] = 32'b00000000000000010110000001100101;
assign LUT_3[38138] = 32'b00000000000000010001011101101100;
assign LUT_3[38139] = 32'b00000000000000011000001001001001;
assign LUT_3[38140] = 32'b00000000000000001100100011111110;
assign LUT_3[38141] = 32'b00000000000000010011001111011011;
assign LUT_3[38142] = 32'b00000000000000001110101011100010;
assign LUT_3[38143] = 32'b00000000000000010101010110111111;
assign LUT_3[38144] = 32'b11111111111111111111100111010111;
assign LUT_3[38145] = 32'b00000000000000000110010010110100;
assign LUT_3[38146] = 32'b00000000000000000001101110111011;
assign LUT_3[38147] = 32'b00000000000000001000011010011000;
assign LUT_3[38148] = 32'b11111111111111111100110101001101;
assign LUT_3[38149] = 32'b00000000000000000011100000101010;
assign LUT_3[38150] = 32'b11111111111111111110111100110001;
assign LUT_3[38151] = 32'b00000000000000000101101000001110;
assign LUT_3[38152] = 32'b00000000000000000101000000011101;
assign LUT_3[38153] = 32'b00000000000000001011101011111010;
assign LUT_3[38154] = 32'b00000000000000000111001000000001;
assign LUT_3[38155] = 32'b00000000000000001101110011011110;
assign LUT_3[38156] = 32'b00000000000000000010001110010011;
assign LUT_3[38157] = 32'b00000000000000001000111001110000;
assign LUT_3[38158] = 32'b00000000000000000100010101110111;
assign LUT_3[38159] = 32'b00000000000000001011000001010100;
assign LUT_3[38160] = 32'b00000000000000000010111010011010;
assign LUT_3[38161] = 32'b00000000000000001001100101110111;
assign LUT_3[38162] = 32'b00000000000000000101000001111110;
assign LUT_3[38163] = 32'b00000000000000001011101101011011;
assign LUT_3[38164] = 32'b00000000000000000000001000010000;
assign LUT_3[38165] = 32'b00000000000000000110110011101101;
assign LUT_3[38166] = 32'b00000000000000000010001111110100;
assign LUT_3[38167] = 32'b00000000000000001000111011010001;
assign LUT_3[38168] = 32'b00000000000000001000010011100000;
assign LUT_3[38169] = 32'b00000000000000001110111110111101;
assign LUT_3[38170] = 32'b00000000000000001010011011000100;
assign LUT_3[38171] = 32'b00000000000000010001000110100001;
assign LUT_3[38172] = 32'b00000000000000000101100001010110;
assign LUT_3[38173] = 32'b00000000000000001100001100110011;
assign LUT_3[38174] = 32'b00000000000000000111101000111010;
assign LUT_3[38175] = 32'b00000000000000001110010100010111;
assign LUT_3[38176] = 32'b00000000000000000000110101110111;
assign LUT_3[38177] = 32'b00000000000000000111100001010100;
assign LUT_3[38178] = 32'b00000000000000000010111101011011;
assign LUT_3[38179] = 32'b00000000000000001001101000111000;
assign LUT_3[38180] = 32'b11111111111111111110000011101101;
assign LUT_3[38181] = 32'b00000000000000000100101111001010;
assign LUT_3[38182] = 32'b00000000000000000000001011010001;
assign LUT_3[38183] = 32'b00000000000000000110110110101110;
assign LUT_3[38184] = 32'b00000000000000000110001110111101;
assign LUT_3[38185] = 32'b00000000000000001100111010011010;
assign LUT_3[38186] = 32'b00000000000000001000010110100001;
assign LUT_3[38187] = 32'b00000000000000001111000001111110;
assign LUT_3[38188] = 32'b00000000000000000011011100110011;
assign LUT_3[38189] = 32'b00000000000000001010001000010000;
assign LUT_3[38190] = 32'b00000000000000000101100100010111;
assign LUT_3[38191] = 32'b00000000000000001100001111110100;
assign LUT_3[38192] = 32'b00000000000000000100001000111010;
assign LUT_3[38193] = 32'b00000000000000001010110100010111;
assign LUT_3[38194] = 32'b00000000000000000110010000011110;
assign LUT_3[38195] = 32'b00000000000000001100111011111011;
assign LUT_3[38196] = 32'b00000000000000000001010110110000;
assign LUT_3[38197] = 32'b00000000000000001000000010001101;
assign LUT_3[38198] = 32'b00000000000000000011011110010100;
assign LUT_3[38199] = 32'b00000000000000001010001001110001;
assign LUT_3[38200] = 32'b00000000000000001001100010000000;
assign LUT_3[38201] = 32'b00000000000000010000001101011101;
assign LUT_3[38202] = 32'b00000000000000001011101001100100;
assign LUT_3[38203] = 32'b00000000000000010010010101000001;
assign LUT_3[38204] = 32'b00000000000000000110101111110110;
assign LUT_3[38205] = 32'b00000000000000001101011011010011;
assign LUT_3[38206] = 32'b00000000000000001000110111011010;
assign LUT_3[38207] = 32'b00000000000000001111100010110111;
assign LUT_3[38208] = 32'b11111111111111111111100000000010;
assign LUT_3[38209] = 32'b00000000000000000110001011011111;
assign LUT_3[38210] = 32'b00000000000000000001100111100110;
assign LUT_3[38211] = 32'b00000000000000001000010011000011;
assign LUT_3[38212] = 32'b11111111111111111100101101111000;
assign LUT_3[38213] = 32'b00000000000000000011011001010101;
assign LUT_3[38214] = 32'b11111111111111111110110101011100;
assign LUT_3[38215] = 32'b00000000000000000101100000111001;
assign LUT_3[38216] = 32'b00000000000000000100111001001000;
assign LUT_3[38217] = 32'b00000000000000001011100100100101;
assign LUT_3[38218] = 32'b00000000000000000111000000101100;
assign LUT_3[38219] = 32'b00000000000000001101101100001001;
assign LUT_3[38220] = 32'b00000000000000000010000110111110;
assign LUT_3[38221] = 32'b00000000000000001000110010011011;
assign LUT_3[38222] = 32'b00000000000000000100001110100010;
assign LUT_3[38223] = 32'b00000000000000001010111001111111;
assign LUT_3[38224] = 32'b00000000000000000010110011000101;
assign LUT_3[38225] = 32'b00000000000000001001011110100010;
assign LUT_3[38226] = 32'b00000000000000000100111010101001;
assign LUT_3[38227] = 32'b00000000000000001011100110000110;
assign LUT_3[38228] = 32'b00000000000000000000000000111011;
assign LUT_3[38229] = 32'b00000000000000000110101100011000;
assign LUT_3[38230] = 32'b00000000000000000010001000011111;
assign LUT_3[38231] = 32'b00000000000000001000110011111100;
assign LUT_3[38232] = 32'b00000000000000001000001100001011;
assign LUT_3[38233] = 32'b00000000000000001110110111101000;
assign LUT_3[38234] = 32'b00000000000000001010010011101111;
assign LUT_3[38235] = 32'b00000000000000010000111111001100;
assign LUT_3[38236] = 32'b00000000000000000101011010000001;
assign LUT_3[38237] = 32'b00000000000000001100000101011110;
assign LUT_3[38238] = 32'b00000000000000000111100001100101;
assign LUT_3[38239] = 32'b00000000000000001110001101000010;
assign LUT_3[38240] = 32'b00000000000000000000101110100010;
assign LUT_3[38241] = 32'b00000000000000000111011001111111;
assign LUT_3[38242] = 32'b00000000000000000010110110000110;
assign LUT_3[38243] = 32'b00000000000000001001100001100011;
assign LUT_3[38244] = 32'b11111111111111111101111100011000;
assign LUT_3[38245] = 32'b00000000000000000100100111110101;
assign LUT_3[38246] = 32'b00000000000000000000000011111100;
assign LUT_3[38247] = 32'b00000000000000000110101111011001;
assign LUT_3[38248] = 32'b00000000000000000110000111101000;
assign LUT_3[38249] = 32'b00000000000000001100110011000101;
assign LUT_3[38250] = 32'b00000000000000001000001111001100;
assign LUT_3[38251] = 32'b00000000000000001110111010101001;
assign LUT_3[38252] = 32'b00000000000000000011010101011110;
assign LUT_3[38253] = 32'b00000000000000001010000000111011;
assign LUT_3[38254] = 32'b00000000000000000101011101000010;
assign LUT_3[38255] = 32'b00000000000000001100001000011111;
assign LUT_3[38256] = 32'b00000000000000000100000001100101;
assign LUT_3[38257] = 32'b00000000000000001010101101000010;
assign LUT_3[38258] = 32'b00000000000000000110001001001001;
assign LUT_3[38259] = 32'b00000000000000001100110100100110;
assign LUT_3[38260] = 32'b00000000000000000001001111011011;
assign LUT_3[38261] = 32'b00000000000000000111111010111000;
assign LUT_3[38262] = 32'b00000000000000000011010110111111;
assign LUT_3[38263] = 32'b00000000000000001010000010011100;
assign LUT_3[38264] = 32'b00000000000000001001011010101011;
assign LUT_3[38265] = 32'b00000000000000010000000110001000;
assign LUT_3[38266] = 32'b00000000000000001011100010001111;
assign LUT_3[38267] = 32'b00000000000000010010001101101100;
assign LUT_3[38268] = 32'b00000000000000000110101000100001;
assign LUT_3[38269] = 32'b00000000000000001101010011111110;
assign LUT_3[38270] = 32'b00000000000000001000110000000101;
assign LUT_3[38271] = 32'b00000000000000001111011011100010;
assign LUT_3[38272] = 32'b00000000000000000001110010010101;
assign LUT_3[38273] = 32'b00000000000000001000011101110010;
assign LUT_3[38274] = 32'b00000000000000000011111001111001;
assign LUT_3[38275] = 32'b00000000000000001010100101010110;
assign LUT_3[38276] = 32'b11111111111111111111000000001011;
assign LUT_3[38277] = 32'b00000000000000000101101011101000;
assign LUT_3[38278] = 32'b00000000000000000001000111101111;
assign LUT_3[38279] = 32'b00000000000000000111110011001100;
assign LUT_3[38280] = 32'b00000000000000000111001011011011;
assign LUT_3[38281] = 32'b00000000000000001101110110111000;
assign LUT_3[38282] = 32'b00000000000000001001010010111111;
assign LUT_3[38283] = 32'b00000000000000001111111110011100;
assign LUT_3[38284] = 32'b00000000000000000100011001010001;
assign LUT_3[38285] = 32'b00000000000000001011000100101110;
assign LUT_3[38286] = 32'b00000000000000000110100000110101;
assign LUT_3[38287] = 32'b00000000000000001101001100010010;
assign LUT_3[38288] = 32'b00000000000000000101000101011000;
assign LUT_3[38289] = 32'b00000000000000001011110000110101;
assign LUT_3[38290] = 32'b00000000000000000111001100111100;
assign LUT_3[38291] = 32'b00000000000000001101111000011001;
assign LUT_3[38292] = 32'b00000000000000000010010011001110;
assign LUT_3[38293] = 32'b00000000000000001000111110101011;
assign LUT_3[38294] = 32'b00000000000000000100011010110010;
assign LUT_3[38295] = 32'b00000000000000001011000110001111;
assign LUT_3[38296] = 32'b00000000000000001010011110011110;
assign LUT_3[38297] = 32'b00000000000000010001001001111011;
assign LUT_3[38298] = 32'b00000000000000001100100110000010;
assign LUT_3[38299] = 32'b00000000000000010011010001011111;
assign LUT_3[38300] = 32'b00000000000000000111101100010100;
assign LUT_3[38301] = 32'b00000000000000001110010111110001;
assign LUT_3[38302] = 32'b00000000000000001001110011111000;
assign LUT_3[38303] = 32'b00000000000000010000011111010101;
assign LUT_3[38304] = 32'b00000000000000000011000000110101;
assign LUT_3[38305] = 32'b00000000000000001001101100010010;
assign LUT_3[38306] = 32'b00000000000000000101001000011001;
assign LUT_3[38307] = 32'b00000000000000001011110011110110;
assign LUT_3[38308] = 32'b00000000000000000000001110101011;
assign LUT_3[38309] = 32'b00000000000000000110111010001000;
assign LUT_3[38310] = 32'b00000000000000000010010110001111;
assign LUT_3[38311] = 32'b00000000000000001001000001101100;
assign LUT_3[38312] = 32'b00000000000000001000011001111011;
assign LUT_3[38313] = 32'b00000000000000001111000101011000;
assign LUT_3[38314] = 32'b00000000000000001010100001011111;
assign LUT_3[38315] = 32'b00000000000000010001001100111100;
assign LUT_3[38316] = 32'b00000000000000000101100111110001;
assign LUT_3[38317] = 32'b00000000000000001100010011001110;
assign LUT_3[38318] = 32'b00000000000000000111101111010101;
assign LUT_3[38319] = 32'b00000000000000001110011010110010;
assign LUT_3[38320] = 32'b00000000000000000110010011111000;
assign LUT_3[38321] = 32'b00000000000000001100111111010101;
assign LUT_3[38322] = 32'b00000000000000001000011011011100;
assign LUT_3[38323] = 32'b00000000000000001111000110111001;
assign LUT_3[38324] = 32'b00000000000000000011100001101110;
assign LUT_3[38325] = 32'b00000000000000001010001101001011;
assign LUT_3[38326] = 32'b00000000000000000101101001010010;
assign LUT_3[38327] = 32'b00000000000000001100010100101111;
assign LUT_3[38328] = 32'b00000000000000001011101100111110;
assign LUT_3[38329] = 32'b00000000000000010010011000011011;
assign LUT_3[38330] = 32'b00000000000000001101110100100010;
assign LUT_3[38331] = 32'b00000000000000010100011111111111;
assign LUT_3[38332] = 32'b00000000000000001000111010110100;
assign LUT_3[38333] = 32'b00000000000000001111100110010001;
assign LUT_3[38334] = 32'b00000000000000001011000010011000;
assign LUT_3[38335] = 32'b00000000000000010001101101110101;
assign LUT_3[38336] = 32'b00000000000000000001101011000000;
assign LUT_3[38337] = 32'b00000000000000001000010110011101;
assign LUT_3[38338] = 32'b00000000000000000011110010100100;
assign LUT_3[38339] = 32'b00000000000000001010011110000001;
assign LUT_3[38340] = 32'b11111111111111111110111000110110;
assign LUT_3[38341] = 32'b00000000000000000101100100010011;
assign LUT_3[38342] = 32'b00000000000000000001000000011010;
assign LUT_3[38343] = 32'b00000000000000000111101011110111;
assign LUT_3[38344] = 32'b00000000000000000111000100000110;
assign LUT_3[38345] = 32'b00000000000000001101101111100011;
assign LUT_3[38346] = 32'b00000000000000001001001011101010;
assign LUT_3[38347] = 32'b00000000000000001111110111000111;
assign LUT_3[38348] = 32'b00000000000000000100010001111100;
assign LUT_3[38349] = 32'b00000000000000001010111101011001;
assign LUT_3[38350] = 32'b00000000000000000110011001100000;
assign LUT_3[38351] = 32'b00000000000000001101000100111101;
assign LUT_3[38352] = 32'b00000000000000000100111110000011;
assign LUT_3[38353] = 32'b00000000000000001011101001100000;
assign LUT_3[38354] = 32'b00000000000000000111000101100111;
assign LUT_3[38355] = 32'b00000000000000001101110001000100;
assign LUT_3[38356] = 32'b00000000000000000010001011111001;
assign LUT_3[38357] = 32'b00000000000000001000110111010110;
assign LUT_3[38358] = 32'b00000000000000000100010011011101;
assign LUT_3[38359] = 32'b00000000000000001010111110111010;
assign LUT_3[38360] = 32'b00000000000000001010010111001001;
assign LUT_3[38361] = 32'b00000000000000010001000010100110;
assign LUT_3[38362] = 32'b00000000000000001100011110101101;
assign LUT_3[38363] = 32'b00000000000000010011001010001010;
assign LUT_3[38364] = 32'b00000000000000000111100100111111;
assign LUT_3[38365] = 32'b00000000000000001110010000011100;
assign LUT_3[38366] = 32'b00000000000000001001101100100011;
assign LUT_3[38367] = 32'b00000000000000010000011000000000;
assign LUT_3[38368] = 32'b00000000000000000010111001100000;
assign LUT_3[38369] = 32'b00000000000000001001100100111101;
assign LUT_3[38370] = 32'b00000000000000000101000001000100;
assign LUT_3[38371] = 32'b00000000000000001011101100100001;
assign LUT_3[38372] = 32'b00000000000000000000000111010110;
assign LUT_3[38373] = 32'b00000000000000000110110010110011;
assign LUT_3[38374] = 32'b00000000000000000010001110111010;
assign LUT_3[38375] = 32'b00000000000000001000111010010111;
assign LUT_3[38376] = 32'b00000000000000001000010010100110;
assign LUT_3[38377] = 32'b00000000000000001110111110000011;
assign LUT_3[38378] = 32'b00000000000000001010011010001010;
assign LUT_3[38379] = 32'b00000000000000010001000101100111;
assign LUT_3[38380] = 32'b00000000000000000101100000011100;
assign LUT_3[38381] = 32'b00000000000000001100001011111001;
assign LUT_3[38382] = 32'b00000000000000000111101000000000;
assign LUT_3[38383] = 32'b00000000000000001110010011011101;
assign LUT_3[38384] = 32'b00000000000000000110001100100011;
assign LUT_3[38385] = 32'b00000000000000001100111000000000;
assign LUT_3[38386] = 32'b00000000000000001000010100000111;
assign LUT_3[38387] = 32'b00000000000000001110111111100100;
assign LUT_3[38388] = 32'b00000000000000000011011010011001;
assign LUT_3[38389] = 32'b00000000000000001010000101110110;
assign LUT_3[38390] = 32'b00000000000000000101100001111101;
assign LUT_3[38391] = 32'b00000000000000001100001101011010;
assign LUT_3[38392] = 32'b00000000000000001011100101101001;
assign LUT_3[38393] = 32'b00000000000000010010010001000110;
assign LUT_3[38394] = 32'b00000000000000001101101101001101;
assign LUT_3[38395] = 32'b00000000000000010100011000101010;
assign LUT_3[38396] = 32'b00000000000000001000110011011111;
assign LUT_3[38397] = 32'b00000000000000001111011110111100;
assign LUT_3[38398] = 32'b00000000000000001010111011000011;
assign LUT_3[38399] = 32'b00000000000000010001100110100000;
assign LUT_3[38400] = 32'b00000000000000000110101101000010;
assign LUT_3[38401] = 32'b00000000000000001101011000011111;
assign LUT_3[38402] = 32'b00000000000000001000110100100110;
assign LUT_3[38403] = 32'b00000000000000001111100000000011;
assign LUT_3[38404] = 32'b00000000000000000011111010111000;
assign LUT_3[38405] = 32'b00000000000000001010100110010101;
assign LUT_3[38406] = 32'b00000000000000000110000010011100;
assign LUT_3[38407] = 32'b00000000000000001100101101111001;
assign LUT_3[38408] = 32'b00000000000000001100000110001000;
assign LUT_3[38409] = 32'b00000000000000010010110001100101;
assign LUT_3[38410] = 32'b00000000000000001110001101101100;
assign LUT_3[38411] = 32'b00000000000000010100111001001001;
assign LUT_3[38412] = 32'b00000000000000001001010011111110;
assign LUT_3[38413] = 32'b00000000000000001111111111011011;
assign LUT_3[38414] = 32'b00000000000000001011011011100010;
assign LUT_3[38415] = 32'b00000000000000010010000110111111;
assign LUT_3[38416] = 32'b00000000000000001010000000000101;
assign LUT_3[38417] = 32'b00000000000000010000101011100010;
assign LUT_3[38418] = 32'b00000000000000001100000111101001;
assign LUT_3[38419] = 32'b00000000000000010010110011000110;
assign LUT_3[38420] = 32'b00000000000000000111001101111011;
assign LUT_3[38421] = 32'b00000000000000001101111001011000;
assign LUT_3[38422] = 32'b00000000000000001001010101011111;
assign LUT_3[38423] = 32'b00000000000000010000000000111100;
assign LUT_3[38424] = 32'b00000000000000001111011001001011;
assign LUT_3[38425] = 32'b00000000000000010110000100101000;
assign LUT_3[38426] = 32'b00000000000000010001100000101111;
assign LUT_3[38427] = 32'b00000000000000011000001100001100;
assign LUT_3[38428] = 32'b00000000000000001100100111000001;
assign LUT_3[38429] = 32'b00000000000000010011010010011110;
assign LUT_3[38430] = 32'b00000000000000001110101110100101;
assign LUT_3[38431] = 32'b00000000000000010101011010000010;
assign LUT_3[38432] = 32'b00000000000000000111111011100010;
assign LUT_3[38433] = 32'b00000000000000001110100110111111;
assign LUT_3[38434] = 32'b00000000000000001010000011000110;
assign LUT_3[38435] = 32'b00000000000000010000101110100011;
assign LUT_3[38436] = 32'b00000000000000000101001001011000;
assign LUT_3[38437] = 32'b00000000000000001011110100110101;
assign LUT_3[38438] = 32'b00000000000000000111010000111100;
assign LUT_3[38439] = 32'b00000000000000001101111100011001;
assign LUT_3[38440] = 32'b00000000000000001101010100101000;
assign LUT_3[38441] = 32'b00000000000000010100000000000101;
assign LUT_3[38442] = 32'b00000000000000001111011100001100;
assign LUT_3[38443] = 32'b00000000000000010110000111101001;
assign LUT_3[38444] = 32'b00000000000000001010100010011110;
assign LUT_3[38445] = 32'b00000000000000010001001101111011;
assign LUT_3[38446] = 32'b00000000000000001100101010000010;
assign LUT_3[38447] = 32'b00000000000000010011010101011111;
assign LUT_3[38448] = 32'b00000000000000001011001110100101;
assign LUT_3[38449] = 32'b00000000000000010001111010000010;
assign LUT_3[38450] = 32'b00000000000000001101010110001001;
assign LUT_3[38451] = 32'b00000000000000010100000001100110;
assign LUT_3[38452] = 32'b00000000000000001000011100011011;
assign LUT_3[38453] = 32'b00000000000000001111000111111000;
assign LUT_3[38454] = 32'b00000000000000001010100011111111;
assign LUT_3[38455] = 32'b00000000000000010001001111011100;
assign LUT_3[38456] = 32'b00000000000000010000100111101011;
assign LUT_3[38457] = 32'b00000000000000010111010011001000;
assign LUT_3[38458] = 32'b00000000000000010010101111001111;
assign LUT_3[38459] = 32'b00000000000000011001011010101100;
assign LUT_3[38460] = 32'b00000000000000001101110101100001;
assign LUT_3[38461] = 32'b00000000000000010100100000111110;
assign LUT_3[38462] = 32'b00000000000000001111111101000101;
assign LUT_3[38463] = 32'b00000000000000010110101000100010;
assign LUT_3[38464] = 32'b00000000000000000110100101101101;
assign LUT_3[38465] = 32'b00000000000000001101010001001010;
assign LUT_3[38466] = 32'b00000000000000001000101101010001;
assign LUT_3[38467] = 32'b00000000000000001111011000101110;
assign LUT_3[38468] = 32'b00000000000000000011110011100011;
assign LUT_3[38469] = 32'b00000000000000001010011111000000;
assign LUT_3[38470] = 32'b00000000000000000101111011000111;
assign LUT_3[38471] = 32'b00000000000000001100100110100100;
assign LUT_3[38472] = 32'b00000000000000001011111110110011;
assign LUT_3[38473] = 32'b00000000000000010010101010010000;
assign LUT_3[38474] = 32'b00000000000000001110000110010111;
assign LUT_3[38475] = 32'b00000000000000010100110001110100;
assign LUT_3[38476] = 32'b00000000000000001001001100101001;
assign LUT_3[38477] = 32'b00000000000000001111111000000110;
assign LUT_3[38478] = 32'b00000000000000001011010100001101;
assign LUT_3[38479] = 32'b00000000000000010001111111101010;
assign LUT_3[38480] = 32'b00000000000000001001111000110000;
assign LUT_3[38481] = 32'b00000000000000010000100100001101;
assign LUT_3[38482] = 32'b00000000000000001100000000010100;
assign LUT_3[38483] = 32'b00000000000000010010101011110001;
assign LUT_3[38484] = 32'b00000000000000000111000110100110;
assign LUT_3[38485] = 32'b00000000000000001101110010000011;
assign LUT_3[38486] = 32'b00000000000000001001001110001010;
assign LUT_3[38487] = 32'b00000000000000001111111001100111;
assign LUT_3[38488] = 32'b00000000000000001111010001110110;
assign LUT_3[38489] = 32'b00000000000000010101111101010011;
assign LUT_3[38490] = 32'b00000000000000010001011001011010;
assign LUT_3[38491] = 32'b00000000000000011000000100110111;
assign LUT_3[38492] = 32'b00000000000000001100011111101100;
assign LUT_3[38493] = 32'b00000000000000010011001011001001;
assign LUT_3[38494] = 32'b00000000000000001110100111010000;
assign LUT_3[38495] = 32'b00000000000000010101010010101101;
assign LUT_3[38496] = 32'b00000000000000000111110100001101;
assign LUT_3[38497] = 32'b00000000000000001110011111101010;
assign LUT_3[38498] = 32'b00000000000000001001111011110001;
assign LUT_3[38499] = 32'b00000000000000010000100111001110;
assign LUT_3[38500] = 32'b00000000000000000101000010000011;
assign LUT_3[38501] = 32'b00000000000000001011101101100000;
assign LUT_3[38502] = 32'b00000000000000000111001001100111;
assign LUT_3[38503] = 32'b00000000000000001101110101000100;
assign LUT_3[38504] = 32'b00000000000000001101001101010011;
assign LUT_3[38505] = 32'b00000000000000010011111000110000;
assign LUT_3[38506] = 32'b00000000000000001111010100110111;
assign LUT_3[38507] = 32'b00000000000000010110000000010100;
assign LUT_3[38508] = 32'b00000000000000001010011011001001;
assign LUT_3[38509] = 32'b00000000000000010001000110100110;
assign LUT_3[38510] = 32'b00000000000000001100100010101101;
assign LUT_3[38511] = 32'b00000000000000010011001110001010;
assign LUT_3[38512] = 32'b00000000000000001011000111010000;
assign LUT_3[38513] = 32'b00000000000000010001110010101101;
assign LUT_3[38514] = 32'b00000000000000001101001110110100;
assign LUT_3[38515] = 32'b00000000000000010011111010010001;
assign LUT_3[38516] = 32'b00000000000000001000010101000110;
assign LUT_3[38517] = 32'b00000000000000001111000000100011;
assign LUT_3[38518] = 32'b00000000000000001010011100101010;
assign LUT_3[38519] = 32'b00000000000000010001001000000111;
assign LUT_3[38520] = 32'b00000000000000010000100000010110;
assign LUT_3[38521] = 32'b00000000000000010111001011110011;
assign LUT_3[38522] = 32'b00000000000000010010100111111010;
assign LUT_3[38523] = 32'b00000000000000011001010011010111;
assign LUT_3[38524] = 32'b00000000000000001101101110001100;
assign LUT_3[38525] = 32'b00000000000000010100011001101001;
assign LUT_3[38526] = 32'b00000000000000001111110101110000;
assign LUT_3[38527] = 32'b00000000000000010110100001001101;
assign LUT_3[38528] = 32'b00000000000000001000111000000000;
assign LUT_3[38529] = 32'b00000000000000001111100011011101;
assign LUT_3[38530] = 32'b00000000000000001010111111100100;
assign LUT_3[38531] = 32'b00000000000000010001101011000001;
assign LUT_3[38532] = 32'b00000000000000000110000101110110;
assign LUT_3[38533] = 32'b00000000000000001100110001010011;
assign LUT_3[38534] = 32'b00000000000000001000001101011010;
assign LUT_3[38535] = 32'b00000000000000001110111000110111;
assign LUT_3[38536] = 32'b00000000000000001110010001000110;
assign LUT_3[38537] = 32'b00000000000000010100111100100011;
assign LUT_3[38538] = 32'b00000000000000010000011000101010;
assign LUT_3[38539] = 32'b00000000000000010111000100000111;
assign LUT_3[38540] = 32'b00000000000000001011011110111100;
assign LUT_3[38541] = 32'b00000000000000010010001010011001;
assign LUT_3[38542] = 32'b00000000000000001101100110100000;
assign LUT_3[38543] = 32'b00000000000000010100010001111101;
assign LUT_3[38544] = 32'b00000000000000001100001011000011;
assign LUT_3[38545] = 32'b00000000000000010010110110100000;
assign LUT_3[38546] = 32'b00000000000000001110010010100111;
assign LUT_3[38547] = 32'b00000000000000010100111110000100;
assign LUT_3[38548] = 32'b00000000000000001001011000111001;
assign LUT_3[38549] = 32'b00000000000000010000000100010110;
assign LUT_3[38550] = 32'b00000000000000001011100000011101;
assign LUT_3[38551] = 32'b00000000000000010010001011111010;
assign LUT_3[38552] = 32'b00000000000000010001100100001001;
assign LUT_3[38553] = 32'b00000000000000011000001111100110;
assign LUT_3[38554] = 32'b00000000000000010011101011101101;
assign LUT_3[38555] = 32'b00000000000000011010010111001010;
assign LUT_3[38556] = 32'b00000000000000001110110001111111;
assign LUT_3[38557] = 32'b00000000000000010101011101011100;
assign LUT_3[38558] = 32'b00000000000000010000111001100011;
assign LUT_3[38559] = 32'b00000000000000010111100101000000;
assign LUT_3[38560] = 32'b00000000000000001010000110100000;
assign LUT_3[38561] = 32'b00000000000000010000110001111101;
assign LUT_3[38562] = 32'b00000000000000001100001110000100;
assign LUT_3[38563] = 32'b00000000000000010010111001100001;
assign LUT_3[38564] = 32'b00000000000000000111010100010110;
assign LUT_3[38565] = 32'b00000000000000001101111111110011;
assign LUT_3[38566] = 32'b00000000000000001001011011111010;
assign LUT_3[38567] = 32'b00000000000000010000000111010111;
assign LUT_3[38568] = 32'b00000000000000001111011111100110;
assign LUT_3[38569] = 32'b00000000000000010110001011000011;
assign LUT_3[38570] = 32'b00000000000000010001100111001010;
assign LUT_3[38571] = 32'b00000000000000011000010010100111;
assign LUT_3[38572] = 32'b00000000000000001100101101011100;
assign LUT_3[38573] = 32'b00000000000000010011011000111001;
assign LUT_3[38574] = 32'b00000000000000001110110101000000;
assign LUT_3[38575] = 32'b00000000000000010101100000011101;
assign LUT_3[38576] = 32'b00000000000000001101011001100011;
assign LUT_3[38577] = 32'b00000000000000010100000101000000;
assign LUT_3[38578] = 32'b00000000000000001111100001000111;
assign LUT_3[38579] = 32'b00000000000000010110001100100100;
assign LUT_3[38580] = 32'b00000000000000001010100111011001;
assign LUT_3[38581] = 32'b00000000000000010001010010110110;
assign LUT_3[38582] = 32'b00000000000000001100101110111101;
assign LUT_3[38583] = 32'b00000000000000010011011010011010;
assign LUT_3[38584] = 32'b00000000000000010010110010101001;
assign LUT_3[38585] = 32'b00000000000000011001011110000110;
assign LUT_3[38586] = 32'b00000000000000010100111010001101;
assign LUT_3[38587] = 32'b00000000000000011011100101101010;
assign LUT_3[38588] = 32'b00000000000000010000000000011111;
assign LUT_3[38589] = 32'b00000000000000010110101011111100;
assign LUT_3[38590] = 32'b00000000000000010010001000000011;
assign LUT_3[38591] = 32'b00000000000000011000110011100000;
assign LUT_3[38592] = 32'b00000000000000001000110000101011;
assign LUT_3[38593] = 32'b00000000000000001111011100001000;
assign LUT_3[38594] = 32'b00000000000000001010111000001111;
assign LUT_3[38595] = 32'b00000000000000010001100011101100;
assign LUT_3[38596] = 32'b00000000000000000101111110100001;
assign LUT_3[38597] = 32'b00000000000000001100101001111110;
assign LUT_3[38598] = 32'b00000000000000001000000110000101;
assign LUT_3[38599] = 32'b00000000000000001110110001100010;
assign LUT_3[38600] = 32'b00000000000000001110001001110001;
assign LUT_3[38601] = 32'b00000000000000010100110101001110;
assign LUT_3[38602] = 32'b00000000000000010000010001010101;
assign LUT_3[38603] = 32'b00000000000000010110111100110010;
assign LUT_3[38604] = 32'b00000000000000001011010111100111;
assign LUT_3[38605] = 32'b00000000000000010010000011000100;
assign LUT_3[38606] = 32'b00000000000000001101011111001011;
assign LUT_3[38607] = 32'b00000000000000010100001010101000;
assign LUT_3[38608] = 32'b00000000000000001100000011101110;
assign LUT_3[38609] = 32'b00000000000000010010101111001011;
assign LUT_3[38610] = 32'b00000000000000001110001011010010;
assign LUT_3[38611] = 32'b00000000000000010100110110101111;
assign LUT_3[38612] = 32'b00000000000000001001010001100100;
assign LUT_3[38613] = 32'b00000000000000001111111101000001;
assign LUT_3[38614] = 32'b00000000000000001011011001001000;
assign LUT_3[38615] = 32'b00000000000000010010000100100101;
assign LUT_3[38616] = 32'b00000000000000010001011100110100;
assign LUT_3[38617] = 32'b00000000000000011000001000010001;
assign LUT_3[38618] = 32'b00000000000000010011100100011000;
assign LUT_3[38619] = 32'b00000000000000011010001111110101;
assign LUT_3[38620] = 32'b00000000000000001110101010101010;
assign LUT_3[38621] = 32'b00000000000000010101010110000111;
assign LUT_3[38622] = 32'b00000000000000010000110010001110;
assign LUT_3[38623] = 32'b00000000000000010111011101101011;
assign LUT_3[38624] = 32'b00000000000000001001111111001011;
assign LUT_3[38625] = 32'b00000000000000010000101010101000;
assign LUT_3[38626] = 32'b00000000000000001100000110101111;
assign LUT_3[38627] = 32'b00000000000000010010110010001100;
assign LUT_3[38628] = 32'b00000000000000000111001101000001;
assign LUT_3[38629] = 32'b00000000000000001101111000011110;
assign LUT_3[38630] = 32'b00000000000000001001010100100101;
assign LUT_3[38631] = 32'b00000000000000010000000000000010;
assign LUT_3[38632] = 32'b00000000000000001111011000010001;
assign LUT_3[38633] = 32'b00000000000000010110000011101110;
assign LUT_3[38634] = 32'b00000000000000010001011111110101;
assign LUT_3[38635] = 32'b00000000000000011000001011010010;
assign LUT_3[38636] = 32'b00000000000000001100100110000111;
assign LUT_3[38637] = 32'b00000000000000010011010001100100;
assign LUT_3[38638] = 32'b00000000000000001110101101101011;
assign LUT_3[38639] = 32'b00000000000000010101011001001000;
assign LUT_3[38640] = 32'b00000000000000001101010010001110;
assign LUT_3[38641] = 32'b00000000000000010011111101101011;
assign LUT_3[38642] = 32'b00000000000000001111011001110010;
assign LUT_3[38643] = 32'b00000000000000010110000101001111;
assign LUT_3[38644] = 32'b00000000000000001010100000000100;
assign LUT_3[38645] = 32'b00000000000000010001001011100001;
assign LUT_3[38646] = 32'b00000000000000001100100111101000;
assign LUT_3[38647] = 32'b00000000000000010011010011000101;
assign LUT_3[38648] = 32'b00000000000000010010101011010100;
assign LUT_3[38649] = 32'b00000000000000011001010110110001;
assign LUT_3[38650] = 32'b00000000000000010100110010111000;
assign LUT_3[38651] = 32'b00000000000000011011011110010101;
assign LUT_3[38652] = 32'b00000000000000001111111001001010;
assign LUT_3[38653] = 32'b00000000000000010110100100100111;
assign LUT_3[38654] = 32'b00000000000000010010000000101110;
assign LUT_3[38655] = 32'b00000000000000011000101100001011;
assign LUT_3[38656] = 32'b00000000000000000010111100100011;
assign LUT_3[38657] = 32'b00000000000000001001101000000000;
assign LUT_3[38658] = 32'b00000000000000000101000100000111;
assign LUT_3[38659] = 32'b00000000000000001011101111100100;
assign LUT_3[38660] = 32'b00000000000000000000001010011001;
assign LUT_3[38661] = 32'b00000000000000000110110101110110;
assign LUT_3[38662] = 32'b00000000000000000010010001111101;
assign LUT_3[38663] = 32'b00000000000000001000111101011010;
assign LUT_3[38664] = 32'b00000000000000001000010101101001;
assign LUT_3[38665] = 32'b00000000000000001111000001000110;
assign LUT_3[38666] = 32'b00000000000000001010011101001101;
assign LUT_3[38667] = 32'b00000000000000010001001000101010;
assign LUT_3[38668] = 32'b00000000000000000101100011011111;
assign LUT_3[38669] = 32'b00000000000000001100001110111100;
assign LUT_3[38670] = 32'b00000000000000000111101011000011;
assign LUT_3[38671] = 32'b00000000000000001110010110100000;
assign LUT_3[38672] = 32'b00000000000000000110001111100110;
assign LUT_3[38673] = 32'b00000000000000001100111011000011;
assign LUT_3[38674] = 32'b00000000000000001000010111001010;
assign LUT_3[38675] = 32'b00000000000000001111000010100111;
assign LUT_3[38676] = 32'b00000000000000000011011101011100;
assign LUT_3[38677] = 32'b00000000000000001010001000111001;
assign LUT_3[38678] = 32'b00000000000000000101100101000000;
assign LUT_3[38679] = 32'b00000000000000001100010000011101;
assign LUT_3[38680] = 32'b00000000000000001011101000101100;
assign LUT_3[38681] = 32'b00000000000000010010010100001001;
assign LUT_3[38682] = 32'b00000000000000001101110000010000;
assign LUT_3[38683] = 32'b00000000000000010100011011101101;
assign LUT_3[38684] = 32'b00000000000000001000110110100010;
assign LUT_3[38685] = 32'b00000000000000001111100001111111;
assign LUT_3[38686] = 32'b00000000000000001010111110000110;
assign LUT_3[38687] = 32'b00000000000000010001101001100011;
assign LUT_3[38688] = 32'b00000000000000000100001011000011;
assign LUT_3[38689] = 32'b00000000000000001010110110100000;
assign LUT_3[38690] = 32'b00000000000000000110010010100111;
assign LUT_3[38691] = 32'b00000000000000001100111110000100;
assign LUT_3[38692] = 32'b00000000000000000001011000111001;
assign LUT_3[38693] = 32'b00000000000000001000000100010110;
assign LUT_3[38694] = 32'b00000000000000000011100000011101;
assign LUT_3[38695] = 32'b00000000000000001010001011111010;
assign LUT_3[38696] = 32'b00000000000000001001100100001001;
assign LUT_3[38697] = 32'b00000000000000010000001111100110;
assign LUT_3[38698] = 32'b00000000000000001011101011101101;
assign LUT_3[38699] = 32'b00000000000000010010010111001010;
assign LUT_3[38700] = 32'b00000000000000000110110001111111;
assign LUT_3[38701] = 32'b00000000000000001101011101011100;
assign LUT_3[38702] = 32'b00000000000000001000111001100011;
assign LUT_3[38703] = 32'b00000000000000001111100101000000;
assign LUT_3[38704] = 32'b00000000000000000111011110000110;
assign LUT_3[38705] = 32'b00000000000000001110001001100011;
assign LUT_3[38706] = 32'b00000000000000001001100101101010;
assign LUT_3[38707] = 32'b00000000000000010000010001000111;
assign LUT_3[38708] = 32'b00000000000000000100101011111100;
assign LUT_3[38709] = 32'b00000000000000001011010111011001;
assign LUT_3[38710] = 32'b00000000000000000110110011100000;
assign LUT_3[38711] = 32'b00000000000000001101011110111101;
assign LUT_3[38712] = 32'b00000000000000001100110111001100;
assign LUT_3[38713] = 32'b00000000000000010011100010101001;
assign LUT_3[38714] = 32'b00000000000000001110111110110000;
assign LUT_3[38715] = 32'b00000000000000010101101010001101;
assign LUT_3[38716] = 32'b00000000000000001010000101000010;
assign LUT_3[38717] = 32'b00000000000000010000110000011111;
assign LUT_3[38718] = 32'b00000000000000001100001100100110;
assign LUT_3[38719] = 32'b00000000000000010010111000000011;
assign LUT_3[38720] = 32'b00000000000000000010110101001110;
assign LUT_3[38721] = 32'b00000000000000001001100000101011;
assign LUT_3[38722] = 32'b00000000000000000100111100110010;
assign LUT_3[38723] = 32'b00000000000000001011101000001111;
assign LUT_3[38724] = 32'b00000000000000000000000011000100;
assign LUT_3[38725] = 32'b00000000000000000110101110100001;
assign LUT_3[38726] = 32'b00000000000000000010001010101000;
assign LUT_3[38727] = 32'b00000000000000001000110110000101;
assign LUT_3[38728] = 32'b00000000000000001000001110010100;
assign LUT_3[38729] = 32'b00000000000000001110111001110001;
assign LUT_3[38730] = 32'b00000000000000001010010101111000;
assign LUT_3[38731] = 32'b00000000000000010001000001010101;
assign LUT_3[38732] = 32'b00000000000000000101011100001010;
assign LUT_3[38733] = 32'b00000000000000001100000111100111;
assign LUT_3[38734] = 32'b00000000000000000111100011101110;
assign LUT_3[38735] = 32'b00000000000000001110001111001011;
assign LUT_3[38736] = 32'b00000000000000000110001000010001;
assign LUT_3[38737] = 32'b00000000000000001100110011101110;
assign LUT_3[38738] = 32'b00000000000000001000001111110101;
assign LUT_3[38739] = 32'b00000000000000001110111011010010;
assign LUT_3[38740] = 32'b00000000000000000011010110000111;
assign LUT_3[38741] = 32'b00000000000000001010000001100100;
assign LUT_3[38742] = 32'b00000000000000000101011101101011;
assign LUT_3[38743] = 32'b00000000000000001100001001001000;
assign LUT_3[38744] = 32'b00000000000000001011100001010111;
assign LUT_3[38745] = 32'b00000000000000010010001100110100;
assign LUT_3[38746] = 32'b00000000000000001101101000111011;
assign LUT_3[38747] = 32'b00000000000000010100010100011000;
assign LUT_3[38748] = 32'b00000000000000001000101111001101;
assign LUT_3[38749] = 32'b00000000000000001111011010101010;
assign LUT_3[38750] = 32'b00000000000000001010110110110001;
assign LUT_3[38751] = 32'b00000000000000010001100010001110;
assign LUT_3[38752] = 32'b00000000000000000100000011101110;
assign LUT_3[38753] = 32'b00000000000000001010101111001011;
assign LUT_3[38754] = 32'b00000000000000000110001011010010;
assign LUT_3[38755] = 32'b00000000000000001100110110101111;
assign LUT_3[38756] = 32'b00000000000000000001010001100100;
assign LUT_3[38757] = 32'b00000000000000000111111101000001;
assign LUT_3[38758] = 32'b00000000000000000011011001001000;
assign LUT_3[38759] = 32'b00000000000000001010000100100101;
assign LUT_3[38760] = 32'b00000000000000001001011100110100;
assign LUT_3[38761] = 32'b00000000000000010000001000010001;
assign LUT_3[38762] = 32'b00000000000000001011100100011000;
assign LUT_3[38763] = 32'b00000000000000010010001111110101;
assign LUT_3[38764] = 32'b00000000000000000110101010101010;
assign LUT_3[38765] = 32'b00000000000000001101010110000111;
assign LUT_3[38766] = 32'b00000000000000001000110010001110;
assign LUT_3[38767] = 32'b00000000000000001111011101101011;
assign LUT_3[38768] = 32'b00000000000000000111010110110001;
assign LUT_3[38769] = 32'b00000000000000001110000010001110;
assign LUT_3[38770] = 32'b00000000000000001001011110010101;
assign LUT_3[38771] = 32'b00000000000000010000001001110010;
assign LUT_3[38772] = 32'b00000000000000000100100100100111;
assign LUT_3[38773] = 32'b00000000000000001011010000000100;
assign LUT_3[38774] = 32'b00000000000000000110101100001011;
assign LUT_3[38775] = 32'b00000000000000001101010111101000;
assign LUT_3[38776] = 32'b00000000000000001100101111110111;
assign LUT_3[38777] = 32'b00000000000000010011011011010100;
assign LUT_3[38778] = 32'b00000000000000001110110111011011;
assign LUT_3[38779] = 32'b00000000000000010101100010111000;
assign LUT_3[38780] = 32'b00000000000000001001111101101101;
assign LUT_3[38781] = 32'b00000000000000010000101001001010;
assign LUT_3[38782] = 32'b00000000000000001100000101010001;
assign LUT_3[38783] = 32'b00000000000000010010110000101110;
assign LUT_3[38784] = 32'b00000000000000000101000111100001;
assign LUT_3[38785] = 32'b00000000000000001011110010111110;
assign LUT_3[38786] = 32'b00000000000000000111001111000101;
assign LUT_3[38787] = 32'b00000000000000001101111010100010;
assign LUT_3[38788] = 32'b00000000000000000010010101010111;
assign LUT_3[38789] = 32'b00000000000000001001000000110100;
assign LUT_3[38790] = 32'b00000000000000000100011100111011;
assign LUT_3[38791] = 32'b00000000000000001011001000011000;
assign LUT_3[38792] = 32'b00000000000000001010100000100111;
assign LUT_3[38793] = 32'b00000000000000010001001100000100;
assign LUT_3[38794] = 32'b00000000000000001100101000001011;
assign LUT_3[38795] = 32'b00000000000000010011010011101000;
assign LUT_3[38796] = 32'b00000000000000000111101110011101;
assign LUT_3[38797] = 32'b00000000000000001110011001111010;
assign LUT_3[38798] = 32'b00000000000000001001110110000001;
assign LUT_3[38799] = 32'b00000000000000010000100001011110;
assign LUT_3[38800] = 32'b00000000000000001000011010100100;
assign LUT_3[38801] = 32'b00000000000000001111000110000001;
assign LUT_3[38802] = 32'b00000000000000001010100010001000;
assign LUT_3[38803] = 32'b00000000000000010001001101100101;
assign LUT_3[38804] = 32'b00000000000000000101101000011010;
assign LUT_3[38805] = 32'b00000000000000001100010011110111;
assign LUT_3[38806] = 32'b00000000000000000111101111111110;
assign LUT_3[38807] = 32'b00000000000000001110011011011011;
assign LUT_3[38808] = 32'b00000000000000001101110011101010;
assign LUT_3[38809] = 32'b00000000000000010100011111000111;
assign LUT_3[38810] = 32'b00000000000000001111111011001110;
assign LUT_3[38811] = 32'b00000000000000010110100110101011;
assign LUT_3[38812] = 32'b00000000000000001011000001100000;
assign LUT_3[38813] = 32'b00000000000000010001101100111101;
assign LUT_3[38814] = 32'b00000000000000001101001001000100;
assign LUT_3[38815] = 32'b00000000000000010011110100100001;
assign LUT_3[38816] = 32'b00000000000000000110010110000001;
assign LUT_3[38817] = 32'b00000000000000001101000001011110;
assign LUT_3[38818] = 32'b00000000000000001000011101100101;
assign LUT_3[38819] = 32'b00000000000000001111001001000010;
assign LUT_3[38820] = 32'b00000000000000000011100011110111;
assign LUT_3[38821] = 32'b00000000000000001010001111010100;
assign LUT_3[38822] = 32'b00000000000000000101101011011011;
assign LUT_3[38823] = 32'b00000000000000001100010110111000;
assign LUT_3[38824] = 32'b00000000000000001011101111000111;
assign LUT_3[38825] = 32'b00000000000000010010011010100100;
assign LUT_3[38826] = 32'b00000000000000001101110110101011;
assign LUT_3[38827] = 32'b00000000000000010100100010001000;
assign LUT_3[38828] = 32'b00000000000000001000111100111101;
assign LUT_3[38829] = 32'b00000000000000001111101000011010;
assign LUT_3[38830] = 32'b00000000000000001011000100100001;
assign LUT_3[38831] = 32'b00000000000000010001101111111110;
assign LUT_3[38832] = 32'b00000000000000001001101001000100;
assign LUT_3[38833] = 32'b00000000000000010000010100100001;
assign LUT_3[38834] = 32'b00000000000000001011110000101000;
assign LUT_3[38835] = 32'b00000000000000010010011100000101;
assign LUT_3[38836] = 32'b00000000000000000110110110111010;
assign LUT_3[38837] = 32'b00000000000000001101100010010111;
assign LUT_3[38838] = 32'b00000000000000001000111110011110;
assign LUT_3[38839] = 32'b00000000000000001111101001111011;
assign LUT_3[38840] = 32'b00000000000000001111000010001010;
assign LUT_3[38841] = 32'b00000000000000010101101101100111;
assign LUT_3[38842] = 32'b00000000000000010001001001101110;
assign LUT_3[38843] = 32'b00000000000000010111110101001011;
assign LUT_3[38844] = 32'b00000000000000001100010000000000;
assign LUT_3[38845] = 32'b00000000000000010010111011011101;
assign LUT_3[38846] = 32'b00000000000000001110010111100100;
assign LUT_3[38847] = 32'b00000000000000010101000011000001;
assign LUT_3[38848] = 32'b00000000000000000101000000001100;
assign LUT_3[38849] = 32'b00000000000000001011101011101001;
assign LUT_3[38850] = 32'b00000000000000000111000111110000;
assign LUT_3[38851] = 32'b00000000000000001101110011001101;
assign LUT_3[38852] = 32'b00000000000000000010001110000010;
assign LUT_3[38853] = 32'b00000000000000001000111001011111;
assign LUT_3[38854] = 32'b00000000000000000100010101100110;
assign LUT_3[38855] = 32'b00000000000000001011000001000011;
assign LUT_3[38856] = 32'b00000000000000001010011001010010;
assign LUT_3[38857] = 32'b00000000000000010001000100101111;
assign LUT_3[38858] = 32'b00000000000000001100100000110110;
assign LUT_3[38859] = 32'b00000000000000010011001100010011;
assign LUT_3[38860] = 32'b00000000000000000111100111001000;
assign LUT_3[38861] = 32'b00000000000000001110010010100101;
assign LUT_3[38862] = 32'b00000000000000001001101110101100;
assign LUT_3[38863] = 32'b00000000000000010000011010001001;
assign LUT_3[38864] = 32'b00000000000000001000010011001111;
assign LUT_3[38865] = 32'b00000000000000001110111110101100;
assign LUT_3[38866] = 32'b00000000000000001010011010110011;
assign LUT_3[38867] = 32'b00000000000000010001000110010000;
assign LUT_3[38868] = 32'b00000000000000000101100001000101;
assign LUT_3[38869] = 32'b00000000000000001100001100100010;
assign LUT_3[38870] = 32'b00000000000000000111101000101001;
assign LUT_3[38871] = 32'b00000000000000001110010100000110;
assign LUT_3[38872] = 32'b00000000000000001101101100010101;
assign LUT_3[38873] = 32'b00000000000000010100010111110010;
assign LUT_3[38874] = 32'b00000000000000001111110011111001;
assign LUT_3[38875] = 32'b00000000000000010110011111010110;
assign LUT_3[38876] = 32'b00000000000000001010111010001011;
assign LUT_3[38877] = 32'b00000000000000010001100101101000;
assign LUT_3[38878] = 32'b00000000000000001101000001101111;
assign LUT_3[38879] = 32'b00000000000000010011101101001100;
assign LUT_3[38880] = 32'b00000000000000000110001110101100;
assign LUT_3[38881] = 32'b00000000000000001100111010001001;
assign LUT_3[38882] = 32'b00000000000000001000010110010000;
assign LUT_3[38883] = 32'b00000000000000001111000001101101;
assign LUT_3[38884] = 32'b00000000000000000011011100100010;
assign LUT_3[38885] = 32'b00000000000000001010000111111111;
assign LUT_3[38886] = 32'b00000000000000000101100100000110;
assign LUT_3[38887] = 32'b00000000000000001100001111100011;
assign LUT_3[38888] = 32'b00000000000000001011100111110010;
assign LUT_3[38889] = 32'b00000000000000010010010011001111;
assign LUT_3[38890] = 32'b00000000000000001101101111010110;
assign LUT_3[38891] = 32'b00000000000000010100011010110011;
assign LUT_3[38892] = 32'b00000000000000001000110101101000;
assign LUT_3[38893] = 32'b00000000000000001111100001000101;
assign LUT_3[38894] = 32'b00000000000000001010111101001100;
assign LUT_3[38895] = 32'b00000000000000010001101000101001;
assign LUT_3[38896] = 32'b00000000000000001001100001101111;
assign LUT_3[38897] = 32'b00000000000000010000001101001100;
assign LUT_3[38898] = 32'b00000000000000001011101001010011;
assign LUT_3[38899] = 32'b00000000000000010010010100110000;
assign LUT_3[38900] = 32'b00000000000000000110101111100101;
assign LUT_3[38901] = 32'b00000000000000001101011011000010;
assign LUT_3[38902] = 32'b00000000000000001000110111001001;
assign LUT_3[38903] = 32'b00000000000000001111100010100110;
assign LUT_3[38904] = 32'b00000000000000001110111010110101;
assign LUT_3[38905] = 32'b00000000000000010101100110010010;
assign LUT_3[38906] = 32'b00000000000000010001000010011001;
assign LUT_3[38907] = 32'b00000000000000010111101101110110;
assign LUT_3[38908] = 32'b00000000000000001100001000101011;
assign LUT_3[38909] = 32'b00000000000000010010110100001000;
assign LUT_3[38910] = 32'b00000000000000001110010000001111;
assign LUT_3[38911] = 32'b00000000000000010100111011101100;
assign LUT_3[38912] = 32'b11111111111111111110101001000111;
assign LUT_3[38913] = 32'b00000000000000000101010100100100;
assign LUT_3[38914] = 32'b00000000000000000000110000101011;
assign LUT_3[38915] = 32'b00000000000000000111011100001000;
assign LUT_3[38916] = 32'b11111111111111111011110110111101;
assign LUT_3[38917] = 32'b00000000000000000010100010011010;
assign LUT_3[38918] = 32'b11111111111111111101111110100001;
assign LUT_3[38919] = 32'b00000000000000000100101001111110;
assign LUT_3[38920] = 32'b00000000000000000100000010001101;
assign LUT_3[38921] = 32'b00000000000000001010101101101010;
assign LUT_3[38922] = 32'b00000000000000000110001001110001;
assign LUT_3[38923] = 32'b00000000000000001100110101001110;
assign LUT_3[38924] = 32'b00000000000000000001010000000011;
assign LUT_3[38925] = 32'b00000000000000000111111011100000;
assign LUT_3[38926] = 32'b00000000000000000011010111100111;
assign LUT_3[38927] = 32'b00000000000000001010000011000100;
assign LUT_3[38928] = 32'b00000000000000000001111100001010;
assign LUT_3[38929] = 32'b00000000000000001000100111100111;
assign LUT_3[38930] = 32'b00000000000000000100000011101110;
assign LUT_3[38931] = 32'b00000000000000001010101111001011;
assign LUT_3[38932] = 32'b11111111111111111111001010000000;
assign LUT_3[38933] = 32'b00000000000000000101110101011101;
assign LUT_3[38934] = 32'b00000000000000000001010001100100;
assign LUT_3[38935] = 32'b00000000000000000111111101000001;
assign LUT_3[38936] = 32'b00000000000000000111010101010000;
assign LUT_3[38937] = 32'b00000000000000001110000000101101;
assign LUT_3[38938] = 32'b00000000000000001001011100110100;
assign LUT_3[38939] = 32'b00000000000000010000001000010001;
assign LUT_3[38940] = 32'b00000000000000000100100011000110;
assign LUT_3[38941] = 32'b00000000000000001011001110100011;
assign LUT_3[38942] = 32'b00000000000000000110101010101010;
assign LUT_3[38943] = 32'b00000000000000001101010110000111;
assign LUT_3[38944] = 32'b11111111111111111111110111100111;
assign LUT_3[38945] = 32'b00000000000000000110100011000100;
assign LUT_3[38946] = 32'b00000000000000000001111111001011;
assign LUT_3[38947] = 32'b00000000000000001000101010101000;
assign LUT_3[38948] = 32'b11111111111111111101000101011101;
assign LUT_3[38949] = 32'b00000000000000000011110000111010;
assign LUT_3[38950] = 32'b11111111111111111111001101000001;
assign LUT_3[38951] = 32'b00000000000000000101111000011110;
assign LUT_3[38952] = 32'b00000000000000000101010000101101;
assign LUT_3[38953] = 32'b00000000000000001011111100001010;
assign LUT_3[38954] = 32'b00000000000000000111011000010001;
assign LUT_3[38955] = 32'b00000000000000001110000011101110;
assign LUT_3[38956] = 32'b00000000000000000010011110100011;
assign LUT_3[38957] = 32'b00000000000000001001001010000000;
assign LUT_3[38958] = 32'b00000000000000000100100110000111;
assign LUT_3[38959] = 32'b00000000000000001011010001100100;
assign LUT_3[38960] = 32'b00000000000000000011001010101010;
assign LUT_3[38961] = 32'b00000000000000001001110110000111;
assign LUT_3[38962] = 32'b00000000000000000101010010001110;
assign LUT_3[38963] = 32'b00000000000000001011111101101011;
assign LUT_3[38964] = 32'b00000000000000000000011000100000;
assign LUT_3[38965] = 32'b00000000000000000111000011111101;
assign LUT_3[38966] = 32'b00000000000000000010100000000100;
assign LUT_3[38967] = 32'b00000000000000001001001011100001;
assign LUT_3[38968] = 32'b00000000000000001000100011110000;
assign LUT_3[38969] = 32'b00000000000000001111001111001101;
assign LUT_3[38970] = 32'b00000000000000001010101011010100;
assign LUT_3[38971] = 32'b00000000000000010001010110110001;
assign LUT_3[38972] = 32'b00000000000000000101110001100110;
assign LUT_3[38973] = 32'b00000000000000001100011101000011;
assign LUT_3[38974] = 32'b00000000000000000111111001001010;
assign LUT_3[38975] = 32'b00000000000000001110100100100111;
assign LUT_3[38976] = 32'b11111111111111111110100001110010;
assign LUT_3[38977] = 32'b00000000000000000101001101001111;
assign LUT_3[38978] = 32'b00000000000000000000101001010110;
assign LUT_3[38979] = 32'b00000000000000000111010100110011;
assign LUT_3[38980] = 32'b11111111111111111011101111101000;
assign LUT_3[38981] = 32'b00000000000000000010011011000101;
assign LUT_3[38982] = 32'b11111111111111111101110111001100;
assign LUT_3[38983] = 32'b00000000000000000100100010101001;
assign LUT_3[38984] = 32'b00000000000000000011111010111000;
assign LUT_3[38985] = 32'b00000000000000001010100110010101;
assign LUT_3[38986] = 32'b00000000000000000110000010011100;
assign LUT_3[38987] = 32'b00000000000000001100101101111001;
assign LUT_3[38988] = 32'b00000000000000000001001000101110;
assign LUT_3[38989] = 32'b00000000000000000111110100001011;
assign LUT_3[38990] = 32'b00000000000000000011010000010010;
assign LUT_3[38991] = 32'b00000000000000001001111011101111;
assign LUT_3[38992] = 32'b00000000000000000001110100110101;
assign LUT_3[38993] = 32'b00000000000000001000100000010010;
assign LUT_3[38994] = 32'b00000000000000000011111100011001;
assign LUT_3[38995] = 32'b00000000000000001010100111110110;
assign LUT_3[38996] = 32'b11111111111111111111000010101011;
assign LUT_3[38997] = 32'b00000000000000000101101110001000;
assign LUT_3[38998] = 32'b00000000000000000001001010001111;
assign LUT_3[38999] = 32'b00000000000000000111110101101100;
assign LUT_3[39000] = 32'b00000000000000000111001101111011;
assign LUT_3[39001] = 32'b00000000000000001101111001011000;
assign LUT_3[39002] = 32'b00000000000000001001010101011111;
assign LUT_3[39003] = 32'b00000000000000010000000000111100;
assign LUT_3[39004] = 32'b00000000000000000100011011110001;
assign LUT_3[39005] = 32'b00000000000000001011000111001110;
assign LUT_3[39006] = 32'b00000000000000000110100011010101;
assign LUT_3[39007] = 32'b00000000000000001101001110110010;
assign LUT_3[39008] = 32'b11111111111111111111110000010010;
assign LUT_3[39009] = 32'b00000000000000000110011011101111;
assign LUT_3[39010] = 32'b00000000000000000001110111110110;
assign LUT_3[39011] = 32'b00000000000000001000100011010011;
assign LUT_3[39012] = 32'b11111111111111111100111110001000;
assign LUT_3[39013] = 32'b00000000000000000011101001100101;
assign LUT_3[39014] = 32'b11111111111111111111000101101100;
assign LUT_3[39015] = 32'b00000000000000000101110001001001;
assign LUT_3[39016] = 32'b00000000000000000101001001011000;
assign LUT_3[39017] = 32'b00000000000000001011110100110101;
assign LUT_3[39018] = 32'b00000000000000000111010000111100;
assign LUT_3[39019] = 32'b00000000000000001101111100011001;
assign LUT_3[39020] = 32'b00000000000000000010010111001110;
assign LUT_3[39021] = 32'b00000000000000001001000010101011;
assign LUT_3[39022] = 32'b00000000000000000100011110110010;
assign LUT_3[39023] = 32'b00000000000000001011001010001111;
assign LUT_3[39024] = 32'b00000000000000000011000011010101;
assign LUT_3[39025] = 32'b00000000000000001001101110110010;
assign LUT_3[39026] = 32'b00000000000000000101001010111001;
assign LUT_3[39027] = 32'b00000000000000001011110110010110;
assign LUT_3[39028] = 32'b00000000000000000000010001001011;
assign LUT_3[39029] = 32'b00000000000000000110111100101000;
assign LUT_3[39030] = 32'b00000000000000000010011000101111;
assign LUT_3[39031] = 32'b00000000000000001001000100001100;
assign LUT_3[39032] = 32'b00000000000000001000011100011011;
assign LUT_3[39033] = 32'b00000000000000001111000111111000;
assign LUT_3[39034] = 32'b00000000000000001010100011111111;
assign LUT_3[39035] = 32'b00000000000000010001001111011100;
assign LUT_3[39036] = 32'b00000000000000000101101010010001;
assign LUT_3[39037] = 32'b00000000000000001100010101101110;
assign LUT_3[39038] = 32'b00000000000000000111110001110101;
assign LUT_3[39039] = 32'b00000000000000001110011101010010;
assign LUT_3[39040] = 32'b00000000000000000000110100000101;
assign LUT_3[39041] = 32'b00000000000000000111011111100010;
assign LUT_3[39042] = 32'b00000000000000000010111011101001;
assign LUT_3[39043] = 32'b00000000000000001001100111000110;
assign LUT_3[39044] = 32'b11111111111111111110000001111011;
assign LUT_3[39045] = 32'b00000000000000000100101101011000;
assign LUT_3[39046] = 32'b00000000000000000000001001011111;
assign LUT_3[39047] = 32'b00000000000000000110110100111100;
assign LUT_3[39048] = 32'b00000000000000000110001101001011;
assign LUT_3[39049] = 32'b00000000000000001100111000101000;
assign LUT_3[39050] = 32'b00000000000000001000010100101111;
assign LUT_3[39051] = 32'b00000000000000001111000000001100;
assign LUT_3[39052] = 32'b00000000000000000011011011000001;
assign LUT_3[39053] = 32'b00000000000000001010000110011110;
assign LUT_3[39054] = 32'b00000000000000000101100010100101;
assign LUT_3[39055] = 32'b00000000000000001100001110000010;
assign LUT_3[39056] = 32'b00000000000000000100000111001000;
assign LUT_3[39057] = 32'b00000000000000001010110010100101;
assign LUT_3[39058] = 32'b00000000000000000110001110101100;
assign LUT_3[39059] = 32'b00000000000000001100111010001001;
assign LUT_3[39060] = 32'b00000000000000000001010100111110;
assign LUT_3[39061] = 32'b00000000000000001000000000011011;
assign LUT_3[39062] = 32'b00000000000000000011011100100010;
assign LUT_3[39063] = 32'b00000000000000001010000111111111;
assign LUT_3[39064] = 32'b00000000000000001001100000001110;
assign LUT_3[39065] = 32'b00000000000000010000001011101011;
assign LUT_3[39066] = 32'b00000000000000001011100111110010;
assign LUT_3[39067] = 32'b00000000000000010010010011001111;
assign LUT_3[39068] = 32'b00000000000000000110101110000100;
assign LUT_3[39069] = 32'b00000000000000001101011001100001;
assign LUT_3[39070] = 32'b00000000000000001000110101101000;
assign LUT_3[39071] = 32'b00000000000000001111100001000101;
assign LUT_3[39072] = 32'b00000000000000000010000010100101;
assign LUT_3[39073] = 32'b00000000000000001000101110000010;
assign LUT_3[39074] = 32'b00000000000000000100001010001001;
assign LUT_3[39075] = 32'b00000000000000001010110101100110;
assign LUT_3[39076] = 32'b11111111111111111111010000011011;
assign LUT_3[39077] = 32'b00000000000000000101111011111000;
assign LUT_3[39078] = 32'b00000000000000000001010111111111;
assign LUT_3[39079] = 32'b00000000000000001000000011011100;
assign LUT_3[39080] = 32'b00000000000000000111011011101011;
assign LUT_3[39081] = 32'b00000000000000001110000111001000;
assign LUT_3[39082] = 32'b00000000000000001001100011001111;
assign LUT_3[39083] = 32'b00000000000000010000001110101100;
assign LUT_3[39084] = 32'b00000000000000000100101001100001;
assign LUT_3[39085] = 32'b00000000000000001011010100111110;
assign LUT_3[39086] = 32'b00000000000000000110110001000101;
assign LUT_3[39087] = 32'b00000000000000001101011100100010;
assign LUT_3[39088] = 32'b00000000000000000101010101101000;
assign LUT_3[39089] = 32'b00000000000000001100000001000101;
assign LUT_3[39090] = 32'b00000000000000000111011101001100;
assign LUT_3[39091] = 32'b00000000000000001110001000101001;
assign LUT_3[39092] = 32'b00000000000000000010100011011110;
assign LUT_3[39093] = 32'b00000000000000001001001110111011;
assign LUT_3[39094] = 32'b00000000000000000100101011000010;
assign LUT_3[39095] = 32'b00000000000000001011010110011111;
assign LUT_3[39096] = 32'b00000000000000001010101110101110;
assign LUT_3[39097] = 32'b00000000000000010001011010001011;
assign LUT_3[39098] = 32'b00000000000000001100110110010010;
assign LUT_3[39099] = 32'b00000000000000010011100001101111;
assign LUT_3[39100] = 32'b00000000000000000111111100100100;
assign LUT_3[39101] = 32'b00000000000000001110101000000001;
assign LUT_3[39102] = 32'b00000000000000001010000100001000;
assign LUT_3[39103] = 32'b00000000000000010000101111100101;
assign LUT_3[39104] = 32'b00000000000000000000101100110000;
assign LUT_3[39105] = 32'b00000000000000000111011000001101;
assign LUT_3[39106] = 32'b00000000000000000010110100010100;
assign LUT_3[39107] = 32'b00000000000000001001011111110001;
assign LUT_3[39108] = 32'b11111111111111111101111010100110;
assign LUT_3[39109] = 32'b00000000000000000100100110000011;
assign LUT_3[39110] = 32'b00000000000000000000000010001010;
assign LUT_3[39111] = 32'b00000000000000000110101101100111;
assign LUT_3[39112] = 32'b00000000000000000110000101110110;
assign LUT_3[39113] = 32'b00000000000000001100110001010011;
assign LUT_3[39114] = 32'b00000000000000001000001101011010;
assign LUT_3[39115] = 32'b00000000000000001110111000110111;
assign LUT_3[39116] = 32'b00000000000000000011010011101100;
assign LUT_3[39117] = 32'b00000000000000001001111111001001;
assign LUT_3[39118] = 32'b00000000000000000101011011010000;
assign LUT_3[39119] = 32'b00000000000000001100000110101101;
assign LUT_3[39120] = 32'b00000000000000000011111111110011;
assign LUT_3[39121] = 32'b00000000000000001010101011010000;
assign LUT_3[39122] = 32'b00000000000000000110000111010111;
assign LUT_3[39123] = 32'b00000000000000001100110010110100;
assign LUT_3[39124] = 32'b00000000000000000001001101101001;
assign LUT_3[39125] = 32'b00000000000000000111111001000110;
assign LUT_3[39126] = 32'b00000000000000000011010101001101;
assign LUT_3[39127] = 32'b00000000000000001010000000101010;
assign LUT_3[39128] = 32'b00000000000000001001011000111001;
assign LUT_3[39129] = 32'b00000000000000010000000100010110;
assign LUT_3[39130] = 32'b00000000000000001011100000011101;
assign LUT_3[39131] = 32'b00000000000000010010001011111010;
assign LUT_3[39132] = 32'b00000000000000000110100110101111;
assign LUT_3[39133] = 32'b00000000000000001101010010001100;
assign LUT_3[39134] = 32'b00000000000000001000101110010011;
assign LUT_3[39135] = 32'b00000000000000001111011001110000;
assign LUT_3[39136] = 32'b00000000000000000001111011010000;
assign LUT_3[39137] = 32'b00000000000000001000100110101101;
assign LUT_3[39138] = 32'b00000000000000000100000010110100;
assign LUT_3[39139] = 32'b00000000000000001010101110010001;
assign LUT_3[39140] = 32'b11111111111111111111001001000110;
assign LUT_3[39141] = 32'b00000000000000000101110100100011;
assign LUT_3[39142] = 32'b00000000000000000001010000101010;
assign LUT_3[39143] = 32'b00000000000000000111111100000111;
assign LUT_3[39144] = 32'b00000000000000000111010100010110;
assign LUT_3[39145] = 32'b00000000000000001101111111110011;
assign LUT_3[39146] = 32'b00000000000000001001011011111010;
assign LUT_3[39147] = 32'b00000000000000010000000111010111;
assign LUT_3[39148] = 32'b00000000000000000100100010001100;
assign LUT_3[39149] = 32'b00000000000000001011001101101001;
assign LUT_3[39150] = 32'b00000000000000000110101001110000;
assign LUT_3[39151] = 32'b00000000000000001101010101001101;
assign LUT_3[39152] = 32'b00000000000000000101001110010011;
assign LUT_3[39153] = 32'b00000000000000001011111001110000;
assign LUT_3[39154] = 32'b00000000000000000111010101110111;
assign LUT_3[39155] = 32'b00000000000000001110000001010100;
assign LUT_3[39156] = 32'b00000000000000000010011100001001;
assign LUT_3[39157] = 32'b00000000000000001001000111100110;
assign LUT_3[39158] = 32'b00000000000000000100100011101101;
assign LUT_3[39159] = 32'b00000000000000001011001111001010;
assign LUT_3[39160] = 32'b00000000000000001010100111011001;
assign LUT_3[39161] = 32'b00000000000000010001010010110110;
assign LUT_3[39162] = 32'b00000000000000001100101110111101;
assign LUT_3[39163] = 32'b00000000000000010011011010011010;
assign LUT_3[39164] = 32'b00000000000000000111110101001111;
assign LUT_3[39165] = 32'b00000000000000001110100000101100;
assign LUT_3[39166] = 32'b00000000000000001001111100110011;
assign LUT_3[39167] = 32'b00000000000000010000101000010000;
assign LUT_3[39168] = 32'b11111111111111111010111000101000;
assign LUT_3[39169] = 32'b00000000000000000001100100000101;
assign LUT_3[39170] = 32'b11111111111111111101000000001100;
assign LUT_3[39171] = 32'b00000000000000000011101011101001;
assign LUT_3[39172] = 32'b11111111111111111000000110011110;
assign LUT_3[39173] = 32'b11111111111111111110110001111011;
assign LUT_3[39174] = 32'b11111111111111111010001110000010;
assign LUT_3[39175] = 32'b00000000000000000000111001011111;
assign LUT_3[39176] = 32'b00000000000000000000010001101110;
assign LUT_3[39177] = 32'b00000000000000000110111101001011;
assign LUT_3[39178] = 32'b00000000000000000010011001010010;
assign LUT_3[39179] = 32'b00000000000000001001000100101111;
assign LUT_3[39180] = 32'b11111111111111111101011111100100;
assign LUT_3[39181] = 32'b00000000000000000100001011000001;
assign LUT_3[39182] = 32'b11111111111111111111100111001000;
assign LUT_3[39183] = 32'b00000000000000000110010010100101;
assign LUT_3[39184] = 32'b11111111111111111110001011101011;
assign LUT_3[39185] = 32'b00000000000000000100110111001000;
assign LUT_3[39186] = 32'b00000000000000000000010011001111;
assign LUT_3[39187] = 32'b00000000000000000110111110101100;
assign LUT_3[39188] = 32'b11111111111111111011011001100001;
assign LUT_3[39189] = 32'b00000000000000000010000100111110;
assign LUT_3[39190] = 32'b11111111111111111101100001000101;
assign LUT_3[39191] = 32'b00000000000000000100001100100010;
assign LUT_3[39192] = 32'b00000000000000000011100100110001;
assign LUT_3[39193] = 32'b00000000000000001010010000001110;
assign LUT_3[39194] = 32'b00000000000000000101101100010101;
assign LUT_3[39195] = 32'b00000000000000001100010111110010;
assign LUT_3[39196] = 32'b00000000000000000000110010100111;
assign LUT_3[39197] = 32'b00000000000000000111011110000100;
assign LUT_3[39198] = 32'b00000000000000000010111010001011;
assign LUT_3[39199] = 32'b00000000000000001001100101101000;
assign LUT_3[39200] = 32'b11111111111111111100000111001000;
assign LUT_3[39201] = 32'b00000000000000000010110010100101;
assign LUT_3[39202] = 32'b11111111111111111110001110101100;
assign LUT_3[39203] = 32'b00000000000000000100111010001001;
assign LUT_3[39204] = 32'b11111111111111111001010100111110;
assign LUT_3[39205] = 32'b00000000000000000000000000011011;
assign LUT_3[39206] = 32'b11111111111111111011011100100010;
assign LUT_3[39207] = 32'b00000000000000000010000111111111;
assign LUT_3[39208] = 32'b00000000000000000001100000001110;
assign LUT_3[39209] = 32'b00000000000000001000001011101011;
assign LUT_3[39210] = 32'b00000000000000000011100111110010;
assign LUT_3[39211] = 32'b00000000000000001010010011001111;
assign LUT_3[39212] = 32'b11111111111111111110101110000100;
assign LUT_3[39213] = 32'b00000000000000000101011001100001;
assign LUT_3[39214] = 32'b00000000000000000000110101101000;
assign LUT_3[39215] = 32'b00000000000000000111100001000101;
assign LUT_3[39216] = 32'b11111111111111111111011010001011;
assign LUT_3[39217] = 32'b00000000000000000110000101101000;
assign LUT_3[39218] = 32'b00000000000000000001100001101111;
assign LUT_3[39219] = 32'b00000000000000001000001101001100;
assign LUT_3[39220] = 32'b11111111111111111100101000000001;
assign LUT_3[39221] = 32'b00000000000000000011010011011110;
assign LUT_3[39222] = 32'b11111111111111111110101111100101;
assign LUT_3[39223] = 32'b00000000000000000101011011000010;
assign LUT_3[39224] = 32'b00000000000000000100110011010001;
assign LUT_3[39225] = 32'b00000000000000001011011110101110;
assign LUT_3[39226] = 32'b00000000000000000110111010110101;
assign LUT_3[39227] = 32'b00000000000000001101100110010010;
assign LUT_3[39228] = 32'b00000000000000000010000001000111;
assign LUT_3[39229] = 32'b00000000000000001000101100100100;
assign LUT_3[39230] = 32'b00000000000000000100001000101011;
assign LUT_3[39231] = 32'b00000000000000001010110100001000;
assign LUT_3[39232] = 32'b11111111111111111010110001010011;
assign LUT_3[39233] = 32'b00000000000000000001011100110000;
assign LUT_3[39234] = 32'b11111111111111111100111000110111;
assign LUT_3[39235] = 32'b00000000000000000011100100010100;
assign LUT_3[39236] = 32'b11111111111111110111111111001001;
assign LUT_3[39237] = 32'b11111111111111111110101010100110;
assign LUT_3[39238] = 32'b11111111111111111010000110101101;
assign LUT_3[39239] = 32'b00000000000000000000110010001010;
assign LUT_3[39240] = 32'b00000000000000000000001010011001;
assign LUT_3[39241] = 32'b00000000000000000110110101110110;
assign LUT_3[39242] = 32'b00000000000000000010010001111101;
assign LUT_3[39243] = 32'b00000000000000001000111101011010;
assign LUT_3[39244] = 32'b11111111111111111101011000001111;
assign LUT_3[39245] = 32'b00000000000000000100000011101100;
assign LUT_3[39246] = 32'b11111111111111111111011111110011;
assign LUT_3[39247] = 32'b00000000000000000110001011010000;
assign LUT_3[39248] = 32'b11111111111111111110000100010110;
assign LUT_3[39249] = 32'b00000000000000000100101111110011;
assign LUT_3[39250] = 32'b00000000000000000000001011111010;
assign LUT_3[39251] = 32'b00000000000000000110110111010111;
assign LUT_3[39252] = 32'b11111111111111111011010010001100;
assign LUT_3[39253] = 32'b00000000000000000001111101101001;
assign LUT_3[39254] = 32'b11111111111111111101011001110000;
assign LUT_3[39255] = 32'b00000000000000000100000101001101;
assign LUT_3[39256] = 32'b00000000000000000011011101011100;
assign LUT_3[39257] = 32'b00000000000000001010001000111001;
assign LUT_3[39258] = 32'b00000000000000000101100101000000;
assign LUT_3[39259] = 32'b00000000000000001100010000011101;
assign LUT_3[39260] = 32'b00000000000000000000101011010010;
assign LUT_3[39261] = 32'b00000000000000000111010110101111;
assign LUT_3[39262] = 32'b00000000000000000010110010110110;
assign LUT_3[39263] = 32'b00000000000000001001011110010011;
assign LUT_3[39264] = 32'b11111111111111111011111111110011;
assign LUT_3[39265] = 32'b00000000000000000010101011010000;
assign LUT_3[39266] = 32'b11111111111111111110000111010111;
assign LUT_3[39267] = 32'b00000000000000000100110010110100;
assign LUT_3[39268] = 32'b11111111111111111001001101101001;
assign LUT_3[39269] = 32'b11111111111111111111111001000110;
assign LUT_3[39270] = 32'b11111111111111111011010101001101;
assign LUT_3[39271] = 32'b00000000000000000010000000101010;
assign LUT_3[39272] = 32'b00000000000000000001011000111001;
assign LUT_3[39273] = 32'b00000000000000001000000100010110;
assign LUT_3[39274] = 32'b00000000000000000011100000011101;
assign LUT_3[39275] = 32'b00000000000000001010001011111010;
assign LUT_3[39276] = 32'b11111111111111111110100110101111;
assign LUT_3[39277] = 32'b00000000000000000101010010001100;
assign LUT_3[39278] = 32'b00000000000000000000101110010011;
assign LUT_3[39279] = 32'b00000000000000000111011001110000;
assign LUT_3[39280] = 32'b11111111111111111111010010110110;
assign LUT_3[39281] = 32'b00000000000000000101111110010011;
assign LUT_3[39282] = 32'b00000000000000000001011010011010;
assign LUT_3[39283] = 32'b00000000000000001000000101110111;
assign LUT_3[39284] = 32'b11111111111111111100100000101100;
assign LUT_3[39285] = 32'b00000000000000000011001100001001;
assign LUT_3[39286] = 32'b11111111111111111110101000010000;
assign LUT_3[39287] = 32'b00000000000000000101010011101101;
assign LUT_3[39288] = 32'b00000000000000000100101011111100;
assign LUT_3[39289] = 32'b00000000000000001011010111011001;
assign LUT_3[39290] = 32'b00000000000000000110110011100000;
assign LUT_3[39291] = 32'b00000000000000001101011110111101;
assign LUT_3[39292] = 32'b00000000000000000001111001110010;
assign LUT_3[39293] = 32'b00000000000000001000100101001111;
assign LUT_3[39294] = 32'b00000000000000000100000001010110;
assign LUT_3[39295] = 32'b00000000000000001010101100110011;
assign LUT_3[39296] = 32'b11111111111111111101000011100110;
assign LUT_3[39297] = 32'b00000000000000000011101111000011;
assign LUT_3[39298] = 32'b11111111111111111111001011001010;
assign LUT_3[39299] = 32'b00000000000000000101110110100111;
assign LUT_3[39300] = 32'b11111111111111111010010001011100;
assign LUT_3[39301] = 32'b00000000000000000000111100111001;
assign LUT_3[39302] = 32'b11111111111111111100011001000000;
assign LUT_3[39303] = 32'b00000000000000000011000100011101;
assign LUT_3[39304] = 32'b00000000000000000010011100101100;
assign LUT_3[39305] = 32'b00000000000000001001001000001001;
assign LUT_3[39306] = 32'b00000000000000000100100100010000;
assign LUT_3[39307] = 32'b00000000000000001011001111101101;
assign LUT_3[39308] = 32'b11111111111111111111101010100010;
assign LUT_3[39309] = 32'b00000000000000000110010101111111;
assign LUT_3[39310] = 32'b00000000000000000001110010000110;
assign LUT_3[39311] = 32'b00000000000000001000011101100011;
assign LUT_3[39312] = 32'b00000000000000000000010110101001;
assign LUT_3[39313] = 32'b00000000000000000111000010000110;
assign LUT_3[39314] = 32'b00000000000000000010011110001101;
assign LUT_3[39315] = 32'b00000000000000001001001001101010;
assign LUT_3[39316] = 32'b11111111111111111101100100011111;
assign LUT_3[39317] = 32'b00000000000000000100001111111100;
assign LUT_3[39318] = 32'b11111111111111111111101100000011;
assign LUT_3[39319] = 32'b00000000000000000110010111100000;
assign LUT_3[39320] = 32'b00000000000000000101101111101111;
assign LUT_3[39321] = 32'b00000000000000001100011011001100;
assign LUT_3[39322] = 32'b00000000000000000111110111010011;
assign LUT_3[39323] = 32'b00000000000000001110100010110000;
assign LUT_3[39324] = 32'b00000000000000000010111101100101;
assign LUT_3[39325] = 32'b00000000000000001001101001000010;
assign LUT_3[39326] = 32'b00000000000000000101000101001001;
assign LUT_3[39327] = 32'b00000000000000001011110000100110;
assign LUT_3[39328] = 32'b11111111111111111110010010000110;
assign LUT_3[39329] = 32'b00000000000000000100111101100011;
assign LUT_3[39330] = 32'b00000000000000000000011001101010;
assign LUT_3[39331] = 32'b00000000000000000111000101000111;
assign LUT_3[39332] = 32'b11111111111111111011011111111100;
assign LUT_3[39333] = 32'b00000000000000000010001011011001;
assign LUT_3[39334] = 32'b11111111111111111101100111100000;
assign LUT_3[39335] = 32'b00000000000000000100010010111101;
assign LUT_3[39336] = 32'b00000000000000000011101011001100;
assign LUT_3[39337] = 32'b00000000000000001010010110101001;
assign LUT_3[39338] = 32'b00000000000000000101110010110000;
assign LUT_3[39339] = 32'b00000000000000001100011110001101;
assign LUT_3[39340] = 32'b00000000000000000000111001000010;
assign LUT_3[39341] = 32'b00000000000000000111100100011111;
assign LUT_3[39342] = 32'b00000000000000000011000000100110;
assign LUT_3[39343] = 32'b00000000000000001001101100000011;
assign LUT_3[39344] = 32'b00000000000000000001100101001001;
assign LUT_3[39345] = 32'b00000000000000001000010000100110;
assign LUT_3[39346] = 32'b00000000000000000011101100101101;
assign LUT_3[39347] = 32'b00000000000000001010011000001010;
assign LUT_3[39348] = 32'b11111111111111111110110010111111;
assign LUT_3[39349] = 32'b00000000000000000101011110011100;
assign LUT_3[39350] = 32'b00000000000000000000111010100011;
assign LUT_3[39351] = 32'b00000000000000000111100110000000;
assign LUT_3[39352] = 32'b00000000000000000110111110001111;
assign LUT_3[39353] = 32'b00000000000000001101101001101100;
assign LUT_3[39354] = 32'b00000000000000001001000101110011;
assign LUT_3[39355] = 32'b00000000000000001111110001010000;
assign LUT_3[39356] = 32'b00000000000000000100001100000101;
assign LUT_3[39357] = 32'b00000000000000001010110111100010;
assign LUT_3[39358] = 32'b00000000000000000110010011101001;
assign LUT_3[39359] = 32'b00000000000000001100111111000110;
assign LUT_3[39360] = 32'b11111111111111111100111100010001;
assign LUT_3[39361] = 32'b00000000000000000011100111101110;
assign LUT_3[39362] = 32'b11111111111111111111000011110101;
assign LUT_3[39363] = 32'b00000000000000000101101111010010;
assign LUT_3[39364] = 32'b11111111111111111010001010000111;
assign LUT_3[39365] = 32'b00000000000000000000110101100100;
assign LUT_3[39366] = 32'b11111111111111111100010001101011;
assign LUT_3[39367] = 32'b00000000000000000010111101001000;
assign LUT_3[39368] = 32'b00000000000000000010010101010111;
assign LUT_3[39369] = 32'b00000000000000001001000000110100;
assign LUT_3[39370] = 32'b00000000000000000100011100111011;
assign LUT_3[39371] = 32'b00000000000000001011001000011000;
assign LUT_3[39372] = 32'b11111111111111111111100011001101;
assign LUT_3[39373] = 32'b00000000000000000110001110101010;
assign LUT_3[39374] = 32'b00000000000000000001101010110001;
assign LUT_3[39375] = 32'b00000000000000001000010110001110;
assign LUT_3[39376] = 32'b00000000000000000000001111010100;
assign LUT_3[39377] = 32'b00000000000000000110111010110001;
assign LUT_3[39378] = 32'b00000000000000000010010110111000;
assign LUT_3[39379] = 32'b00000000000000001001000010010101;
assign LUT_3[39380] = 32'b11111111111111111101011101001010;
assign LUT_3[39381] = 32'b00000000000000000100001000100111;
assign LUT_3[39382] = 32'b11111111111111111111100100101110;
assign LUT_3[39383] = 32'b00000000000000000110010000001011;
assign LUT_3[39384] = 32'b00000000000000000101101000011010;
assign LUT_3[39385] = 32'b00000000000000001100010011110111;
assign LUT_3[39386] = 32'b00000000000000000111101111111110;
assign LUT_3[39387] = 32'b00000000000000001110011011011011;
assign LUT_3[39388] = 32'b00000000000000000010110110010000;
assign LUT_3[39389] = 32'b00000000000000001001100001101101;
assign LUT_3[39390] = 32'b00000000000000000100111101110100;
assign LUT_3[39391] = 32'b00000000000000001011101001010001;
assign LUT_3[39392] = 32'b11111111111111111110001010110001;
assign LUT_3[39393] = 32'b00000000000000000100110110001110;
assign LUT_3[39394] = 32'b00000000000000000000010010010101;
assign LUT_3[39395] = 32'b00000000000000000110111101110010;
assign LUT_3[39396] = 32'b11111111111111111011011000100111;
assign LUT_3[39397] = 32'b00000000000000000010000100000100;
assign LUT_3[39398] = 32'b11111111111111111101100000001011;
assign LUT_3[39399] = 32'b00000000000000000100001011101000;
assign LUT_3[39400] = 32'b00000000000000000011100011110111;
assign LUT_3[39401] = 32'b00000000000000001010001111010100;
assign LUT_3[39402] = 32'b00000000000000000101101011011011;
assign LUT_3[39403] = 32'b00000000000000001100010110111000;
assign LUT_3[39404] = 32'b00000000000000000000110001101101;
assign LUT_3[39405] = 32'b00000000000000000111011101001010;
assign LUT_3[39406] = 32'b00000000000000000010111001010001;
assign LUT_3[39407] = 32'b00000000000000001001100100101110;
assign LUT_3[39408] = 32'b00000000000000000001011101110100;
assign LUT_3[39409] = 32'b00000000000000001000001001010001;
assign LUT_3[39410] = 32'b00000000000000000011100101011000;
assign LUT_3[39411] = 32'b00000000000000001010010000110101;
assign LUT_3[39412] = 32'b11111111111111111110101011101010;
assign LUT_3[39413] = 32'b00000000000000000101010111000111;
assign LUT_3[39414] = 32'b00000000000000000000110011001110;
assign LUT_3[39415] = 32'b00000000000000000111011110101011;
assign LUT_3[39416] = 32'b00000000000000000110110110111010;
assign LUT_3[39417] = 32'b00000000000000001101100010010111;
assign LUT_3[39418] = 32'b00000000000000001000111110011110;
assign LUT_3[39419] = 32'b00000000000000001111101001111011;
assign LUT_3[39420] = 32'b00000000000000000100000100110000;
assign LUT_3[39421] = 32'b00000000000000001010110000001101;
assign LUT_3[39422] = 32'b00000000000000000110001100010100;
assign LUT_3[39423] = 32'b00000000000000001100110111110001;
assign LUT_3[39424] = 32'b00000000000000000001111110010011;
assign LUT_3[39425] = 32'b00000000000000001000101001110000;
assign LUT_3[39426] = 32'b00000000000000000100000101110111;
assign LUT_3[39427] = 32'b00000000000000001010110001010100;
assign LUT_3[39428] = 32'b11111111111111111111001100001001;
assign LUT_3[39429] = 32'b00000000000000000101110111100110;
assign LUT_3[39430] = 32'b00000000000000000001010011101101;
assign LUT_3[39431] = 32'b00000000000000000111111111001010;
assign LUT_3[39432] = 32'b00000000000000000111010111011001;
assign LUT_3[39433] = 32'b00000000000000001110000010110110;
assign LUT_3[39434] = 32'b00000000000000001001011110111101;
assign LUT_3[39435] = 32'b00000000000000010000001010011010;
assign LUT_3[39436] = 32'b00000000000000000100100101001111;
assign LUT_3[39437] = 32'b00000000000000001011010000101100;
assign LUT_3[39438] = 32'b00000000000000000110101100110011;
assign LUT_3[39439] = 32'b00000000000000001101011000010000;
assign LUT_3[39440] = 32'b00000000000000000101010001010110;
assign LUT_3[39441] = 32'b00000000000000001011111100110011;
assign LUT_3[39442] = 32'b00000000000000000111011000111010;
assign LUT_3[39443] = 32'b00000000000000001110000100010111;
assign LUT_3[39444] = 32'b00000000000000000010011111001100;
assign LUT_3[39445] = 32'b00000000000000001001001010101001;
assign LUT_3[39446] = 32'b00000000000000000100100110110000;
assign LUT_3[39447] = 32'b00000000000000001011010010001101;
assign LUT_3[39448] = 32'b00000000000000001010101010011100;
assign LUT_3[39449] = 32'b00000000000000010001010101111001;
assign LUT_3[39450] = 32'b00000000000000001100110010000000;
assign LUT_3[39451] = 32'b00000000000000010011011101011101;
assign LUT_3[39452] = 32'b00000000000000000111111000010010;
assign LUT_3[39453] = 32'b00000000000000001110100011101111;
assign LUT_3[39454] = 32'b00000000000000001001111111110110;
assign LUT_3[39455] = 32'b00000000000000010000101011010011;
assign LUT_3[39456] = 32'b00000000000000000011001100110011;
assign LUT_3[39457] = 32'b00000000000000001001111000010000;
assign LUT_3[39458] = 32'b00000000000000000101010100010111;
assign LUT_3[39459] = 32'b00000000000000001011111111110100;
assign LUT_3[39460] = 32'b00000000000000000000011010101001;
assign LUT_3[39461] = 32'b00000000000000000111000110000110;
assign LUT_3[39462] = 32'b00000000000000000010100010001101;
assign LUT_3[39463] = 32'b00000000000000001001001101101010;
assign LUT_3[39464] = 32'b00000000000000001000100101111001;
assign LUT_3[39465] = 32'b00000000000000001111010001010110;
assign LUT_3[39466] = 32'b00000000000000001010101101011101;
assign LUT_3[39467] = 32'b00000000000000010001011000111010;
assign LUT_3[39468] = 32'b00000000000000000101110011101111;
assign LUT_3[39469] = 32'b00000000000000001100011111001100;
assign LUT_3[39470] = 32'b00000000000000000111111011010011;
assign LUT_3[39471] = 32'b00000000000000001110100110110000;
assign LUT_3[39472] = 32'b00000000000000000110011111110110;
assign LUT_3[39473] = 32'b00000000000000001101001011010011;
assign LUT_3[39474] = 32'b00000000000000001000100111011010;
assign LUT_3[39475] = 32'b00000000000000001111010010110111;
assign LUT_3[39476] = 32'b00000000000000000011101101101100;
assign LUT_3[39477] = 32'b00000000000000001010011001001001;
assign LUT_3[39478] = 32'b00000000000000000101110101010000;
assign LUT_3[39479] = 32'b00000000000000001100100000101101;
assign LUT_3[39480] = 32'b00000000000000001011111000111100;
assign LUT_3[39481] = 32'b00000000000000010010100100011001;
assign LUT_3[39482] = 32'b00000000000000001110000000100000;
assign LUT_3[39483] = 32'b00000000000000010100101011111101;
assign LUT_3[39484] = 32'b00000000000000001001000110110010;
assign LUT_3[39485] = 32'b00000000000000001111110010001111;
assign LUT_3[39486] = 32'b00000000000000001011001110010110;
assign LUT_3[39487] = 32'b00000000000000010001111001110011;
assign LUT_3[39488] = 32'b00000000000000000001110110111110;
assign LUT_3[39489] = 32'b00000000000000001000100010011011;
assign LUT_3[39490] = 32'b00000000000000000011111110100010;
assign LUT_3[39491] = 32'b00000000000000001010101001111111;
assign LUT_3[39492] = 32'b11111111111111111111000100110100;
assign LUT_3[39493] = 32'b00000000000000000101110000010001;
assign LUT_3[39494] = 32'b00000000000000000001001100011000;
assign LUT_3[39495] = 32'b00000000000000000111110111110101;
assign LUT_3[39496] = 32'b00000000000000000111010000000100;
assign LUT_3[39497] = 32'b00000000000000001101111011100001;
assign LUT_3[39498] = 32'b00000000000000001001010111101000;
assign LUT_3[39499] = 32'b00000000000000010000000011000101;
assign LUT_3[39500] = 32'b00000000000000000100011101111010;
assign LUT_3[39501] = 32'b00000000000000001011001001010111;
assign LUT_3[39502] = 32'b00000000000000000110100101011110;
assign LUT_3[39503] = 32'b00000000000000001101010000111011;
assign LUT_3[39504] = 32'b00000000000000000101001010000001;
assign LUT_3[39505] = 32'b00000000000000001011110101011110;
assign LUT_3[39506] = 32'b00000000000000000111010001100101;
assign LUT_3[39507] = 32'b00000000000000001101111101000010;
assign LUT_3[39508] = 32'b00000000000000000010010111110111;
assign LUT_3[39509] = 32'b00000000000000001001000011010100;
assign LUT_3[39510] = 32'b00000000000000000100011111011011;
assign LUT_3[39511] = 32'b00000000000000001011001010111000;
assign LUT_3[39512] = 32'b00000000000000001010100011000111;
assign LUT_3[39513] = 32'b00000000000000010001001110100100;
assign LUT_3[39514] = 32'b00000000000000001100101010101011;
assign LUT_3[39515] = 32'b00000000000000010011010110001000;
assign LUT_3[39516] = 32'b00000000000000000111110000111101;
assign LUT_3[39517] = 32'b00000000000000001110011100011010;
assign LUT_3[39518] = 32'b00000000000000001001111000100001;
assign LUT_3[39519] = 32'b00000000000000010000100011111110;
assign LUT_3[39520] = 32'b00000000000000000011000101011110;
assign LUT_3[39521] = 32'b00000000000000001001110000111011;
assign LUT_3[39522] = 32'b00000000000000000101001101000010;
assign LUT_3[39523] = 32'b00000000000000001011111000011111;
assign LUT_3[39524] = 32'b00000000000000000000010011010100;
assign LUT_3[39525] = 32'b00000000000000000110111110110001;
assign LUT_3[39526] = 32'b00000000000000000010011010111000;
assign LUT_3[39527] = 32'b00000000000000001001000110010101;
assign LUT_3[39528] = 32'b00000000000000001000011110100100;
assign LUT_3[39529] = 32'b00000000000000001111001010000001;
assign LUT_3[39530] = 32'b00000000000000001010100110001000;
assign LUT_3[39531] = 32'b00000000000000010001010001100101;
assign LUT_3[39532] = 32'b00000000000000000101101100011010;
assign LUT_3[39533] = 32'b00000000000000001100010111110111;
assign LUT_3[39534] = 32'b00000000000000000111110011111110;
assign LUT_3[39535] = 32'b00000000000000001110011111011011;
assign LUT_3[39536] = 32'b00000000000000000110011000100001;
assign LUT_3[39537] = 32'b00000000000000001101000011111110;
assign LUT_3[39538] = 32'b00000000000000001000100000000101;
assign LUT_3[39539] = 32'b00000000000000001111001011100010;
assign LUT_3[39540] = 32'b00000000000000000011100110010111;
assign LUT_3[39541] = 32'b00000000000000001010010001110100;
assign LUT_3[39542] = 32'b00000000000000000101101101111011;
assign LUT_3[39543] = 32'b00000000000000001100011001011000;
assign LUT_3[39544] = 32'b00000000000000001011110001100111;
assign LUT_3[39545] = 32'b00000000000000010010011101000100;
assign LUT_3[39546] = 32'b00000000000000001101111001001011;
assign LUT_3[39547] = 32'b00000000000000010100100100101000;
assign LUT_3[39548] = 32'b00000000000000001000111111011101;
assign LUT_3[39549] = 32'b00000000000000001111101010111010;
assign LUT_3[39550] = 32'b00000000000000001011000111000001;
assign LUT_3[39551] = 32'b00000000000000010001110010011110;
assign LUT_3[39552] = 32'b00000000000000000100001001010001;
assign LUT_3[39553] = 32'b00000000000000001010110100101110;
assign LUT_3[39554] = 32'b00000000000000000110010000110101;
assign LUT_3[39555] = 32'b00000000000000001100111100010010;
assign LUT_3[39556] = 32'b00000000000000000001010111000111;
assign LUT_3[39557] = 32'b00000000000000001000000010100100;
assign LUT_3[39558] = 32'b00000000000000000011011110101011;
assign LUT_3[39559] = 32'b00000000000000001010001010001000;
assign LUT_3[39560] = 32'b00000000000000001001100010010111;
assign LUT_3[39561] = 32'b00000000000000010000001101110100;
assign LUT_3[39562] = 32'b00000000000000001011101001111011;
assign LUT_3[39563] = 32'b00000000000000010010010101011000;
assign LUT_3[39564] = 32'b00000000000000000110110000001101;
assign LUT_3[39565] = 32'b00000000000000001101011011101010;
assign LUT_3[39566] = 32'b00000000000000001000110111110001;
assign LUT_3[39567] = 32'b00000000000000001111100011001110;
assign LUT_3[39568] = 32'b00000000000000000111011100010100;
assign LUT_3[39569] = 32'b00000000000000001110000111110001;
assign LUT_3[39570] = 32'b00000000000000001001100011111000;
assign LUT_3[39571] = 32'b00000000000000010000001111010101;
assign LUT_3[39572] = 32'b00000000000000000100101010001010;
assign LUT_3[39573] = 32'b00000000000000001011010101100111;
assign LUT_3[39574] = 32'b00000000000000000110110001101110;
assign LUT_3[39575] = 32'b00000000000000001101011101001011;
assign LUT_3[39576] = 32'b00000000000000001100110101011010;
assign LUT_3[39577] = 32'b00000000000000010011100000110111;
assign LUT_3[39578] = 32'b00000000000000001110111100111110;
assign LUT_3[39579] = 32'b00000000000000010101101000011011;
assign LUT_3[39580] = 32'b00000000000000001010000011010000;
assign LUT_3[39581] = 32'b00000000000000010000101110101101;
assign LUT_3[39582] = 32'b00000000000000001100001010110100;
assign LUT_3[39583] = 32'b00000000000000010010110110010001;
assign LUT_3[39584] = 32'b00000000000000000101010111110001;
assign LUT_3[39585] = 32'b00000000000000001100000011001110;
assign LUT_3[39586] = 32'b00000000000000000111011111010101;
assign LUT_3[39587] = 32'b00000000000000001110001010110010;
assign LUT_3[39588] = 32'b00000000000000000010100101100111;
assign LUT_3[39589] = 32'b00000000000000001001010001000100;
assign LUT_3[39590] = 32'b00000000000000000100101101001011;
assign LUT_3[39591] = 32'b00000000000000001011011000101000;
assign LUT_3[39592] = 32'b00000000000000001010110000110111;
assign LUT_3[39593] = 32'b00000000000000010001011100010100;
assign LUT_3[39594] = 32'b00000000000000001100111000011011;
assign LUT_3[39595] = 32'b00000000000000010011100011111000;
assign LUT_3[39596] = 32'b00000000000000000111111110101101;
assign LUT_3[39597] = 32'b00000000000000001110101010001010;
assign LUT_3[39598] = 32'b00000000000000001010000110010001;
assign LUT_3[39599] = 32'b00000000000000010000110001101110;
assign LUT_3[39600] = 32'b00000000000000001000101010110100;
assign LUT_3[39601] = 32'b00000000000000001111010110010001;
assign LUT_3[39602] = 32'b00000000000000001010110010011000;
assign LUT_3[39603] = 32'b00000000000000010001011101110101;
assign LUT_3[39604] = 32'b00000000000000000101111000101010;
assign LUT_3[39605] = 32'b00000000000000001100100100000111;
assign LUT_3[39606] = 32'b00000000000000001000000000001110;
assign LUT_3[39607] = 32'b00000000000000001110101011101011;
assign LUT_3[39608] = 32'b00000000000000001110000011111010;
assign LUT_3[39609] = 32'b00000000000000010100101111010111;
assign LUT_3[39610] = 32'b00000000000000010000001011011110;
assign LUT_3[39611] = 32'b00000000000000010110110110111011;
assign LUT_3[39612] = 32'b00000000000000001011010001110000;
assign LUT_3[39613] = 32'b00000000000000010001111101001101;
assign LUT_3[39614] = 32'b00000000000000001101011001010100;
assign LUT_3[39615] = 32'b00000000000000010100000100110001;
assign LUT_3[39616] = 32'b00000000000000000100000001111100;
assign LUT_3[39617] = 32'b00000000000000001010101101011001;
assign LUT_3[39618] = 32'b00000000000000000110001001100000;
assign LUT_3[39619] = 32'b00000000000000001100110100111101;
assign LUT_3[39620] = 32'b00000000000000000001001111110010;
assign LUT_3[39621] = 32'b00000000000000000111111011001111;
assign LUT_3[39622] = 32'b00000000000000000011010111010110;
assign LUT_3[39623] = 32'b00000000000000001010000010110011;
assign LUT_3[39624] = 32'b00000000000000001001011011000010;
assign LUT_3[39625] = 32'b00000000000000010000000110011111;
assign LUT_3[39626] = 32'b00000000000000001011100010100110;
assign LUT_3[39627] = 32'b00000000000000010010001110000011;
assign LUT_3[39628] = 32'b00000000000000000110101000111000;
assign LUT_3[39629] = 32'b00000000000000001101010100010101;
assign LUT_3[39630] = 32'b00000000000000001000110000011100;
assign LUT_3[39631] = 32'b00000000000000001111011011111001;
assign LUT_3[39632] = 32'b00000000000000000111010100111111;
assign LUT_3[39633] = 32'b00000000000000001110000000011100;
assign LUT_3[39634] = 32'b00000000000000001001011100100011;
assign LUT_3[39635] = 32'b00000000000000010000001000000000;
assign LUT_3[39636] = 32'b00000000000000000100100010110101;
assign LUT_3[39637] = 32'b00000000000000001011001110010010;
assign LUT_3[39638] = 32'b00000000000000000110101010011001;
assign LUT_3[39639] = 32'b00000000000000001101010101110110;
assign LUT_3[39640] = 32'b00000000000000001100101110000101;
assign LUT_3[39641] = 32'b00000000000000010011011001100010;
assign LUT_3[39642] = 32'b00000000000000001110110101101001;
assign LUT_3[39643] = 32'b00000000000000010101100001000110;
assign LUT_3[39644] = 32'b00000000000000001001111011111011;
assign LUT_3[39645] = 32'b00000000000000010000100111011000;
assign LUT_3[39646] = 32'b00000000000000001100000011011111;
assign LUT_3[39647] = 32'b00000000000000010010101110111100;
assign LUT_3[39648] = 32'b00000000000000000101010000011100;
assign LUT_3[39649] = 32'b00000000000000001011111011111001;
assign LUT_3[39650] = 32'b00000000000000000111011000000000;
assign LUT_3[39651] = 32'b00000000000000001110000011011101;
assign LUT_3[39652] = 32'b00000000000000000010011110010010;
assign LUT_3[39653] = 32'b00000000000000001001001001101111;
assign LUT_3[39654] = 32'b00000000000000000100100101110110;
assign LUT_3[39655] = 32'b00000000000000001011010001010011;
assign LUT_3[39656] = 32'b00000000000000001010101001100010;
assign LUT_3[39657] = 32'b00000000000000010001010100111111;
assign LUT_3[39658] = 32'b00000000000000001100110001000110;
assign LUT_3[39659] = 32'b00000000000000010011011100100011;
assign LUT_3[39660] = 32'b00000000000000000111110111011000;
assign LUT_3[39661] = 32'b00000000000000001110100010110101;
assign LUT_3[39662] = 32'b00000000000000001001111110111100;
assign LUT_3[39663] = 32'b00000000000000010000101010011001;
assign LUT_3[39664] = 32'b00000000000000001000100011011111;
assign LUT_3[39665] = 32'b00000000000000001111001110111100;
assign LUT_3[39666] = 32'b00000000000000001010101011000011;
assign LUT_3[39667] = 32'b00000000000000010001010110100000;
assign LUT_3[39668] = 32'b00000000000000000101110001010101;
assign LUT_3[39669] = 32'b00000000000000001100011100110010;
assign LUT_3[39670] = 32'b00000000000000000111111000111001;
assign LUT_3[39671] = 32'b00000000000000001110100100010110;
assign LUT_3[39672] = 32'b00000000000000001101111100100101;
assign LUT_3[39673] = 32'b00000000000000010100101000000010;
assign LUT_3[39674] = 32'b00000000000000010000000100001001;
assign LUT_3[39675] = 32'b00000000000000010110101111100110;
assign LUT_3[39676] = 32'b00000000000000001011001010011011;
assign LUT_3[39677] = 32'b00000000000000010001110101111000;
assign LUT_3[39678] = 32'b00000000000000001101010001111111;
assign LUT_3[39679] = 32'b00000000000000010011111101011100;
assign LUT_3[39680] = 32'b11111111111111111110001101110100;
assign LUT_3[39681] = 32'b00000000000000000100111001010001;
assign LUT_3[39682] = 32'b00000000000000000000010101011000;
assign LUT_3[39683] = 32'b00000000000000000111000000110101;
assign LUT_3[39684] = 32'b11111111111111111011011011101010;
assign LUT_3[39685] = 32'b00000000000000000010000111000111;
assign LUT_3[39686] = 32'b11111111111111111101100011001110;
assign LUT_3[39687] = 32'b00000000000000000100001110101011;
assign LUT_3[39688] = 32'b00000000000000000011100110111010;
assign LUT_3[39689] = 32'b00000000000000001010010010010111;
assign LUT_3[39690] = 32'b00000000000000000101101110011110;
assign LUT_3[39691] = 32'b00000000000000001100011001111011;
assign LUT_3[39692] = 32'b00000000000000000000110100110000;
assign LUT_3[39693] = 32'b00000000000000000111100000001101;
assign LUT_3[39694] = 32'b00000000000000000010111100010100;
assign LUT_3[39695] = 32'b00000000000000001001100111110001;
assign LUT_3[39696] = 32'b00000000000000000001100000110111;
assign LUT_3[39697] = 32'b00000000000000001000001100010100;
assign LUT_3[39698] = 32'b00000000000000000011101000011011;
assign LUT_3[39699] = 32'b00000000000000001010010011111000;
assign LUT_3[39700] = 32'b11111111111111111110101110101101;
assign LUT_3[39701] = 32'b00000000000000000101011010001010;
assign LUT_3[39702] = 32'b00000000000000000000110110010001;
assign LUT_3[39703] = 32'b00000000000000000111100001101110;
assign LUT_3[39704] = 32'b00000000000000000110111001111101;
assign LUT_3[39705] = 32'b00000000000000001101100101011010;
assign LUT_3[39706] = 32'b00000000000000001001000001100001;
assign LUT_3[39707] = 32'b00000000000000001111101100111110;
assign LUT_3[39708] = 32'b00000000000000000100000111110011;
assign LUT_3[39709] = 32'b00000000000000001010110011010000;
assign LUT_3[39710] = 32'b00000000000000000110001111010111;
assign LUT_3[39711] = 32'b00000000000000001100111010110100;
assign LUT_3[39712] = 32'b11111111111111111111011100010100;
assign LUT_3[39713] = 32'b00000000000000000110000111110001;
assign LUT_3[39714] = 32'b00000000000000000001100011111000;
assign LUT_3[39715] = 32'b00000000000000001000001111010101;
assign LUT_3[39716] = 32'b11111111111111111100101010001010;
assign LUT_3[39717] = 32'b00000000000000000011010101100111;
assign LUT_3[39718] = 32'b11111111111111111110110001101110;
assign LUT_3[39719] = 32'b00000000000000000101011101001011;
assign LUT_3[39720] = 32'b00000000000000000100110101011010;
assign LUT_3[39721] = 32'b00000000000000001011100000110111;
assign LUT_3[39722] = 32'b00000000000000000110111100111110;
assign LUT_3[39723] = 32'b00000000000000001101101000011011;
assign LUT_3[39724] = 32'b00000000000000000010000011010000;
assign LUT_3[39725] = 32'b00000000000000001000101110101101;
assign LUT_3[39726] = 32'b00000000000000000100001010110100;
assign LUT_3[39727] = 32'b00000000000000001010110110010001;
assign LUT_3[39728] = 32'b00000000000000000010101111010111;
assign LUT_3[39729] = 32'b00000000000000001001011010110100;
assign LUT_3[39730] = 32'b00000000000000000100110110111011;
assign LUT_3[39731] = 32'b00000000000000001011100010011000;
assign LUT_3[39732] = 32'b11111111111111111111111101001101;
assign LUT_3[39733] = 32'b00000000000000000110101000101010;
assign LUT_3[39734] = 32'b00000000000000000010000100110001;
assign LUT_3[39735] = 32'b00000000000000001000110000001110;
assign LUT_3[39736] = 32'b00000000000000001000001000011101;
assign LUT_3[39737] = 32'b00000000000000001110110011111010;
assign LUT_3[39738] = 32'b00000000000000001010010000000001;
assign LUT_3[39739] = 32'b00000000000000010000111011011110;
assign LUT_3[39740] = 32'b00000000000000000101010110010011;
assign LUT_3[39741] = 32'b00000000000000001100000001110000;
assign LUT_3[39742] = 32'b00000000000000000111011101110111;
assign LUT_3[39743] = 32'b00000000000000001110001001010100;
assign LUT_3[39744] = 32'b11111111111111111110000110011111;
assign LUT_3[39745] = 32'b00000000000000000100110001111100;
assign LUT_3[39746] = 32'b00000000000000000000001110000011;
assign LUT_3[39747] = 32'b00000000000000000110111001100000;
assign LUT_3[39748] = 32'b11111111111111111011010100010101;
assign LUT_3[39749] = 32'b00000000000000000001111111110010;
assign LUT_3[39750] = 32'b11111111111111111101011011111001;
assign LUT_3[39751] = 32'b00000000000000000100000111010110;
assign LUT_3[39752] = 32'b00000000000000000011011111100101;
assign LUT_3[39753] = 32'b00000000000000001010001011000010;
assign LUT_3[39754] = 32'b00000000000000000101100111001001;
assign LUT_3[39755] = 32'b00000000000000001100010010100110;
assign LUT_3[39756] = 32'b00000000000000000000101101011011;
assign LUT_3[39757] = 32'b00000000000000000111011000111000;
assign LUT_3[39758] = 32'b00000000000000000010110100111111;
assign LUT_3[39759] = 32'b00000000000000001001100000011100;
assign LUT_3[39760] = 32'b00000000000000000001011001100010;
assign LUT_3[39761] = 32'b00000000000000001000000100111111;
assign LUT_3[39762] = 32'b00000000000000000011100001000110;
assign LUT_3[39763] = 32'b00000000000000001010001100100011;
assign LUT_3[39764] = 32'b11111111111111111110100111011000;
assign LUT_3[39765] = 32'b00000000000000000101010010110101;
assign LUT_3[39766] = 32'b00000000000000000000101110111100;
assign LUT_3[39767] = 32'b00000000000000000111011010011001;
assign LUT_3[39768] = 32'b00000000000000000110110010101000;
assign LUT_3[39769] = 32'b00000000000000001101011110000101;
assign LUT_3[39770] = 32'b00000000000000001000111010001100;
assign LUT_3[39771] = 32'b00000000000000001111100101101001;
assign LUT_3[39772] = 32'b00000000000000000100000000011110;
assign LUT_3[39773] = 32'b00000000000000001010101011111011;
assign LUT_3[39774] = 32'b00000000000000000110001000000010;
assign LUT_3[39775] = 32'b00000000000000001100110011011111;
assign LUT_3[39776] = 32'b11111111111111111111010100111111;
assign LUT_3[39777] = 32'b00000000000000000110000000011100;
assign LUT_3[39778] = 32'b00000000000000000001011100100011;
assign LUT_3[39779] = 32'b00000000000000001000001000000000;
assign LUT_3[39780] = 32'b11111111111111111100100010110101;
assign LUT_3[39781] = 32'b00000000000000000011001110010010;
assign LUT_3[39782] = 32'b11111111111111111110101010011001;
assign LUT_3[39783] = 32'b00000000000000000101010101110110;
assign LUT_3[39784] = 32'b00000000000000000100101110000101;
assign LUT_3[39785] = 32'b00000000000000001011011001100010;
assign LUT_3[39786] = 32'b00000000000000000110110101101001;
assign LUT_3[39787] = 32'b00000000000000001101100001000110;
assign LUT_3[39788] = 32'b00000000000000000001111011111011;
assign LUT_3[39789] = 32'b00000000000000001000100111011000;
assign LUT_3[39790] = 32'b00000000000000000100000011011111;
assign LUT_3[39791] = 32'b00000000000000001010101110111100;
assign LUT_3[39792] = 32'b00000000000000000010101000000010;
assign LUT_3[39793] = 32'b00000000000000001001010011011111;
assign LUT_3[39794] = 32'b00000000000000000100101111100110;
assign LUT_3[39795] = 32'b00000000000000001011011011000011;
assign LUT_3[39796] = 32'b11111111111111111111110101111000;
assign LUT_3[39797] = 32'b00000000000000000110100001010101;
assign LUT_3[39798] = 32'b00000000000000000001111101011100;
assign LUT_3[39799] = 32'b00000000000000001000101000111001;
assign LUT_3[39800] = 32'b00000000000000001000000001001000;
assign LUT_3[39801] = 32'b00000000000000001110101100100101;
assign LUT_3[39802] = 32'b00000000000000001010001000101100;
assign LUT_3[39803] = 32'b00000000000000010000110100001001;
assign LUT_3[39804] = 32'b00000000000000000101001110111110;
assign LUT_3[39805] = 32'b00000000000000001011111010011011;
assign LUT_3[39806] = 32'b00000000000000000111010110100010;
assign LUT_3[39807] = 32'b00000000000000001110000001111111;
assign LUT_3[39808] = 32'b00000000000000000000011000110010;
assign LUT_3[39809] = 32'b00000000000000000111000100001111;
assign LUT_3[39810] = 32'b00000000000000000010100000010110;
assign LUT_3[39811] = 32'b00000000000000001001001011110011;
assign LUT_3[39812] = 32'b11111111111111111101100110101000;
assign LUT_3[39813] = 32'b00000000000000000100010010000101;
assign LUT_3[39814] = 32'b11111111111111111111101110001100;
assign LUT_3[39815] = 32'b00000000000000000110011001101001;
assign LUT_3[39816] = 32'b00000000000000000101110001111000;
assign LUT_3[39817] = 32'b00000000000000001100011101010101;
assign LUT_3[39818] = 32'b00000000000000000111111001011100;
assign LUT_3[39819] = 32'b00000000000000001110100100111001;
assign LUT_3[39820] = 32'b00000000000000000010111111101110;
assign LUT_3[39821] = 32'b00000000000000001001101011001011;
assign LUT_3[39822] = 32'b00000000000000000101000111010010;
assign LUT_3[39823] = 32'b00000000000000001011110010101111;
assign LUT_3[39824] = 32'b00000000000000000011101011110101;
assign LUT_3[39825] = 32'b00000000000000001010010111010010;
assign LUT_3[39826] = 32'b00000000000000000101110011011001;
assign LUT_3[39827] = 32'b00000000000000001100011110110110;
assign LUT_3[39828] = 32'b00000000000000000000111001101011;
assign LUT_3[39829] = 32'b00000000000000000111100101001000;
assign LUT_3[39830] = 32'b00000000000000000011000001001111;
assign LUT_3[39831] = 32'b00000000000000001001101100101100;
assign LUT_3[39832] = 32'b00000000000000001001000100111011;
assign LUT_3[39833] = 32'b00000000000000001111110000011000;
assign LUT_3[39834] = 32'b00000000000000001011001100011111;
assign LUT_3[39835] = 32'b00000000000000010001110111111100;
assign LUT_3[39836] = 32'b00000000000000000110010010110001;
assign LUT_3[39837] = 32'b00000000000000001100111110001110;
assign LUT_3[39838] = 32'b00000000000000001000011010010101;
assign LUT_3[39839] = 32'b00000000000000001111000101110010;
assign LUT_3[39840] = 32'b00000000000000000001100111010010;
assign LUT_3[39841] = 32'b00000000000000001000010010101111;
assign LUT_3[39842] = 32'b00000000000000000011101110110110;
assign LUT_3[39843] = 32'b00000000000000001010011010010011;
assign LUT_3[39844] = 32'b11111111111111111110110101001000;
assign LUT_3[39845] = 32'b00000000000000000101100000100101;
assign LUT_3[39846] = 32'b00000000000000000000111100101100;
assign LUT_3[39847] = 32'b00000000000000000111101000001001;
assign LUT_3[39848] = 32'b00000000000000000111000000011000;
assign LUT_3[39849] = 32'b00000000000000001101101011110101;
assign LUT_3[39850] = 32'b00000000000000001001000111111100;
assign LUT_3[39851] = 32'b00000000000000001111110011011001;
assign LUT_3[39852] = 32'b00000000000000000100001110001110;
assign LUT_3[39853] = 32'b00000000000000001010111001101011;
assign LUT_3[39854] = 32'b00000000000000000110010101110010;
assign LUT_3[39855] = 32'b00000000000000001101000001001111;
assign LUT_3[39856] = 32'b00000000000000000100111010010101;
assign LUT_3[39857] = 32'b00000000000000001011100101110010;
assign LUT_3[39858] = 32'b00000000000000000111000001111001;
assign LUT_3[39859] = 32'b00000000000000001101101101010110;
assign LUT_3[39860] = 32'b00000000000000000010001000001011;
assign LUT_3[39861] = 32'b00000000000000001000110011101000;
assign LUT_3[39862] = 32'b00000000000000000100001111101111;
assign LUT_3[39863] = 32'b00000000000000001010111011001100;
assign LUT_3[39864] = 32'b00000000000000001010010011011011;
assign LUT_3[39865] = 32'b00000000000000010000111110111000;
assign LUT_3[39866] = 32'b00000000000000001100011010111111;
assign LUT_3[39867] = 32'b00000000000000010011000110011100;
assign LUT_3[39868] = 32'b00000000000000000111100001010001;
assign LUT_3[39869] = 32'b00000000000000001110001100101110;
assign LUT_3[39870] = 32'b00000000000000001001101000110101;
assign LUT_3[39871] = 32'b00000000000000010000010100010010;
assign LUT_3[39872] = 32'b00000000000000000000010001011101;
assign LUT_3[39873] = 32'b00000000000000000110111100111010;
assign LUT_3[39874] = 32'b00000000000000000010011001000001;
assign LUT_3[39875] = 32'b00000000000000001001000100011110;
assign LUT_3[39876] = 32'b11111111111111111101011111010011;
assign LUT_3[39877] = 32'b00000000000000000100001010110000;
assign LUT_3[39878] = 32'b11111111111111111111100110110111;
assign LUT_3[39879] = 32'b00000000000000000110010010010100;
assign LUT_3[39880] = 32'b00000000000000000101101010100011;
assign LUT_3[39881] = 32'b00000000000000001100010110000000;
assign LUT_3[39882] = 32'b00000000000000000111110010000111;
assign LUT_3[39883] = 32'b00000000000000001110011101100100;
assign LUT_3[39884] = 32'b00000000000000000010111000011001;
assign LUT_3[39885] = 32'b00000000000000001001100011110110;
assign LUT_3[39886] = 32'b00000000000000000100111111111101;
assign LUT_3[39887] = 32'b00000000000000001011101011011010;
assign LUT_3[39888] = 32'b00000000000000000011100100100000;
assign LUT_3[39889] = 32'b00000000000000001010001111111101;
assign LUT_3[39890] = 32'b00000000000000000101101100000100;
assign LUT_3[39891] = 32'b00000000000000001100010111100001;
assign LUT_3[39892] = 32'b00000000000000000000110010010110;
assign LUT_3[39893] = 32'b00000000000000000111011101110011;
assign LUT_3[39894] = 32'b00000000000000000010111001111010;
assign LUT_3[39895] = 32'b00000000000000001001100101010111;
assign LUT_3[39896] = 32'b00000000000000001000111101100110;
assign LUT_3[39897] = 32'b00000000000000001111101001000011;
assign LUT_3[39898] = 32'b00000000000000001011000101001010;
assign LUT_3[39899] = 32'b00000000000000010001110000100111;
assign LUT_3[39900] = 32'b00000000000000000110001011011100;
assign LUT_3[39901] = 32'b00000000000000001100110110111001;
assign LUT_3[39902] = 32'b00000000000000001000010011000000;
assign LUT_3[39903] = 32'b00000000000000001110111110011101;
assign LUT_3[39904] = 32'b00000000000000000001011111111101;
assign LUT_3[39905] = 32'b00000000000000001000001011011010;
assign LUT_3[39906] = 32'b00000000000000000011100111100001;
assign LUT_3[39907] = 32'b00000000000000001010010010111110;
assign LUT_3[39908] = 32'b11111111111111111110101101110011;
assign LUT_3[39909] = 32'b00000000000000000101011001010000;
assign LUT_3[39910] = 32'b00000000000000000000110101010111;
assign LUT_3[39911] = 32'b00000000000000000111100000110100;
assign LUT_3[39912] = 32'b00000000000000000110111001000011;
assign LUT_3[39913] = 32'b00000000000000001101100100100000;
assign LUT_3[39914] = 32'b00000000000000001001000000100111;
assign LUT_3[39915] = 32'b00000000000000001111101100000100;
assign LUT_3[39916] = 32'b00000000000000000100000110111001;
assign LUT_3[39917] = 32'b00000000000000001010110010010110;
assign LUT_3[39918] = 32'b00000000000000000110001110011101;
assign LUT_3[39919] = 32'b00000000000000001100111001111010;
assign LUT_3[39920] = 32'b00000000000000000100110011000000;
assign LUT_3[39921] = 32'b00000000000000001011011110011101;
assign LUT_3[39922] = 32'b00000000000000000110111010100100;
assign LUT_3[39923] = 32'b00000000000000001101100110000001;
assign LUT_3[39924] = 32'b00000000000000000010000000110110;
assign LUT_3[39925] = 32'b00000000000000001000101100010011;
assign LUT_3[39926] = 32'b00000000000000000100001000011010;
assign LUT_3[39927] = 32'b00000000000000001010110011110111;
assign LUT_3[39928] = 32'b00000000000000001010001100000110;
assign LUT_3[39929] = 32'b00000000000000010000110111100011;
assign LUT_3[39930] = 32'b00000000000000001100010011101010;
assign LUT_3[39931] = 32'b00000000000000010010111111000111;
assign LUT_3[39932] = 32'b00000000000000000111011001111100;
assign LUT_3[39933] = 32'b00000000000000001110000101011001;
assign LUT_3[39934] = 32'b00000000000000001001100001100000;
assign LUT_3[39935] = 32'b00000000000000010000001100111101;
assign LUT_3[39936] = 32'b00000000000000000101001110000100;
assign LUT_3[39937] = 32'b00000000000000001011111001100001;
assign LUT_3[39938] = 32'b00000000000000000111010101101000;
assign LUT_3[39939] = 32'b00000000000000001110000001000101;
assign LUT_3[39940] = 32'b00000000000000000010011011111010;
assign LUT_3[39941] = 32'b00000000000000001001000111010111;
assign LUT_3[39942] = 32'b00000000000000000100100011011110;
assign LUT_3[39943] = 32'b00000000000000001011001110111011;
assign LUT_3[39944] = 32'b00000000000000001010100111001010;
assign LUT_3[39945] = 32'b00000000000000010001010010100111;
assign LUT_3[39946] = 32'b00000000000000001100101110101110;
assign LUT_3[39947] = 32'b00000000000000010011011010001011;
assign LUT_3[39948] = 32'b00000000000000000111110101000000;
assign LUT_3[39949] = 32'b00000000000000001110100000011101;
assign LUT_3[39950] = 32'b00000000000000001001111100100100;
assign LUT_3[39951] = 32'b00000000000000010000101000000001;
assign LUT_3[39952] = 32'b00000000000000001000100001000111;
assign LUT_3[39953] = 32'b00000000000000001111001100100100;
assign LUT_3[39954] = 32'b00000000000000001010101000101011;
assign LUT_3[39955] = 32'b00000000000000010001010100001000;
assign LUT_3[39956] = 32'b00000000000000000101101110111101;
assign LUT_3[39957] = 32'b00000000000000001100011010011010;
assign LUT_3[39958] = 32'b00000000000000000111110110100001;
assign LUT_3[39959] = 32'b00000000000000001110100001111110;
assign LUT_3[39960] = 32'b00000000000000001101111010001101;
assign LUT_3[39961] = 32'b00000000000000010100100101101010;
assign LUT_3[39962] = 32'b00000000000000010000000001110001;
assign LUT_3[39963] = 32'b00000000000000010110101101001110;
assign LUT_3[39964] = 32'b00000000000000001011001000000011;
assign LUT_3[39965] = 32'b00000000000000010001110011100000;
assign LUT_3[39966] = 32'b00000000000000001101001111100111;
assign LUT_3[39967] = 32'b00000000000000010011111011000100;
assign LUT_3[39968] = 32'b00000000000000000110011100100100;
assign LUT_3[39969] = 32'b00000000000000001101001000000001;
assign LUT_3[39970] = 32'b00000000000000001000100100001000;
assign LUT_3[39971] = 32'b00000000000000001111001111100101;
assign LUT_3[39972] = 32'b00000000000000000011101010011010;
assign LUT_3[39973] = 32'b00000000000000001010010101110111;
assign LUT_3[39974] = 32'b00000000000000000101110001111110;
assign LUT_3[39975] = 32'b00000000000000001100011101011011;
assign LUT_3[39976] = 32'b00000000000000001011110101101010;
assign LUT_3[39977] = 32'b00000000000000010010100001000111;
assign LUT_3[39978] = 32'b00000000000000001101111101001110;
assign LUT_3[39979] = 32'b00000000000000010100101000101011;
assign LUT_3[39980] = 32'b00000000000000001001000011100000;
assign LUT_3[39981] = 32'b00000000000000001111101110111101;
assign LUT_3[39982] = 32'b00000000000000001011001011000100;
assign LUT_3[39983] = 32'b00000000000000010001110110100001;
assign LUT_3[39984] = 32'b00000000000000001001101111100111;
assign LUT_3[39985] = 32'b00000000000000010000011011000100;
assign LUT_3[39986] = 32'b00000000000000001011110111001011;
assign LUT_3[39987] = 32'b00000000000000010010100010101000;
assign LUT_3[39988] = 32'b00000000000000000110111101011101;
assign LUT_3[39989] = 32'b00000000000000001101101000111010;
assign LUT_3[39990] = 32'b00000000000000001001000101000001;
assign LUT_3[39991] = 32'b00000000000000001111110000011110;
assign LUT_3[39992] = 32'b00000000000000001111001000101101;
assign LUT_3[39993] = 32'b00000000000000010101110100001010;
assign LUT_3[39994] = 32'b00000000000000010001010000010001;
assign LUT_3[39995] = 32'b00000000000000010111111011101110;
assign LUT_3[39996] = 32'b00000000000000001100010110100011;
assign LUT_3[39997] = 32'b00000000000000010011000010000000;
assign LUT_3[39998] = 32'b00000000000000001110011110000111;
assign LUT_3[39999] = 32'b00000000000000010101001001100100;
assign LUT_3[40000] = 32'b00000000000000000101000110101111;
assign LUT_3[40001] = 32'b00000000000000001011110010001100;
assign LUT_3[40002] = 32'b00000000000000000111001110010011;
assign LUT_3[40003] = 32'b00000000000000001101111001110000;
assign LUT_3[40004] = 32'b00000000000000000010010100100101;
assign LUT_3[40005] = 32'b00000000000000001001000000000010;
assign LUT_3[40006] = 32'b00000000000000000100011100001001;
assign LUT_3[40007] = 32'b00000000000000001011000111100110;
assign LUT_3[40008] = 32'b00000000000000001010011111110101;
assign LUT_3[40009] = 32'b00000000000000010001001011010010;
assign LUT_3[40010] = 32'b00000000000000001100100111011001;
assign LUT_3[40011] = 32'b00000000000000010011010010110110;
assign LUT_3[40012] = 32'b00000000000000000111101101101011;
assign LUT_3[40013] = 32'b00000000000000001110011001001000;
assign LUT_3[40014] = 32'b00000000000000001001110101001111;
assign LUT_3[40015] = 32'b00000000000000010000100000101100;
assign LUT_3[40016] = 32'b00000000000000001000011001110010;
assign LUT_3[40017] = 32'b00000000000000001111000101001111;
assign LUT_3[40018] = 32'b00000000000000001010100001010110;
assign LUT_3[40019] = 32'b00000000000000010001001100110011;
assign LUT_3[40020] = 32'b00000000000000000101100111101000;
assign LUT_3[40021] = 32'b00000000000000001100010011000101;
assign LUT_3[40022] = 32'b00000000000000000111101111001100;
assign LUT_3[40023] = 32'b00000000000000001110011010101001;
assign LUT_3[40024] = 32'b00000000000000001101110010111000;
assign LUT_3[40025] = 32'b00000000000000010100011110010101;
assign LUT_3[40026] = 32'b00000000000000001111111010011100;
assign LUT_3[40027] = 32'b00000000000000010110100101111001;
assign LUT_3[40028] = 32'b00000000000000001011000000101110;
assign LUT_3[40029] = 32'b00000000000000010001101100001011;
assign LUT_3[40030] = 32'b00000000000000001101001000010010;
assign LUT_3[40031] = 32'b00000000000000010011110011101111;
assign LUT_3[40032] = 32'b00000000000000000110010101001111;
assign LUT_3[40033] = 32'b00000000000000001101000000101100;
assign LUT_3[40034] = 32'b00000000000000001000011100110011;
assign LUT_3[40035] = 32'b00000000000000001111001000010000;
assign LUT_3[40036] = 32'b00000000000000000011100011000101;
assign LUT_3[40037] = 32'b00000000000000001010001110100010;
assign LUT_3[40038] = 32'b00000000000000000101101010101001;
assign LUT_3[40039] = 32'b00000000000000001100010110000110;
assign LUT_3[40040] = 32'b00000000000000001011101110010101;
assign LUT_3[40041] = 32'b00000000000000010010011001110010;
assign LUT_3[40042] = 32'b00000000000000001101110101111001;
assign LUT_3[40043] = 32'b00000000000000010100100001010110;
assign LUT_3[40044] = 32'b00000000000000001000111100001011;
assign LUT_3[40045] = 32'b00000000000000001111100111101000;
assign LUT_3[40046] = 32'b00000000000000001011000011101111;
assign LUT_3[40047] = 32'b00000000000000010001101111001100;
assign LUT_3[40048] = 32'b00000000000000001001101000010010;
assign LUT_3[40049] = 32'b00000000000000010000010011101111;
assign LUT_3[40050] = 32'b00000000000000001011101111110110;
assign LUT_3[40051] = 32'b00000000000000010010011011010011;
assign LUT_3[40052] = 32'b00000000000000000110110110001000;
assign LUT_3[40053] = 32'b00000000000000001101100001100101;
assign LUT_3[40054] = 32'b00000000000000001000111101101100;
assign LUT_3[40055] = 32'b00000000000000001111101001001001;
assign LUT_3[40056] = 32'b00000000000000001111000001011000;
assign LUT_3[40057] = 32'b00000000000000010101101100110101;
assign LUT_3[40058] = 32'b00000000000000010001001000111100;
assign LUT_3[40059] = 32'b00000000000000010111110100011001;
assign LUT_3[40060] = 32'b00000000000000001100001111001110;
assign LUT_3[40061] = 32'b00000000000000010010111010101011;
assign LUT_3[40062] = 32'b00000000000000001110010110110010;
assign LUT_3[40063] = 32'b00000000000000010101000010001111;
assign LUT_3[40064] = 32'b00000000000000000111011001000010;
assign LUT_3[40065] = 32'b00000000000000001110000100011111;
assign LUT_3[40066] = 32'b00000000000000001001100000100110;
assign LUT_3[40067] = 32'b00000000000000010000001100000011;
assign LUT_3[40068] = 32'b00000000000000000100100110111000;
assign LUT_3[40069] = 32'b00000000000000001011010010010101;
assign LUT_3[40070] = 32'b00000000000000000110101110011100;
assign LUT_3[40071] = 32'b00000000000000001101011001111001;
assign LUT_3[40072] = 32'b00000000000000001100110010001000;
assign LUT_3[40073] = 32'b00000000000000010011011101100101;
assign LUT_3[40074] = 32'b00000000000000001110111001101100;
assign LUT_3[40075] = 32'b00000000000000010101100101001001;
assign LUT_3[40076] = 32'b00000000000000001001111111111110;
assign LUT_3[40077] = 32'b00000000000000010000101011011011;
assign LUT_3[40078] = 32'b00000000000000001100000111100010;
assign LUT_3[40079] = 32'b00000000000000010010110010111111;
assign LUT_3[40080] = 32'b00000000000000001010101100000101;
assign LUT_3[40081] = 32'b00000000000000010001010111100010;
assign LUT_3[40082] = 32'b00000000000000001100110011101001;
assign LUT_3[40083] = 32'b00000000000000010011011111000110;
assign LUT_3[40084] = 32'b00000000000000000111111001111011;
assign LUT_3[40085] = 32'b00000000000000001110100101011000;
assign LUT_3[40086] = 32'b00000000000000001010000001011111;
assign LUT_3[40087] = 32'b00000000000000010000101100111100;
assign LUT_3[40088] = 32'b00000000000000010000000101001011;
assign LUT_3[40089] = 32'b00000000000000010110110000101000;
assign LUT_3[40090] = 32'b00000000000000010010001100101111;
assign LUT_3[40091] = 32'b00000000000000011000111000001100;
assign LUT_3[40092] = 32'b00000000000000001101010011000001;
assign LUT_3[40093] = 32'b00000000000000010011111110011110;
assign LUT_3[40094] = 32'b00000000000000001111011010100101;
assign LUT_3[40095] = 32'b00000000000000010110000110000010;
assign LUT_3[40096] = 32'b00000000000000001000100111100010;
assign LUT_3[40097] = 32'b00000000000000001111010010111111;
assign LUT_3[40098] = 32'b00000000000000001010101111000110;
assign LUT_3[40099] = 32'b00000000000000010001011010100011;
assign LUT_3[40100] = 32'b00000000000000000101110101011000;
assign LUT_3[40101] = 32'b00000000000000001100100000110101;
assign LUT_3[40102] = 32'b00000000000000000111111100111100;
assign LUT_3[40103] = 32'b00000000000000001110101000011001;
assign LUT_3[40104] = 32'b00000000000000001110000000101000;
assign LUT_3[40105] = 32'b00000000000000010100101100000101;
assign LUT_3[40106] = 32'b00000000000000010000001000001100;
assign LUT_3[40107] = 32'b00000000000000010110110011101001;
assign LUT_3[40108] = 32'b00000000000000001011001110011110;
assign LUT_3[40109] = 32'b00000000000000010001111001111011;
assign LUT_3[40110] = 32'b00000000000000001101010110000010;
assign LUT_3[40111] = 32'b00000000000000010100000001011111;
assign LUT_3[40112] = 32'b00000000000000001011111010100101;
assign LUT_3[40113] = 32'b00000000000000010010100110000010;
assign LUT_3[40114] = 32'b00000000000000001110000010001001;
assign LUT_3[40115] = 32'b00000000000000010100101101100110;
assign LUT_3[40116] = 32'b00000000000000001001001000011011;
assign LUT_3[40117] = 32'b00000000000000001111110011111000;
assign LUT_3[40118] = 32'b00000000000000001011001111111111;
assign LUT_3[40119] = 32'b00000000000000010001111011011100;
assign LUT_3[40120] = 32'b00000000000000010001010011101011;
assign LUT_3[40121] = 32'b00000000000000010111111111001000;
assign LUT_3[40122] = 32'b00000000000000010011011011001111;
assign LUT_3[40123] = 32'b00000000000000011010000110101100;
assign LUT_3[40124] = 32'b00000000000000001110100001100001;
assign LUT_3[40125] = 32'b00000000000000010101001100111110;
assign LUT_3[40126] = 32'b00000000000000010000101001000101;
assign LUT_3[40127] = 32'b00000000000000010111010100100010;
assign LUT_3[40128] = 32'b00000000000000000111010001101101;
assign LUT_3[40129] = 32'b00000000000000001101111101001010;
assign LUT_3[40130] = 32'b00000000000000001001011001010001;
assign LUT_3[40131] = 32'b00000000000000010000000100101110;
assign LUT_3[40132] = 32'b00000000000000000100011111100011;
assign LUT_3[40133] = 32'b00000000000000001011001011000000;
assign LUT_3[40134] = 32'b00000000000000000110100111000111;
assign LUT_3[40135] = 32'b00000000000000001101010010100100;
assign LUT_3[40136] = 32'b00000000000000001100101010110011;
assign LUT_3[40137] = 32'b00000000000000010011010110010000;
assign LUT_3[40138] = 32'b00000000000000001110110010010111;
assign LUT_3[40139] = 32'b00000000000000010101011101110100;
assign LUT_3[40140] = 32'b00000000000000001001111000101001;
assign LUT_3[40141] = 32'b00000000000000010000100100000110;
assign LUT_3[40142] = 32'b00000000000000001100000000001101;
assign LUT_3[40143] = 32'b00000000000000010010101011101010;
assign LUT_3[40144] = 32'b00000000000000001010100100110000;
assign LUT_3[40145] = 32'b00000000000000010001010000001101;
assign LUT_3[40146] = 32'b00000000000000001100101100010100;
assign LUT_3[40147] = 32'b00000000000000010011010111110001;
assign LUT_3[40148] = 32'b00000000000000000111110010100110;
assign LUT_3[40149] = 32'b00000000000000001110011110000011;
assign LUT_3[40150] = 32'b00000000000000001001111010001010;
assign LUT_3[40151] = 32'b00000000000000010000100101100111;
assign LUT_3[40152] = 32'b00000000000000001111111101110110;
assign LUT_3[40153] = 32'b00000000000000010110101001010011;
assign LUT_3[40154] = 32'b00000000000000010010000101011010;
assign LUT_3[40155] = 32'b00000000000000011000110000110111;
assign LUT_3[40156] = 32'b00000000000000001101001011101100;
assign LUT_3[40157] = 32'b00000000000000010011110111001001;
assign LUT_3[40158] = 32'b00000000000000001111010011010000;
assign LUT_3[40159] = 32'b00000000000000010101111110101101;
assign LUT_3[40160] = 32'b00000000000000001000100000001101;
assign LUT_3[40161] = 32'b00000000000000001111001011101010;
assign LUT_3[40162] = 32'b00000000000000001010100111110001;
assign LUT_3[40163] = 32'b00000000000000010001010011001110;
assign LUT_3[40164] = 32'b00000000000000000101101110000011;
assign LUT_3[40165] = 32'b00000000000000001100011001100000;
assign LUT_3[40166] = 32'b00000000000000000111110101100111;
assign LUT_3[40167] = 32'b00000000000000001110100001000100;
assign LUT_3[40168] = 32'b00000000000000001101111001010011;
assign LUT_3[40169] = 32'b00000000000000010100100100110000;
assign LUT_3[40170] = 32'b00000000000000010000000000110111;
assign LUT_3[40171] = 32'b00000000000000010110101100010100;
assign LUT_3[40172] = 32'b00000000000000001011000111001001;
assign LUT_3[40173] = 32'b00000000000000010001110010100110;
assign LUT_3[40174] = 32'b00000000000000001101001110101101;
assign LUT_3[40175] = 32'b00000000000000010011111010001010;
assign LUT_3[40176] = 32'b00000000000000001011110011010000;
assign LUT_3[40177] = 32'b00000000000000010010011110101101;
assign LUT_3[40178] = 32'b00000000000000001101111010110100;
assign LUT_3[40179] = 32'b00000000000000010100100110010001;
assign LUT_3[40180] = 32'b00000000000000001001000001000110;
assign LUT_3[40181] = 32'b00000000000000001111101100100011;
assign LUT_3[40182] = 32'b00000000000000001011001000101010;
assign LUT_3[40183] = 32'b00000000000000010001110100000111;
assign LUT_3[40184] = 32'b00000000000000010001001100010110;
assign LUT_3[40185] = 32'b00000000000000010111110111110011;
assign LUT_3[40186] = 32'b00000000000000010011010011111010;
assign LUT_3[40187] = 32'b00000000000000011001111111010111;
assign LUT_3[40188] = 32'b00000000000000001110011010001100;
assign LUT_3[40189] = 32'b00000000000000010101000101101001;
assign LUT_3[40190] = 32'b00000000000000010000100001110000;
assign LUT_3[40191] = 32'b00000000000000010111001101001101;
assign LUT_3[40192] = 32'b00000000000000000001011101100101;
assign LUT_3[40193] = 32'b00000000000000001000001001000010;
assign LUT_3[40194] = 32'b00000000000000000011100101001001;
assign LUT_3[40195] = 32'b00000000000000001010010000100110;
assign LUT_3[40196] = 32'b11111111111111111110101011011011;
assign LUT_3[40197] = 32'b00000000000000000101010110111000;
assign LUT_3[40198] = 32'b00000000000000000000110010111111;
assign LUT_3[40199] = 32'b00000000000000000111011110011100;
assign LUT_3[40200] = 32'b00000000000000000110110110101011;
assign LUT_3[40201] = 32'b00000000000000001101100010001000;
assign LUT_3[40202] = 32'b00000000000000001000111110001111;
assign LUT_3[40203] = 32'b00000000000000001111101001101100;
assign LUT_3[40204] = 32'b00000000000000000100000100100001;
assign LUT_3[40205] = 32'b00000000000000001010101111111110;
assign LUT_3[40206] = 32'b00000000000000000110001100000101;
assign LUT_3[40207] = 32'b00000000000000001100110111100010;
assign LUT_3[40208] = 32'b00000000000000000100110000101000;
assign LUT_3[40209] = 32'b00000000000000001011011100000101;
assign LUT_3[40210] = 32'b00000000000000000110111000001100;
assign LUT_3[40211] = 32'b00000000000000001101100011101001;
assign LUT_3[40212] = 32'b00000000000000000001111110011110;
assign LUT_3[40213] = 32'b00000000000000001000101001111011;
assign LUT_3[40214] = 32'b00000000000000000100000110000010;
assign LUT_3[40215] = 32'b00000000000000001010110001011111;
assign LUT_3[40216] = 32'b00000000000000001010001001101110;
assign LUT_3[40217] = 32'b00000000000000010000110101001011;
assign LUT_3[40218] = 32'b00000000000000001100010001010010;
assign LUT_3[40219] = 32'b00000000000000010010111100101111;
assign LUT_3[40220] = 32'b00000000000000000111010111100100;
assign LUT_3[40221] = 32'b00000000000000001110000011000001;
assign LUT_3[40222] = 32'b00000000000000001001011111001000;
assign LUT_3[40223] = 32'b00000000000000010000001010100101;
assign LUT_3[40224] = 32'b00000000000000000010101100000101;
assign LUT_3[40225] = 32'b00000000000000001001010111100010;
assign LUT_3[40226] = 32'b00000000000000000100110011101001;
assign LUT_3[40227] = 32'b00000000000000001011011111000110;
assign LUT_3[40228] = 32'b11111111111111111111111001111011;
assign LUT_3[40229] = 32'b00000000000000000110100101011000;
assign LUT_3[40230] = 32'b00000000000000000010000001011111;
assign LUT_3[40231] = 32'b00000000000000001000101100111100;
assign LUT_3[40232] = 32'b00000000000000001000000101001011;
assign LUT_3[40233] = 32'b00000000000000001110110000101000;
assign LUT_3[40234] = 32'b00000000000000001010001100101111;
assign LUT_3[40235] = 32'b00000000000000010000111000001100;
assign LUT_3[40236] = 32'b00000000000000000101010011000001;
assign LUT_3[40237] = 32'b00000000000000001011111110011110;
assign LUT_3[40238] = 32'b00000000000000000111011010100101;
assign LUT_3[40239] = 32'b00000000000000001110000110000010;
assign LUT_3[40240] = 32'b00000000000000000101111111001000;
assign LUT_3[40241] = 32'b00000000000000001100101010100101;
assign LUT_3[40242] = 32'b00000000000000001000000110101100;
assign LUT_3[40243] = 32'b00000000000000001110110010001001;
assign LUT_3[40244] = 32'b00000000000000000011001100111110;
assign LUT_3[40245] = 32'b00000000000000001001111000011011;
assign LUT_3[40246] = 32'b00000000000000000101010100100010;
assign LUT_3[40247] = 32'b00000000000000001011111111111111;
assign LUT_3[40248] = 32'b00000000000000001011011000001110;
assign LUT_3[40249] = 32'b00000000000000010010000011101011;
assign LUT_3[40250] = 32'b00000000000000001101011111110010;
assign LUT_3[40251] = 32'b00000000000000010100001011001111;
assign LUT_3[40252] = 32'b00000000000000001000100110000100;
assign LUT_3[40253] = 32'b00000000000000001111010001100001;
assign LUT_3[40254] = 32'b00000000000000001010101101101000;
assign LUT_3[40255] = 32'b00000000000000010001011001000101;
assign LUT_3[40256] = 32'b00000000000000000001010110010000;
assign LUT_3[40257] = 32'b00000000000000001000000001101101;
assign LUT_3[40258] = 32'b00000000000000000011011101110100;
assign LUT_3[40259] = 32'b00000000000000001010001001010001;
assign LUT_3[40260] = 32'b11111111111111111110100100000110;
assign LUT_3[40261] = 32'b00000000000000000101001111100011;
assign LUT_3[40262] = 32'b00000000000000000000101011101010;
assign LUT_3[40263] = 32'b00000000000000000111010111000111;
assign LUT_3[40264] = 32'b00000000000000000110101111010110;
assign LUT_3[40265] = 32'b00000000000000001101011010110011;
assign LUT_3[40266] = 32'b00000000000000001000110110111010;
assign LUT_3[40267] = 32'b00000000000000001111100010010111;
assign LUT_3[40268] = 32'b00000000000000000011111101001100;
assign LUT_3[40269] = 32'b00000000000000001010101000101001;
assign LUT_3[40270] = 32'b00000000000000000110000100110000;
assign LUT_3[40271] = 32'b00000000000000001100110000001101;
assign LUT_3[40272] = 32'b00000000000000000100101001010011;
assign LUT_3[40273] = 32'b00000000000000001011010100110000;
assign LUT_3[40274] = 32'b00000000000000000110110000110111;
assign LUT_3[40275] = 32'b00000000000000001101011100010100;
assign LUT_3[40276] = 32'b00000000000000000001110111001001;
assign LUT_3[40277] = 32'b00000000000000001000100010100110;
assign LUT_3[40278] = 32'b00000000000000000011111110101101;
assign LUT_3[40279] = 32'b00000000000000001010101010001010;
assign LUT_3[40280] = 32'b00000000000000001010000010011001;
assign LUT_3[40281] = 32'b00000000000000010000101101110110;
assign LUT_3[40282] = 32'b00000000000000001100001001111101;
assign LUT_3[40283] = 32'b00000000000000010010110101011010;
assign LUT_3[40284] = 32'b00000000000000000111010000001111;
assign LUT_3[40285] = 32'b00000000000000001101111011101100;
assign LUT_3[40286] = 32'b00000000000000001001010111110011;
assign LUT_3[40287] = 32'b00000000000000010000000011010000;
assign LUT_3[40288] = 32'b00000000000000000010100100110000;
assign LUT_3[40289] = 32'b00000000000000001001010000001101;
assign LUT_3[40290] = 32'b00000000000000000100101100010100;
assign LUT_3[40291] = 32'b00000000000000001011010111110001;
assign LUT_3[40292] = 32'b11111111111111111111110010100110;
assign LUT_3[40293] = 32'b00000000000000000110011110000011;
assign LUT_3[40294] = 32'b00000000000000000001111010001010;
assign LUT_3[40295] = 32'b00000000000000001000100101100111;
assign LUT_3[40296] = 32'b00000000000000000111111101110110;
assign LUT_3[40297] = 32'b00000000000000001110101001010011;
assign LUT_3[40298] = 32'b00000000000000001010000101011010;
assign LUT_3[40299] = 32'b00000000000000010000110000110111;
assign LUT_3[40300] = 32'b00000000000000000101001011101100;
assign LUT_3[40301] = 32'b00000000000000001011110111001001;
assign LUT_3[40302] = 32'b00000000000000000111010011010000;
assign LUT_3[40303] = 32'b00000000000000001101111110101101;
assign LUT_3[40304] = 32'b00000000000000000101110111110011;
assign LUT_3[40305] = 32'b00000000000000001100100011010000;
assign LUT_3[40306] = 32'b00000000000000000111111111010111;
assign LUT_3[40307] = 32'b00000000000000001110101010110100;
assign LUT_3[40308] = 32'b00000000000000000011000101101001;
assign LUT_3[40309] = 32'b00000000000000001001110001000110;
assign LUT_3[40310] = 32'b00000000000000000101001101001101;
assign LUT_3[40311] = 32'b00000000000000001011111000101010;
assign LUT_3[40312] = 32'b00000000000000001011010000111001;
assign LUT_3[40313] = 32'b00000000000000010001111100010110;
assign LUT_3[40314] = 32'b00000000000000001101011000011101;
assign LUT_3[40315] = 32'b00000000000000010100000011111010;
assign LUT_3[40316] = 32'b00000000000000001000011110101111;
assign LUT_3[40317] = 32'b00000000000000001111001010001100;
assign LUT_3[40318] = 32'b00000000000000001010100110010011;
assign LUT_3[40319] = 32'b00000000000000010001010001110000;
assign LUT_3[40320] = 32'b00000000000000000011101000100011;
assign LUT_3[40321] = 32'b00000000000000001010010100000000;
assign LUT_3[40322] = 32'b00000000000000000101110000000111;
assign LUT_3[40323] = 32'b00000000000000001100011011100100;
assign LUT_3[40324] = 32'b00000000000000000000110110011001;
assign LUT_3[40325] = 32'b00000000000000000111100001110110;
assign LUT_3[40326] = 32'b00000000000000000010111101111101;
assign LUT_3[40327] = 32'b00000000000000001001101001011010;
assign LUT_3[40328] = 32'b00000000000000001001000001101001;
assign LUT_3[40329] = 32'b00000000000000001111101101000110;
assign LUT_3[40330] = 32'b00000000000000001011001001001101;
assign LUT_3[40331] = 32'b00000000000000010001110100101010;
assign LUT_3[40332] = 32'b00000000000000000110001111011111;
assign LUT_3[40333] = 32'b00000000000000001100111010111100;
assign LUT_3[40334] = 32'b00000000000000001000010111000011;
assign LUT_3[40335] = 32'b00000000000000001111000010100000;
assign LUT_3[40336] = 32'b00000000000000000110111011100110;
assign LUT_3[40337] = 32'b00000000000000001101100111000011;
assign LUT_3[40338] = 32'b00000000000000001001000011001010;
assign LUT_3[40339] = 32'b00000000000000001111101110100111;
assign LUT_3[40340] = 32'b00000000000000000100001001011100;
assign LUT_3[40341] = 32'b00000000000000001010110100111001;
assign LUT_3[40342] = 32'b00000000000000000110010001000000;
assign LUT_3[40343] = 32'b00000000000000001100111100011101;
assign LUT_3[40344] = 32'b00000000000000001100010100101100;
assign LUT_3[40345] = 32'b00000000000000010011000000001001;
assign LUT_3[40346] = 32'b00000000000000001110011100010000;
assign LUT_3[40347] = 32'b00000000000000010101000111101101;
assign LUT_3[40348] = 32'b00000000000000001001100010100010;
assign LUT_3[40349] = 32'b00000000000000010000001101111111;
assign LUT_3[40350] = 32'b00000000000000001011101010000110;
assign LUT_3[40351] = 32'b00000000000000010010010101100011;
assign LUT_3[40352] = 32'b00000000000000000100110111000011;
assign LUT_3[40353] = 32'b00000000000000001011100010100000;
assign LUT_3[40354] = 32'b00000000000000000110111110100111;
assign LUT_3[40355] = 32'b00000000000000001101101010000100;
assign LUT_3[40356] = 32'b00000000000000000010000100111001;
assign LUT_3[40357] = 32'b00000000000000001000110000010110;
assign LUT_3[40358] = 32'b00000000000000000100001100011101;
assign LUT_3[40359] = 32'b00000000000000001010110111111010;
assign LUT_3[40360] = 32'b00000000000000001010010000001001;
assign LUT_3[40361] = 32'b00000000000000010000111011100110;
assign LUT_3[40362] = 32'b00000000000000001100010111101101;
assign LUT_3[40363] = 32'b00000000000000010011000011001010;
assign LUT_3[40364] = 32'b00000000000000000111011101111111;
assign LUT_3[40365] = 32'b00000000000000001110001001011100;
assign LUT_3[40366] = 32'b00000000000000001001100101100011;
assign LUT_3[40367] = 32'b00000000000000010000010001000000;
assign LUT_3[40368] = 32'b00000000000000001000001010000110;
assign LUT_3[40369] = 32'b00000000000000001110110101100011;
assign LUT_3[40370] = 32'b00000000000000001010010001101010;
assign LUT_3[40371] = 32'b00000000000000010000111101000111;
assign LUT_3[40372] = 32'b00000000000000000101010111111100;
assign LUT_3[40373] = 32'b00000000000000001100000011011001;
assign LUT_3[40374] = 32'b00000000000000000111011111100000;
assign LUT_3[40375] = 32'b00000000000000001110001010111101;
assign LUT_3[40376] = 32'b00000000000000001101100011001100;
assign LUT_3[40377] = 32'b00000000000000010100001110101001;
assign LUT_3[40378] = 32'b00000000000000001111101010110000;
assign LUT_3[40379] = 32'b00000000000000010110010110001101;
assign LUT_3[40380] = 32'b00000000000000001010110001000010;
assign LUT_3[40381] = 32'b00000000000000010001011100011111;
assign LUT_3[40382] = 32'b00000000000000001100111000100110;
assign LUT_3[40383] = 32'b00000000000000010011100100000011;
assign LUT_3[40384] = 32'b00000000000000000011100001001110;
assign LUT_3[40385] = 32'b00000000000000001010001100101011;
assign LUT_3[40386] = 32'b00000000000000000101101000110010;
assign LUT_3[40387] = 32'b00000000000000001100010100001111;
assign LUT_3[40388] = 32'b00000000000000000000101111000100;
assign LUT_3[40389] = 32'b00000000000000000111011010100001;
assign LUT_3[40390] = 32'b00000000000000000010110110101000;
assign LUT_3[40391] = 32'b00000000000000001001100010000101;
assign LUT_3[40392] = 32'b00000000000000001000111010010100;
assign LUT_3[40393] = 32'b00000000000000001111100101110001;
assign LUT_3[40394] = 32'b00000000000000001011000001111000;
assign LUT_3[40395] = 32'b00000000000000010001101101010101;
assign LUT_3[40396] = 32'b00000000000000000110001000001010;
assign LUT_3[40397] = 32'b00000000000000001100110011100111;
assign LUT_3[40398] = 32'b00000000000000001000001111101110;
assign LUT_3[40399] = 32'b00000000000000001110111011001011;
assign LUT_3[40400] = 32'b00000000000000000110110100010001;
assign LUT_3[40401] = 32'b00000000000000001101011111101110;
assign LUT_3[40402] = 32'b00000000000000001000111011110101;
assign LUT_3[40403] = 32'b00000000000000001111100111010010;
assign LUT_3[40404] = 32'b00000000000000000100000010000111;
assign LUT_3[40405] = 32'b00000000000000001010101101100100;
assign LUT_3[40406] = 32'b00000000000000000110001001101011;
assign LUT_3[40407] = 32'b00000000000000001100110101001000;
assign LUT_3[40408] = 32'b00000000000000001100001101010111;
assign LUT_3[40409] = 32'b00000000000000010010111000110100;
assign LUT_3[40410] = 32'b00000000000000001110010100111011;
assign LUT_3[40411] = 32'b00000000000000010101000000011000;
assign LUT_3[40412] = 32'b00000000000000001001011011001101;
assign LUT_3[40413] = 32'b00000000000000010000000110101010;
assign LUT_3[40414] = 32'b00000000000000001011100010110001;
assign LUT_3[40415] = 32'b00000000000000010010001110001110;
assign LUT_3[40416] = 32'b00000000000000000100101111101110;
assign LUT_3[40417] = 32'b00000000000000001011011011001011;
assign LUT_3[40418] = 32'b00000000000000000110110111010010;
assign LUT_3[40419] = 32'b00000000000000001101100010101111;
assign LUT_3[40420] = 32'b00000000000000000001111101100100;
assign LUT_3[40421] = 32'b00000000000000001000101001000001;
assign LUT_3[40422] = 32'b00000000000000000100000101001000;
assign LUT_3[40423] = 32'b00000000000000001010110000100101;
assign LUT_3[40424] = 32'b00000000000000001010001000110100;
assign LUT_3[40425] = 32'b00000000000000010000110100010001;
assign LUT_3[40426] = 32'b00000000000000001100010000011000;
assign LUT_3[40427] = 32'b00000000000000010010111011110101;
assign LUT_3[40428] = 32'b00000000000000000111010110101010;
assign LUT_3[40429] = 32'b00000000000000001110000010000111;
assign LUT_3[40430] = 32'b00000000000000001001011110001110;
assign LUT_3[40431] = 32'b00000000000000010000001001101011;
assign LUT_3[40432] = 32'b00000000000000001000000010110001;
assign LUT_3[40433] = 32'b00000000000000001110101110001110;
assign LUT_3[40434] = 32'b00000000000000001010001010010101;
assign LUT_3[40435] = 32'b00000000000000010000110101110010;
assign LUT_3[40436] = 32'b00000000000000000101010000100111;
assign LUT_3[40437] = 32'b00000000000000001011111100000100;
assign LUT_3[40438] = 32'b00000000000000000111011000001011;
assign LUT_3[40439] = 32'b00000000000000001110000011101000;
assign LUT_3[40440] = 32'b00000000000000001101011011110111;
assign LUT_3[40441] = 32'b00000000000000010100000111010100;
assign LUT_3[40442] = 32'b00000000000000001111100011011011;
assign LUT_3[40443] = 32'b00000000000000010110001110111000;
assign LUT_3[40444] = 32'b00000000000000001010101001101101;
assign LUT_3[40445] = 32'b00000000000000010001010101001010;
assign LUT_3[40446] = 32'b00000000000000001100110001010001;
assign LUT_3[40447] = 32'b00000000000000010011011100101110;
assign LUT_3[40448] = 32'b00000000000000001000100011010000;
assign LUT_3[40449] = 32'b00000000000000001111001110101101;
assign LUT_3[40450] = 32'b00000000000000001010101010110100;
assign LUT_3[40451] = 32'b00000000000000010001010110010001;
assign LUT_3[40452] = 32'b00000000000000000101110001000110;
assign LUT_3[40453] = 32'b00000000000000001100011100100011;
assign LUT_3[40454] = 32'b00000000000000000111111000101010;
assign LUT_3[40455] = 32'b00000000000000001110100100000111;
assign LUT_3[40456] = 32'b00000000000000001101111100010110;
assign LUT_3[40457] = 32'b00000000000000010100100111110011;
assign LUT_3[40458] = 32'b00000000000000010000000011111010;
assign LUT_3[40459] = 32'b00000000000000010110101111010111;
assign LUT_3[40460] = 32'b00000000000000001011001010001100;
assign LUT_3[40461] = 32'b00000000000000010001110101101001;
assign LUT_3[40462] = 32'b00000000000000001101010001110000;
assign LUT_3[40463] = 32'b00000000000000010011111101001101;
assign LUT_3[40464] = 32'b00000000000000001011110110010011;
assign LUT_3[40465] = 32'b00000000000000010010100001110000;
assign LUT_3[40466] = 32'b00000000000000001101111101110111;
assign LUT_3[40467] = 32'b00000000000000010100101001010100;
assign LUT_3[40468] = 32'b00000000000000001001000100001001;
assign LUT_3[40469] = 32'b00000000000000001111101111100110;
assign LUT_3[40470] = 32'b00000000000000001011001011101101;
assign LUT_3[40471] = 32'b00000000000000010001110111001010;
assign LUT_3[40472] = 32'b00000000000000010001001111011001;
assign LUT_3[40473] = 32'b00000000000000010111111010110110;
assign LUT_3[40474] = 32'b00000000000000010011010110111101;
assign LUT_3[40475] = 32'b00000000000000011010000010011010;
assign LUT_3[40476] = 32'b00000000000000001110011101001111;
assign LUT_3[40477] = 32'b00000000000000010101001000101100;
assign LUT_3[40478] = 32'b00000000000000010000100100110011;
assign LUT_3[40479] = 32'b00000000000000010111010000010000;
assign LUT_3[40480] = 32'b00000000000000001001110001110000;
assign LUT_3[40481] = 32'b00000000000000010000011101001101;
assign LUT_3[40482] = 32'b00000000000000001011111001010100;
assign LUT_3[40483] = 32'b00000000000000010010100100110001;
assign LUT_3[40484] = 32'b00000000000000000110111111100110;
assign LUT_3[40485] = 32'b00000000000000001101101011000011;
assign LUT_3[40486] = 32'b00000000000000001001000111001010;
assign LUT_3[40487] = 32'b00000000000000001111110010100111;
assign LUT_3[40488] = 32'b00000000000000001111001010110110;
assign LUT_3[40489] = 32'b00000000000000010101110110010011;
assign LUT_3[40490] = 32'b00000000000000010001010010011010;
assign LUT_3[40491] = 32'b00000000000000010111111101110111;
assign LUT_3[40492] = 32'b00000000000000001100011000101100;
assign LUT_3[40493] = 32'b00000000000000010011000100001001;
assign LUT_3[40494] = 32'b00000000000000001110100000010000;
assign LUT_3[40495] = 32'b00000000000000010101001011101101;
assign LUT_3[40496] = 32'b00000000000000001101000100110011;
assign LUT_3[40497] = 32'b00000000000000010011110000010000;
assign LUT_3[40498] = 32'b00000000000000001111001100010111;
assign LUT_3[40499] = 32'b00000000000000010101110111110100;
assign LUT_3[40500] = 32'b00000000000000001010010010101001;
assign LUT_3[40501] = 32'b00000000000000010000111110000110;
assign LUT_3[40502] = 32'b00000000000000001100011010001101;
assign LUT_3[40503] = 32'b00000000000000010011000101101010;
assign LUT_3[40504] = 32'b00000000000000010010011101111001;
assign LUT_3[40505] = 32'b00000000000000011001001001010110;
assign LUT_3[40506] = 32'b00000000000000010100100101011101;
assign LUT_3[40507] = 32'b00000000000000011011010000111010;
assign LUT_3[40508] = 32'b00000000000000001111101011101111;
assign LUT_3[40509] = 32'b00000000000000010110010111001100;
assign LUT_3[40510] = 32'b00000000000000010001110011010011;
assign LUT_3[40511] = 32'b00000000000000011000011110110000;
assign LUT_3[40512] = 32'b00000000000000001000011011111011;
assign LUT_3[40513] = 32'b00000000000000001111000111011000;
assign LUT_3[40514] = 32'b00000000000000001010100011011111;
assign LUT_3[40515] = 32'b00000000000000010001001110111100;
assign LUT_3[40516] = 32'b00000000000000000101101001110001;
assign LUT_3[40517] = 32'b00000000000000001100010101001110;
assign LUT_3[40518] = 32'b00000000000000000111110001010101;
assign LUT_3[40519] = 32'b00000000000000001110011100110010;
assign LUT_3[40520] = 32'b00000000000000001101110101000001;
assign LUT_3[40521] = 32'b00000000000000010100100000011110;
assign LUT_3[40522] = 32'b00000000000000001111111100100101;
assign LUT_3[40523] = 32'b00000000000000010110101000000010;
assign LUT_3[40524] = 32'b00000000000000001011000010110111;
assign LUT_3[40525] = 32'b00000000000000010001101110010100;
assign LUT_3[40526] = 32'b00000000000000001101001010011011;
assign LUT_3[40527] = 32'b00000000000000010011110101111000;
assign LUT_3[40528] = 32'b00000000000000001011101110111110;
assign LUT_3[40529] = 32'b00000000000000010010011010011011;
assign LUT_3[40530] = 32'b00000000000000001101110110100010;
assign LUT_3[40531] = 32'b00000000000000010100100001111111;
assign LUT_3[40532] = 32'b00000000000000001000111100110100;
assign LUT_3[40533] = 32'b00000000000000001111101000010001;
assign LUT_3[40534] = 32'b00000000000000001011000100011000;
assign LUT_3[40535] = 32'b00000000000000010001101111110101;
assign LUT_3[40536] = 32'b00000000000000010001001000000100;
assign LUT_3[40537] = 32'b00000000000000010111110011100001;
assign LUT_3[40538] = 32'b00000000000000010011001111101000;
assign LUT_3[40539] = 32'b00000000000000011001111011000101;
assign LUT_3[40540] = 32'b00000000000000001110010101111010;
assign LUT_3[40541] = 32'b00000000000000010101000001010111;
assign LUT_3[40542] = 32'b00000000000000010000011101011110;
assign LUT_3[40543] = 32'b00000000000000010111001000111011;
assign LUT_3[40544] = 32'b00000000000000001001101010011011;
assign LUT_3[40545] = 32'b00000000000000010000010101111000;
assign LUT_3[40546] = 32'b00000000000000001011110001111111;
assign LUT_3[40547] = 32'b00000000000000010010011101011100;
assign LUT_3[40548] = 32'b00000000000000000110111000010001;
assign LUT_3[40549] = 32'b00000000000000001101100011101110;
assign LUT_3[40550] = 32'b00000000000000001000111111110101;
assign LUT_3[40551] = 32'b00000000000000001111101011010010;
assign LUT_3[40552] = 32'b00000000000000001111000011100001;
assign LUT_3[40553] = 32'b00000000000000010101101110111110;
assign LUT_3[40554] = 32'b00000000000000010001001011000101;
assign LUT_3[40555] = 32'b00000000000000010111110110100010;
assign LUT_3[40556] = 32'b00000000000000001100010001010111;
assign LUT_3[40557] = 32'b00000000000000010010111100110100;
assign LUT_3[40558] = 32'b00000000000000001110011000111011;
assign LUT_3[40559] = 32'b00000000000000010101000100011000;
assign LUT_3[40560] = 32'b00000000000000001100111101011110;
assign LUT_3[40561] = 32'b00000000000000010011101000111011;
assign LUT_3[40562] = 32'b00000000000000001111000101000010;
assign LUT_3[40563] = 32'b00000000000000010101110000011111;
assign LUT_3[40564] = 32'b00000000000000001010001011010100;
assign LUT_3[40565] = 32'b00000000000000010000110110110001;
assign LUT_3[40566] = 32'b00000000000000001100010010111000;
assign LUT_3[40567] = 32'b00000000000000010010111110010101;
assign LUT_3[40568] = 32'b00000000000000010010010110100100;
assign LUT_3[40569] = 32'b00000000000000011001000010000001;
assign LUT_3[40570] = 32'b00000000000000010100011110001000;
assign LUT_3[40571] = 32'b00000000000000011011001001100101;
assign LUT_3[40572] = 32'b00000000000000001111100100011010;
assign LUT_3[40573] = 32'b00000000000000010110001111110111;
assign LUT_3[40574] = 32'b00000000000000010001101011111110;
assign LUT_3[40575] = 32'b00000000000000011000010111011011;
assign LUT_3[40576] = 32'b00000000000000001010101110001110;
assign LUT_3[40577] = 32'b00000000000000010001011001101011;
assign LUT_3[40578] = 32'b00000000000000001100110101110010;
assign LUT_3[40579] = 32'b00000000000000010011100001001111;
assign LUT_3[40580] = 32'b00000000000000000111111100000100;
assign LUT_3[40581] = 32'b00000000000000001110100111100001;
assign LUT_3[40582] = 32'b00000000000000001010000011101000;
assign LUT_3[40583] = 32'b00000000000000010000101111000101;
assign LUT_3[40584] = 32'b00000000000000010000000111010100;
assign LUT_3[40585] = 32'b00000000000000010110110010110001;
assign LUT_3[40586] = 32'b00000000000000010010001110111000;
assign LUT_3[40587] = 32'b00000000000000011000111010010101;
assign LUT_3[40588] = 32'b00000000000000001101010101001010;
assign LUT_3[40589] = 32'b00000000000000010100000000100111;
assign LUT_3[40590] = 32'b00000000000000001111011100101110;
assign LUT_3[40591] = 32'b00000000000000010110001000001011;
assign LUT_3[40592] = 32'b00000000000000001110000001010001;
assign LUT_3[40593] = 32'b00000000000000010100101100101110;
assign LUT_3[40594] = 32'b00000000000000010000001000110101;
assign LUT_3[40595] = 32'b00000000000000010110110100010010;
assign LUT_3[40596] = 32'b00000000000000001011001111000111;
assign LUT_3[40597] = 32'b00000000000000010001111010100100;
assign LUT_3[40598] = 32'b00000000000000001101010110101011;
assign LUT_3[40599] = 32'b00000000000000010100000010001000;
assign LUT_3[40600] = 32'b00000000000000010011011010010111;
assign LUT_3[40601] = 32'b00000000000000011010000101110100;
assign LUT_3[40602] = 32'b00000000000000010101100001111011;
assign LUT_3[40603] = 32'b00000000000000011100001101011000;
assign LUT_3[40604] = 32'b00000000000000010000101000001101;
assign LUT_3[40605] = 32'b00000000000000010111010011101010;
assign LUT_3[40606] = 32'b00000000000000010010101111110001;
assign LUT_3[40607] = 32'b00000000000000011001011011001110;
assign LUT_3[40608] = 32'b00000000000000001011111100101110;
assign LUT_3[40609] = 32'b00000000000000010010101000001011;
assign LUT_3[40610] = 32'b00000000000000001110000100010010;
assign LUT_3[40611] = 32'b00000000000000010100101111101111;
assign LUT_3[40612] = 32'b00000000000000001001001010100100;
assign LUT_3[40613] = 32'b00000000000000001111110110000001;
assign LUT_3[40614] = 32'b00000000000000001011010010001000;
assign LUT_3[40615] = 32'b00000000000000010001111101100101;
assign LUT_3[40616] = 32'b00000000000000010001010101110100;
assign LUT_3[40617] = 32'b00000000000000011000000001010001;
assign LUT_3[40618] = 32'b00000000000000010011011101011000;
assign LUT_3[40619] = 32'b00000000000000011010001000110101;
assign LUT_3[40620] = 32'b00000000000000001110100011101010;
assign LUT_3[40621] = 32'b00000000000000010101001111000111;
assign LUT_3[40622] = 32'b00000000000000010000101011001110;
assign LUT_3[40623] = 32'b00000000000000010111010110101011;
assign LUT_3[40624] = 32'b00000000000000001111001111110001;
assign LUT_3[40625] = 32'b00000000000000010101111011001110;
assign LUT_3[40626] = 32'b00000000000000010001010111010101;
assign LUT_3[40627] = 32'b00000000000000011000000010110010;
assign LUT_3[40628] = 32'b00000000000000001100011101100111;
assign LUT_3[40629] = 32'b00000000000000010011001001000100;
assign LUT_3[40630] = 32'b00000000000000001110100101001011;
assign LUT_3[40631] = 32'b00000000000000010101010000101000;
assign LUT_3[40632] = 32'b00000000000000010100101000110111;
assign LUT_3[40633] = 32'b00000000000000011011010100010100;
assign LUT_3[40634] = 32'b00000000000000010110110000011011;
assign LUT_3[40635] = 32'b00000000000000011101011011111000;
assign LUT_3[40636] = 32'b00000000000000010001110110101101;
assign LUT_3[40637] = 32'b00000000000000011000100010001010;
assign LUT_3[40638] = 32'b00000000000000010011111110010001;
assign LUT_3[40639] = 32'b00000000000000011010101001101110;
assign LUT_3[40640] = 32'b00000000000000001010100110111001;
assign LUT_3[40641] = 32'b00000000000000010001010010010110;
assign LUT_3[40642] = 32'b00000000000000001100101110011101;
assign LUT_3[40643] = 32'b00000000000000010011011001111010;
assign LUT_3[40644] = 32'b00000000000000000111110100101111;
assign LUT_3[40645] = 32'b00000000000000001110100000001100;
assign LUT_3[40646] = 32'b00000000000000001001111100010011;
assign LUT_3[40647] = 32'b00000000000000010000100111110000;
assign LUT_3[40648] = 32'b00000000000000001111111111111111;
assign LUT_3[40649] = 32'b00000000000000010110101011011100;
assign LUT_3[40650] = 32'b00000000000000010010000111100011;
assign LUT_3[40651] = 32'b00000000000000011000110011000000;
assign LUT_3[40652] = 32'b00000000000000001101001101110101;
assign LUT_3[40653] = 32'b00000000000000010011111001010010;
assign LUT_3[40654] = 32'b00000000000000001111010101011001;
assign LUT_3[40655] = 32'b00000000000000010110000000110110;
assign LUT_3[40656] = 32'b00000000000000001101111001111100;
assign LUT_3[40657] = 32'b00000000000000010100100101011001;
assign LUT_3[40658] = 32'b00000000000000010000000001100000;
assign LUT_3[40659] = 32'b00000000000000010110101100111101;
assign LUT_3[40660] = 32'b00000000000000001011000111110010;
assign LUT_3[40661] = 32'b00000000000000010001110011001111;
assign LUT_3[40662] = 32'b00000000000000001101001111010110;
assign LUT_3[40663] = 32'b00000000000000010011111010110011;
assign LUT_3[40664] = 32'b00000000000000010011010011000010;
assign LUT_3[40665] = 32'b00000000000000011001111110011111;
assign LUT_3[40666] = 32'b00000000000000010101011010100110;
assign LUT_3[40667] = 32'b00000000000000011100000110000011;
assign LUT_3[40668] = 32'b00000000000000010000100000111000;
assign LUT_3[40669] = 32'b00000000000000010111001100010101;
assign LUT_3[40670] = 32'b00000000000000010010101000011100;
assign LUT_3[40671] = 32'b00000000000000011001010011111001;
assign LUT_3[40672] = 32'b00000000000000001011110101011001;
assign LUT_3[40673] = 32'b00000000000000010010100000110110;
assign LUT_3[40674] = 32'b00000000000000001101111100111101;
assign LUT_3[40675] = 32'b00000000000000010100101000011010;
assign LUT_3[40676] = 32'b00000000000000001001000011001111;
assign LUT_3[40677] = 32'b00000000000000001111101110101100;
assign LUT_3[40678] = 32'b00000000000000001011001010110011;
assign LUT_3[40679] = 32'b00000000000000010001110110010000;
assign LUT_3[40680] = 32'b00000000000000010001001110011111;
assign LUT_3[40681] = 32'b00000000000000010111111001111100;
assign LUT_3[40682] = 32'b00000000000000010011010110000011;
assign LUT_3[40683] = 32'b00000000000000011010000001100000;
assign LUT_3[40684] = 32'b00000000000000001110011100010101;
assign LUT_3[40685] = 32'b00000000000000010101000111110010;
assign LUT_3[40686] = 32'b00000000000000010000100011111001;
assign LUT_3[40687] = 32'b00000000000000010111001111010110;
assign LUT_3[40688] = 32'b00000000000000001111001000011100;
assign LUT_3[40689] = 32'b00000000000000010101110011111001;
assign LUT_3[40690] = 32'b00000000000000010001010000000000;
assign LUT_3[40691] = 32'b00000000000000010111111011011101;
assign LUT_3[40692] = 32'b00000000000000001100010110010010;
assign LUT_3[40693] = 32'b00000000000000010011000001101111;
assign LUT_3[40694] = 32'b00000000000000001110011101110110;
assign LUT_3[40695] = 32'b00000000000000010101001001010011;
assign LUT_3[40696] = 32'b00000000000000010100100001100010;
assign LUT_3[40697] = 32'b00000000000000011011001100111111;
assign LUT_3[40698] = 32'b00000000000000010110101001000110;
assign LUT_3[40699] = 32'b00000000000000011101010100100011;
assign LUT_3[40700] = 32'b00000000000000010001101111011000;
assign LUT_3[40701] = 32'b00000000000000011000011010110101;
assign LUT_3[40702] = 32'b00000000000000010011110110111100;
assign LUT_3[40703] = 32'b00000000000000011010100010011001;
assign LUT_3[40704] = 32'b00000000000000000100110010110001;
assign LUT_3[40705] = 32'b00000000000000001011011110001110;
assign LUT_3[40706] = 32'b00000000000000000110111010010101;
assign LUT_3[40707] = 32'b00000000000000001101100101110010;
assign LUT_3[40708] = 32'b00000000000000000010000000100111;
assign LUT_3[40709] = 32'b00000000000000001000101100000100;
assign LUT_3[40710] = 32'b00000000000000000100001000001011;
assign LUT_3[40711] = 32'b00000000000000001010110011101000;
assign LUT_3[40712] = 32'b00000000000000001010001011110111;
assign LUT_3[40713] = 32'b00000000000000010000110111010100;
assign LUT_3[40714] = 32'b00000000000000001100010011011011;
assign LUT_3[40715] = 32'b00000000000000010010111110111000;
assign LUT_3[40716] = 32'b00000000000000000111011001101101;
assign LUT_3[40717] = 32'b00000000000000001110000101001010;
assign LUT_3[40718] = 32'b00000000000000001001100001010001;
assign LUT_3[40719] = 32'b00000000000000010000001100101110;
assign LUT_3[40720] = 32'b00000000000000001000000101110100;
assign LUT_3[40721] = 32'b00000000000000001110110001010001;
assign LUT_3[40722] = 32'b00000000000000001010001101011000;
assign LUT_3[40723] = 32'b00000000000000010000111000110101;
assign LUT_3[40724] = 32'b00000000000000000101010011101010;
assign LUT_3[40725] = 32'b00000000000000001011111111000111;
assign LUT_3[40726] = 32'b00000000000000000111011011001110;
assign LUT_3[40727] = 32'b00000000000000001110000110101011;
assign LUT_3[40728] = 32'b00000000000000001101011110111010;
assign LUT_3[40729] = 32'b00000000000000010100001010010111;
assign LUT_3[40730] = 32'b00000000000000001111100110011110;
assign LUT_3[40731] = 32'b00000000000000010110010001111011;
assign LUT_3[40732] = 32'b00000000000000001010101100110000;
assign LUT_3[40733] = 32'b00000000000000010001011000001101;
assign LUT_3[40734] = 32'b00000000000000001100110100010100;
assign LUT_3[40735] = 32'b00000000000000010011011111110001;
assign LUT_3[40736] = 32'b00000000000000000110000001010001;
assign LUT_3[40737] = 32'b00000000000000001100101100101110;
assign LUT_3[40738] = 32'b00000000000000001000001000110101;
assign LUT_3[40739] = 32'b00000000000000001110110100010010;
assign LUT_3[40740] = 32'b00000000000000000011001111000111;
assign LUT_3[40741] = 32'b00000000000000001001111010100100;
assign LUT_3[40742] = 32'b00000000000000000101010110101011;
assign LUT_3[40743] = 32'b00000000000000001100000010001000;
assign LUT_3[40744] = 32'b00000000000000001011011010010111;
assign LUT_3[40745] = 32'b00000000000000010010000101110100;
assign LUT_3[40746] = 32'b00000000000000001101100001111011;
assign LUT_3[40747] = 32'b00000000000000010100001101011000;
assign LUT_3[40748] = 32'b00000000000000001000101000001101;
assign LUT_3[40749] = 32'b00000000000000001111010011101010;
assign LUT_3[40750] = 32'b00000000000000001010101111110001;
assign LUT_3[40751] = 32'b00000000000000010001011011001110;
assign LUT_3[40752] = 32'b00000000000000001001010100010100;
assign LUT_3[40753] = 32'b00000000000000001111111111110001;
assign LUT_3[40754] = 32'b00000000000000001011011011111000;
assign LUT_3[40755] = 32'b00000000000000010010000111010101;
assign LUT_3[40756] = 32'b00000000000000000110100010001010;
assign LUT_3[40757] = 32'b00000000000000001101001101100111;
assign LUT_3[40758] = 32'b00000000000000001000101001101110;
assign LUT_3[40759] = 32'b00000000000000001111010101001011;
assign LUT_3[40760] = 32'b00000000000000001110101101011010;
assign LUT_3[40761] = 32'b00000000000000010101011000110111;
assign LUT_3[40762] = 32'b00000000000000010000110100111110;
assign LUT_3[40763] = 32'b00000000000000010111100000011011;
assign LUT_3[40764] = 32'b00000000000000001011111011010000;
assign LUT_3[40765] = 32'b00000000000000010010100110101101;
assign LUT_3[40766] = 32'b00000000000000001110000010110100;
assign LUT_3[40767] = 32'b00000000000000010100101110010001;
assign LUT_3[40768] = 32'b00000000000000000100101011011100;
assign LUT_3[40769] = 32'b00000000000000001011010110111001;
assign LUT_3[40770] = 32'b00000000000000000110110011000000;
assign LUT_3[40771] = 32'b00000000000000001101011110011101;
assign LUT_3[40772] = 32'b00000000000000000001111001010010;
assign LUT_3[40773] = 32'b00000000000000001000100100101111;
assign LUT_3[40774] = 32'b00000000000000000100000000110110;
assign LUT_3[40775] = 32'b00000000000000001010101100010011;
assign LUT_3[40776] = 32'b00000000000000001010000100100010;
assign LUT_3[40777] = 32'b00000000000000010000101111111111;
assign LUT_3[40778] = 32'b00000000000000001100001100000110;
assign LUT_3[40779] = 32'b00000000000000010010110111100011;
assign LUT_3[40780] = 32'b00000000000000000111010010011000;
assign LUT_3[40781] = 32'b00000000000000001101111101110101;
assign LUT_3[40782] = 32'b00000000000000001001011001111100;
assign LUT_3[40783] = 32'b00000000000000010000000101011001;
assign LUT_3[40784] = 32'b00000000000000000111111110011111;
assign LUT_3[40785] = 32'b00000000000000001110101001111100;
assign LUT_3[40786] = 32'b00000000000000001010000110000011;
assign LUT_3[40787] = 32'b00000000000000010000110001100000;
assign LUT_3[40788] = 32'b00000000000000000101001100010101;
assign LUT_3[40789] = 32'b00000000000000001011110111110010;
assign LUT_3[40790] = 32'b00000000000000000111010011111001;
assign LUT_3[40791] = 32'b00000000000000001101111111010110;
assign LUT_3[40792] = 32'b00000000000000001101010111100101;
assign LUT_3[40793] = 32'b00000000000000010100000011000010;
assign LUT_3[40794] = 32'b00000000000000001111011111001001;
assign LUT_3[40795] = 32'b00000000000000010110001010100110;
assign LUT_3[40796] = 32'b00000000000000001010100101011011;
assign LUT_3[40797] = 32'b00000000000000010001010000111000;
assign LUT_3[40798] = 32'b00000000000000001100101100111111;
assign LUT_3[40799] = 32'b00000000000000010011011000011100;
assign LUT_3[40800] = 32'b00000000000000000101111001111100;
assign LUT_3[40801] = 32'b00000000000000001100100101011001;
assign LUT_3[40802] = 32'b00000000000000001000000001100000;
assign LUT_3[40803] = 32'b00000000000000001110101100111101;
assign LUT_3[40804] = 32'b00000000000000000011000111110010;
assign LUT_3[40805] = 32'b00000000000000001001110011001111;
assign LUT_3[40806] = 32'b00000000000000000101001111010110;
assign LUT_3[40807] = 32'b00000000000000001011111010110011;
assign LUT_3[40808] = 32'b00000000000000001011010011000010;
assign LUT_3[40809] = 32'b00000000000000010001111110011111;
assign LUT_3[40810] = 32'b00000000000000001101011010100110;
assign LUT_3[40811] = 32'b00000000000000010100000110000011;
assign LUT_3[40812] = 32'b00000000000000001000100000111000;
assign LUT_3[40813] = 32'b00000000000000001111001100010101;
assign LUT_3[40814] = 32'b00000000000000001010101000011100;
assign LUT_3[40815] = 32'b00000000000000010001010011111001;
assign LUT_3[40816] = 32'b00000000000000001001001100111111;
assign LUT_3[40817] = 32'b00000000000000001111111000011100;
assign LUT_3[40818] = 32'b00000000000000001011010100100011;
assign LUT_3[40819] = 32'b00000000000000010010000000000000;
assign LUT_3[40820] = 32'b00000000000000000110011010110101;
assign LUT_3[40821] = 32'b00000000000000001101000110010010;
assign LUT_3[40822] = 32'b00000000000000001000100010011001;
assign LUT_3[40823] = 32'b00000000000000001111001101110110;
assign LUT_3[40824] = 32'b00000000000000001110100110000101;
assign LUT_3[40825] = 32'b00000000000000010101010001100010;
assign LUT_3[40826] = 32'b00000000000000010000101101101001;
assign LUT_3[40827] = 32'b00000000000000010111011001000110;
assign LUT_3[40828] = 32'b00000000000000001011110011111011;
assign LUT_3[40829] = 32'b00000000000000010010011111011000;
assign LUT_3[40830] = 32'b00000000000000001101111011011111;
assign LUT_3[40831] = 32'b00000000000000010100100110111100;
assign LUT_3[40832] = 32'b00000000000000000110111101101111;
assign LUT_3[40833] = 32'b00000000000000001101101001001100;
assign LUT_3[40834] = 32'b00000000000000001001000101010011;
assign LUT_3[40835] = 32'b00000000000000001111110000110000;
assign LUT_3[40836] = 32'b00000000000000000100001011100101;
assign LUT_3[40837] = 32'b00000000000000001010110111000010;
assign LUT_3[40838] = 32'b00000000000000000110010011001001;
assign LUT_3[40839] = 32'b00000000000000001100111110100110;
assign LUT_3[40840] = 32'b00000000000000001100010110110101;
assign LUT_3[40841] = 32'b00000000000000010011000010010010;
assign LUT_3[40842] = 32'b00000000000000001110011110011001;
assign LUT_3[40843] = 32'b00000000000000010101001001110110;
assign LUT_3[40844] = 32'b00000000000000001001100100101011;
assign LUT_3[40845] = 32'b00000000000000010000010000001000;
assign LUT_3[40846] = 32'b00000000000000001011101100001111;
assign LUT_3[40847] = 32'b00000000000000010010010111101100;
assign LUT_3[40848] = 32'b00000000000000001010010000110010;
assign LUT_3[40849] = 32'b00000000000000010000111100001111;
assign LUT_3[40850] = 32'b00000000000000001100011000010110;
assign LUT_3[40851] = 32'b00000000000000010011000011110011;
assign LUT_3[40852] = 32'b00000000000000000111011110101000;
assign LUT_3[40853] = 32'b00000000000000001110001010000101;
assign LUT_3[40854] = 32'b00000000000000001001100110001100;
assign LUT_3[40855] = 32'b00000000000000010000010001101001;
assign LUT_3[40856] = 32'b00000000000000001111101001111000;
assign LUT_3[40857] = 32'b00000000000000010110010101010101;
assign LUT_3[40858] = 32'b00000000000000010001110001011100;
assign LUT_3[40859] = 32'b00000000000000011000011100111001;
assign LUT_3[40860] = 32'b00000000000000001100110111101110;
assign LUT_3[40861] = 32'b00000000000000010011100011001011;
assign LUT_3[40862] = 32'b00000000000000001110111111010010;
assign LUT_3[40863] = 32'b00000000000000010101101010101111;
assign LUT_3[40864] = 32'b00000000000000001000001100001111;
assign LUT_3[40865] = 32'b00000000000000001110110111101100;
assign LUT_3[40866] = 32'b00000000000000001010010011110011;
assign LUT_3[40867] = 32'b00000000000000010000111111010000;
assign LUT_3[40868] = 32'b00000000000000000101011010000101;
assign LUT_3[40869] = 32'b00000000000000001100000101100010;
assign LUT_3[40870] = 32'b00000000000000000111100001101001;
assign LUT_3[40871] = 32'b00000000000000001110001101000110;
assign LUT_3[40872] = 32'b00000000000000001101100101010101;
assign LUT_3[40873] = 32'b00000000000000010100010000110010;
assign LUT_3[40874] = 32'b00000000000000001111101100111001;
assign LUT_3[40875] = 32'b00000000000000010110011000010110;
assign LUT_3[40876] = 32'b00000000000000001010110011001011;
assign LUT_3[40877] = 32'b00000000000000010001011110101000;
assign LUT_3[40878] = 32'b00000000000000001100111010101111;
assign LUT_3[40879] = 32'b00000000000000010011100110001100;
assign LUT_3[40880] = 32'b00000000000000001011011111010010;
assign LUT_3[40881] = 32'b00000000000000010010001010101111;
assign LUT_3[40882] = 32'b00000000000000001101100110110110;
assign LUT_3[40883] = 32'b00000000000000010100010010010011;
assign LUT_3[40884] = 32'b00000000000000001000101101001000;
assign LUT_3[40885] = 32'b00000000000000001111011000100101;
assign LUT_3[40886] = 32'b00000000000000001010110100101100;
assign LUT_3[40887] = 32'b00000000000000010001100000001001;
assign LUT_3[40888] = 32'b00000000000000010000111000011000;
assign LUT_3[40889] = 32'b00000000000000010111100011110101;
assign LUT_3[40890] = 32'b00000000000000010010111111111100;
assign LUT_3[40891] = 32'b00000000000000011001101011011001;
assign LUT_3[40892] = 32'b00000000000000001110000110001110;
assign LUT_3[40893] = 32'b00000000000000010100110001101011;
assign LUT_3[40894] = 32'b00000000000000010000001101110010;
assign LUT_3[40895] = 32'b00000000000000010110111001001111;
assign LUT_3[40896] = 32'b00000000000000000110110110011010;
assign LUT_3[40897] = 32'b00000000000000001101100001110111;
assign LUT_3[40898] = 32'b00000000000000001000111101111110;
assign LUT_3[40899] = 32'b00000000000000001111101001011011;
assign LUT_3[40900] = 32'b00000000000000000100000100010000;
assign LUT_3[40901] = 32'b00000000000000001010101111101101;
assign LUT_3[40902] = 32'b00000000000000000110001011110100;
assign LUT_3[40903] = 32'b00000000000000001100110111010001;
assign LUT_3[40904] = 32'b00000000000000001100001111100000;
assign LUT_3[40905] = 32'b00000000000000010010111010111101;
assign LUT_3[40906] = 32'b00000000000000001110010111000100;
assign LUT_3[40907] = 32'b00000000000000010101000010100001;
assign LUT_3[40908] = 32'b00000000000000001001011101010110;
assign LUT_3[40909] = 32'b00000000000000010000001000110011;
assign LUT_3[40910] = 32'b00000000000000001011100100111010;
assign LUT_3[40911] = 32'b00000000000000010010010000010111;
assign LUT_3[40912] = 32'b00000000000000001010001001011101;
assign LUT_3[40913] = 32'b00000000000000010000110100111010;
assign LUT_3[40914] = 32'b00000000000000001100010001000001;
assign LUT_3[40915] = 32'b00000000000000010010111100011110;
assign LUT_3[40916] = 32'b00000000000000000111010111010011;
assign LUT_3[40917] = 32'b00000000000000001110000010110000;
assign LUT_3[40918] = 32'b00000000000000001001011110110111;
assign LUT_3[40919] = 32'b00000000000000010000001010010100;
assign LUT_3[40920] = 32'b00000000000000001111100010100011;
assign LUT_3[40921] = 32'b00000000000000010110001110000000;
assign LUT_3[40922] = 32'b00000000000000010001101010000111;
assign LUT_3[40923] = 32'b00000000000000011000010101100100;
assign LUT_3[40924] = 32'b00000000000000001100110000011001;
assign LUT_3[40925] = 32'b00000000000000010011011011110110;
assign LUT_3[40926] = 32'b00000000000000001110110111111101;
assign LUT_3[40927] = 32'b00000000000000010101100011011010;
assign LUT_3[40928] = 32'b00000000000000001000000100111010;
assign LUT_3[40929] = 32'b00000000000000001110110000010111;
assign LUT_3[40930] = 32'b00000000000000001010001100011110;
assign LUT_3[40931] = 32'b00000000000000010000110111111011;
assign LUT_3[40932] = 32'b00000000000000000101010010110000;
assign LUT_3[40933] = 32'b00000000000000001011111110001101;
assign LUT_3[40934] = 32'b00000000000000000111011010010100;
assign LUT_3[40935] = 32'b00000000000000001110000101110001;
assign LUT_3[40936] = 32'b00000000000000001101011110000000;
assign LUT_3[40937] = 32'b00000000000000010100001001011101;
assign LUT_3[40938] = 32'b00000000000000001111100101100100;
assign LUT_3[40939] = 32'b00000000000000010110010001000001;
assign LUT_3[40940] = 32'b00000000000000001010101011110110;
assign LUT_3[40941] = 32'b00000000000000010001010111010011;
assign LUT_3[40942] = 32'b00000000000000001100110011011010;
assign LUT_3[40943] = 32'b00000000000000010011011110110111;
assign LUT_3[40944] = 32'b00000000000000001011010111111101;
assign LUT_3[40945] = 32'b00000000000000010010000011011010;
assign LUT_3[40946] = 32'b00000000000000001101011111100001;
assign LUT_3[40947] = 32'b00000000000000010100001010111110;
assign LUT_3[40948] = 32'b00000000000000001000100101110011;
assign LUT_3[40949] = 32'b00000000000000001111010001010000;
assign LUT_3[40950] = 32'b00000000000000001010101101010111;
assign LUT_3[40951] = 32'b00000000000000010001011000110100;
assign LUT_3[40952] = 32'b00000000000000010000110001000011;
assign LUT_3[40953] = 32'b00000000000000010111011100100000;
assign LUT_3[40954] = 32'b00000000000000010010111000100111;
assign LUT_3[40955] = 32'b00000000000000011001100100000100;
assign LUT_3[40956] = 32'b00000000000000001101111110111001;
assign LUT_3[40957] = 32'b00000000000000010100101010010110;
assign LUT_3[40958] = 32'b00000000000000010000000110011101;
assign LUT_3[40959] = 32'b00000000000000010110110001111010;
assign LUT_3[40960] = 32'b11111111111111111110110110111001;
assign LUT_3[40961] = 32'b00000000000000000101100010010110;
assign LUT_3[40962] = 32'b00000000000000000000111110011101;
assign LUT_3[40963] = 32'b00000000000000000111101001111010;
assign LUT_3[40964] = 32'b11111111111111111100000100101111;
assign LUT_3[40965] = 32'b00000000000000000010110000001100;
assign LUT_3[40966] = 32'b11111111111111111110001100010011;
assign LUT_3[40967] = 32'b00000000000000000100110111110000;
assign LUT_3[40968] = 32'b00000000000000000100001111111111;
assign LUT_3[40969] = 32'b00000000000000001010111011011100;
assign LUT_3[40970] = 32'b00000000000000000110010111100011;
assign LUT_3[40971] = 32'b00000000000000001101000011000000;
assign LUT_3[40972] = 32'b00000000000000000001011101110101;
assign LUT_3[40973] = 32'b00000000000000001000001001010010;
assign LUT_3[40974] = 32'b00000000000000000011100101011001;
assign LUT_3[40975] = 32'b00000000000000001010010000110110;
assign LUT_3[40976] = 32'b00000000000000000010001001111100;
assign LUT_3[40977] = 32'b00000000000000001000110101011001;
assign LUT_3[40978] = 32'b00000000000000000100010001100000;
assign LUT_3[40979] = 32'b00000000000000001010111100111101;
assign LUT_3[40980] = 32'b11111111111111111111010111110010;
assign LUT_3[40981] = 32'b00000000000000000110000011001111;
assign LUT_3[40982] = 32'b00000000000000000001011111010110;
assign LUT_3[40983] = 32'b00000000000000001000001010110011;
assign LUT_3[40984] = 32'b00000000000000000111100011000010;
assign LUT_3[40985] = 32'b00000000000000001110001110011111;
assign LUT_3[40986] = 32'b00000000000000001001101010100110;
assign LUT_3[40987] = 32'b00000000000000010000010110000011;
assign LUT_3[40988] = 32'b00000000000000000100110000111000;
assign LUT_3[40989] = 32'b00000000000000001011011100010101;
assign LUT_3[40990] = 32'b00000000000000000110111000011100;
assign LUT_3[40991] = 32'b00000000000000001101100011111001;
assign LUT_3[40992] = 32'b00000000000000000000000101011001;
assign LUT_3[40993] = 32'b00000000000000000110110000110110;
assign LUT_3[40994] = 32'b00000000000000000010001100111101;
assign LUT_3[40995] = 32'b00000000000000001000111000011010;
assign LUT_3[40996] = 32'b11111111111111111101010011001111;
assign LUT_3[40997] = 32'b00000000000000000011111110101100;
assign LUT_3[40998] = 32'b11111111111111111111011010110011;
assign LUT_3[40999] = 32'b00000000000000000110000110010000;
assign LUT_3[41000] = 32'b00000000000000000101011110011111;
assign LUT_3[41001] = 32'b00000000000000001100001001111100;
assign LUT_3[41002] = 32'b00000000000000000111100110000011;
assign LUT_3[41003] = 32'b00000000000000001110010001100000;
assign LUT_3[41004] = 32'b00000000000000000010101100010101;
assign LUT_3[41005] = 32'b00000000000000001001010111110010;
assign LUT_3[41006] = 32'b00000000000000000100110011111001;
assign LUT_3[41007] = 32'b00000000000000001011011111010110;
assign LUT_3[41008] = 32'b00000000000000000011011000011100;
assign LUT_3[41009] = 32'b00000000000000001010000011111001;
assign LUT_3[41010] = 32'b00000000000000000101100000000000;
assign LUT_3[41011] = 32'b00000000000000001100001011011101;
assign LUT_3[41012] = 32'b00000000000000000000100110010010;
assign LUT_3[41013] = 32'b00000000000000000111010001101111;
assign LUT_3[41014] = 32'b00000000000000000010101101110110;
assign LUT_3[41015] = 32'b00000000000000001001011001010011;
assign LUT_3[41016] = 32'b00000000000000001000110001100010;
assign LUT_3[41017] = 32'b00000000000000001111011100111111;
assign LUT_3[41018] = 32'b00000000000000001010111001000110;
assign LUT_3[41019] = 32'b00000000000000010001100100100011;
assign LUT_3[41020] = 32'b00000000000000000101111111011000;
assign LUT_3[41021] = 32'b00000000000000001100101010110101;
assign LUT_3[41022] = 32'b00000000000000001000000110111100;
assign LUT_3[41023] = 32'b00000000000000001110110010011001;
assign LUT_3[41024] = 32'b11111111111111111110101111100100;
assign LUT_3[41025] = 32'b00000000000000000101011011000001;
assign LUT_3[41026] = 32'b00000000000000000000110111001000;
assign LUT_3[41027] = 32'b00000000000000000111100010100101;
assign LUT_3[41028] = 32'b11111111111111111011111101011010;
assign LUT_3[41029] = 32'b00000000000000000010101000110111;
assign LUT_3[41030] = 32'b11111111111111111110000100111110;
assign LUT_3[41031] = 32'b00000000000000000100110000011011;
assign LUT_3[41032] = 32'b00000000000000000100001000101010;
assign LUT_3[41033] = 32'b00000000000000001010110100000111;
assign LUT_3[41034] = 32'b00000000000000000110010000001110;
assign LUT_3[41035] = 32'b00000000000000001100111011101011;
assign LUT_3[41036] = 32'b00000000000000000001010110100000;
assign LUT_3[41037] = 32'b00000000000000001000000001111101;
assign LUT_3[41038] = 32'b00000000000000000011011110000100;
assign LUT_3[41039] = 32'b00000000000000001010001001100001;
assign LUT_3[41040] = 32'b00000000000000000010000010100111;
assign LUT_3[41041] = 32'b00000000000000001000101110000100;
assign LUT_3[41042] = 32'b00000000000000000100001010001011;
assign LUT_3[41043] = 32'b00000000000000001010110101101000;
assign LUT_3[41044] = 32'b11111111111111111111010000011101;
assign LUT_3[41045] = 32'b00000000000000000101111011111010;
assign LUT_3[41046] = 32'b00000000000000000001011000000001;
assign LUT_3[41047] = 32'b00000000000000001000000011011110;
assign LUT_3[41048] = 32'b00000000000000000111011011101101;
assign LUT_3[41049] = 32'b00000000000000001110000111001010;
assign LUT_3[41050] = 32'b00000000000000001001100011010001;
assign LUT_3[41051] = 32'b00000000000000010000001110101110;
assign LUT_3[41052] = 32'b00000000000000000100101001100011;
assign LUT_3[41053] = 32'b00000000000000001011010101000000;
assign LUT_3[41054] = 32'b00000000000000000110110001000111;
assign LUT_3[41055] = 32'b00000000000000001101011100100100;
assign LUT_3[41056] = 32'b11111111111111111111111110000100;
assign LUT_3[41057] = 32'b00000000000000000110101001100001;
assign LUT_3[41058] = 32'b00000000000000000010000101101000;
assign LUT_3[41059] = 32'b00000000000000001000110001000101;
assign LUT_3[41060] = 32'b11111111111111111101001011111010;
assign LUT_3[41061] = 32'b00000000000000000011110111010111;
assign LUT_3[41062] = 32'b11111111111111111111010011011110;
assign LUT_3[41063] = 32'b00000000000000000101111110111011;
assign LUT_3[41064] = 32'b00000000000000000101010111001010;
assign LUT_3[41065] = 32'b00000000000000001100000010100111;
assign LUT_3[41066] = 32'b00000000000000000111011110101110;
assign LUT_3[41067] = 32'b00000000000000001110001010001011;
assign LUT_3[41068] = 32'b00000000000000000010100101000000;
assign LUT_3[41069] = 32'b00000000000000001001010000011101;
assign LUT_3[41070] = 32'b00000000000000000100101100100100;
assign LUT_3[41071] = 32'b00000000000000001011011000000001;
assign LUT_3[41072] = 32'b00000000000000000011010001000111;
assign LUT_3[41073] = 32'b00000000000000001001111100100100;
assign LUT_3[41074] = 32'b00000000000000000101011000101011;
assign LUT_3[41075] = 32'b00000000000000001100000100001000;
assign LUT_3[41076] = 32'b00000000000000000000011110111101;
assign LUT_3[41077] = 32'b00000000000000000111001010011010;
assign LUT_3[41078] = 32'b00000000000000000010100110100001;
assign LUT_3[41079] = 32'b00000000000000001001010001111110;
assign LUT_3[41080] = 32'b00000000000000001000101010001101;
assign LUT_3[41081] = 32'b00000000000000001111010101101010;
assign LUT_3[41082] = 32'b00000000000000001010110001110001;
assign LUT_3[41083] = 32'b00000000000000010001011101001110;
assign LUT_3[41084] = 32'b00000000000000000101111000000011;
assign LUT_3[41085] = 32'b00000000000000001100100011100000;
assign LUT_3[41086] = 32'b00000000000000000111111111100111;
assign LUT_3[41087] = 32'b00000000000000001110101011000100;
assign LUT_3[41088] = 32'b00000000000000000001000001110111;
assign LUT_3[41089] = 32'b00000000000000000111101101010100;
assign LUT_3[41090] = 32'b00000000000000000011001001011011;
assign LUT_3[41091] = 32'b00000000000000001001110100111000;
assign LUT_3[41092] = 32'b11111111111111111110001111101101;
assign LUT_3[41093] = 32'b00000000000000000100111011001010;
assign LUT_3[41094] = 32'b00000000000000000000010111010001;
assign LUT_3[41095] = 32'b00000000000000000111000010101110;
assign LUT_3[41096] = 32'b00000000000000000110011010111101;
assign LUT_3[41097] = 32'b00000000000000001101000110011010;
assign LUT_3[41098] = 32'b00000000000000001000100010100001;
assign LUT_3[41099] = 32'b00000000000000001111001101111110;
assign LUT_3[41100] = 32'b00000000000000000011101000110011;
assign LUT_3[41101] = 32'b00000000000000001010010100010000;
assign LUT_3[41102] = 32'b00000000000000000101110000010111;
assign LUT_3[41103] = 32'b00000000000000001100011011110100;
assign LUT_3[41104] = 32'b00000000000000000100010100111010;
assign LUT_3[41105] = 32'b00000000000000001011000000010111;
assign LUT_3[41106] = 32'b00000000000000000110011100011110;
assign LUT_3[41107] = 32'b00000000000000001101000111111011;
assign LUT_3[41108] = 32'b00000000000000000001100010110000;
assign LUT_3[41109] = 32'b00000000000000001000001110001101;
assign LUT_3[41110] = 32'b00000000000000000011101010010100;
assign LUT_3[41111] = 32'b00000000000000001010010101110001;
assign LUT_3[41112] = 32'b00000000000000001001101110000000;
assign LUT_3[41113] = 32'b00000000000000010000011001011101;
assign LUT_3[41114] = 32'b00000000000000001011110101100100;
assign LUT_3[41115] = 32'b00000000000000010010100001000001;
assign LUT_3[41116] = 32'b00000000000000000110111011110110;
assign LUT_3[41117] = 32'b00000000000000001101100111010011;
assign LUT_3[41118] = 32'b00000000000000001001000011011010;
assign LUT_3[41119] = 32'b00000000000000001111101110110111;
assign LUT_3[41120] = 32'b00000000000000000010010000010111;
assign LUT_3[41121] = 32'b00000000000000001000111011110100;
assign LUT_3[41122] = 32'b00000000000000000100010111111011;
assign LUT_3[41123] = 32'b00000000000000001011000011011000;
assign LUT_3[41124] = 32'b11111111111111111111011110001101;
assign LUT_3[41125] = 32'b00000000000000000110001001101010;
assign LUT_3[41126] = 32'b00000000000000000001100101110001;
assign LUT_3[41127] = 32'b00000000000000001000010001001110;
assign LUT_3[41128] = 32'b00000000000000000111101001011101;
assign LUT_3[41129] = 32'b00000000000000001110010100111010;
assign LUT_3[41130] = 32'b00000000000000001001110001000001;
assign LUT_3[41131] = 32'b00000000000000010000011100011110;
assign LUT_3[41132] = 32'b00000000000000000100110111010011;
assign LUT_3[41133] = 32'b00000000000000001011100010110000;
assign LUT_3[41134] = 32'b00000000000000000110111110110111;
assign LUT_3[41135] = 32'b00000000000000001101101010010100;
assign LUT_3[41136] = 32'b00000000000000000101100011011010;
assign LUT_3[41137] = 32'b00000000000000001100001110110111;
assign LUT_3[41138] = 32'b00000000000000000111101010111110;
assign LUT_3[41139] = 32'b00000000000000001110010110011011;
assign LUT_3[41140] = 32'b00000000000000000010110001010000;
assign LUT_3[41141] = 32'b00000000000000001001011100101101;
assign LUT_3[41142] = 32'b00000000000000000100111000110100;
assign LUT_3[41143] = 32'b00000000000000001011100100010001;
assign LUT_3[41144] = 32'b00000000000000001010111100100000;
assign LUT_3[41145] = 32'b00000000000000010001100111111101;
assign LUT_3[41146] = 32'b00000000000000001101000100000100;
assign LUT_3[41147] = 32'b00000000000000010011101111100001;
assign LUT_3[41148] = 32'b00000000000000001000001010010110;
assign LUT_3[41149] = 32'b00000000000000001110110101110011;
assign LUT_3[41150] = 32'b00000000000000001010010001111010;
assign LUT_3[41151] = 32'b00000000000000010000111101010111;
assign LUT_3[41152] = 32'b00000000000000000000111010100010;
assign LUT_3[41153] = 32'b00000000000000000111100101111111;
assign LUT_3[41154] = 32'b00000000000000000011000010000110;
assign LUT_3[41155] = 32'b00000000000000001001101101100011;
assign LUT_3[41156] = 32'b11111111111111111110001000011000;
assign LUT_3[41157] = 32'b00000000000000000100110011110101;
assign LUT_3[41158] = 32'b00000000000000000000001111111100;
assign LUT_3[41159] = 32'b00000000000000000110111011011001;
assign LUT_3[41160] = 32'b00000000000000000110010011101000;
assign LUT_3[41161] = 32'b00000000000000001100111111000101;
assign LUT_3[41162] = 32'b00000000000000001000011011001100;
assign LUT_3[41163] = 32'b00000000000000001111000110101001;
assign LUT_3[41164] = 32'b00000000000000000011100001011110;
assign LUT_3[41165] = 32'b00000000000000001010001100111011;
assign LUT_3[41166] = 32'b00000000000000000101101001000010;
assign LUT_3[41167] = 32'b00000000000000001100010100011111;
assign LUT_3[41168] = 32'b00000000000000000100001101100101;
assign LUT_3[41169] = 32'b00000000000000001010111001000010;
assign LUT_3[41170] = 32'b00000000000000000110010101001001;
assign LUT_3[41171] = 32'b00000000000000001101000000100110;
assign LUT_3[41172] = 32'b00000000000000000001011011011011;
assign LUT_3[41173] = 32'b00000000000000001000000110111000;
assign LUT_3[41174] = 32'b00000000000000000011100010111111;
assign LUT_3[41175] = 32'b00000000000000001010001110011100;
assign LUT_3[41176] = 32'b00000000000000001001100110101011;
assign LUT_3[41177] = 32'b00000000000000010000010010001000;
assign LUT_3[41178] = 32'b00000000000000001011101110001111;
assign LUT_3[41179] = 32'b00000000000000010010011001101100;
assign LUT_3[41180] = 32'b00000000000000000110110100100001;
assign LUT_3[41181] = 32'b00000000000000001101011111111110;
assign LUT_3[41182] = 32'b00000000000000001000111100000101;
assign LUT_3[41183] = 32'b00000000000000001111100111100010;
assign LUT_3[41184] = 32'b00000000000000000010001001000010;
assign LUT_3[41185] = 32'b00000000000000001000110100011111;
assign LUT_3[41186] = 32'b00000000000000000100010000100110;
assign LUT_3[41187] = 32'b00000000000000001010111100000011;
assign LUT_3[41188] = 32'b11111111111111111111010110111000;
assign LUT_3[41189] = 32'b00000000000000000110000010010101;
assign LUT_3[41190] = 32'b00000000000000000001011110011100;
assign LUT_3[41191] = 32'b00000000000000001000001001111001;
assign LUT_3[41192] = 32'b00000000000000000111100010001000;
assign LUT_3[41193] = 32'b00000000000000001110001101100101;
assign LUT_3[41194] = 32'b00000000000000001001101001101100;
assign LUT_3[41195] = 32'b00000000000000010000010101001001;
assign LUT_3[41196] = 32'b00000000000000000100101111111110;
assign LUT_3[41197] = 32'b00000000000000001011011011011011;
assign LUT_3[41198] = 32'b00000000000000000110110111100010;
assign LUT_3[41199] = 32'b00000000000000001101100010111111;
assign LUT_3[41200] = 32'b00000000000000000101011100000101;
assign LUT_3[41201] = 32'b00000000000000001100000111100010;
assign LUT_3[41202] = 32'b00000000000000000111100011101001;
assign LUT_3[41203] = 32'b00000000000000001110001111000110;
assign LUT_3[41204] = 32'b00000000000000000010101001111011;
assign LUT_3[41205] = 32'b00000000000000001001010101011000;
assign LUT_3[41206] = 32'b00000000000000000100110001011111;
assign LUT_3[41207] = 32'b00000000000000001011011100111100;
assign LUT_3[41208] = 32'b00000000000000001010110101001011;
assign LUT_3[41209] = 32'b00000000000000010001100000101000;
assign LUT_3[41210] = 32'b00000000000000001100111100101111;
assign LUT_3[41211] = 32'b00000000000000010011101000001100;
assign LUT_3[41212] = 32'b00000000000000001000000011000001;
assign LUT_3[41213] = 32'b00000000000000001110101110011110;
assign LUT_3[41214] = 32'b00000000000000001010001010100101;
assign LUT_3[41215] = 32'b00000000000000010000110110000010;
assign LUT_3[41216] = 32'b11111111111111111011000110011010;
assign LUT_3[41217] = 32'b00000000000000000001110001110111;
assign LUT_3[41218] = 32'b11111111111111111101001101111110;
assign LUT_3[41219] = 32'b00000000000000000011111001011011;
assign LUT_3[41220] = 32'b11111111111111111000010100010000;
assign LUT_3[41221] = 32'b11111111111111111110111111101101;
assign LUT_3[41222] = 32'b11111111111111111010011011110100;
assign LUT_3[41223] = 32'b00000000000000000001000111010001;
assign LUT_3[41224] = 32'b00000000000000000000011111100000;
assign LUT_3[41225] = 32'b00000000000000000111001010111101;
assign LUT_3[41226] = 32'b00000000000000000010100111000100;
assign LUT_3[41227] = 32'b00000000000000001001010010100001;
assign LUT_3[41228] = 32'b11111111111111111101101101010110;
assign LUT_3[41229] = 32'b00000000000000000100011000110011;
assign LUT_3[41230] = 32'b11111111111111111111110100111010;
assign LUT_3[41231] = 32'b00000000000000000110100000010111;
assign LUT_3[41232] = 32'b11111111111111111110011001011101;
assign LUT_3[41233] = 32'b00000000000000000101000100111010;
assign LUT_3[41234] = 32'b00000000000000000000100001000001;
assign LUT_3[41235] = 32'b00000000000000000111001100011110;
assign LUT_3[41236] = 32'b11111111111111111011100111010011;
assign LUT_3[41237] = 32'b00000000000000000010010010110000;
assign LUT_3[41238] = 32'b11111111111111111101101110110111;
assign LUT_3[41239] = 32'b00000000000000000100011010010100;
assign LUT_3[41240] = 32'b00000000000000000011110010100011;
assign LUT_3[41241] = 32'b00000000000000001010011110000000;
assign LUT_3[41242] = 32'b00000000000000000101111010000111;
assign LUT_3[41243] = 32'b00000000000000001100100101100100;
assign LUT_3[41244] = 32'b00000000000000000001000000011001;
assign LUT_3[41245] = 32'b00000000000000000111101011110110;
assign LUT_3[41246] = 32'b00000000000000000011000111111101;
assign LUT_3[41247] = 32'b00000000000000001001110011011010;
assign LUT_3[41248] = 32'b11111111111111111100010100111010;
assign LUT_3[41249] = 32'b00000000000000000011000000010111;
assign LUT_3[41250] = 32'b11111111111111111110011100011110;
assign LUT_3[41251] = 32'b00000000000000000101000111111011;
assign LUT_3[41252] = 32'b11111111111111111001100010110000;
assign LUT_3[41253] = 32'b00000000000000000000001110001101;
assign LUT_3[41254] = 32'b11111111111111111011101010010100;
assign LUT_3[41255] = 32'b00000000000000000010010101110001;
assign LUT_3[41256] = 32'b00000000000000000001101110000000;
assign LUT_3[41257] = 32'b00000000000000001000011001011101;
assign LUT_3[41258] = 32'b00000000000000000011110101100100;
assign LUT_3[41259] = 32'b00000000000000001010100001000001;
assign LUT_3[41260] = 32'b11111111111111111110111011110110;
assign LUT_3[41261] = 32'b00000000000000000101100111010011;
assign LUT_3[41262] = 32'b00000000000000000001000011011010;
assign LUT_3[41263] = 32'b00000000000000000111101110110111;
assign LUT_3[41264] = 32'b11111111111111111111100111111101;
assign LUT_3[41265] = 32'b00000000000000000110010011011010;
assign LUT_3[41266] = 32'b00000000000000000001101111100001;
assign LUT_3[41267] = 32'b00000000000000001000011010111110;
assign LUT_3[41268] = 32'b11111111111111111100110101110011;
assign LUT_3[41269] = 32'b00000000000000000011100001010000;
assign LUT_3[41270] = 32'b11111111111111111110111101010111;
assign LUT_3[41271] = 32'b00000000000000000101101000110100;
assign LUT_3[41272] = 32'b00000000000000000101000001000011;
assign LUT_3[41273] = 32'b00000000000000001011101100100000;
assign LUT_3[41274] = 32'b00000000000000000111001000100111;
assign LUT_3[41275] = 32'b00000000000000001101110100000100;
assign LUT_3[41276] = 32'b00000000000000000010001110111001;
assign LUT_3[41277] = 32'b00000000000000001000111010010110;
assign LUT_3[41278] = 32'b00000000000000000100010110011101;
assign LUT_3[41279] = 32'b00000000000000001011000001111010;
assign LUT_3[41280] = 32'b11111111111111111010111111000101;
assign LUT_3[41281] = 32'b00000000000000000001101010100010;
assign LUT_3[41282] = 32'b11111111111111111101000110101001;
assign LUT_3[41283] = 32'b00000000000000000011110010000110;
assign LUT_3[41284] = 32'b11111111111111111000001100111011;
assign LUT_3[41285] = 32'b11111111111111111110111000011000;
assign LUT_3[41286] = 32'b11111111111111111010010100011111;
assign LUT_3[41287] = 32'b00000000000000000000111111111100;
assign LUT_3[41288] = 32'b00000000000000000000011000001011;
assign LUT_3[41289] = 32'b00000000000000000111000011101000;
assign LUT_3[41290] = 32'b00000000000000000010011111101111;
assign LUT_3[41291] = 32'b00000000000000001001001011001100;
assign LUT_3[41292] = 32'b11111111111111111101100110000001;
assign LUT_3[41293] = 32'b00000000000000000100010001011110;
assign LUT_3[41294] = 32'b11111111111111111111101101100101;
assign LUT_3[41295] = 32'b00000000000000000110011001000010;
assign LUT_3[41296] = 32'b11111111111111111110010010001000;
assign LUT_3[41297] = 32'b00000000000000000100111101100101;
assign LUT_3[41298] = 32'b00000000000000000000011001101100;
assign LUT_3[41299] = 32'b00000000000000000111000101001001;
assign LUT_3[41300] = 32'b11111111111111111011011111111110;
assign LUT_3[41301] = 32'b00000000000000000010001011011011;
assign LUT_3[41302] = 32'b11111111111111111101100111100010;
assign LUT_3[41303] = 32'b00000000000000000100010010111111;
assign LUT_3[41304] = 32'b00000000000000000011101011001110;
assign LUT_3[41305] = 32'b00000000000000001010010110101011;
assign LUT_3[41306] = 32'b00000000000000000101110010110010;
assign LUT_3[41307] = 32'b00000000000000001100011110001111;
assign LUT_3[41308] = 32'b00000000000000000000111001000100;
assign LUT_3[41309] = 32'b00000000000000000111100100100001;
assign LUT_3[41310] = 32'b00000000000000000011000000101000;
assign LUT_3[41311] = 32'b00000000000000001001101100000101;
assign LUT_3[41312] = 32'b11111111111111111100001101100101;
assign LUT_3[41313] = 32'b00000000000000000010111001000010;
assign LUT_3[41314] = 32'b11111111111111111110010101001001;
assign LUT_3[41315] = 32'b00000000000000000101000000100110;
assign LUT_3[41316] = 32'b11111111111111111001011011011011;
assign LUT_3[41317] = 32'b00000000000000000000000110111000;
assign LUT_3[41318] = 32'b11111111111111111011100010111111;
assign LUT_3[41319] = 32'b00000000000000000010001110011100;
assign LUT_3[41320] = 32'b00000000000000000001100110101011;
assign LUT_3[41321] = 32'b00000000000000001000010010001000;
assign LUT_3[41322] = 32'b00000000000000000011101110001111;
assign LUT_3[41323] = 32'b00000000000000001010011001101100;
assign LUT_3[41324] = 32'b11111111111111111110110100100001;
assign LUT_3[41325] = 32'b00000000000000000101011111111110;
assign LUT_3[41326] = 32'b00000000000000000000111100000101;
assign LUT_3[41327] = 32'b00000000000000000111100111100010;
assign LUT_3[41328] = 32'b11111111111111111111100000101000;
assign LUT_3[41329] = 32'b00000000000000000110001100000101;
assign LUT_3[41330] = 32'b00000000000000000001101000001100;
assign LUT_3[41331] = 32'b00000000000000001000010011101001;
assign LUT_3[41332] = 32'b11111111111111111100101110011110;
assign LUT_3[41333] = 32'b00000000000000000011011001111011;
assign LUT_3[41334] = 32'b11111111111111111110110110000010;
assign LUT_3[41335] = 32'b00000000000000000101100001011111;
assign LUT_3[41336] = 32'b00000000000000000100111001101110;
assign LUT_3[41337] = 32'b00000000000000001011100101001011;
assign LUT_3[41338] = 32'b00000000000000000111000001010010;
assign LUT_3[41339] = 32'b00000000000000001101101100101111;
assign LUT_3[41340] = 32'b00000000000000000010000111100100;
assign LUT_3[41341] = 32'b00000000000000001000110011000001;
assign LUT_3[41342] = 32'b00000000000000000100001111001000;
assign LUT_3[41343] = 32'b00000000000000001010111010100101;
assign LUT_3[41344] = 32'b11111111111111111101010001011000;
assign LUT_3[41345] = 32'b00000000000000000011111100110101;
assign LUT_3[41346] = 32'b11111111111111111111011000111100;
assign LUT_3[41347] = 32'b00000000000000000110000100011001;
assign LUT_3[41348] = 32'b11111111111111111010011111001110;
assign LUT_3[41349] = 32'b00000000000000000001001010101011;
assign LUT_3[41350] = 32'b11111111111111111100100110110010;
assign LUT_3[41351] = 32'b00000000000000000011010010001111;
assign LUT_3[41352] = 32'b00000000000000000010101010011110;
assign LUT_3[41353] = 32'b00000000000000001001010101111011;
assign LUT_3[41354] = 32'b00000000000000000100110010000010;
assign LUT_3[41355] = 32'b00000000000000001011011101011111;
assign LUT_3[41356] = 32'b11111111111111111111111000010100;
assign LUT_3[41357] = 32'b00000000000000000110100011110001;
assign LUT_3[41358] = 32'b00000000000000000001111111111000;
assign LUT_3[41359] = 32'b00000000000000001000101011010101;
assign LUT_3[41360] = 32'b00000000000000000000100100011011;
assign LUT_3[41361] = 32'b00000000000000000111001111111000;
assign LUT_3[41362] = 32'b00000000000000000010101011111111;
assign LUT_3[41363] = 32'b00000000000000001001010111011100;
assign LUT_3[41364] = 32'b11111111111111111101110010010001;
assign LUT_3[41365] = 32'b00000000000000000100011101101110;
assign LUT_3[41366] = 32'b11111111111111111111111001110101;
assign LUT_3[41367] = 32'b00000000000000000110100101010010;
assign LUT_3[41368] = 32'b00000000000000000101111101100001;
assign LUT_3[41369] = 32'b00000000000000001100101000111110;
assign LUT_3[41370] = 32'b00000000000000001000000101000101;
assign LUT_3[41371] = 32'b00000000000000001110110000100010;
assign LUT_3[41372] = 32'b00000000000000000011001011010111;
assign LUT_3[41373] = 32'b00000000000000001001110110110100;
assign LUT_3[41374] = 32'b00000000000000000101010010111011;
assign LUT_3[41375] = 32'b00000000000000001011111110011000;
assign LUT_3[41376] = 32'b11111111111111111110011111111000;
assign LUT_3[41377] = 32'b00000000000000000101001011010101;
assign LUT_3[41378] = 32'b00000000000000000000100111011100;
assign LUT_3[41379] = 32'b00000000000000000111010010111001;
assign LUT_3[41380] = 32'b11111111111111111011101101101110;
assign LUT_3[41381] = 32'b00000000000000000010011001001011;
assign LUT_3[41382] = 32'b11111111111111111101110101010010;
assign LUT_3[41383] = 32'b00000000000000000100100000101111;
assign LUT_3[41384] = 32'b00000000000000000011111000111110;
assign LUT_3[41385] = 32'b00000000000000001010100100011011;
assign LUT_3[41386] = 32'b00000000000000000110000000100010;
assign LUT_3[41387] = 32'b00000000000000001100101011111111;
assign LUT_3[41388] = 32'b00000000000000000001000110110100;
assign LUT_3[41389] = 32'b00000000000000000111110010010001;
assign LUT_3[41390] = 32'b00000000000000000011001110011000;
assign LUT_3[41391] = 32'b00000000000000001001111001110101;
assign LUT_3[41392] = 32'b00000000000000000001110010111011;
assign LUT_3[41393] = 32'b00000000000000001000011110011000;
assign LUT_3[41394] = 32'b00000000000000000011111010011111;
assign LUT_3[41395] = 32'b00000000000000001010100101111100;
assign LUT_3[41396] = 32'b11111111111111111111000000110001;
assign LUT_3[41397] = 32'b00000000000000000101101100001110;
assign LUT_3[41398] = 32'b00000000000000000001001000010101;
assign LUT_3[41399] = 32'b00000000000000000111110011110010;
assign LUT_3[41400] = 32'b00000000000000000111001100000001;
assign LUT_3[41401] = 32'b00000000000000001101110111011110;
assign LUT_3[41402] = 32'b00000000000000001001010011100101;
assign LUT_3[41403] = 32'b00000000000000001111111111000010;
assign LUT_3[41404] = 32'b00000000000000000100011001110111;
assign LUT_3[41405] = 32'b00000000000000001011000101010100;
assign LUT_3[41406] = 32'b00000000000000000110100001011011;
assign LUT_3[41407] = 32'b00000000000000001101001100111000;
assign LUT_3[41408] = 32'b11111111111111111101001010000011;
assign LUT_3[41409] = 32'b00000000000000000011110101100000;
assign LUT_3[41410] = 32'b11111111111111111111010001100111;
assign LUT_3[41411] = 32'b00000000000000000101111101000100;
assign LUT_3[41412] = 32'b11111111111111111010010111111001;
assign LUT_3[41413] = 32'b00000000000000000001000011010110;
assign LUT_3[41414] = 32'b11111111111111111100011111011101;
assign LUT_3[41415] = 32'b00000000000000000011001010111010;
assign LUT_3[41416] = 32'b00000000000000000010100011001001;
assign LUT_3[41417] = 32'b00000000000000001001001110100110;
assign LUT_3[41418] = 32'b00000000000000000100101010101101;
assign LUT_3[41419] = 32'b00000000000000001011010110001010;
assign LUT_3[41420] = 32'b11111111111111111111110000111111;
assign LUT_3[41421] = 32'b00000000000000000110011100011100;
assign LUT_3[41422] = 32'b00000000000000000001111000100011;
assign LUT_3[41423] = 32'b00000000000000001000100100000000;
assign LUT_3[41424] = 32'b00000000000000000000011101000110;
assign LUT_3[41425] = 32'b00000000000000000111001000100011;
assign LUT_3[41426] = 32'b00000000000000000010100100101010;
assign LUT_3[41427] = 32'b00000000000000001001010000000111;
assign LUT_3[41428] = 32'b11111111111111111101101010111100;
assign LUT_3[41429] = 32'b00000000000000000100010110011001;
assign LUT_3[41430] = 32'b11111111111111111111110010100000;
assign LUT_3[41431] = 32'b00000000000000000110011101111101;
assign LUT_3[41432] = 32'b00000000000000000101110110001100;
assign LUT_3[41433] = 32'b00000000000000001100100001101001;
assign LUT_3[41434] = 32'b00000000000000000111111101110000;
assign LUT_3[41435] = 32'b00000000000000001110101001001101;
assign LUT_3[41436] = 32'b00000000000000000011000100000010;
assign LUT_3[41437] = 32'b00000000000000001001101111011111;
assign LUT_3[41438] = 32'b00000000000000000101001011100110;
assign LUT_3[41439] = 32'b00000000000000001011110111000011;
assign LUT_3[41440] = 32'b11111111111111111110011000100011;
assign LUT_3[41441] = 32'b00000000000000000101000100000000;
assign LUT_3[41442] = 32'b00000000000000000000100000000111;
assign LUT_3[41443] = 32'b00000000000000000111001011100100;
assign LUT_3[41444] = 32'b11111111111111111011100110011001;
assign LUT_3[41445] = 32'b00000000000000000010010001110110;
assign LUT_3[41446] = 32'b11111111111111111101101101111101;
assign LUT_3[41447] = 32'b00000000000000000100011001011010;
assign LUT_3[41448] = 32'b00000000000000000011110001101001;
assign LUT_3[41449] = 32'b00000000000000001010011101000110;
assign LUT_3[41450] = 32'b00000000000000000101111001001101;
assign LUT_3[41451] = 32'b00000000000000001100100100101010;
assign LUT_3[41452] = 32'b00000000000000000000111111011111;
assign LUT_3[41453] = 32'b00000000000000000111101010111100;
assign LUT_3[41454] = 32'b00000000000000000011000111000011;
assign LUT_3[41455] = 32'b00000000000000001001110010100000;
assign LUT_3[41456] = 32'b00000000000000000001101011100110;
assign LUT_3[41457] = 32'b00000000000000001000010111000011;
assign LUT_3[41458] = 32'b00000000000000000011110011001010;
assign LUT_3[41459] = 32'b00000000000000001010011110100111;
assign LUT_3[41460] = 32'b11111111111111111110111001011100;
assign LUT_3[41461] = 32'b00000000000000000101100100111001;
assign LUT_3[41462] = 32'b00000000000000000001000001000000;
assign LUT_3[41463] = 32'b00000000000000000111101100011101;
assign LUT_3[41464] = 32'b00000000000000000111000100101100;
assign LUT_3[41465] = 32'b00000000000000001101110000001001;
assign LUT_3[41466] = 32'b00000000000000001001001100010000;
assign LUT_3[41467] = 32'b00000000000000001111110111101101;
assign LUT_3[41468] = 32'b00000000000000000100010010100010;
assign LUT_3[41469] = 32'b00000000000000001010111101111111;
assign LUT_3[41470] = 32'b00000000000000000110011010000110;
assign LUT_3[41471] = 32'b00000000000000001101000101100011;
assign LUT_3[41472] = 32'b00000000000000000010001100000101;
assign LUT_3[41473] = 32'b00000000000000001000110111100010;
assign LUT_3[41474] = 32'b00000000000000000100010011101001;
assign LUT_3[41475] = 32'b00000000000000001010111111000110;
assign LUT_3[41476] = 32'b11111111111111111111011001111011;
assign LUT_3[41477] = 32'b00000000000000000110000101011000;
assign LUT_3[41478] = 32'b00000000000000000001100001011111;
assign LUT_3[41479] = 32'b00000000000000001000001100111100;
assign LUT_3[41480] = 32'b00000000000000000111100101001011;
assign LUT_3[41481] = 32'b00000000000000001110010000101000;
assign LUT_3[41482] = 32'b00000000000000001001101100101111;
assign LUT_3[41483] = 32'b00000000000000010000011000001100;
assign LUT_3[41484] = 32'b00000000000000000100110011000001;
assign LUT_3[41485] = 32'b00000000000000001011011110011110;
assign LUT_3[41486] = 32'b00000000000000000110111010100101;
assign LUT_3[41487] = 32'b00000000000000001101100110000010;
assign LUT_3[41488] = 32'b00000000000000000101011111001000;
assign LUT_3[41489] = 32'b00000000000000001100001010100101;
assign LUT_3[41490] = 32'b00000000000000000111100110101100;
assign LUT_3[41491] = 32'b00000000000000001110010010001001;
assign LUT_3[41492] = 32'b00000000000000000010101100111110;
assign LUT_3[41493] = 32'b00000000000000001001011000011011;
assign LUT_3[41494] = 32'b00000000000000000100110100100010;
assign LUT_3[41495] = 32'b00000000000000001011011111111111;
assign LUT_3[41496] = 32'b00000000000000001010111000001110;
assign LUT_3[41497] = 32'b00000000000000010001100011101011;
assign LUT_3[41498] = 32'b00000000000000001100111111110010;
assign LUT_3[41499] = 32'b00000000000000010011101011001111;
assign LUT_3[41500] = 32'b00000000000000001000000110000100;
assign LUT_3[41501] = 32'b00000000000000001110110001100001;
assign LUT_3[41502] = 32'b00000000000000001010001101101000;
assign LUT_3[41503] = 32'b00000000000000010000111001000101;
assign LUT_3[41504] = 32'b00000000000000000011011010100101;
assign LUT_3[41505] = 32'b00000000000000001010000110000010;
assign LUT_3[41506] = 32'b00000000000000000101100010001001;
assign LUT_3[41507] = 32'b00000000000000001100001101100110;
assign LUT_3[41508] = 32'b00000000000000000000101000011011;
assign LUT_3[41509] = 32'b00000000000000000111010011111000;
assign LUT_3[41510] = 32'b00000000000000000010101111111111;
assign LUT_3[41511] = 32'b00000000000000001001011011011100;
assign LUT_3[41512] = 32'b00000000000000001000110011101011;
assign LUT_3[41513] = 32'b00000000000000001111011111001000;
assign LUT_3[41514] = 32'b00000000000000001010111011001111;
assign LUT_3[41515] = 32'b00000000000000010001100110101100;
assign LUT_3[41516] = 32'b00000000000000000110000001100001;
assign LUT_3[41517] = 32'b00000000000000001100101100111110;
assign LUT_3[41518] = 32'b00000000000000001000001001000101;
assign LUT_3[41519] = 32'b00000000000000001110110100100010;
assign LUT_3[41520] = 32'b00000000000000000110101101101000;
assign LUT_3[41521] = 32'b00000000000000001101011001000101;
assign LUT_3[41522] = 32'b00000000000000001000110101001100;
assign LUT_3[41523] = 32'b00000000000000001111100000101001;
assign LUT_3[41524] = 32'b00000000000000000011111011011110;
assign LUT_3[41525] = 32'b00000000000000001010100110111011;
assign LUT_3[41526] = 32'b00000000000000000110000011000010;
assign LUT_3[41527] = 32'b00000000000000001100101110011111;
assign LUT_3[41528] = 32'b00000000000000001100000110101110;
assign LUT_3[41529] = 32'b00000000000000010010110010001011;
assign LUT_3[41530] = 32'b00000000000000001110001110010010;
assign LUT_3[41531] = 32'b00000000000000010100111001101111;
assign LUT_3[41532] = 32'b00000000000000001001010100100100;
assign LUT_3[41533] = 32'b00000000000000010000000000000001;
assign LUT_3[41534] = 32'b00000000000000001011011100001000;
assign LUT_3[41535] = 32'b00000000000000010010000111100101;
assign LUT_3[41536] = 32'b00000000000000000010000100110000;
assign LUT_3[41537] = 32'b00000000000000001000110000001101;
assign LUT_3[41538] = 32'b00000000000000000100001100010100;
assign LUT_3[41539] = 32'b00000000000000001010110111110001;
assign LUT_3[41540] = 32'b11111111111111111111010010100110;
assign LUT_3[41541] = 32'b00000000000000000101111110000011;
assign LUT_3[41542] = 32'b00000000000000000001011010001010;
assign LUT_3[41543] = 32'b00000000000000001000000101100111;
assign LUT_3[41544] = 32'b00000000000000000111011101110110;
assign LUT_3[41545] = 32'b00000000000000001110001001010011;
assign LUT_3[41546] = 32'b00000000000000001001100101011010;
assign LUT_3[41547] = 32'b00000000000000010000010000110111;
assign LUT_3[41548] = 32'b00000000000000000100101011101100;
assign LUT_3[41549] = 32'b00000000000000001011010111001001;
assign LUT_3[41550] = 32'b00000000000000000110110011010000;
assign LUT_3[41551] = 32'b00000000000000001101011110101101;
assign LUT_3[41552] = 32'b00000000000000000101010111110011;
assign LUT_3[41553] = 32'b00000000000000001100000011010000;
assign LUT_3[41554] = 32'b00000000000000000111011111010111;
assign LUT_3[41555] = 32'b00000000000000001110001010110100;
assign LUT_3[41556] = 32'b00000000000000000010100101101001;
assign LUT_3[41557] = 32'b00000000000000001001010001000110;
assign LUT_3[41558] = 32'b00000000000000000100101101001101;
assign LUT_3[41559] = 32'b00000000000000001011011000101010;
assign LUT_3[41560] = 32'b00000000000000001010110000111001;
assign LUT_3[41561] = 32'b00000000000000010001011100010110;
assign LUT_3[41562] = 32'b00000000000000001100111000011101;
assign LUT_3[41563] = 32'b00000000000000010011100011111010;
assign LUT_3[41564] = 32'b00000000000000000111111110101111;
assign LUT_3[41565] = 32'b00000000000000001110101010001100;
assign LUT_3[41566] = 32'b00000000000000001010000110010011;
assign LUT_3[41567] = 32'b00000000000000010000110001110000;
assign LUT_3[41568] = 32'b00000000000000000011010011010000;
assign LUT_3[41569] = 32'b00000000000000001001111110101101;
assign LUT_3[41570] = 32'b00000000000000000101011010110100;
assign LUT_3[41571] = 32'b00000000000000001100000110010001;
assign LUT_3[41572] = 32'b00000000000000000000100001000110;
assign LUT_3[41573] = 32'b00000000000000000111001100100011;
assign LUT_3[41574] = 32'b00000000000000000010101000101010;
assign LUT_3[41575] = 32'b00000000000000001001010100000111;
assign LUT_3[41576] = 32'b00000000000000001000101100010110;
assign LUT_3[41577] = 32'b00000000000000001111010111110011;
assign LUT_3[41578] = 32'b00000000000000001010110011111010;
assign LUT_3[41579] = 32'b00000000000000010001011111010111;
assign LUT_3[41580] = 32'b00000000000000000101111010001100;
assign LUT_3[41581] = 32'b00000000000000001100100101101001;
assign LUT_3[41582] = 32'b00000000000000001000000001110000;
assign LUT_3[41583] = 32'b00000000000000001110101101001101;
assign LUT_3[41584] = 32'b00000000000000000110100110010011;
assign LUT_3[41585] = 32'b00000000000000001101010001110000;
assign LUT_3[41586] = 32'b00000000000000001000101101110111;
assign LUT_3[41587] = 32'b00000000000000001111011001010100;
assign LUT_3[41588] = 32'b00000000000000000011110100001001;
assign LUT_3[41589] = 32'b00000000000000001010011111100110;
assign LUT_3[41590] = 32'b00000000000000000101111011101101;
assign LUT_3[41591] = 32'b00000000000000001100100111001010;
assign LUT_3[41592] = 32'b00000000000000001011111111011001;
assign LUT_3[41593] = 32'b00000000000000010010101010110110;
assign LUT_3[41594] = 32'b00000000000000001110000110111101;
assign LUT_3[41595] = 32'b00000000000000010100110010011010;
assign LUT_3[41596] = 32'b00000000000000001001001101001111;
assign LUT_3[41597] = 32'b00000000000000001111111000101100;
assign LUT_3[41598] = 32'b00000000000000001011010100110011;
assign LUT_3[41599] = 32'b00000000000000010010000000010000;
assign LUT_3[41600] = 32'b00000000000000000100010111000011;
assign LUT_3[41601] = 32'b00000000000000001011000010100000;
assign LUT_3[41602] = 32'b00000000000000000110011110100111;
assign LUT_3[41603] = 32'b00000000000000001101001010000100;
assign LUT_3[41604] = 32'b00000000000000000001100100111001;
assign LUT_3[41605] = 32'b00000000000000001000010000010110;
assign LUT_3[41606] = 32'b00000000000000000011101100011101;
assign LUT_3[41607] = 32'b00000000000000001010010111111010;
assign LUT_3[41608] = 32'b00000000000000001001110000001001;
assign LUT_3[41609] = 32'b00000000000000010000011011100110;
assign LUT_3[41610] = 32'b00000000000000001011110111101101;
assign LUT_3[41611] = 32'b00000000000000010010100011001010;
assign LUT_3[41612] = 32'b00000000000000000110111101111111;
assign LUT_3[41613] = 32'b00000000000000001101101001011100;
assign LUT_3[41614] = 32'b00000000000000001001000101100011;
assign LUT_3[41615] = 32'b00000000000000001111110001000000;
assign LUT_3[41616] = 32'b00000000000000000111101010000110;
assign LUT_3[41617] = 32'b00000000000000001110010101100011;
assign LUT_3[41618] = 32'b00000000000000001001110001101010;
assign LUT_3[41619] = 32'b00000000000000010000011101000111;
assign LUT_3[41620] = 32'b00000000000000000100110111111100;
assign LUT_3[41621] = 32'b00000000000000001011100011011001;
assign LUT_3[41622] = 32'b00000000000000000110111111100000;
assign LUT_3[41623] = 32'b00000000000000001101101010111101;
assign LUT_3[41624] = 32'b00000000000000001101000011001100;
assign LUT_3[41625] = 32'b00000000000000010011101110101001;
assign LUT_3[41626] = 32'b00000000000000001111001010110000;
assign LUT_3[41627] = 32'b00000000000000010101110110001101;
assign LUT_3[41628] = 32'b00000000000000001010010001000010;
assign LUT_3[41629] = 32'b00000000000000010000111100011111;
assign LUT_3[41630] = 32'b00000000000000001100011000100110;
assign LUT_3[41631] = 32'b00000000000000010011000100000011;
assign LUT_3[41632] = 32'b00000000000000000101100101100011;
assign LUT_3[41633] = 32'b00000000000000001100010001000000;
assign LUT_3[41634] = 32'b00000000000000000111101101000111;
assign LUT_3[41635] = 32'b00000000000000001110011000100100;
assign LUT_3[41636] = 32'b00000000000000000010110011011001;
assign LUT_3[41637] = 32'b00000000000000001001011110110110;
assign LUT_3[41638] = 32'b00000000000000000100111010111101;
assign LUT_3[41639] = 32'b00000000000000001011100110011010;
assign LUT_3[41640] = 32'b00000000000000001010111110101001;
assign LUT_3[41641] = 32'b00000000000000010001101010000110;
assign LUT_3[41642] = 32'b00000000000000001101000110001101;
assign LUT_3[41643] = 32'b00000000000000010011110001101010;
assign LUT_3[41644] = 32'b00000000000000001000001100011111;
assign LUT_3[41645] = 32'b00000000000000001110110111111100;
assign LUT_3[41646] = 32'b00000000000000001010010100000011;
assign LUT_3[41647] = 32'b00000000000000010000111111100000;
assign LUT_3[41648] = 32'b00000000000000001000111000100110;
assign LUT_3[41649] = 32'b00000000000000001111100100000011;
assign LUT_3[41650] = 32'b00000000000000001011000000001010;
assign LUT_3[41651] = 32'b00000000000000010001101011100111;
assign LUT_3[41652] = 32'b00000000000000000110000110011100;
assign LUT_3[41653] = 32'b00000000000000001100110001111001;
assign LUT_3[41654] = 32'b00000000000000001000001110000000;
assign LUT_3[41655] = 32'b00000000000000001110111001011101;
assign LUT_3[41656] = 32'b00000000000000001110010001101100;
assign LUT_3[41657] = 32'b00000000000000010100111101001001;
assign LUT_3[41658] = 32'b00000000000000010000011001010000;
assign LUT_3[41659] = 32'b00000000000000010111000100101101;
assign LUT_3[41660] = 32'b00000000000000001011011111100010;
assign LUT_3[41661] = 32'b00000000000000010010001010111111;
assign LUT_3[41662] = 32'b00000000000000001101100111000110;
assign LUT_3[41663] = 32'b00000000000000010100010010100011;
assign LUT_3[41664] = 32'b00000000000000000100001111101110;
assign LUT_3[41665] = 32'b00000000000000001010111011001011;
assign LUT_3[41666] = 32'b00000000000000000110010111010010;
assign LUT_3[41667] = 32'b00000000000000001101000010101111;
assign LUT_3[41668] = 32'b00000000000000000001011101100100;
assign LUT_3[41669] = 32'b00000000000000001000001001000001;
assign LUT_3[41670] = 32'b00000000000000000011100101001000;
assign LUT_3[41671] = 32'b00000000000000001010010000100101;
assign LUT_3[41672] = 32'b00000000000000001001101000110100;
assign LUT_3[41673] = 32'b00000000000000010000010100010001;
assign LUT_3[41674] = 32'b00000000000000001011110000011000;
assign LUT_3[41675] = 32'b00000000000000010010011011110101;
assign LUT_3[41676] = 32'b00000000000000000110110110101010;
assign LUT_3[41677] = 32'b00000000000000001101100010000111;
assign LUT_3[41678] = 32'b00000000000000001000111110001110;
assign LUT_3[41679] = 32'b00000000000000001111101001101011;
assign LUT_3[41680] = 32'b00000000000000000111100010110001;
assign LUT_3[41681] = 32'b00000000000000001110001110001110;
assign LUT_3[41682] = 32'b00000000000000001001101010010101;
assign LUT_3[41683] = 32'b00000000000000010000010101110010;
assign LUT_3[41684] = 32'b00000000000000000100110000100111;
assign LUT_3[41685] = 32'b00000000000000001011011100000100;
assign LUT_3[41686] = 32'b00000000000000000110111000001011;
assign LUT_3[41687] = 32'b00000000000000001101100011101000;
assign LUT_3[41688] = 32'b00000000000000001100111011110111;
assign LUT_3[41689] = 32'b00000000000000010011100111010100;
assign LUT_3[41690] = 32'b00000000000000001111000011011011;
assign LUT_3[41691] = 32'b00000000000000010101101110111000;
assign LUT_3[41692] = 32'b00000000000000001010001001101101;
assign LUT_3[41693] = 32'b00000000000000010000110101001010;
assign LUT_3[41694] = 32'b00000000000000001100010001010001;
assign LUT_3[41695] = 32'b00000000000000010010111100101110;
assign LUT_3[41696] = 32'b00000000000000000101011110001110;
assign LUT_3[41697] = 32'b00000000000000001100001001101011;
assign LUT_3[41698] = 32'b00000000000000000111100101110010;
assign LUT_3[41699] = 32'b00000000000000001110010001001111;
assign LUT_3[41700] = 32'b00000000000000000010101100000100;
assign LUT_3[41701] = 32'b00000000000000001001010111100001;
assign LUT_3[41702] = 32'b00000000000000000100110011101000;
assign LUT_3[41703] = 32'b00000000000000001011011111000101;
assign LUT_3[41704] = 32'b00000000000000001010110111010100;
assign LUT_3[41705] = 32'b00000000000000010001100010110001;
assign LUT_3[41706] = 32'b00000000000000001100111110111000;
assign LUT_3[41707] = 32'b00000000000000010011101010010101;
assign LUT_3[41708] = 32'b00000000000000001000000101001010;
assign LUT_3[41709] = 32'b00000000000000001110110000100111;
assign LUT_3[41710] = 32'b00000000000000001010001100101110;
assign LUT_3[41711] = 32'b00000000000000010000111000001011;
assign LUT_3[41712] = 32'b00000000000000001000110001010001;
assign LUT_3[41713] = 32'b00000000000000001111011100101110;
assign LUT_3[41714] = 32'b00000000000000001010111000110101;
assign LUT_3[41715] = 32'b00000000000000010001100100010010;
assign LUT_3[41716] = 32'b00000000000000000101111111000111;
assign LUT_3[41717] = 32'b00000000000000001100101010100100;
assign LUT_3[41718] = 32'b00000000000000001000000110101011;
assign LUT_3[41719] = 32'b00000000000000001110110010001000;
assign LUT_3[41720] = 32'b00000000000000001110001010010111;
assign LUT_3[41721] = 32'b00000000000000010100110101110100;
assign LUT_3[41722] = 32'b00000000000000010000010001111011;
assign LUT_3[41723] = 32'b00000000000000010110111101011000;
assign LUT_3[41724] = 32'b00000000000000001011011000001101;
assign LUT_3[41725] = 32'b00000000000000010010000011101010;
assign LUT_3[41726] = 32'b00000000000000001101011111110001;
assign LUT_3[41727] = 32'b00000000000000010100001011001110;
assign LUT_3[41728] = 32'b11111111111111111110011011100110;
assign LUT_3[41729] = 32'b00000000000000000101000111000011;
assign LUT_3[41730] = 32'b00000000000000000000100011001010;
assign LUT_3[41731] = 32'b00000000000000000111001110100111;
assign LUT_3[41732] = 32'b11111111111111111011101001011100;
assign LUT_3[41733] = 32'b00000000000000000010010100111001;
assign LUT_3[41734] = 32'b11111111111111111101110001000000;
assign LUT_3[41735] = 32'b00000000000000000100011100011101;
assign LUT_3[41736] = 32'b00000000000000000011110100101100;
assign LUT_3[41737] = 32'b00000000000000001010100000001001;
assign LUT_3[41738] = 32'b00000000000000000101111100010000;
assign LUT_3[41739] = 32'b00000000000000001100100111101101;
assign LUT_3[41740] = 32'b00000000000000000001000010100010;
assign LUT_3[41741] = 32'b00000000000000000111101101111111;
assign LUT_3[41742] = 32'b00000000000000000011001010000110;
assign LUT_3[41743] = 32'b00000000000000001001110101100011;
assign LUT_3[41744] = 32'b00000000000000000001101110101001;
assign LUT_3[41745] = 32'b00000000000000001000011010000110;
assign LUT_3[41746] = 32'b00000000000000000011110110001101;
assign LUT_3[41747] = 32'b00000000000000001010100001101010;
assign LUT_3[41748] = 32'b11111111111111111110111100011111;
assign LUT_3[41749] = 32'b00000000000000000101100111111100;
assign LUT_3[41750] = 32'b00000000000000000001000100000011;
assign LUT_3[41751] = 32'b00000000000000000111101111100000;
assign LUT_3[41752] = 32'b00000000000000000111000111101111;
assign LUT_3[41753] = 32'b00000000000000001101110011001100;
assign LUT_3[41754] = 32'b00000000000000001001001111010011;
assign LUT_3[41755] = 32'b00000000000000001111111010110000;
assign LUT_3[41756] = 32'b00000000000000000100010101100101;
assign LUT_3[41757] = 32'b00000000000000001011000001000010;
assign LUT_3[41758] = 32'b00000000000000000110011101001001;
assign LUT_3[41759] = 32'b00000000000000001101001000100110;
assign LUT_3[41760] = 32'b11111111111111111111101010000110;
assign LUT_3[41761] = 32'b00000000000000000110010101100011;
assign LUT_3[41762] = 32'b00000000000000000001110001101010;
assign LUT_3[41763] = 32'b00000000000000001000011101000111;
assign LUT_3[41764] = 32'b11111111111111111100110111111100;
assign LUT_3[41765] = 32'b00000000000000000011100011011001;
assign LUT_3[41766] = 32'b11111111111111111110111111100000;
assign LUT_3[41767] = 32'b00000000000000000101101010111101;
assign LUT_3[41768] = 32'b00000000000000000101000011001100;
assign LUT_3[41769] = 32'b00000000000000001011101110101001;
assign LUT_3[41770] = 32'b00000000000000000111001010110000;
assign LUT_3[41771] = 32'b00000000000000001101110110001101;
assign LUT_3[41772] = 32'b00000000000000000010010001000010;
assign LUT_3[41773] = 32'b00000000000000001000111100011111;
assign LUT_3[41774] = 32'b00000000000000000100011000100110;
assign LUT_3[41775] = 32'b00000000000000001011000100000011;
assign LUT_3[41776] = 32'b00000000000000000010111101001001;
assign LUT_3[41777] = 32'b00000000000000001001101000100110;
assign LUT_3[41778] = 32'b00000000000000000101000100101101;
assign LUT_3[41779] = 32'b00000000000000001011110000001010;
assign LUT_3[41780] = 32'b00000000000000000000001010111111;
assign LUT_3[41781] = 32'b00000000000000000110110110011100;
assign LUT_3[41782] = 32'b00000000000000000010010010100011;
assign LUT_3[41783] = 32'b00000000000000001000111110000000;
assign LUT_3[41784] = 32'b00000000000000001000010110001111;
assign LUT_3[41785] = 32'b00000000000000001111000001101100;
assign LUT_3[41786] = 32'b00000000000000001010011101110011;
assign LUT_3[41787] = 32'b00000000000000010001001001010000;
assign LUT_3[41788] = 32'b00000000000000000101100100000101;
assign LUT_3[41789] = 32'b00000000000000001100001111100010;
assign LUT_3[41790] = 32'b00000000000000000111101011101001;
assign LUT_3[41791] = 32'b00000000000000001110010111000110;
assign LUT_3[41792] = 32'b11111111111111111110010100010001;
assign LUT_3[41793] = 32'b00000000000000000100111111101110;
assign LUT_3[41794] = 32'b00000000000000000000011011110101;
assign LUT_3[41795] = 32'b00000000000000000111000111010010;
assign LUT_3[41796] = 32'b11111111111111111011100010000111;
assign LUT_3[41797] = 32'b00000000000000000010001101100100;
assign LUT_3[41798] = 32'b11111111111111111101101001101011;
assign LUT_3[41799] = 32'b00000000000000000100010101001000;
assign LUT_3[41800] = 32'b00000000000000000011101101010111;
assign LUT_3[41801] = 32'b00000000000000001010011000110100;
assign LUT_3[41802] = 32'b00000000000000000101110100111011;
assign LUT_3[41803] = 32'b00000000000000001100100000011000;
assign LUT_3[41804] = 32'b00000000000000000000111011001101;
assign LUT_3[41805] = 32'b00000000000000000111100110101010;
assign LUT_3[41806] = 32'b00000000000000000011000010110001;
assign LUT_3[41807] = 32'b00000000000000001001101110001110;
assign LUT_3[41808] = 32'b00000000000000000001100111010100;
assign LUT_3[41809] = 32'b00000000000000001000010010110001;
assign LUT_3[41810] = 32'b00000000000000000011101110111000;
assign LUT_3[41811] = 32'b00000000000000001010011010010101;
assign LUT_3[41812] = 32'b11111111111111111110110101001010;
assign LUT_3[41813] = 32'b00000000000000000101100000100111;
assign LUT_3[41814] = 32'b00000000000000000000111100101110;
assign LUT_3[41815] = 32'b00000000000000000111101000001011;
assign LUT_3[41816] = 32'b00000000000000000111000000011010;
assign LUT_3[41817] = 32'b00000000000000001101101011110111;
assign LUT_3[41818] = 32'b00000000000000001001000111111110;
assign LUT_3[41819] = 32'b00000000000000001111110011011011;
assign LUT_3[41820] = 32'b00000000000000000100001110010000;
assign LUT_3[41821] = 32'b00000000000000001010111001101101;
assign LUT_3[41822] = 32'b00000000000000000110010101110100;
assign LUT_3[41823] = 32'b00000000000000001101000001010001;
assign LUT_3[41824] = 32'b11111111111111111111100010110001;
assign LUT_3[41825] = 32'b00000000000000000110001110001110;
assign LUT_3[41826] = 32'b00000000000000000001101010010101;
assign LUT_3[41827] = 32'b00000000000000001000010101110010;
assign LUT_3[41828] = 32'b11111111111111111100110000100111;
assign LUT_3[41829] = 32'b00000000000000000011011100000100;
assign LUT_3[41830] = 32'b11111111111111111110111000001011;
assign LUT_3[41831] = 32'b00000000000000000101100011101000;
assign LUT_3[41832] = 32'b00000000000000000100111011110111;
assign LUT_3[41833] = 32'b00000000000000001011100111010100;
assign LUT_3[41834] = 32'b00000000000000000111000011011011;
assign LUT_3[41835] = 32'b00000000000000001101101110111000;
assign LUT_3[41836] = 32'b00000000000000000010001001101101;
assign LUT_3[41837] = 32'b00000000000000001000110101001010;
assign LUT_3[41838] = 32'b00000000000000000100010001010001;
assign LUT_3[41839] = 32'b00000000000000001010111100101110;
assign LUT_3[41840] = 32'b00000000000000000010110101110100;
assign LUT_3[41841] = 32'b00000000000000001001100001010001;
assign LUT_3[41842] = 32'b00000000000000000100111101011000;
assign LUT_3[41843] = 32'b00000000000000001011101000110101;
assign LUT_3[41844] = 32'b00000000000000000000000011101010;
assign LUT_3[41845] = 32'b00000000000000000110101111000111;
assign LUT_3[41846] = 32'b00000000000000000010001011001110;
assign LUT_3[41847] = 32'b00000000000000001000110110101011;
assign LUT_3[41848] = 32'b00000000000000001000001110111010;
assign LUT_3[41849] = 32'b00000000000000001110111010010111;
assign LUT_3[41850] = 32'b00000000000000001010010110011110;
assign LUT_3[41851] = 32'b00000000000000010001000001111011;
assign LUT_3[41852] = 32'b00000000000000000101011100110000;
assign LUT_3[41853] = 32'b00000000000000001100001000001101;
assign LUT_3[41854] = 32'b00000000000000000111100100010100;
assign LUT_3[41855] = 32'b00000000000000001110001111110001;
assign LUT_3[41856] = 32'b00000000000000000000100110100100;
assign LUT_3[41857] = 32'b00000000000000000111010010000001;
assign LUT_3[41858] = 32'b00000000000000000010101110001000;
assign LUT_3[41859] = 32'b00000000000000001001011001100101;
assign LUT_3[41860] = 32'b11111111111111111101110100011010;
assign LUT_3[41861] = 32'b00000000000000000100011111110111;
assign LUT_3[41862] = 32'b11111111111111111111111011111110;
assign LUT_3[41863] = 32'b00000000000000000110100111011011;
assign LUT_3[41864] = 32'b00000000000000000101111111101010;
assign LUT_3[41865] = 32'b00000000000000001100101011000111;
assign LUT_3[41866] = 32'b00000000000000001000000111001110;
assign LUT_3[41867] = 32'b00000000000000001110110010101011;
assign LUT_3[41868] = 32'b00000000000000000011001101100000;
assign LUT_3[41869] = 32'b00000000000000001001111000111101;
assign LUT_3[41870] = 32'b00000000000000000101010101000100;
assign LUT_3[41871] = 32'b00000000000000001100000000100001;
assign LUT_3[41872] = 32'b00000000000000000011111001100111;
assign LUT_3[41873] = 32'b00000000000000001010100101000100;
assign LUT_3[41874] = 32'b00000000000000000110000001001011;
assign LUT_3[41875] = 32'b00000000000000001100101100101000;
assign LUT_3[41876] = 32'b00000000000000000001000111011101;
assign LUT_3[41877] = 32'b00000000000000000111110010111010;
assign LUT_3[41878] = 32'b00000000000000000011001111000001;
assign LUT_3[41879] = 32'b00000000000000001001111010011110;
assign LUT_3[41880] = 32'b00000000000000001001010010101101;
assign LUT_3[41881] = 32'b00000000000000001111111110001010;
assign LUT_3[41882] = 32'b00000000000000001011011010010001;
assign LUT_3[41883] = 32'b00000000000000010010000101101110;
assign LUT_3[41884] = 32'b00000000000000000110100000100011;
assign LUT_3[41885] = 32'b00000000000000001101001100000000;
assign LUT_3[41886] = 32'b00000000000000001000101000000111;
assign LUT_3[41887] = 32'b00000000000000001111010011100100;
assign LUT_3[41888] = 32'b00000000000000000001110101000100;
assign LUT_3[41889] = 32'b00000000000000001000100000100001;
assign LUT_3[41890] = 32'b00000000000000000011111100101000;
assign LUT_3[41891] = 32'b00000000000000001010101000000101;
assign LUT_3[41892] = 32'b11111111111111111111000010111010;
assign LUT_3[41893] = 32'b00000000000000000101101110010111;
assign LUT_3[41894] = 32'b00000000000000000001001010011110;
assign LUT_3[41895] = 32'b00000000000000000111110101111011;
assign LUT_3[41896] = 32'b00000000000000000111001110001010;
assign LUT_3[41897] = 32'b00000000000000001101111001100111;
assign LUT_3[41898] = 32'b00000000000000001001010101101110;
assign LUT_3[41899] = 32'b00000000000000010000000001001011;
assign LUT_3[41900] = 32'b00000000000000000100011100000000;
assign LUT_3[41901] = 32'b00000000000000001011000111011101;
assign LUT_3[41902] = 32'b00000000000000000110100011100100;
assign LUT_3[41903] = 32'b00000000000000001101001111000001;
assign LUT_3[41904] = 32'b00000000000000000101001000000111;
assign LUT_3[41905] = 32'b00000000000000001011110011100100;
assign LUT_3[41906] = 32'b00000000000000000111001111101011;
assign LUT_3[41907] = 32'b00000000000000001101111011001000;
assign LUT_3[41908] = 32'b00000000000000000010010101111101;
assign LUT_3[41909] = 32'b00000000000000001001000001011010;
assign LUT_3[41910] = 32'b00000000000000000100011101100001;
assign LUT_3[41911] = 32'b00000000000000001011001000111110;
assign LUT_3[41912] = 32'b00000000000000001010100001001101;
assign LUT_3[41913] = 32'b00000000000000010001001100101010;
assign LUT_3[41914] = 32'b00000000000000001100101000110001;
assign LUT_3[41915] = 32'b00000000000000010011010100001110;
assign LUT_3[41916] = 32'b00000000000000000111101111000011;
assign LUT_3[41917] = 32'b00000000000000001110011010100000;
assign LUT_3[41918] = 32'b00000000000000001001110110100111;
assign LUT_3[41919] = 32'b00000000000000010000100010000100;
assign LUT_3[41920] = 32'b00000000000000000000011111001111;
assign LUT_3[41921] = 32'b00000000000000000111001010101100;
assign LUT_3[41922] = 32'b00000000000000000010100110110011;
assign LUT_3[41923] = 32'b00000000000000001001010010010000;
assign LUT_3[41924] = 32'b11111111111111111101101101000101;
assign LUT_3[41925] = 32'b00000000000000000100011000100010;
assign LUT_3[41926] = 32'b11111111111111111111110100101001;
assign LUT_3[41927] = 32'b00000000000000000110100000000110;
assign LUT_3[41928] = 32'b00000000000000000101111000010101;
assign LUT_3[41929] = 32'b00000000000000001100100011110010;
assign LUT_3[41930] = 32'b00000000000000000111111111111001;
assign LUT_3[41931] = 32'b00000000000000001110101011010110;
assign LUT_3[41932] = 32'b00000000000000000011000110001011;
assign LUT_3[41933] = 32'b00000000000000001001110001101000;
assign LUT_3[41934] = 32'b00000000000000000101001101101111;
assign LUT_3[41935] = 32'b00000000000000001011111001001100;
assign LUT_3[41936] = 32'b00000000000000000011110010010010;
assign LUT_3[41937] = 32'b00000000000000001010011101101111;
assign LUT_3[41938] = 32'b00000000000000000101111001110110;
assign LUT_3[41939] = 32'b00000000000000001100100101010011;
assign LUT_3[41940] = 32'b00000000000000000001000000001000;
assign LUT_3[41941] = 32'b00000000000000000111101011100101;
assign LUT_3[41942] = 32'b00000000000000000011000111101100;
assign LUT_3[41943] = 32'b00000000000000001001110011001001;
assign LUT_3[41944] = 32'b00000000000000001001001011011000;
assign LUT_3[41945] = 32'b00000000000000001111110110110101;
assign LUT_3[41946] = 32'b00000000000000001011010010111100;
assign LUT_3[41947] = 32'b00000000000000010001111110011001;
assign LUT_3[41948] = 32'b00000000000000000110011001001110;
assign LUT_3[41949] = 32'b00000000000000001101000100101011;
assign LUT_3[41950] = 32'b00000000000000001000100000110010;
assign LUT_3[41951] = 32'b00000000000000001111001100001111;
assign LUT_3[41952] = 32'b00000000000000000001101101101111;
assign LUT_3[41953] = 32'b00000000000000001000011001001100;
assign LUT_3[41954] = 32'b00000000000000000011110101010011;
assign LUT_3[41955] = 32'b00000000000000001010100000110000;
assign LUT_3[41956] = 32'b11111111111111111110111011100101;
assign LUT_3[41957] = 32'b00000000000000000101100111000010;
assign LUT_3[41958] = 32'b00000000000000000001000011001001;
assign LUT_3[41959] = 32'b00000000000000000111101110100110;
assign LUT_3[41960] = 32'b00000000000000000111000110110101;
assign LUT_3[41961] = 32'b00000000000000001101110010010010;
assign LUT_3[41962] = 32'b00000000000000001001001110011001;
assign LUT_3[41963] = 32'b00000000000000001111111001110110;
assign LUT_3[41964] = 32'b00000000000000000100010100101011;
assign LUT_3[41965] = 32'b00000000000000001011000000001000;
assign LUT_3[41966] = 32'b00000000000000000110011100001111;
assign LUT_3[41967] = 32'b00000000000000001101000111101100;
assign LUT_3[41968] = 32'b00000000000000000101000000110010;
assign LUT_3[41969] = 32'b00000000000000001011101100001111;
assign LUT_3[41970] = 32'b00000000000000000111001000010110;
assign LUT_3[41971] = 32'b00000000000000001101110011110011;
assign LUT_3[41972] = 32'b00000000000000000010001110101000;
assign LUT_3[41973] = 32'b00000000000000001000111010000101;
assign LUT_3[41974] = 32'b00000000000000000100010110001100;
assign LUT_3[41975] = 32'b00000000000000001011000001101001;
assign LUT_3[41976] = 32'b00000000000000001010011001111000;
assign LUT_3[41977] = 32'b00000000000000010001000101010101;
assign LUT_3[41978] = 32'b00000000000000001100100001011100;
assign LUT_3[41979] = 32'b00000000000000010011001100111001;
assign LUT_3[41980] = 32'b00000000000000000111100111101110;
assign LUT_3[41981] = 32'b00000000000000001110010011001011;
assign LUT_3[41982] = 32'b00000000000000001001101111010010;
assign LUT_3[41983] = 32'b00000000000000010000011010101111;
assign LUT_3[41984] = 32'b00000000000000000101011011110110;
assign LUT_3[41985] = 32'b00000000000000001100000111010011;
assign LUT_3[41986] = 32'b00000000000000000111100011011010;
assign LUT_3[41987] = 32'b00000000000000001110001110110111;
assign LUT_3[41988] = 32'b00000000000000000010101001101100;
assign LUT_3[41989] = 32'b00000000000000001001010101001001;
assign LUT_3[41990] = 32'b00000000000000000100110001010000;
assign LUT_3[41991] = 32'b00000000000000001011011100101101;
assign LUT_3[41992] = 32'b00000000000000001010110100111100;
assign LUT_3[41993] = 32'b00000000000000010001100000011001;
assign LUT_3[41994] = 32'b00000000000000001100111100100000;
assign LUT_3[41995] = 32'b00000000000000010011100111111101;
assign LUT_3[41996] = 32'b00000000000000001000000010110010;
assign LUT_3[41997] = 32'b00000000000000001110101110001111;
assign LUT_3[41998] = 32'b00000000000000001010001010010110;
assign LUT_3[41999] = 32'b00000000000000010000110101110011;
assign LUT_3[42000] = 32'b00000000000000001000101110111001;
assign LUT_3[42001] = 32'b00000000000000001111011010010110;
assign LUT_3[42002] = 32'b00000000000000001010110110011101;
assign LUT_3[42003] = 32'b00000000000000010001100001111010;
assign LUT_3[42004] = 32'b00000000000000000101111100101111;
assign LUT_3[42005] = 32'b00000000000000001100101000001100;
assign LUT_3[42006] = 32'b00000000000000001000000100010011;
assign LUT_3[42007] = 32'b00000000000000001110101111110000;
assign LUT_3[42008] = 32'b00000000000000001110000111111111;
assign LUT_3[42009] = 32'b00000000000000010100110011011100;
assign LUT_3[42010] = 32'b00000000000000010000001111100011;
assign LUT_3[42011] = 32'b00000000000000010110111011000000;
assign LUT_3[42012] = 32'b00000000000000001011010101110101;
assign LUT_3[42013] = 32'b00000000000000010010000001010010;
assign LUT_3[42014] = 32'b00000000000000001101011101011001;
assign LUT_3[42015] = 32'b00000000000000010100001000110110;
assign LUT_3[42016] = 32'b00000000000000000110101010010110;
assign LUT_3[42017] = 32'b00000000000000001101010101110011;
assign LUT_3[42018] = 32'b00000000000000001000110001111010;
assign LUT_3[42019] = 32'b00000000000000001111011101010111;
assign LUT_3[42020] = 32'b00000000000000000011111000001100;
assign LUT_3[42021] = 32'b00000000000000001010100011101001;
assign LUT_3[42022] = 32'b00000000000000000101111111110000;
assign LUT_3[42023] = 32'b00000000000000001100101011001101;
assign LUT_3[42024] = 32'b00000000000000001100000011011100;
assign LUT_3[42025] = 32'b00000000000000010010101110111001;
assign LUT_3[42026] = 32'b00000000000000001110001011000000;
assign LUT_3[42027] = 32'b00000000000000010100110110011101;
assign LUT_3[42028] = 32'b00000000000000001001010001010010;
assign LUT_3[42029] = 32'b00000000000000001111111100101111;
assign LUT_3[42030] = 32'b00000000000000001011011000110110;
assign LUT_3[42031] = 32'b00000000000000010010000100010011;
assign LUT_3[42032] = 32'b00000000000000001001111101011001;
assign LUT_3[42033] = 32'b00000000000000010000101000110110;
assign LUT_3[42034] = 32'b00000000000000001100000100111101;
assign LUT_3[42035] = 32'b00000000000000010010110000011010;
assign LUT_3[42036] = 32'b00000000000000000111001011001111;
assign LUT_3[42037] = 32'b00000000000000001101110110101100;
assign LUT_3[42038] = 32'b00000000000000001001010010110011;
assign LUT_3[42039] = 32'b00000000000000001111111110010000;
assign LUT_3[42040] = 32'b00000000000000001111010110011111;
assign LUT_3[42041] = 32'b00000000000000010110000001111100;
assign LUT_3[42042] = 32'b00000000000000010001011110000011;
assign LUT_3[42043] = 32'b00000000000000011000001001100000;
assign LUT_3[42044] = 32'b00000000000000001100100100010101;
assign LUT_3[42045] = 32'b00000000000000010011001111110010;
assign LUT_3[42046] = 32'b00000000000000001110101011111001;
assign LUT_3[42047] = 32'b00000000000000010101010111010110;
assign LUT_3[42048] = 32'b00000000000000000101010100100001;
assign LUT_3[42049] = 32'b00000000000000001011111111111110;
assign LUT_3[42050] = 32'b00000000000000000111011100000101;
assign LUT_3[42051] = 32'b00000000000000001110000111100010;
assign LUT_3[42052] = 32'b00000000000000000010100010010111;
assign LUT_3[42053] = 32'b00000000000000001001001101110100;
assign LUT_3[42054] = 32'b00000000000000000100101001111011;
assign LUT_3[42055] = 32'b00000000000000001011010101011000;
assign LUT_3[42056] = 32'b00000000000000001010101101100111;
assign LUT_3[42057] = 32'b00000000000000010001011001000100;
assign LUT_3[42058] = 32'b00000000000000001100110101001011;
assign LUT_3[42059] = 32'b00000000000000010011100000101000;
assign LUT_3[42060] = 32'b00000000000000000111111011011101;
assign LUT_3[42061] = 32'b00000000000000001110100110111010;
assign LUT_3[42062] = 32'b00000000000000001010000011000001;
assign LUT_3[42063] = 32'b00000000000000010000101110011110;
assign LUT_3[42064] = 32'b00000000000000001000100111100100;
assign LUT_3[42065] = 32'b00000000000000001111010011000001;
assign LUT_3[42066] = 32'b00000000000000001010101111001000;
assign LUT_3[42067] = 32'b00000000000000010001011010100101;
assign LUT_3[42068] = 32'b00000000000000000101110101011010;
assign LUT_3[42069] = 32'b00000000000000001100100000110111;
assign LUT_3[42070] = 32'b00000000000000000111111100111110;
assign LUT_3[42071] = 32'b00000000000000001110101000011011;
assign LUT_3[42072] = 32'b00000000000000001110000000101010;
assign LUT_3[42073] = 32'b00000000000000010100101100000111;
assign LUT_3[42074] = 32'b00000000000000010000001000001110;
assign LUT_3[42075] = 32'b00000000000000010110110011101011;
assign LUT_3[42076] = 32'b00000000000000001011001110100000;
assign LUT_3[42077] = 32'b00000000000000010001111001111101;
assign LUT_3[42078] = 32'b00000000000000001101010110000100;
assign LUT_3[42079] = 32'b00000000000000010100000001100001;
assign LUT_3[42080] = 32'b00000000000000000110100011000001;
assign LUT_3[42081] = 32'b00000000000000001101001110011110;
assign LUT_3[42082] = 32'b00000000000000001000101010100101;
assign LUT_3[42083] = 32'b00000000000000001111010110000010;
assign LUT_3[42084] = 32'b00000000000000000011110000110111;
assign LUT_3[42085] = 32'b00000000000000001010011100010100;
assign LUT_3[42086] = 32'b00000000000000000101111000011011;
assign LUT_3[42087] = 32'b00000000000000001100100011111000;
assign LUT_3[42088] = 32'b00000000000000001011111100000111;
assign LUT_3[42089] = 32'b00000000000000010010100111100100;
assign LUT_3[42090] = 32'b00000000000000001110000011101011;
assign LUT_3[42091] = 32'b00000000000000010100101111001000;
assign LUT_3[42092] = 32'b00000000000000001001001001111101;
assign LUT_3[42093] = 32'b00000000000000001111110101011010;
assign LUT_3[42094] = 32'b00000000000000001011010001100001;
assign LUT_3[42095] = 32'b00000000000000010001111100111110;
assign LUT_3[42096] = 32'b00000000000000001001110110000100;
assign LUT_3[42097] = 32'b00000000000000010000100001100001;
assign LUT_3[42098] = 32'b00000000000000001011111101101000;
assign LUT_3[42099] = 32'b00000000000000010010101001000101;
assign LUT_3[42100] = 32'b00000000000000000111000011111010;
assign LUT_3[42101] = 32'b00000000000000001101101111010111;
assign LUT_3[42102] = 32'b00000000000000001001001011011110;
assign LUT_3[42103] = 32'b00000000000000001111110110111011;
assign LUT_3[42104] = 32'b00000000000000001111001111001010;
assign LUT_3[42105] = 32'b00000000000000010101111010100111;
assign LUT_3[42106] = 32'b00000000000000010001010110101110;
assign LUT_3[42107] = 32'b00000000000000011000000010001011;
assign LUT_3[42108] = 32'b00000000000000001100011101000000;
assign LUT_3[42109] = 32'b00000000000000010011001000011101;
assign LUT_3[42110] = 32'b00000000000000001110100100100100;
assign LUT_3[42111] = 32'b00000000000000010101010000000001;
assign LUT_3[42112] = 32'b00000000000000000111100110110100;
assign LUT_3[42113] = 32'b00000000000000001110010010010001;
assign LUT_3[42114] = 32'b00000000000000001001101110011000;
assign LUT_3[42115] = 32'b00000000000000010000011001110101;
assign LUT_3[42116] = 32'b00000000000000000100110100101010;
assign LUT_3[42117] = 32'b00000000000000001011100000000111;
assign LUT_3[42118] = 32'b00000000000000000110111100001110;
assign LUT_3[42119] = 32'b00000000000000001101100111101011;
assign LUT_3[42120] = 32'b00000000000000001100111111111010;
assign LUT_3[42121] = 32'b00000000000000010011101011010111;
assign LUT_3[42122] = 32'b00000000000000001111000111011110;
assign LUT_3[42123] = 32'b00000000000000010101110010111011;
assign LUT_3[42124] = 32'b00000000000000001010001101110000;
assign LUT_3[42125] = 32'b00000000000000010000111001001101;
assign LUT_3[42126] = 32'b00000000000000001100010101010100;
assign LUT_3[42127] = 32'b00000000000000010011000000110001;
assign LUT_3[42128] = 32'b00000000000000001010111001110111;
assign LUT_3[42129] = 32'b00000000000000010001100101010100;
assign LUT_3[42130] = 32'b00000000000000001101000001011011;
assign LUT_3[42131] = 32'b00000000000000010011101100111000;
assign LUT_3[42132] = 32'b00000000000000001000000111101101;
assign LUT_3[42133] = 32'b00000000000000001110110011001010;
assign LUT_3[42134] = 32'b00000000000000001010001111010001;
assign LUT_3[42135] = 32'b00000000000000010000111010101110;
assign LUT_3[42136] = 32'b00000000000000010000010010111101;
assign LUT_3[42137] = 32'b00000000000000010110111110011010;
assign LUT_3[42138] = 32'b00000000000000010010011010100001;
assign LUT_3[42139] = 32'b00000000000000011001000101111110;
assign LUT_3[42140] = 32'b00000000000000001101100000110011;
assign LUT_3[42141] = 32'b00000000000000010100001100010000;
assign LUT_3[42142] = 32'b00000000000000001111101000010111;
assign LUT_3[42143] = 32'b00000000000000010110010011110100;
assign LUT_3[42144] = 32'b00000000000000001000110101010100;
assign LUT_3[42145] = 32'b00000000000000001111100000110001;
assign LUT_3[42146] = 32'b00000000000000001010111100111000;
assign LUT_3[42147] = 32'b00000000000000010001101000010101;
assign LUT_3[42148] = 32'b00000000000000000110000011001010;
assign LUT_3[42149] = 32'b00000000000000001100101110100111;
assign LUT_3[42150] = 32'b00000000000000001000001010101110;
assign LUT_3[42151] = 32'b00000000000000001110110110001011;
assign LUT_3[42152] = 32'b00000000000000001110001110011010;
assign LUT_3[42153] = 32'b00000000000000010100111001110111;
assign LUT_3[42154] = 32'b00000000000000010000010101111110;
assign LUT_3[42155] = 32'b00000000000000010111000001011011;
assign LUT_3[42156] = 32'b00000000000000001011011100010000;
assign LUT_3[42157] = 32'b00000000000000010010000111101101;
assign LUT_3[42158] = 32'b00000000000000001101100011110100;
assign LUT_3[42159] = 32'b00000000000000010100001111010001;
assign LUT_3[42160] = 32'b00000000000000001100001000010111;
assign LUT_3[42161] = 32'b00000000000000010010110011110100;
assign LUT_3[42162] = 32'b00000000000000001110001111111011;
assign LUT_3[42163] = 32'b00000000000000010100111011011000;
assign LUT_3[42164] = 32'b00000000000000001001010110001101;
assign LUT_3[42165] = 32'b00000000000000010000000001101010;
assign LUT_3[42166] = 32'b00000000000000001011011101110001;
assign LUT_3[42167] = 32'b00000000000000010010001001001110;
assign LUT_3[42168] = 32'b00000000000000010001100001011101;
assign LUT_3[42169] = 32'b00000000000000011000001100111010;
assign LUT_3[42170] = 32'b00000000000000010011101001000001;
assign LUT_3[42171] = 32'b00000000000000011010010100011110;
assign LUT_3[42172] = 32'b00000000000000001110101111010011;
assign LUT_3[42173] = 32'b00000000000000010101011010110000;
assign LUT_3[42174] = 32'b00000000000000010000110110110111;
assign LUT_3[42175] = 32'b00000000000000010111100010010100;
assign LUT_3[42176] = 32'b00000000000000000111011111011111;
assign LUT_3[42177] = 32'b00000000000000001110001010111100;
assign LUT_3[42178] = 32'b00000000000000001001100111000011;
assign LUT_3[42179] = 32'b00000000000000010000010010100000;
assign LUT_3[42180] = 32'b00000000000000000100101101010101;
assign LUT_3[42181] = 32'b00000000000000001011011000110010;
assign LUT_3[42182] = 32'b00000000000000000110110100111001;
assign LUT_3[42183] = 32'b00000000000000001101100000010110;
assign LUT_3[42184] = 32'b00000000000000001100111000100101;
assign LUT_3[42185] = 32'b00000000000000010011100100000010;
assign LUT_3[42186] = 32'b00000000000000001111000000001001;
assign LUT_3[42187] = 32'b00000000000000010101101011100110;
assign LUT_3[42188] = 32'b00000000000000001010000110011011;
assign LUT_3[42189] = 32'b00000000000000010000110001111000;
assign LUT_3[42190] = 32'b00000000000000001100001101111111;
assign LUT_3[42191] = 32'b00000000000000010010111001011100;
assign LUT_3[42192] = 32'b00000000000000001010110010100010;
assign LUT_3[42193] = 32'b00000000000000010001011101111111;
assign LUT_3[42194] = 32'b00000000000000001100111010000110;
assign LUT_3[42195] = 32'b00000000000000010011100101100011;
assign LUT_3[42196] = 32'b00000000000000001000000000011000;
assign LUT_3[42197] = 32'b00000000000000001110101011110101;
assign LUT_3[42198] = 32'b00000000000000001010000111111100;
assign LUT_3[42199] = 32'b00000000000000010000110011011001;
assign LUT_3[42200] = 32'b00000000000000010000001011101000;
assign LUT_3[42201] = 32'b00000000000000010110110111000101;
assign LUT_3[42202] = 32'b00000000000000010010010011001100;
assign LUT_3[42203] = 32'b00000000000000011000111110101001;
assign LUT_3[42204] = 32'b00000000000000001101011001011110;
assign LUT_3[42205] = 32'b00000000000000010100000100111011;
assign LUT_3[42206] = 32'b00000000000000001111100001000010;
assign LUT_3[42207] = 32'b00000000000000010110001100011111;
assign LUT_3[42208] = 32'b00000000000000001000101101111111;
assign LUT_3[42209] = 32'b00000000000000001111011001011100;
assign LUT_3[42210] = 32'b00000000000000001010110101100011;
assign LUT_3[42211] = 32'b00000000000000010001100001000000;
assign LUT_3[42212] = 32'b00000000000000000101111011110101;
assign LUT_3[42213] = 32'b00000000000000001100100111010010;
assign LUT_3[42214] = 32'b00000000000000001000000011011001;
assign LUT_3[42215] = 32'b00000000000000001110101110110110;
assign LUT_3[42216] = 32'b00000000000000001110000111000101;
assign LUT_3[42217] = 32'b00000000000000010100110010100010;
assign LUT_3[42218] = 32'b00000000000000010000001110101001;
assign LUT_3[42219] = 32'b00000000000000010110111010000110;
assign LUT_3[42220] = 32'b00000000000000001011010100111011;
assign LUT_3[42221] = 32'b00000000000000010010000000011000;
assign LUT_3[42222] = 32'b00000000000000001101011100011111;
assign LUT_3[42223] = 32'b00000000000000010100000111111100;
assign LUT_3[42224] = 32'b00000000000000001100000001000010;
assign LUT_3[42225] = 32'b00000000000000010010101100011111;
assign LUT_3[42226] = 32'b00000000000000001110001000100110;
assign LUT_3[42227] = 32'b00000000000000010100110100000011;
assign LUT_3[42228] = 32'b00000000000000001001001110111000;
assign LUT_3[42229] = 32'b00000000000000001111111010010101;
assign LUT_3[42230] = 32'b00000000000000001011010110011100;
assign LUT_3[42231] = 32'b00000000000000010010000001111001;
assign LUT_3[42232] = 32'b00000000000000010001011010001000;
assign LUT_3[42233] = 32'b00000000000000011000000101100101;
assign LUT_3[42234] = 32'b00000000000000010011100001101100;
assign LUT_3[42235] = 32'b00000000000000011010001101001001;
assign LUT_3[42236] = 32'b00000000000000001110100111111110;
assign LUT_3[42237] = 32'b00000000000000010101010011011011;
assign LUT_3[42238] = 32'b00000000000000010000101111100010;
assign LUT_3[42239] = 32'b00000000000000010111011010111111;
assign LUT_3[42240] = 32'b00000000000000000001101011010111;
assign LUT_3[42241] = 32'b00000000000000001000010110110100;
assign LUT_3[42242] = 32'b00000000000000000011110010111011;
assign LUT_3[42243] = 32'b00000000000000001010011110011000;
assign LUT_3[42244] = 32'b11111111111111111110111001001101;
assign LUT_3[42245] = 32'b00000000000000000101100100101010;
assign LUT_3[42246] = 32'b00000000000000000001000000110001;
assign LUT_3[42247] = 32'b00000000000000000111101100001110;
assign LUT_3[42248] = 32'b00000000000000000111000100011101;
assign LUT_3[42249] = 32'b00000000000000001101101111111010;
assign LUT_3[42250] = 32'b00000000000000001001001100000001;
assign LUT_3[42251] = 32'b00000000000000001111110111011110;
assign LUT_3[42252] = 32'b00000000000000000100010010010011;
assign LUT_3[42253] = 32'b00000000000000001010111101110000;
assign LUT_3[42254] = 32'b00000000000000000110011001110111;
assign LUT_3[42255] = 32'b00000000000000001101000101010100;
assign LUT_3[42256] = 32'b00000000000000000100111110011010;
assign LUT_3[42257] = 32'b00000000000000001011101001110111;
assign LUT_3[42258] = 32'b00000000000000000111000101111110;
assign LUT_3[42259] = 32'b00000000000000001101110001011011;
assign LUT_3[42260] = 32'b00000000000000000010001100010000;
assign LUT_3[42261] = 32'b00000000000000001000110111101101;
assign LUT_3[42262] = 32'b00000000000000000100010011110100;
assign LUT_3[42263] = 32'b00000000000000001010111111010001;
assign LUT_3[42264] = 32'b00000000000000001010010111100000;
assign LUT_3[42265] = 32'b00000000000000010001000010111101;
assign LUT_3[42266] = 32'b00000000000000001100011111000100;
assign LUT_3[42267] = 32'b00000000000000010011001010100001;
assign LUT_3[42268] = 32'b00000000000000000111100101010110;
assign LUT_3[42269] = 32'b00000000000000001110010000110011;
assign LUT_3[42270] = 32'b00000000000000001001101100111010;
assign LUT_3[42271] = 32'b00000000000000010000011000010111;
assign LUT_3[42272] = 32'b00000000000000000010111001110111;
assign LUT_3[42273] = 32'b00000000000000001001100101010100;
assign LUT_3[42274] = 32'b00000000000000000101000001011011;
assign LUT_3[42275] = 32'b00000000000000001011101100111000;
assign LUT_3[42276] = 32'b00000000000000000000000111101101;
assign LUT_3[42277] = 32'b00000000000000000110110011001010;
assign LUT_3[42278] = 32'b00000000000000000010001111010001;
assign LUT_3[42279] = 32'b00000000000000001000111010101110;
assign LUT_3[42280] = 32'b00000000000000001000010010111101;
assign LUT_3[42281] = 32'b00000000000000001110111110011010;
assign LUT_3[42282] = 32'b00000000000000001010011010100001;
assign LUT_3[42283] = 32'b00000000000000010001000101111110;
assign LUT_3[42284] = 32'b00000000000000000101100000110011;
assign LUT_3[42285] = 32'b00000000000000001100001100010000;
assign LUT_3[42286] = 32'b00000000000000000111101000010111;
assign LUT_3[42287] = 32'b00000000000000001110010011110100;
assign LUT_3[42288] = 32'b00000000000000000110001100111010;
assign LUT_3[42289] = 32'b00000000000000001100111000010111;
assign LUT_3[42290] = 32'b00000000000000001000010100011110;
assign LUT_3[42291] = 32'b00000000000000001110111111111011;
assign LUT_3[42292] = 32'b00000000000000000011011010110000;
assign LUT_3[42293] = 32'b00000000000000001010000110001101;
assign LUT_3[42294] = 32'b00000000000000000101100010010100;
assign LUT_3[42295] = 32'b00000000000000001100001101110001;
assign LUT_3[42296] = 32'b00000000000000001011100110000000;
assign LUT_3[42297] = 32'b00000000000000010010010001011101;
assign LUT_3[42298] = 32'b00000000000000001101101101100100;
assign LUT_3[42299] = 32'b00000000000000010100011001000001;
assign LUT_3[42300] = 32'b00000000000000001000110011110110;
assign LUT_3[42301] = 32'b00000000000000001111011111010011;
assign LUT_3[42302] = 32'b00000000000000001010111011011010;
assign LUT_3[42303] = 32'b00000000000000010001100110110111;
assign LUT_3[42304] = 32'b00000000000000000001100100000010;
assign LUT_3[42305] = 32'b00000000000000001000001111011111;
assign LUT_3[42306] = 32'b00000000000000000011101011100110;
assign LUT_3[42307] = 32'b00000000000000001010010111000011;
assign LUT_3[42308] = 32'b11111111111111111110110001111000;
assign LUT_3[42309] = 32'b00000000000000000101011101010101;
assign LUT_3[42310] = 32'b00000000000000000000111001011100;
assign LUT_3[42311] = 32'b00000000000000000111100100111001;
assign LUT_3[42312] = 32'b00000000000000000110111101001000;
assign LUT_3[42313] = 32'b00000000000000001101101000100101;
assign LUT_3[42314] = 32'b00000000000000001001000100101100;
assign LUT_3[42315] = 32'b00000000000000001111110000001001;
assign LUT_3[42316] = 32'b00000000000000000100001010111110;
assign LUT_3[42317] = 32'b00000000000000001010110110011011;
assign LUT_3[42318] = 32'b00000000000000000110010010100010;
assign LUT_3[42319] = 32'b00000000000000001100111101111111;
assign LUT_3[42320] = 32'b00000000000000000100110111000101;
assign LUT_3[42321] = 32'b00000000000000001011100010100010;
assign LUT_3[42322] = 32'b00000000000000000110111110101001;
assign LUT_3[42323] = 32'b00000000000000001101101010000110;
assign LUT_3[42324] = 32'b00000000000000000010000100111011;
assign LUT_3[42325] = 32'b00000000000000001000110000011000;
assign LUT_3[42326] = 32'b00000000000000000100001100011111;
assign LUT_3[42327] = 32'b00000000000000001010110111111100;
assign LUT_3[42328] = 32'b00000000000000001010010000001011;
assign LUT_3[42329] = 32'b00000000000000010000111011101000;
assign LUT_3[42330] = 32'b00000000000000001100010111101111;
assign LUT_3[42331] = 32'b00000000000000010011000011001100;
assign LUT_3[42332] = 32'b00000000000000000111011110000001;
assign LUT_3[42333] = 32'b00000000000000001110001001011110;
assign LUT_3[42334] = 32'b00000000000000001001100101100101;
assign LUT_3[42335] = 32'b00000000000000010000010001000010;
assign LUT_3[42336] = 32'b00000000000000000010110010100010;
assign LUT_3[42337] = 32'b00000000000000001001011101111111;
assign LUT_3[42338] = 32'b00000000000000000100111010000110;
assign LUT_3[42339] = 32'b00000000000000001011100101100011;
assign LUT_3[42340] = 32'b00000000000000000000000000011000;
assign LUT_3[42341] = 32'b00000000000000000110101011110101;
assign LUT_3[42342] = 32'b00000000000000000010000111111100;
assign LUT_3[42343] = 32'b00000000000000001000110011011001;
assign LUT_3[42344] = 32'b00000000000000001000001011101000;
assign LUT_3[42345] = 32'b00000000000000001110110111000101;
assign LUT_3[42346] = 32'b00000000000000001010010011001100;
assign LUT_3[42347] = 32'b00000000000000010000111110101001;
assign LUT_3[42348] = 32'b00000000000000000101011001011110;
assign LUT_3[42349] = 32'b00000000000000001100000100111011;
assign LUT_3[42350] = 32'b00000000000000000111100001000010;
assign LUT_3[42351] = 32'b00000000000000001110001100011111;
assign LUT_3[42352] = 32'b00000000000000000110000101100101;
assign LUT_3[42353] = 32'b00000000000000001100110001000010;
assign LUT_3[42354] = 32'b00000000000000001000001101001001;
assign LUT_3[42355] = 32'b00000000000000001110111000100110;
assign LUT_3[42356] = 32'b00000000000000000011010011011011;
assign LUT_3[42357] = 32'b00000000000000001001111110111000;
assign LUT_3[42358] = 32'b00000000000000000101011010111111;
assign LUT_3[42359] = 32'b00000000000000001100000110011100;
assign LUT_3[42360] = 32'b00000000000000001011011110101011;
assign LUT_3[42361] = 32'b00000000000000010010001010001000;
assign LUT_3[42362] = 32'b00000000000000001101100110001111;
assign LUT_3[42363] = 32'b00000000000000010100010001101100;
assign LUT_3[42364] = 32'b00000000000000001000101100100001;
assign LUT_3[42365] = 32'b00000000000000001111010111111110;
assign LUT_3[42366] = 32'b00000000000000001010110100000101;
assign LUT_3[42367] = 32'b00000000000000010001011111100010;
assign LUT_3[42368] = 32'b00000000000000000011110110010101;
assign LUT_3[42369] = 32'b00000000000000001010100001110010;
assign LUT_3[42370] = 32'b00000000000000000101111101111001;
assign LUT_3[42371] = 32'b00000000000000001100101001010110;
assign LUT_3[42372] = 32'b00000000000000000001000100001011;
assign LUT_3[42373] = 32'b00000000000000000111101111101000;
assign LUT_3[42374] = 32'b00000000000000000011001011101111;
assign LUT_3[42375] = 32'b00000000000000001001110111001100;
assign LUT_3[42376] = 32'b00000000000000001001001111011011;
assign LUT_3[42377] = 32'b00000000000000001111111010111000;
assign LUT_3[42378] = 32'b00000000000000001011010110111111;
assign LUT_3[42379] = 32'b00000000000000010010000010011100;
assign LUT_3[42380] = 32'b00000000000000000110011101010001;
assign LUT_3[42381] = 32'b00000000000000001101001000101110;
assign LUT_3[42382] = 32'b00000000000000001000100100110101;
assign LUT_3[42383] = 32'b00000000000000001111010000010010;
assign LUT_3[42384] = 32'b00000000000000000111001001011000;
assign LUT_3[42385] = 32'b00000000000000001101110100110101;
assign LUT_3[42386] = 32'b00000000000000001001010000111100;
assign LUT_3[42387] = 32'b00000000000000001111111100011001;
assign LUT_3[42388] = 32'b00000000000000000100010111001110;
assign LUT_3[42389] = 32'b00000000000000001011000010101011;
assign LUT_3[42390] = 32'b00000000000000000110011110110010;
assign LUT_3[42391] = 32'b00000000000000001101001010001111;
assign LUT_3[42392] = 32'b00000000000000001100100010011110;
assign LUT_3[42393] = 32'b00000000000000010011001101111011;
assign LUT_3[42394] = 32'b00000000000000001110101010000010;
assign LUT_3[42395] = 32'b00000000000000010101010101011111;
assign LUT_3[42396] = 32'b00000000000000001001110000010100;
assign LUT_3[42397] = 32'b00000000000000010000011011110001;
assign LUT_3[42398] = 32'b00000000000000001011110111111000;
assign LUT_3[42399] = 32'b00000000000000010010100011010101;
assign LUT_3[42400] = 32'b00000000000000000101000100110101;
assign LUT_3[42401] = 32'b00000000000000001011110000010010;
assign LUT_3[42402] = 32'b00000000000000000111001100011001;
assign LUT_3[42403] = 32'b00000000000000001101110111110110;
assign LUT_3[42404] = 32'b00000000000000000010010010101011;
assign LUT_3[42405] = 32'b00000000000000001000111110001000;
assign LUT_3[42406] = 32'b00000000000000000100011010001111;
assign LUT_3[42407] = 32'b00000000000000001011000101101100;
assign LUT_3[42408] = 32'b00000000000000001010011101111011;
assign LUT_3[42409] = 32'b00000000000000010001001001011000;
assign LUT_3[42410] = 32'b00000000000000001100100101011111;
assign LUT_3[42411] = 32'b00000000000000010011010000111100;
assign LUT_3[42412] = 32'b00000000000000000111101011110001;
assign LUT_3[42413] = 32'b00000000000000001110010111001110;
assign LUT_3[42414] = 32'b00000000000000001001110011010101;
assign LUT_3[42415] = 32'b00000000000000010000011110110010;
assign LUT_3[42416] = 32'b00000000000000001000010111111000;
assign LUT_3[42417] = 32'b00000000000000001111000011010101;
assign LUT_3[42418] = 32'b00000000000000001010011111011100;
assign LUT_3[42419] = 32'b00000000000000010001001010111001;
assign LUT_3[42420] = 32'b00000000000000000101100101101110;
assign LUT_3[42421] = 32'b00000000000000001100010001001011;
assign LUT_3[42422] = 32'b00000000000000000111101101010010;
assign LUT_3[42423] = 32'b00000000000000001110011000101111;
assign LUT_3[42424] = 32'b00000000000000001101110000111110;
assign LUT_3[42425] = 32'b00000000000000010100011100011011;
assign LUT_3[42426] = 32'b00000000000000001111111000100010;
assign LUT_3[42427] = 32'b00000000000000010110100011111111;
assign LUT_3[42428] = 32'b00000000000000001010111110110100;
assign LUT_3[42429] = 32'b00000000000000010001101010010001;
assign LUT_3[42430] = 32'b00000000000000001101000110011000;
assign LUT_3[42431] = 32'b00000000000000010011110001110101;
assign LUT_3[42432] = 32'b00000000000000000011101111000000;
assign LUT_3[42433] = 32'b00000000000000001010011010011101;
assign LUT_3[42434] = 32'b00000000000000000101110110100100;
assign LUT_3[42435] = 32'b00000000000000001100100010000001;
assign LUT_3[42436] = 32'b00000000000000000000111100110110;
assign LUT_3[42437] = 32'b00000000000000000111101000010011;
assign LUT_3[42438] = 32'b00000000000000000011000100011010;
assign LUT_3[42439] = 32'b00000000000000001001101111110111;
assign LUT_3[42440] = 32'b00000000000000001001001000000110;
assign LUT_3[42441] = 32'b00000000000000001111110011100011;
assign LUT_3[42442] = 32'b00000000000000001011001111101010;
assign LUT_3[42443] = 32'b00000000000000010001111011000111;
assign LUT_3[42444] = 32'b00000000000000000110010101111100;
assign LUT_3[42445] = 32'b00000000000000001101000001011001;
assign LUT_3[42446] = 32'b00000000000000001000011101100000;
assign LUT_3[42447] = 32'b00000000000000001111001000111101;
assign LUT_3[42448] = 32'b00000000000000000111000010000011;
assign LUT_3[42449] = 32'b00000000000000001101101101100000;
assign LUT_3[42450] = 32'b00000000000000001001001001100111;
assign LUT_3[42451] = 32'b00000000000000001111110101000100;
assign LUT_3[42452] = 32'b00000000000000000100001111111001;
assign LUT_3[42453] = 32'b00000000000000001010111011010110;
assign LUT_3[42454] = 32'b00000000000000000110010111011101;
assign LUT_3[42455] = 32'b00000000000000001101000010111010;
assign LUT_3[42456] = 32'b00000000000000001100011011001001;
assign LUT_3[42457] = 32'b00000000000000010011000110100110;
assign LUT_3[42458] = 32'b00000000000000001110100010101101;
assign LUT_3[42459] = 32'b00000000000000010101001110001010;
assign LUT_3[42460] = 32'b00000000000000001001101000111111;
assign LUT_3[42461] = 32'b00000000000000010000010100011100;
assign LUT_3[42462] = 32'b00000000000000001011110000100011;
assign LUT_3[42463] = 32'b00000000000000010010011100000000;
assign LUT_3[42464] = 32'b00000000000000000100111101100000;
assign LUT_3[42465] = 32'b00000000000000001011101000111101;
assign LUT_3[42466] = 32'b00000000000000000111000101000100;
assign LUT_3[42467] = 32'b00000000000000001101110000100001;
assign LUT_3[42468] = 32'b00000000000000000010001011010110;
assign LUT_3[42469] = 32'b00000000000000001000110110110011;
assign LUT_3[42470] = 32'b00000000000000000100010010111010;
assign LUT_3[42471] = 32'b00000000000000001010111110010111;
assign LUT_3[42472] = 32'b00000000000000001010010110100110;
assign LUT_3[42473] = 32'b00000000000000010001000010000011;
assign LUT_3[42474] = 32'b00000000000000001100011110001010;
assign LUT_3[42475] = 32'b00000000000000010011001001100111;
assign LUT_3[42476] = 32'b00000000000000000111100100011100;
assign LUT_3[42477] = 32'b00000000000000001110001111111001;
assign LUT_3[42478] = 32'b00000000000000001001101100000000;
assign LUT_3[42479] = 32'b00000000000000010000010111011101;
assign LUT_3[42480] = 32'b00000000000000001000010000100011;
assign LUT_3[42481] = 32'b00000000000000001110111100000000;
assign LUT_3[42482] = 32'b00000000000000001010011000000111;
assign LUT_3[42483] = 32'b00000000000000010001000011100100;
assign LUT_3[42484] = 32'b00000000000000000101011110011001;
assign LUT_3[42485] = 32'b00000000000000001100001001110110;
assign LUT_3[42486] = 32'b00000000000000000111100101111101;
assign LUT_3[42487] = 32'b00000000000000001110010001011010;
assign LUT_3[42488] = 32'b00000000000000001101101001101001;
assign LUT_3[42489] = 32'b00000000000000010100010101000110;
assign LUT_3[42490] = 32'b00000000000000001111110001001101;
assign LUT_3[42491] = 32'b00000000000000010110011100101010;
assign LUT_3[42492] = 32'b00000000000000001010110111011111;
assign LUT_3[42493] = 32'b00000000000000010001100010111100;
assign LUT_3[42494] = 32'b00000000000000001100111111000011;
assign LUT_3[42495] = 32'b00000000000000010011101010100000;
assign LUT_3[42496] = 32'b00000000000000001000110001000010;
assign LUT_3[42497] = 32'b00000000000000001111011100011111;
assign LUT_3[42498] = 32'b00000000000000001010111000100110;
assign LUT_3[42499] = 32'b00000000000000010001100100000011;
assign LUT_3[42500] = 32'b00000000000000000101111110111000;
assign LUT_3[42501] = 32'b00000000000000001100101010010101;
assign LUT_3[42502] = 32'b00000000000000001000000110011100;
assign LUT_3[42503] = 32'b00000000000000001110110001111001;
assign LUT_3[42504] = 32'b00000000000000001110001010001000;
assign LUT_3[42505] = 32'b00000000000000010100110101100101;
assign LUT_3[42506] = 32'b00000000000000010000010001101100;
assign LUT_3[42507] = 32'b00000000000000010110111101001001;
assign LUT_3[42508] = 32'b00000000000000001011010111111110;
assign LUT_3[42509] = 32'b00000000000000010010000011011011;
assign LUT_3[42510] = 32'b00000000000000001101011111100010;
assign LUT_3[42511] = 32'b00000000000000010100001010111111;
assign LUT_3[42512] = 32'b00000000000000001100000100000101;
assign LUT_3[42513] = 32'b00000000000000010010101111100010;
assign LUT_3[42514] = 32'b00000000000000001110001011101001;
assign LUT_3[42515] = 32'b00000000000000010100110111000110;
assign LUT_3[42516] = 32'b00000000000000001001010001111011;
assign LUT_3[42517] = 32'b00000000000000001111111101011000;
assign LUT_3[42518] = 32'b00000000000000001011011001011111;
assign LUT_3[42519] = 32'b00000000000000010010000100111100;
assign LUT_3[42520] = 32'b00000000000000010001011101001011;
assign LUT_3[42521] = 32'b00000000000000011000001000101000;
assign LUT_3[42522] = 32'b00000000000000010011100100101111;
assign LUT_3[42523] = 32'b00000000000000011010010000001100;
assign LUT_3[42524] = 32'b00000000000000001110101011000001;
assign LUT_3[42525] = 32'b00000000000000010101010110011110;
assign LUT_3[42526] = 32'b00000000000000010000110010100101;
assign LUT_3[42527] = 32'b00000000000000010111011110000010;
assign LUT_3[42528] = 32'b00000000000000001001111111100010;
assign LUT_3[42529] = 32'b00000000000000010000101010111111;
assign LUT_3[42530] = 32'b00000000000000001100000111000110;
assign LUT_3[42531] = 32'b00000000000000010010110010100011;
assign LUT_3[42532] = 32'b00000000000000000111001101011000;
assign LUT_3[42533] = 32'b00000000000000001101111000110101;
assign LUT_3[42534] = 32'b00000000000000001001010100111100;
assign LUT_3[42535] = 32'b00000000000000010000000000011001;
assign LUT_3[42536] = 32'b00000000000000001111011000101000;
assign LUT_3[42537] = 32'b00000000000000010110000100000101;
assign LUT_3[42538] = 32'b00000000000000010001100000001100;
assign LUT_3[42539] = 32'b00000000000000011000001011101001;
assign LUT_3[42540] = 32'b00000000000000001100100110011110;
assign LUT_3[42541] = 32'b00000000000000010011010001111011;
assign LUT_3[42542] = 32'b00000000000000001110101110000010;
assign LUT_3[42543] = 32'b00000000000000010101011001011111;
assign LUT_3[42544] = 32'b00000000000000001101010010100101;
assign LUT_3[42545] = 32'b00000000000000010011111110000010;
assign LUT_3[42546] = 32'b00000000000000001111011010001001;
assign LUT_3[42547] = 32'b00000000000000010110000101100110;
assign LUT_3[42548] = 32'b00000000000000001010100000011011;
assign LUT_3[42549] = 32'b00000000000000010001001011111000;
assign LUT_3[42550] = 32'b00000000000000001100100111111111;
assign LUT_3[42551] = 32'b00000000000000010011010011011100;
assign LUT_3[42552] = 32'b00000000000000010010101011101011;
assign LUT_3[42553] = 32'b00000000000000011001010111001000;
assign LUT_3[42554] = 32'b00000000000000010100110011001111;
assign LUT_3[42555] = 32'b00000000000000011011011110101100;
assign LUT_3[42556] = 32'b00000000000000001111111001100001;
assign LUT_3[42557] = 32'b00000000000000010110100100111110;
assign LUT_3[42558] = 32'b00000000000000010010000001000101;
assign LUT_3[42559] = 32'b00000000000000011000101100100010;
assign LUT_3[42560] = 32'b00000000000000001000101001101101;
assign LUT_3[42561] = 32'b00000000000000001111010101001010;
assign LUT_3[42562] = 32'b00000000000000001010110001010001;
assign LUT_3[42563] = 32'b00000000000000010001011100101110;
assign LUT_3[42564] = 32'b00000000000000000101110111100011;
assign LUT_3[42565] = 32'b00000000000000001100100011000000;
assign LUT_3[42566] = 32'b00000000000000000111111111000111;
assign LUT_3[42567] = 32'b00000000000000001110101010100100;
assign LUT_3[42568] = 32'b00000000000000001110000010110011;
assign LUT_3[42569] = 32'b00000000000000010100101110010000;
assign LUT_3[42570] = 32'b00000000000000010000001010010111;
assign LUT_3[42571] = 32'b00000000000000010110110101110100;
assign LUT_3[42572] = 32'b00000000000000001011010000101001;
assign LUT_3[42573] = 32'b00000000000000010001111100000110;
assign LUT_3[42574] = 32'b00000000000000001101011000001101;
assign LUT_3[42575] = 32'b00000000000000010100000011101010;
assign LUT_3[42576] = 32'b00000000000000001011111100110000;
assign LUT_3[42577] = 32'b00000000000000010010101000001101;
assign LUT_3[42578] = 32'b00000000000000001110000100010100;
assign LUT_3[42579] = 32'b00000000000000010100101111110001;
assign LUT_3[42580] = 32'b00000000000000001001001010100110;
assign LUT_3[42581] = 32'b00000000000000001111110110000011;
assign LUT_3[42582] = 32'b00000000000000001011010010001010;
assign LUT_3[42583] = 32'b00000000000000010001111101100111;
assign LUT_3[42584] = 32'b00000000000000010001010101110110;
assign LUT_3[42585] = 32'b00000000000000011000000001010011;
assign LUT_3[42586] = 32'b00000000000000010011011101011010;
assign LUT_3[42587] = 32'b00000000000000011010001000110111;
assign LUT_3[42588] = 32'b00000000000000001110100011101100;
assign LUT_3[42589] = 32'b00000000000000010101001111001001;
assign LUT_3[42590] = 32'b00000000000000010000101011010000;
assign LUT_3[42591] = 32'b00000000000000010111010110101101;
assign LUT_3[42592] = 32'b00000000000000001001111000001101;
assign LUT_3[42593] = 32'b00000000000000010000100011101010;
assign LUT_3[42594] = 32'b00000000000000001011111111110001;
assign LUT_3[42595] = 32'b00000000000000010010101011001110;
assign LUT_3[42596] = 32'b00000000000000000111000110000011;
assign LUT_3[42597] = 32'b00000000000000001101110001100000;
assign LUT_3[42598] = 32'b00000000000000001001001101100111;
assign LUT_3[42599] = 32'b00000000000000001111111001000100;
assign LUT_3[42600] = 32'b00000000000000001111010001010011;
assign LUT_3[42601] = 32'b00000000000000010101111100110000;
assign LUT_3[42602] = 32'b00000000000000010001011000110111;
assign LUT_3[42603] = 32'b00000000000000011000000100010100;
assign LUT_3[42604] = 32'b00000000000000001100011111001001;
assign LUT_3[42605] = 32'b00000000000000010011001010100110;
assign LUT_3[42606] = 32'b00000000000000001110100110101101;
assign LUT_3[42607] = 32'b00000000000000010101010010001010;
assign LUT_3[42608] = 32'b00000000000000001101001011010000;
assign LUT_3[42609] = 32'b00000000000000010011110110101101;
assign LUT_3[42610] = 32'b00000000000000001111010010110100;
assign LUT_3[42611] = 32'b00000000000000010101111110010001;
assign LUT_3[42612] = 32'b00000000000000001010011001000110;
assign LUT_3[42613] = 32'b00000000000000010001000100100011;
assign LUT_3[42614] = 32'b00000000000000001100100000101010;
assign LUT_3[42615] = 32'b00000000000000010011001100000111;
assign LUT_3[42616] = 32'b00000000000000010010100100010110;
assign LUT_3[42617] = 32'b00000000000000011001001111110011;
assign LUT_3[42618] = 32'b00000000000000010100101011111010;
assign LUT_3[42619] = 32'b00000000000000011011010111010111;
assign LUT_3[42620] = 32'b00000000000000001111110010001100;
assign LUT_3[42621] = 32'b00000000000000010110011101101001;
assign LUT_3[42622] = 32'b00000000000000010001111001110000;
assign LUT_3[42623] = 32'b00000000000000011000100101001101;
assign LUT_3[42624] = 32'b00000000000000001010111100000000;
assign LUT_3[42625] = 32'b00000000000000010001100111011101;
assign LUT_3[42626] = 32'b00000000000000001101000011100100;
assign LUT_3[42627] = 32'b00000000000000010011101111000001;
assign LUT_3[42628] = 32'b00000000000000001000001001110110;
assign LUT_3[42629] = 32'b00000000000000001110110101010011;
assign LUT_3[42630] = 32'b00000000000000001010010001011010;
assign LUT_3[42631] = 32'b00000000000000010000111100110111;
assign LUT_3[42632] = 32'b00000000000000010000010101000110;
assign LUT_3[42633] = 32'b00000000000000010111000000100011;
assign LUT_3[42634] = 32'b00000000000000010010011100101010;
assign LUT_3[42635] = 32'b00000000000000011001001000000111;
assign LUT_3[42636] = 32'b00000000000000001101100010111100;
assign LUT_3[42637] = 32'b00000000000000010100001110011001;
assign LUT_3[42638] = 32'b00000000000000001111101010100000;
assign LUT_3[42639] = 32'b00000000000000010110010101111101;
assign LUT_3[42640] = 32'b00000000000000001110001111000011;
assign LUT_3[42641] = 32'b00000000000000010100111010100000;
assign LUT_3[42642] = 32'b00000000000000010000010110100111;
assign LUT_3[42643] = 32'b00000000000000010111000010000100;
assign LUT_3[42644] = 32'b00000000000000001011011100111001;
assign LUT_3[42645] = 32'b00000000000000010010001000010110;
assign LUT_3[42646] = 32'b00000000000000001101100100011101;
assign LUT_3[42647] = 32'b00000000000000010100001111111010;
assign LUT_3[42648] = 32'b00000000000000010011101000001001;
assign LUT_3[42649] = 32'b00000000000000011010010011100110;
assign LUT_3[42650] = 32'b00000000000000010101101111101101;
assign LUT_3[42651] = 32'b00000000000000011100011011001010;
assign LUT_3[42652] = 32'b00000000000000010000110101111111;
assign LUT_3[42653] = 32'b00000000000000010111100001011100;
assign LUT_3[42654] = 32'b00000000000000010010111101100011;
assign LUT_3[42655] = 32'b00000000000000011001101001000000;
assign LUT_3[42656] = 32'b00000000000000001100001010100000;
assign LUT_3[42657] = 32'b00000000000000010010110101111101;
assign LUT_3[42658] = 32'b00000000000000001110010010000100;
assign LUT_3[42659] = 32'b00000000000000010100111101100001;
assign LUT_3[42660] = 32'b00000000000000001001011000010110;
assign LUT_3[42661] = 32'b00000000000000010000000011110011;
assign LUT_3[42662] = 32'b00000000000000001011011111111010;
assign LUT_3[42663] = 32'b00000000000000010010001011010111;
assign LUT_3[42664] = 32'b00000000000000010001100011100110;
assign LUT_3[42665] = 32'b00000000000000011000001111000011;
assign LUT_3[42666] = 32'b00000000000000010011101011001010;
assign LUT_3[42667] = 32'b00000000000000011010010110100111;
assign LUT_3[42668] = 32'b00000000000000001110110001011100;
assign LUT_3[42669] = 32'b00000000000000010101011100111001;
assign LUT_3[42670] = 32'b00000000000000010000111001000000;
assign LUT_3[42671] = 32'b00000000000000010111100100011101;
assign LUT_3[42672] = 32'b00000000000000001111011101100011;
assign LUT_3[42673] = 32'b00000000000000010110001001000000;
assign LUT_3[42674] = 32'b00000000000000010001100101000111;
assign LUT_3[42675] = 32'b00000000000000011000010000100100;
assign LUT_3[42676] = 32'b00000000000000001100101011011001;
assign LUT_3[42677] = 32'b00000000000000010011010110110110;
assign LUT_3[42678] = 32'b00000000000000001110110010111101;
assign LUT_3[42679] = 32'b00000000000000010101011110011010;
assign LUT_3[42680] = 32'b00000000000000010100110110101001;
assign LUT_3[42681] = 32'b00000000000000011011100010000110;
assign LUT_3[42682] = 32'b00000000000000010110111110001101;
assign LUT_3[42683] = 32'b00000000000000011101101001101010;
assign LUT_3[42684] = 32'b00000000000000010010000100011111;
assign LUT_3[42685] = 32'b00000000000000011000101111111100;
assign LUT_3[42686] = 32'b00000000000000010100001100000011;
assign LUT_3[42687] = 32'b00000000000000011010110111100000;
assign LUT_3[42688] = 32'b00000000000000001010110100101011;
assign LUT_3[42689] = 32'b00000000000000010001100000001000;
assign LUT_3[42690] = 32'b00000000000000001100111100001111;
assign LUT_3[42691] = 32'b00000000000000010011100111101100;
assign LUT_3[42692] = 32'b00000000000000001000000010100001;
assign LUT_3[42693] = 32'b00000000000000001110101101111110;
assign LUT_3[42694] = 32'b00000000000000001010001010000101;
assign LUT_3[42695] = 32'b00000000000000010000110101100010;
assign LUT_3[42696] = 32'b00000000000000010000001101110001;
assign LUT_3[42697] = 32'b00000000000000010110111001001110;
assign LUT_3[42698] = 32'b00000000000000010010010101010101;
assign LUT_3[42699] = 32'b00000000000000011001000000110010;
assign LUT_3[42700] = 32'b00000000000000001101011011100111;
assign LUT_3[42701] = 32'b00000000000000010100000111000100;
assign LUT_3[42702] = 32'b00000000000000001111100011001011;
assign LUT_3[42703] = 32'b00000000000000010110001110101000;
assign LUT_3[42704] = 32'b00000000000000001110000111101110;
assign LUT_3[42705] = 32'b00000000000000010100110011001011;
assign LUT_3[42706] = 32'b00000000000000010000001111010010;
assign LUT_3[42707] = 32'b00000000000000010110111010101111;
assign LUT_3[42708] = 32'b00000000000000001011010101100100;
assign LUT_3[42709] = 32'b00000000000000010010000001000001;
assign LUT_3[42710] = 32'b00000000000000001101011101001000;
assign LUT_3[42711] = 32'b00000000000000010100001000100101;
assign LUT_3[42712] = 32'b00000000000000010011100000110100;
assign LUT_3[42713] = 32'b00000000000000011010001100010001;
assign LUT_3[42714] = 32'b00000000000000010101101000011000;
assign LUT_3[42715] = 32'b00000000000000011100010011110101;
assign LUT_3[42716] = 32'b00000000000000010000101110101010;
assign LUT_3[42717] = 32'b00000000000000010111011010000111;
assign LUT_3[42718] = 32'b00000000000000010010110110001110;
assign LUT_3[42719] = 32'b00000000000000011001100001101011;
assign LUT_3[42720] = 32'b00000000000000001100000011001011;
assign LUT_3[42721] = 32'b00000000000000010010101110101000;
assign LUT_3[42722] = 32'b00000000000000001110001010101111;
assign LUT_3[42723] = 32'b00000000000000010100110110001100;
assign LUT_3[42724] = 32'b00000000000000001001010001000001;
assign LUT_3[42725] = 32'b00000000000000001111111100011110;
assign LUT_3[42726] = 32'b00000000000000001011011000100101;
assign LUT_3[42727] = 32'b00000000000000010010000100000010;
assign LUT_3[42728] = 32'b00000000000000010001011100010001;
assign LUT_3[42729] = 32'b00000000000000011000000111101110;
assign LUT_3[42730] = 32'b00000000000000010011100011110101;
assign LUT_3[42731] = 32'b00000000000000011010001111010010;
assign LUT_3[42732] = 32'b00000000000000001110101010000111;
assign LUT_3[42733] = 32'b00000000000000010101010101100100;
assign LUT_3[42734] = 32'b00000000000000010000110001101011;
assign LUT_3[42735] = 32'b00000000000000010111011101001000;
assign LUT_3[42736] = 32'b00000000000000001111010110001110;
assign LUT_3[42737] = 32'b00000000000000010110000001101011;
assign LUT_3[42738] = 32'b00000000000000010001011101110010;
assign LUT_3[42739] = 32'b00000000000000011000001001001111;
assign LUT_3[42740] = 32'b00000000000000001100100100000100;
assign LUT_3[42741] = 32'b00000000000000010011001111100001;
assign LUT_3[42742] = 32'b00000000000000001110101011101000;
assign LUT_3[42743] = 32'b00000000000000010101010111000101;
assign LUT_3[42744] = 32'b00000000000000010100101111010100;
assign LUT_3[42745] = 32'b00000000000000011011011010110001;
assign LUT_3[42746] = 32'b00000000000000010110110110111000;
assign LUT_3[42747] = 32'b00000000000000011101100010010101;
assign LUT_3[42748] = 32'b00000000000000010001111101001010;
assign LUT_3[42749] = 32'b00000000000000011000101000100111;
assign LUT_3[42750] = 32'b00000000000000010100000100101110;
assign LUT_3[42751] = 32'b00000000000000011010110000001011;
assign LUT_3[42752] = 32'b00000000000000000101000000100011;
assign LUT_3[42753] = 32'b00000000000000001011101100000000;
assign LUT_3[42754] = 32'b00000000000000000111001000000111;
assign LUT_3[42755] = 32'b00000000000000001101110011100100;
assign LUT_3[42756] = 32'b00000000000000000010001110011001;
assign LUT_3[42757] = 32'b00000000000000001000111001110110;
assign LUT_3[42758] = 32'b00000000000000000100010101111101;
assign LUT_3[42759] = 32'b00000000000000001011000001011010;
assign LUT_3[42760] = 32'b00000000000000001010011001101001;
assign LUT_3[42761] = 32'b00000000000000010001000101000110;
assign LUT_3[42762] = 32'b00000000000000001100100001001101;
assign LUT_3[42763] = 32'b00000000000000010011001100101010;
assign LUT_3[42764] = 32'b00000000000000000111100111011111;
assign LUT_3[42765] = 32'b00000000000000001110010010111100;
assign LUT_3[42766] = 32'b00000000000000001001101111000011;
assign LUT_3[42767] = 32'b00000000000000010000011010100000;
assign LUT_3[42768] = 32'b00000000000000001000010011100110;
assign LUT_3[42769] = 32'b00000000000000001110111111000011;
assign LUT_3[42770] = 32'b00000000000000001010011011001010;
assign LUT_3[42771] = 32'b00000000000000010001000110100111;
assign LUT_3[42772] = 32'b00000000000000000101100001011100;
assign LUT_3[42773] = 32'b00000000000000001100001100111001;
assign LUT_3[42774] = 32'b00000000000000000111101001000000;
assign LUT_3[42775] = 32'b00000000000000001110010100011101;
assign LUT_3[42776] = 32'b00000000000000001101101100101100;
assign LUT_3[42777] = 32'b00000000000000010100011000001001;
assign LUT_3[42778] = 32'b00000000000000001111110100010000;
assign LUT_3[42779] = 32'b00000000000000010110011111101101;
assign LUT_3[42780] = 32'b00000000000000001010111010100010;
assign LUT_3[42781] = 32'b00000000000000010001100101111111;
assign LUT_3[42782] = 32'b00000000000000001101000010000110;
assign LUT_3[42783] = 32'b00000000000000010011101101100011;
assign LUT_3[42784] = 32'b00000000000000000110001111000011;
assign LUT_3[42785] = 32'b00000000000000001100111010100000;
assign LUT_3[42786] = 32'b00000000000000001000010110100111;
assign LUT_3[42787] = 32'b00000000000000001111000010000100;
assign LUT_3[42788] = 32'b00000000000000000011011100111001;
assign LUT_3[42789] = 32'b00000000000000001010001000010110;
assign LUT_3[42790] = 32'b00000000000000000101100100011101;
assign LUT_3[42791] = 32'b00000000000000001100001111111010;
assign LUT_3[42792] = 32'b00000000000000001011101000001001;
assign LUT_3[42793] = 32'b00000000000000010010010011100110;
assign LUT_3[42794] = 32'b00000000000000001101101111101101;
assign LUT_3[42795] = 32'b00000000000000010100011011001010;
assign LUT_3[42796] = 32'b00000000000000001000110101111111;
assign LUT_3[42797] = 32'b00000000000000001111100001011100;
assign LUT_3[42798] = 32'b00000000000000001010111101100011;
assign LUT_3[42799] = 32'b00000000000000010001101001000000;
assign LUT_3[42800] = 32'b00000000000000001001100010000110;
assign LUT_3[42801] = 32'b00000000000000010000001101100011;
assign LUT_3[42802] = 32'b00000000000000001011101001101010;
assign LUT_3[42803] = 32'b00000000000000010010010101000111;
assign LUT_3[42804] = 32'b00000000000000000110101111111100;
assign LUT_3[42805] = 32'b00000000000000001101011011011001;
assign LUT_3[42806] = 32'b00000000000000001000110111100000;
assign LUT_3[42807] = 32'b00000000000000001111100010111101;
assign LUT_3[42808] = 32'b00000000000000001110111011001100;
assign LUT_3[42809] = 32'b00000000000000010101100110101001;
assign LUT_3[42810] = 32'b00000000000000010001000010110000;
assign LUT_3[42811] = 32'b00000000000000010111101110001101;
assign LUT_3[42812] = 32'b00000000000000001100001001000010;
assign LUT_3[42813] = 32'b00000000000000010010110100011111;
assign LUT_3[42814] = 32'b00000000000000001110010000100110;
assign LUT_3[42815] = 32'b00000000000000010100111100000011;
assign LUT_3[42816] = 32'b00000000000000000100111001001110;
assign LUT_3[42817] = 32'b00000000000000001011100100101011;
assign LUT_3[42818] = 32'b00000000000000000111000000110010;
assign LUT_3[42819] = 32'b00000000000000001101101100001111;
assign LUT_3[42820] = 32'b00000000000000000010000111000100;
assign LUT_3[42821] = 32'b00000000000000001000110010100001;
assign LUT_3[42822] = 32'b00000000000000000100001110101000;
assign LUT_3[42823] = 32'b00000000000000001010111010000101;
assign LUT_3[42824] = 32'b00000000000000001010010010010100;
assign LUT_3[42825] = 32'b00000000000000010000111101110001;
assign LUT_3[42826] = 32'b00000000000000001100011001111000;
assign LUT_3[42827] = 32'b00000000000000010011000101010101;
assign LUT_3[42828] = 32'b00000000000000000111100000001010;
assign LUT_3[42829] = 32'b00000000000000001110001011100111;
assign LUT_3[42830] = 32'b00000000000000001001100111101110;
assign LUT_3[42831] = 32'b00000000000000010000010011001011;
assign LUT_3[42832] = 32'b00000000000000001000001100010001;
assign LUT_3[42833] = 32'b00000000000000001110110111101110;
assign LUT_3[42834] = 32'b00000000000000001010010011110101;
assign LUT_3[42835] = 32'b00000000000000010000111111010010;
assign LUT_3[42836] = 32'b00000000000000000101011010000111;
assign LUT_3[42837] = 32'b00000000000000001100000101100100;
assign LUT_3[42838] = 32'b00000000000000000111100001101011;
assign LUT_3[42839] = 32'b00000000000000001110001101001000;
assign LUT_3[42840] = 32'b00000000000000001101100101010111;
assign LUT_3[42841] = 32'b00000000000000010100010000110100;
assign LUT_3[42842] = 32'b00000000000000001111101100111011;
assign LUT_3[42843] = 32'b00000000000000010110011000011000;
assign LUT_3[42844] = 32'b00000000000000001010110011001101;
assign LUT_3[42845] = 32'b00000000000000010001011110101010;
assign LUT_3[42846] = 32'b00000000000000001100111010110001;
assign LUT_3[42847] = 32'b00000000000000010011100110001110;
assign LUT_3[42848] = 32'b00000000000000000110000111101110;
assign LUT_3[42849] = 32'b00000000000000001100110011001011;
assign LUT_3[42850] = 32'b00000000000000001000001111010010;
assign LUT_3[42851] = 32'b00000000000000001110111010101111;
assign LUT_3[42852] = 32'b00000000000000000011010101100100;
assign LUT_3[42853] = 32'b00000000000000001010000001000001;
assign LUT_3[42854] = 32'b00000000000000000101011101001000;
assign LUT_3[42855] = 32'b00000000000000001100001000100101;
assign LUT_3[42856] = 32'b00000000000000001011100000110100;
assign LUT_3[42857] = 32'b00000000000000010010001100010001;
assign LUT_3[42858] = 32'b00000000000000001101101000011000;
assign LUT_3[42859] = 32'b00000000000000010100010011110101;
assign LUT_3[42860] = 32'b00000000000000001000101110101010;
assign LUT_3[42861] = 32'b00000000000000001111011010000111;
assign LUT_3[42862] = 32'b00000000000000001010110110001110;
assign LUT_3[42863] = 32'b00000000000000010001100001101011;
assign LUT_3[42864] = 32'b00000000000000001001011010110001;
assign LUT_3[42865] = 32'b00000000000000010000000110001110;
assign LUT_3[42866] = 32'b00000000000000001011100010010101;
assign LUT_3[42867] = 32'b00000000000000010010001101110010;
assign LUT_3[42868] = 32'b00000000000000000110101000100111;
assign LUT_3[42869] = 32'b00000000000000001101010100000100;
assign LUT_3[42870] = 32'b00000000000000001000110000001011;
assign LUT_3[42871] = 32'b00000000000000001111011011101000;
assign LUT_3[42872] = 32'b00000000000000001110110011110111;
assign LUT_3[42873] = 32'b00000000000000010101011111010100;
assign LUT_3[42874] = 32'b00000000000000010000111011011011;
assign LUT_3[42875] = 32'b00000000000000010111100110111000;
assign LUT_3[42876] = 32'b00000000000000001100000001101101;
assign LUT_3[42877] = 32'b00000000000000010010101101001010;
assign LUT_3[42878] = 32'b00000000000000001110001001010001;
assign LUT_3[42879] = 32'b00000000000000010100110100101110;
assign LUT_3[42880] = 32'b00000000000000000111001011100001;
assign LUT_3[42881] = 32'b00000000000000001101110110111110;
assign LUT_3[42882] = 32'b00000000000000001001010011000101;
assign LUT_3[42883] = 32'b00000000000000001111111110100010;
assign LUT_3[42884] = 32'b00000000000000000100011001010111;
assign LUT_3[42885] = 32'b00000000000000001011000100110100;
assign LUT_3[42886] = 32'b00000000000000000110100000111011;
assign LUT_3[42887] = 32'b00000000000000001101001100011000;
assign LUT_3[42888] = 32'b00000000000000001100100100100111;
assign LUT_3[42889] = 32'b00000000000000010011010000000100;
assign LUT_3[42890] = 32'b00000000000000001110101100001011;
assign LUT_3[42891] = 32'b00000000000000010101010111101000;
assign LUT_3[42892] = 32'b00000000000000001001110010011101;
assign LUT_3[42893] = 32'b00000000000000010000011101111010;
assign LUT_3[42894] = 32'b00000000000000001011111010000001;
assign LUT_3[42895] = 32'b00000000000000010010100101011110;
assign LUT_3[42896] = 32'b00000000000000001010011110100100;
assign LUT_3[42897] = 32'b00000000000000010001001010000001;
assign LUT_3[42898] = 32'b00000000000000001100100110001000;
assign LUT_3[42899] = 32'b00000000000000010011010001100101;
assign LUT_3[42900] = 32'b00000000000000000111101100011010;
assign LUT_3[42901] = 32'b00000000000000001110010111110111;
assign LUT_3[42902] = 32'b00000000000000001001110011111110;
assign LUT_3[42903] = 32'b00000000000000010000011111011011;
assign LUT_3[42904] = 32'b00000000000000001111110111101010;
assign LUT_3[42905] = 32'b00000000000000010110100011000111;
assign LUT_3[42906] = 32'b00000000000000010001111111001110;
assign LUT_3[42907] = 32'b00000000000000011000101010101011;
assign LUT_3[42908] = 32'b00000000000000001101000101100000;
assign LUT_3[42909] = 32'b00000000000000010011110000111101;
assign LUT_3[42910] = 32'b00000000000000001111001101000100;
assign LUT_3[42911] = 32'b00000000000000010101111000100001;
assign LUT_3[42912] = 32'b00000000000000001000011010000001;
assign LUT_3[42913] = 32'b00000000000000001111000101011110;
assign LUT_3[42914] = 32'b00000000000000001010100001100101;
assign LUT_3[42915] = 32'b00000000000000010001001101000010;
assign LUT_3[42916] = 32'b00000000000000000101100111110111;
assign LUT_3[42917] = 32'b00000000000000001100010011010100;
assign LUT_3[42918] = 32'b00000000000000000111101111011011;
assign LUT_3[42919] = 32'b00000000000000001110011010111000;
assign LUT_3[42920] = 32'b00000000000000001101110011000111;
assign LUT_3[42921] = 32'b00000000000000010100011110100100;
assign LUT_3[42922] = 32'b00000000000000001111111010101011;
assign LUT_3[42923] = 32'b00000000000000010110100110001000;
assign LUT_3[42924] = 32'b00000000000000001011000000111101;
assign LUT_3[42925] = 32'b00000000000000010001101100011010;
assign LUT_3[42926] = 32'b00000000000000001101001000100001;
assign LUT_3[42927] = 32'b00000000000000010011110011111110;
assign LUT_3[42928] = 32'b00000000000000001011101101000100;
assign LUT_3[42929] = 32'b00000000000000010010011000100001;
assign LUT_3[42930] = 32'b00000000000000001101110100101000;
assign LUT_3[42931] = 32'b00000000000000010100100000000101;
assign LUT_3[42932] = 32'b00000000000000001000111010111010;
assign LUT_3[42933] = 32'b00000000000000001111100110010111;
assign LUT_3[42934] = 32'b00000000000000001011000010011110;
assign LUT_3[42935] = 32'b00000000000000010001101101111011;
assign LUT_3[42936] = 32'b00000000000000010001000110001010;
assign LUT_3[42937] = 32'b00000000000000010111110001100111;
assign LUT_3[42938] = 32'b00000000000000010011001101101110;
assign LUT_3[42939] = 32'b00000000000000011001111001001011;
assign LUT_3[42940] = 32'b00000000000000001110010100000000;
assign LUT_3[42941] = 32'b00000000000000010100111111011101;
assign LUT_3[42942] = 32'b00000000000000010000011011100100;
assign LUT_3[42943] = 32'b00000000000000010111000111000001;
assign LUT_3[42944] = 32'b00000000000000000111000100001100;
assign LUT_3[42945] = 32'b00000000000000001101101111101001;
assign LUT_3[42946] = 32'b00000000000000001001001011110000;
assign LUT_3[42947] = 32'b00000000000000001111110111001101;
assign LUT_3[42948] = 32'b00000000000000000100010010000010;
assign LUT_3[42949] = 32'b00000000000000001010111101011111;
assign LUT_3[42950] = 32'b00000000000000000110011001100110;
assign LUT_3[42951] = 32'b00000000000000001101000101000011;
assign LUT_3[42952] = 32'b00000000000000001100011101010010;
assign LUT_3[42953] = 32'b00000000000000010011001000101111;
assign LUT_3[42954] = 32'b00000000000000001110100100110110;
assign LUT_3[42955] = 32'b00000000000000010101010000010011;
assign LUT_3[42956] = 32'b00000000000000001001101011001000;
assign LUT_3[42957] = 32'b00000000000000010000010110100101;
assign LUT_3[42958] = 32'b00000000000000001011110010101100;
assign LUT_3[42959] = 32'b00000000000000010010011110001001;
assign LUT_3[42960] = 32'b00000000000000001010010111001111;
assign LUT_3[42961] = 32'b00000000000000010001000010101100;
assign LUT_3[42962] = 32'b00000000000000001100011110110011;
assign LUT_3[42963] = 32'b00000000000000010011001010010000;
assign LUT_3[42964] = 32'b00000000000000000111100101000101;
assign LUT_3[42965] = 32'b00000000000000001110010000100010;
assign LUT_3[42966] = 32'b00000000000000001001101100101001;
assign LUT_3[42967] = 32'b00000000000000010000011000000110;
assign LUT_3[42968] = 32'b00000000000000001111110000010101;
assign LUT_3[42969] = 32'b00000000000000010110011011110010;
assign LUT_3[42970] = 32'b00000000000000010001110111111001;
assign LUT_3[42971] = 32'b00000000000000011000100011010110;
assign LUT_3[42972] = 32'b00000000000000001100111110001011;
assign LUT_3[42973] = 32'b00000000000000010011101001101000;
assign LUT_3[42974] = 32'b00000000000000001111000101101111;
assign LUT_3[42975] = 32'b00000000000000010101110001001100;
assign LUT_3[42976] = 32'b00000000000000001000010010101100;
assign LUT_3[42977] = 32'b00000000000000001110111110001001;
assign LUT_3[42978] = 32'b00000000000000001010011010010000;
assign LUT_3[42979] = 32'b00000000000000010001000101101101;
assign LUT_3[42980] = 32'b00000000000000000101100000100010;
assign LUT_3[42981] = 32'b00000000000000001100001011111111;
assign LUT_3[42982] = 32'b00000000000000000111101000000110;
assign LUT_3[42983] = 32'b00000000000000001110010011100011;
assign LUT_3[42984] = 32'b00000000000000001101101011110010;
assign LUT_3[42985] = 32'b00000000000000010100010111001111;
assign LUT_3[42986] = 32'b00000000000000001111110011010110;
assign LUT_3[42987] = 32'b00000000000000010110011110110011;
assign LUT_3[42988] = 32'b00000000000000001010111001101000;
assign LUT_3[42989] = 32'b00000000000000010001100101000101;
assign LUT_3[42990] = 32'b00000000000000001101000001001100;
assign LUT_3[42991] = 32'b00000000000000010011101100101001;
assign LUT_3[42992] = 32'b00000000000000001011100101101111;
assign LUT_3[42993] = 32'b00000000000000010010010001001100;
assign LUT_3[42994] = 32'b00000000000000001101101101010011;
assign LUT_3[42995] = 32'b00000000000000010100011000110000;
assign LUT_3[42996] = 32'b00000000000000001000110011100101;
assign LUT_3[42997] = 32'b00000000000000001111011111000010;
assign LUT_3[42998] = 32'b00000000000000001010111011001001;
assign LUT_3[42999] = 32'b00000000000000010001100110100110;
assign LUT_3[43000] = 32'b00000000000000010000111110110101;
assign LUT_3[43001] = 32'b00000000000000010111101010010010;
assign LUT_3[43002] = 32'b00000000000000010011000110011001;
assign LUT_3[43003] = 32'b00000000000000011001110001110110;
assign LUT_3[43004] = 32'b00000000000000001110001100101011;
assign LUT_3[43005] = 32'b00000000000000010100111000001000;
assign LUT_3[43006] = 32'b00000000000000010000010100001111;
assign LUT_3[43007] = 32'b00000000000000010110111111101100;
assign LUT_3[43008] = 32'b00000000000000000000101101000111;
assign LUT_3[43009] = 32'b00000000000000000111011000100100;
assign LUT_3[43010] = 32'b00000000000000000010110100101011;
assign LUT_3[43011] = 32'b00000000000000001001100000001000;
assign LUT_3[43012] = 32'b11111111111111111101111010111101;
assign LUT_3[43013] = 32'b00000000000000000100100110011010;
assign LUT_3[43014] = 32'b00000000000000000000000010100001;
assign LUT_3[43015] = 32'b00000000000000000110101101111110;
assign LUT_3[43016] = 32'b00000000000000000110000110001101;
assign LUT_3[43017] = 32'b00000000000000001100110001101010;
assign LUT_3[43018] = 32'b00000000000000001000001101110001;
assign LUT_3[43019] = 32'b00000000000000001110111001001110;
assign LUT_3[43020] = 32'b00000000000000000011010100000011;
assign LUT_3[43021] = 32'b00000000000000001001111111100000;
assign LUT_3[43022] = 32'b00000000000000000101011011100111;
assign LUT_3[43023] = 32'b00000000000000001100000111000100;
assign LUT_3[43024] = 32'b00000000000000000100000000001010;
assign LUT_3[43025] = 32'b00000000000000001010101011100111;
assign LUT_3[43026] = 32'b00000000000000000110000111101110;
assign LUT_3[43027] = 32'b00000000000000001100110011001011;
assign LUT_3[43028] = 32'b00000000000000000001001110000000;
assign LUT_3[43029] = 32'b00000000000000000111111001011101;
assign LUT_3[43030] = 32'b00000000000000000011010101100100;
assign LUT_3[43031] = 32'b00000000000000001010000001000001;
assign LUT_3[43032] = 32'b00000000000000001001011001010000;
assign LUT_3[43033] = 32'b00000000000000010000000100101101;
assign LUT_3[43034] = 32'b00000000000000001011100000110100;
assign LUT_3[43035] = 32'b00000000000000010010001100010001;
assign LUT_3[43036] = 32'b00000000000000000110100111000110;
assign LUT_3[43037] = 32'b00000000000000001101010010100011;
assign LUT_3[43038] = 32'b00000000000000001000101110101010;
assign LUT_3[43039] = 32'b00000000000000001111011010000111;
assign LUT_3[43040] = 32'b00000000000000000001111011100111;
assign LUT_3[43041] = 32'b00000000000000001000100111000100;
assign LUT_3[43042] = 32'b00000000000000000100000011001011;
assign LUT_3[43043] = 32'b00000000000000001010101110101000;
assign LUT_3[43044] = 32'b11111111111111111111001001011101;
assign LUT_3[43045] = 32'b00000000000000000101110100111010;
assign LUT_3[43046] = 32'b00000000000000000001010001000001;
assign LUT_3[43047] = 32'b00000000000000000111111100011110;
assign LUT_3[43048] = 32'b00000000000000000111010100101101;
assign LUT_3[43049] = 32'b00000000000000001110000000001010;
assign LUT_3[43050] = 32'b00000000000000001001011100010001;
assign LUT_3[43051] = 32'b00000000000000010000000111101110;
assign LUT_3[43052] = 32'b00000000000000000100100010100011;
assign LUT_3[43053] = 32'b00000000000000001011001110000000;
assign LUT_3[43054] = 32'b00000000000000000110101010000111;
assign LUT_3[43055] = 32'b00000000000000001101010101100100;
assign LUT_3[43056] = 32'b00000000000000000101001110101010;
assign LUT_3[43057] = 32'b00000000000000001011111010000111;
assign LUT_3[43058] = 32'b00000000000000000111010110001110;
assign LUT_3[43059] = 32'b00000000000000001110000001101011;
assign LUT_3[43060] = 32'b00000000000000000010011100100000;
assign LUT_3[43061] = 32'b00000000000000001001000111111101;
assign LUT_3[43062] = 32'b00000000000000000100100100000100;
assign LUT_3[43063] = 32'b00000000000000001011001111100001;
assign LUT_3[43064] = 32'b00000000000000001010100111110000;
assign LUT_3[43065] = 32'b00000000000000010001010011001101;
assign LUT_3[43066] = 32'b00000000000000001100101111010100;
assign LUT_3[43067] = 32'b00000000000000010011011010110001;
assign LUT_3[43068] = 32'b00000000000000000111110101100110;
assign LUT_3[43069] = 32'b00000000000000001110100001000011;
assign LUT_3[43070] = 32'b00000000000000001001111101001010;
assign LUT_3[43071] = 32'b00000000000000010000101000100111;
assign LUT_3[43072] = 32'b00000000000000000000100101110010;
assign LUT_3[43073] = 32'b00000000000000000111010001001111;
assign LUT_3[43074] = 32'b00000000000000000010101101010110;
assign LUT_3[43075] = 32'b00000000000000001001011000110011;
assign LUT_3[43076] = 32'b11111111111111111101110011101000;
assign LUT_3[43077] = 32'b00000000000000000100011111000101;
assign LUT_3[43078] = 32'b11111111111111111111111011001100;
assign LUT_3[43079] = 32'b00000000000000000110100110101001;
assign LUT_3[43080] = 32'b00000000000000000101111110111000;
assign LUT_3[43081] = 32'b00000000000000001100101010010101;
assign LUT_3[43082] = 32'b00000000000000001000000110011100;
assign LUT_3[43083] = 32'b00000000000000001110110001111001;
assign LUT_3[43084] = 32'b00000000000000000011001100101110;
assign LUT_3[43085] = 32'b00000000000000001001111000001011;
assign LUT_3[43086] = 32'b00000000000000000101010100010010;
assign LUT_3[43087] = 32'b00000000000000001011111111101111;
assign LUT_3[43088] = 32'b00000000000000000011111000110101;
assign LUT_3[43089] = 32'b00000000000000001010100100010010;
assign LUT_3[43090] = 32'b00000000000000000110000000011001;
assign LUT_3[43091] = 32'b00000000000000001100101011110110;
assign LUT_3[43092] = 32'b00000000000000000001000110101011;
assign LUT_3[43093] = 32'b00000000000000000111110010001000;
assign LUT_3[43094] = 32'b00000000000000000011001110001111;
assign LUT_3[43095] = 32'b00000000000000001001111001101100;
assign LUT_3[43096] = 32'b00000000000000001001010001111011;
assign LUT_3[43097] = 32'b00000000000000001111111101011000;
assign LUT_3[43098] = 32'b00000000000000001011011001011111;
assign LUT_3[43099] = 32'b00000000000000010010000100111100;
assign LUT_3[43100] = 32'b00000000000000000110011111110001;
assign LUT_3[43101] = 32'b00000000000000001101001011001110;
assign LUT_3[43102] = 32'b00000000000000001000100111010101;
assign LUT_3[43103] = 32'b00000000000000001111010010110010;
assign LUT_3[43104] = 32'b00000000000000000001110100010010;
assign LUT_3[43105] = 32'b00000000000000001000011111101111;
assign LUT_3[43106] = 32'b00000000000000000011111011110110;
assign LUT_3[43107] = 32'b00000000000000001010100111010011;
assign LUT_3[43108] = 32'b11111111111111111111000010001000;
assign LUT_3[43109] = 32'b00000000000000000101101101100101;
assign LUT_3[43110] = 32'b00000000000000000001001001101100;
assign LUT_3[43111] = 32'b00000000000000000111110101001001;
assign LUT_3[43112] = 32'b00000000000000000111001101011000;
assign LUT_3[43113] = 32'b00000000000000001101111000110101;
assign LUT_3[43114] = 32'b00000000000000001001010100111100;
assign LUT_3[43115] = 32'b00000000000000010000000000011001;
assign LUT_3[43116] = 32'b00000000000000000100011011001110;
assign LUT_3[43117] = 32'b00000000000000001011000110101011;
assign LUT_3[43118] = 32'b00000000000000000110100010110010;
assign LUT_3[43119] = 32'b00000000000000001101001110001111;
assign LUT_3[43120] = 32'b00000000000000000101000111010101;
assign LUT_3[43121] = 32'b00000000000000001011110010110010;
assign LUT_3[43122] = 32'b00000000000000000111001110111001;
assign LUT_3[43123] = 32'b00000000000000001101111010010110;
assign LUT_3[43124] = 32'b00000000000000000010010101001011;
assign LUT_3[43125] = 32'b00000000000000001001000000101000;
assign LUT_3[43126] = 32'b00000000000000000100011100101111;
assign LUT_3[43127] = 32'b00000000000000001011001000001100;
assign LUT_3[43128] = 32'b00000000000000001010100000011011;
assign LUT_3[43129] = 32'b00000000000000010001001011111000;
assign LUT_3[43130] = 32'b00000000000000001100100111111111;
assign LUT_3[43131] = 32'b00000000000000010011010011011100;
assign LUT_3[43132] = 32'b00000000000000000111101110010001;
assign LUT_3[43133] = 32'b00000000000000001110011001101110;
assign LUT_3[43134] = 32'b00000000000000001001110101110101;
assign LUT_3[43135] = 32'b00000000000000010000100001010010;
assign LUT_3[43136] = 32'b00000000000000000010111000000101;
assign LUT_3[43137] = 32'b00000000000000001001100011100010;
assign LUT_3[43138] = 32'b00000000000000000100111111101001;
assign LUT_3[43139] = 32'b00000000000000001011101011000110;
assign LUT_3[43140] = 32'b00000000000000000000000101111011;
assign LUT_3[43141] = 32'b00000000000000000110110001011000;
assign LUT_3[43142] = 32'b00000000000000000010001101011111;
assign LUT_3[43143] = 32'b00000000000000001000111000111100;
assign LUT_3[43144] = 32'b00000000000000001000010001001011;
assign LUT_3[43145] = 32'b00000000000000001110111100101000;
assign LUT_3[43146] = 32'b00000000000000001010011000101111;
assign LUT_3[43147] = 32'b00000000000000010001000100001100;
assign LUT_3[43148] = 32'b00000000000000000101011111000001;
assign LUT_3[43149] = 32'b00000000000000001100001010011110;
assign LUT_3[43150] = 32'b00000000000000000111100110100101;
assign LUT_3[43151] = 32'b00000000000000001110010010000010;
assign LUT_3[43152] = 32'b00000000000000000110001011001000;
assign LUT_3[43153] = 32'b00000000000000001100110110100101;
assign LUT_3[43154] = 32'b00000000000000001000010010101100;
assign LUT_3[43155] = 32'b00000000000000001110111110001001;
assign LUT_3[43156] = 32'b00000000000000000011011000111110;
assign LUT_3[43157] = 32'b00000000000000001010000100011011;
assign LUT_3[43158] = 32'b00000000000000000101100000100010;
assign LUT_3[43159] = 32'b00000000000000001100001011111111;
assign LUT_3[43160] = 32'b00000000000000001011100100001110;
assign LUT_3[43161] = 32'b00000000000000010010001111101011;
assign LUT_3[43162] = 32'b00000000000000001101101011110010;
assign LUT_3[43163] = 32'b00000000000000010100010111001111;
assign LUT_3[43164] = 32'b00000000000000001000110010000100;
assign LUT_3[43165] = 32'b00000000000000001111011101100001;
assign LUT_3[43166] = 32'b00000000000000001010111001101000;
assign LUT_3[43167] = 32'b00000000000000010001100101000101;
assign LUT_3[43168] = 32'b00000000000000000100000110100101;
assign LUT_3[43169] = 32'b00000000000000001010110010000010;
assign LUT_3[43170] = 32'b00000000000000000110001110001001;
assign LUT_3[43171] = 32'b00000000000000001100111001100110;
assign LUT_3[43172] = 32'b00000000000000000001010100011011;
assign LUT_3[43173] = 32'b00000000000000000111111111111000;
assign LUT_3[43174] = 32'b00000000000000000011011011111111;
assign LUT_3[43175] = 32'b00000000000000001010000111011100;
assign LUT_3[43176] = 32'b00000000000000001001011111101011;
assign LUT_3[43177] = 32'b00000000000000010000001011001000;
assign LUT_3[43178] = 32'b00000000000000001011100111001111;
assign LUT_3[43179] = 32'b00000000000000010010010010101100;
assign LUT_3[43180] = 32'b00000000000000000110101101100001;
assign LUT_3[43181] = 32'b00000000000000001101011000111110;
assign LUT_3[43182] = 32'b00000000000000001000110101000101;
assign LUT_3[43183] = 32'b00000000000000001111100000100010;
assign LUT_3[43184] = 32'b00000000000000000111011001101000;
assign LUT_3[43185] = 32'b00000000000000001110000101000101;
assign LUT_3[43186] = 32'b00000000000000001001100001001100;
assign LUT_3[43187] = 32'b00000000000000010000001100101001;
assign LUT_3[43188] = 32'b00000000000000000100100111011110;
assign LUT_3[43189] = 32'b00000000000000001011010010111011;
assign LUT_3[43190] = 32'b00000000000000000110101111000010;
assign LUT_3[43191] = 32'b00000000000000001101011010011111;
assign LUT_3[43192] = 32'b00000000000000001100110010101110;
assign LUT_3[43193] = 32'b00000000000000010011011110001011;
assign LUT_3[43194] = 32'b00000000000000001110111010010010;
assign LUT_3[43195] = 32'b00000000000000010101100101101111;
assign LUT_3[43196] = 32'b00000000000000001010000000100100;
assign LUT_3[43197] = 32'b00000000000000010000101100000001;
assign LUT_3[43198] = 32'b00000000000000001100001000001000;
assign LUT_3[43199] = 32'b00000000000000010010110011100101;
assign LUT_3[43200] = 32'b00000000000000000010110000110000;
assign LUT_3[43201] = 32'b00000000000000001001011100001101;
assign LUT_3[43202] = 32'b00000000000000000100111000010100;
assign LUT_3[43203] = 32'b00000000000000001011100011110001;
assign LUT_3[43204] = 32'b11111111111111111111111110100110;
assign LUT_3[43205] = 32'b00000000000000000110101010000011;
assign LUT_3[43206] = 32'b00000000000000000010000110001010;
assign LUT_3[43207] = 32'b00000000000000001000110001100111;
assign LUT_3[43208] = 32'b00000000000000001000001001110110;
assign LUT_3[43209] = 32'b00000000000000001110110101010011;
assign LUT_3[43210] = 32'b00000000000000001010010001011010;
assign LUT_3[43211] = 32'b00000000000000010000111100110111;
assign LUT_3[43212] = 32'b00000000000000000101010111101100;
assign LUT_3[43213] = 32'b00000000000000001100000011001001;
assign LUT_3[43214] = 32'b00000000000000000111011111010000;
assign LUT_3[43215] = 32'b00000000000000001110001010101101;
assign LUT_3[43216] = 32'b00000000000000000110000011110011;
assign LUT_3[43217] = 32'b00000000000000001100101111010000;
assign LUT_3[43218] = 32'b00000000000000001000001011010111;
assign LUT_3[43219] = 32'b00000000000000001110110110110100;
assign LUT_3[43220] = 32'b00000000000000000011010001101001;
assign LUT_3[43221] = 32'b00000000000000001001111101000110;
assign LUT_3[43222] = 32'b00000000000000000101011001001101;
assign LUT_3[43223] = 32'b00000000000000001100000100101010;
assign LUT_3[43224] = 32'b00000000000000001011011100111001;
assign LUT_3[43225] = 32'b00000000000000010010001000010110;
assign LUT_3[43226] = 32'b00000000000000001101100100011101;
assign LUT_3[43227] = 32'b00000000000000010100001111111010;
assign LUT_3[43228] = 32'b00000000000000001000101010101111;
assign LUT_3[43229] = 32'b00000000000000001111010110001100;
assign LUT_3[43230] = 32'b00000000000000001010110010010011;
assign LUT_3[43231] = 32'b00000000000000010001011101110000;
assign LUT_3[43232] = 32'b00000000000000000011111111010000;
assign LUT_3[43233] = 32'b00000000000000001010101010101101;
assign LUT_3[43234] = 32'b00000000000000000110000110110100;
assign LUT_3[43235] = 32'b00000000000000001100110010010001;
assign LUT_3[43236] = 32'b00000000000000000001001101000110;
assign LUT_3[43237] = 32'b00000000000000000111111000100011;
assign LUT_3[43238] = 32'b00000000000000000011010100101010;
assign LUT_3[43239] = 32'b00000000000000001010000000000111;
assign LUT_3[43240] = 32'b00000000000000001001011000010110;
assign LUT_3[43241] = 32'b00000000000000010000000011110011;
assign LUT_3[43242] = 32'b00000000000000001011011111111010;
assign LUT_3[43243] = 32'b00000000000000010010001011010111;
assign LUT_3[43244] = 32'b00000000000000000110100110001100;
assign LUT_3[43245] = 32'b00000000000000001101010001101001;
assign LUT_3[43246] = 32'b00000000000000001000101101110000;
assign LUT_3[43247] = 32'b00000000000000001111011001001101;
assign LUT_3[43248] = 32'b00000000000000000111010010010011;
assign LUT_3[43249] = 32'b00000000000000001101111101110000;
assign LUT_3[43250] = 32'b00000000000000001001011001110111;
assign LUT_3[43251] = 32'b00000000000000010000000101010100;
assign LUT_3[43252] = 32'b00000000000000000100100000001001;
assign LUT_3[43253] = 32'b00000000000000001011001011100110;
assign LUT_3[43254] = 32'b00000000000000000110100111101101;
assign LUT_3[43255] = 32'b00000000000000001101010011001010;
assign LUT_3[43256] = 32'b00000000000000001100101011011001;
assign LUT_3[43257] = 32'b00000000000000010011010110110110;
assign LUT_3[43258] = 32'b00000000000000001110110010111101;
assign LUT_3[43259] = 32'b00000000000000010101011110011010;
assign LUT_3[43260] = 32'b00000000000000001001111001001111;
assign LUT_3[43261] = 32'b00000000000000010000100100101100;
assign LUT_3[43262] = 32'b00000000000000001100000000110011;
assign LUT_3[43263] = 32'b00000000000000010010101100010000;
assign LUT_3[43264] = 32'b11111111111111111100111100101000;
assign LUT_3[43265] = 32'b00000000000000000011101000000101;
assign LUT_3[43266] = 32'b11111111111111111111000100001100;
assign LUT_3[43267] = 32'b00000000000000000101101111101001;
assign LUT_3[43268] = 32'b11111111111111111010001010011110;
assign LUT_3[43269] = 32'b00000000000000000000110101111011;
assign LUT_3[43270] = 32'b11111111111111111100010010000010;
assign LUT_3[43271] = 32'b00000000000000000010111101011111;
assign LUT_3[43272] = 32'b00000000000000000010010101101110;
assign LUT_3[43273] = 32'b00000000000000001001000001001011;
assign LUT_3[43274] = 32'b00000000000000000100011101010010;
assign LUT_3[43275] = 32'b00000000000000001011001000101111;
assign LUT_3[43276] = 32'b11111111111111111111100011100100;
assign LUT_3[43277] = 32'b00000000000000000110001111000001;
assign LUT_3[43278] = 32'b00000000000000000001101011001000;
assign LUT_3[43279] = 32'b00000000000000001000010110100101;
assign LUT_3[43280] = 32'b00000000000000000000001111101011;
assign LUT_3[43281] = 32'b00000000000000000110111011001000;
assign LUT_3[43282] = 32'b00000000000000000010010111001111;
assign LUT_3[43283] = 32'b00000000000000001001000010101100;
assign LUT_3[43284] = 32'b11111111111111111101011101100001;
assign LUT_3[43285] = 32'b00000000000000000100001000111110;
assign LUT_3[43286] = 32'b11111111111111111111100101000101;
assign LUT_3[43287] = 32'b00000000000000000110010000100010;
assign LUT_3[43288] = 32'b00000000000000000101101000110001;
assign LUT_3[43289] = 32'b00000000000000001100010100001110;
assign LUT_3[43290] = 32'b00000000000000000111110000010101;
assign LUT_3[43291] = 32'b00000000000000001110011011110010;
assign LUT_3[43292] = 32'b00000000000000000010110110100111;
assign LUT_3[43293] = 32'b00000000000000001001100010000100;
assign LUT_3[43294] = 32'b00000000000000000100111110001011;
assign LUT_3[43295] = 32'b00000000000000001011101001101000;
assign LUT_3[43296] = 32'b11111111111111111110001011001000;
assign LUT_3[43297] = 32'b00000000000000000100110110100101;
assign LUT_3[43298] = 32'b00000000000000000000010010101100;
assign LUT_3[43299] = 32'b00000000000000000110111110001001;
assign LUT_3[43300] = 32'b11111111111111111011011000111110;
assign LUT_3[43301] = 32'b00000000000000000010000100011011;
assign LUT_3[43302] = 32'b11111111111111111101100000100010;
assign LUT_3[43303] = 32'b00000000000000000100001011111111;
assign LUT_3[43304] = 32'b00000000000000000011100100001110;
assign LUT_3[43305] = 32'b00000000000000001010001111101011;
assign LUT_3[43306] = 32'b00000000000000000101101011110010;
assign LUT_3[43307] = 32'b00000000000000001100010111001111;
assign LUT_3[43308] = 32'b00000000000000000000110010000100;
assign LUT_3[43309] = 32'b00000000000000000111011101100001;
assign LUT_3[43310] = 32'b00000000000000000010111001101000;
assign LUT_3[43311] = 32'b00000000000000001001100101000101;
assign LUT_3[43312] = 32'b00000000000000000001011110001011;
assign LUT_3[43313] = 32'b00000000000000001000001001101000;
assign LUT_3[43314] = 32'b00000000000000000011100101101111;
assign LUT_3[43315] = 32'b00000000000000001010010001001100;
assign LUT_3[43316] = 32'b11111111111111111110101100000001;
assign LUT_3[43317] = 32'b00000000000000000101010111011110;
assign LUT_3[43318] = 32'b00000000000000000000110011100101;
assign LUT_3[43319] = 32'b00000000000000000111011111000010;
assign LUT_3[43320] = 32'b00000000000000000110110111010001;
assign LUT_3[43321] = 32'b00000000000000001101100010101110;
assign LUT_3[43322] = 32'b00000000000000001000111110110101;
assign LUT_3[43323] = 32'b00000000000000001111101010010010;
assign LUT_3[43324] = 32'b00000000000000000100000101000111;
assign LUT_3[43325] = 32'b00000000000000001010110000100100;
assign LUT_3[43326] = 32'b00000000000000000110001100101011;
assign LUT_3[43327] = 32'b00000000000000001100111000001000;
assign LUT_3[43328] = 32'b11111111111111111100110101010011;
assign LUT_3[43329] = 32'b00000000000000000011100000110000;
assign LUT_3[43330] = 32'b11111111111111111110111100110111;
assign LUT_3[43331] = 32'b00000000000000000101101000010100;
assign LUT_3[43332] = 32'b11111111111111111010000011001001;
assign LUT_3[43333] = 32'b00000000000000000000101110100110;
assign LUT_3[43334] = 32'b11111111111111111100001010101101;
assign LUT_3[43335] = 32'b00000000000000000010110110001010;
assign LUT_3[43336] = 32'b00000000000000000010001110011001;
assign LUT_3[43337] = 32'b00000000000000001000111001110110;
assign LUT_3[43338] = 32'b00000000000000000100010101111101;
assign LUT_3[43339] = 32'b00000000000000001011000001011010;
assign LUT_3[43340] = 32'b11111111111111111111011100001111;
assign LUT_3[43341] = 32'b00000000000000000110000111101100;
assign LUT_3[43342] = 32'b00000000000000000001100011110011;
assign LUT_3[43343] = 32'b00000000000000001000001111010000;
assign LUT_3[43344] = 32'b00000000000000000000001000010110;
assign LUT_3[43345] = 32'b00000000000000000110110011110011;
assign LUT_3[43346] = 32'b00000000000000000010001111111010;
assign LUT_3[43347] = 32'b00000000000000001000111011010111;
assign LUT_3[43348] = 32'b11111111111111111101010110001100;
assign LUT_3[43349] = 32'b00000000000000000100000001101001;
assign LUT_3[43350] = 32'b11111111111111111111011101110000;
assign LUT_3[43351] = 32'b00000000000000000110001001001101;
assign LUT_3[43352] = 32'b00000000000000000101100001011100;
assign LUT_3[43353] = 32'b00000000000000001100001100111001;
assign LUT_3[43354] = 32'b00000000000000000111101001000000;
assign LUT_3[43355] = 32'b00000000000000001110010100011101;
assign LUT_3[43356] = 32'b00000000000000000010101111010010;
assign LUT_3[43357] = 32'b00000000000000001001011010101111;
assign LUT_3[43358] = 32'b00000000000000000100110110110110;
assign LUT_3[43359] = 32'b00000000000000001011100010010011;
assign LUT_3[43360] = 32'b11111111111111111110000011110011;
assign LUT_3[43361] = 32'b00000000000000000100101111010000;
assign LUT_3[43362] = 32'b00000000000000000000001011010111;
assign LUT_3[43363] = 32'b00000000000000000110110110110100;
assign LUT_3[43364] = 32'b11111111111111111011010001101001;
assign LUT_3[43365] = 32'b00000000000000000001111101000110;
assign LUT_3[43366] = 32'b11111111111111111101011001001101;
assign LUT_3[43367] = 32'b00000000000000000100000100101010;
assign LUT_3[43368] = 32'b00000000000000000011011100111001;
assign LUT_3[43369] = 32'b00000000000000001010001000010110;
assign LUT_3[43370] = 32'b00000000000000000101100100011101;
assign LUT_3[43371] = 32'b00000000000000001100001111111010;
assign LUT_3[43372] = 32'b00000000000000000000101010101111;
assign LUT_3[43373] = 32'b00000000000000000111010110001100;
assign LUT_3[43374] = 32'b00000000000000000010110010010011;
assign LUT_3[43375] = 32'b00000000000000001001011101110000;
assign LUT_3[43376] = 32'b00000000000000000001010110110110;
assign LUT_3[43377] = 32'b00000000000000001000000010010011;
assign LUT_3[43378] = 32'b00000000000000000011011110011010;
assign LUT_3[43379] = 32'b00000000000000001010001001110111;
assign LUT_3[43380] = 32'b11111111111111111110100100101100;
assign LUT_3[43381] = 32'b00000000000000000101010000001001;
assign LUT_3[43382] = 32'b00000000000000000000101100010000;
assign LUT_3[43383] = 32'b00000000000000000111010111101101;
assign LUT_3[43384] = 32'b00000000000000000110101111111100;
assign LUT_3[43385] = 32'b00000000000000001101011011011001;
assign LUT_3[43386] = 32'b00000000000000001000110111100000;
assign LUT_3[43387] = 32'b00000000000000001111100010111101;
assign LUT_3[43388] = 32'b00000000000000000011111101110010;
assign LUT_3[43389] = 32'b00000000000000001010101001001111;
assign LUT_3[43390] = 32'b00000000000000000110000101010110;
assign LUT_3[43391] = 32'b00000000000000001100110000110011;
assign LUT_3[43392] = 32'b11111111111111111111000111100110;
assign LUT_3[43393] = 32'b00000000000000000101110011000011;
assign LUT_3[43394] = 32'b00000000000000000001001111001010;
assign LUT_3[43395] = 32'b00000000000000000111111010100111;
assign LUT_3[43396] = 32'b11111111111111111100010101011100;
assign LUT_3[43397] = 32'b00000000000000000011000000111001;
assign LUT_3[43398] = 32'b11111111111111111110011101000000;
assign LUT_3[43399] = 32'b00000000000000000101001000011101;
assign LUT_3[43400] = 32'b00000000000000000100100000101100;
assign LUT_3[43401] = 32'b00000000000000001011001100001001;
assign LUT_3[43402] = 32'b00000000000000000110101000010000;
assign LUT_3[43403] = 32'b00000000000000001101010011101101;
assign LUT_3[43404] = 32'b00000000000000000001101110100010;
assign LUT_3[43405] = 32'b00000000000000001000011001111111;
assign LUT_3[43406] = 32'b00000000000000000011110110000110;
assign LUT_3[43407] = 32'b00000000000000001010100001100011;
assign LUT_3[43408] = 32'b00000000000000000010011010101001;
assign LUT_3[43409] = 32'b00000000000000001001000110000110;
assign LUT_3[43410] = 32'b00000000000000000100100010001101;
assign LUT_3[43411] = 32'b00000000000000001011001101101010;
assign LUT_3[43412] = 32'b11111111111111111111101000011111;
assign LUT_3[43413] = 32'b00000000000000000110010011111100;
assign LUT_3[43414] = 32'b00000000000000000001110000000011;
assign LUT_3[43415] = 32'b00000000000000001000011011100000;
assign LUT_3[43416] = 32'b00000000000000000111110011101111;
assign LUT_3[43417] = 32'b00000000000000001110011111001100;
assign LUT_3[43418] = 32'b00000000000000001001111011010011;
assign LUT_3[43419] = 32'b00000000000000010000100110110000;
assign LUT_3[43420] = 32'b00000000000000000101000001100101;
assign LUT_3[43421] = 32'b00000000000000001011101101000010;
assign LUT_3[43422] = 32'b00000000000000000111001001001001;
assign LUT_3[43423] = 32'b00000000000000001101110100100110;
assign LUT_3[43424] = 32'b00000000000000000000010110000110;
assign LUT_3[43425] = 32'b00000000000000000111000001100011;
assign LUT_3[43426] = 32'b00000000000000000010011101101010;
assign LUT_3[43427] = 32'b00000000000000001001001001000111;
assign LUT_3[43428] = 32'b11111111111111111101100011111100;
assign LUT_3[43429] = 32'b00000000000000000100001111011001;
assign LUT_3[43430] = 32'b11111111111111111111101011100000;
assign LUT_3[43431] = 32'b00000000000000000110010110111101;
assign LUT_3[43432] = 32'b00000000000000000101101111001100;
assign LUT_3[43433] = 32'b00000000000000001100011010101001;
assign LUT_3[43434] = 32'b00000000000000000111110110110000;
assign LUT_3[43435] = 32'b00000000000000001110100010001101;
assign LUT_3[43436] = 32'b00000000000000000010111101000010;
assign LUT_3[43437] = 32'b00000000000000001001101000011111;
assign LUT_3[43438] = 32'b00000000000000000101000100100110;
assign LUT_3[43439] = 32'b00000000000000001011110000000011;
assign LUT_3[43440] = 32'b00000000000000000011101001001001;
assign LUT_3[43441] = 32'b00000000000000001010010100100110;
assign LUT_3[43442] = 32'b00000000000000000101110000101101;
assign LUT_3[43443] = 32'b00000000000000001100011100001010;
assign LUT_3[43444] = 32'b00000000000000000000110110111111;
assign LUT_3[43445] = 32'b00000000000000000111100010011100;
assign LUT_3[43446] = 32'b00000000000000000010111110100011;
assign LUT_3[43447] = 32'b00000000000000001001101010000000;
assign LUT_3[43448] = 32'b00000000000000001001000010001111;
assign LUT_3[43449] = 32'b00000000000000001111101101101100;
assign LUT_3[43450] = 32'b00000000000000001011001001110011;
assign LUT_3[43451] = 32'b00000000000000010001110101010000;
assign LUT_3[43452] = 32'b00000000000000000110010000000101;
assign LUT_3[43453] = 32'b00000000000000001100111011100010;
assign LUT_3[43454] = 32'b00000000000000001000010111101001;
assign LUT_3[43455] = 32'b00000000000000001111000011000110;
assign LUT_3[43456] = 32'b11111111111111111111000000010001;
assign LUT_3[43457] = 32'b00000000000000000101101011101110;
assign LUT_3[43458] = 32'b00000000000000000001000111110101;
assign LUT_3[43459] = 32'b00000000000000000111110011010010;
assign LUT_3[43460] = 32'b11111111111111111100001110000111;
assign LUT_3[43461] = 32'b00000000000000000010111001100100;
assign LUT_3[43462] = 32'b11111111111111111110010101101011;
assign LUT_3[43463] = 32'b00000000000000000101000001001000;
assign LUT_3[43464] = 32'b00000000000000000100011001010111;
assign LUT_3[43465] = 32'b00000000000000001011000100110100;
assign LUT_3[43466] = 32'b00000000000000000110100000111011;
assign LUT_3[43467] = 32'b00000000000000001101001100011000;
assign LUT_3[43468] = 32'b00000000000000000001100111001101;
assign LUT_3[43469] = 32'b00000000000000001000010010101010;
assign LUT_3[43470] = 32'b00000000000000000011101110110001;
assign LUT_3[43471] = 32'b00000000000000001010011010001110;
assign LUT_3[43472] = 32'b00000000000000000010010011010100;
assign LUT_3[43473] = 32'b00000000000000001000111110110001;
assign LUT_3[43474] = 32'b00000000000000000100011010111000;
assign LUT_3[43475] = 32'b00000000000000001011000110010101;
assign LUT_3[43476] = 32'b11111111111111111111100001001010;
assign LUT_3[43477] = 32'b00000000000000000110001100100111;
assign LUT_3[43478] = 32'b00000000000000000001101000101110;
assign LUT_3[43479] = 32'b00000000000000001000010100001011;
assign LUT_3[43480] = 32'b00000000000000000111101100011010;
assign LUT_3[43481] = 32'b00000000000000001110010111110111;
assign LUT_3[43482] = 32'b00000000000000001001110011111110;
assign LUT_3[43483] = 32'b00000000000000010000011111011011;
assign LUT_3[43484] = 32'b00000000000000000100111010010000;
assign LUT_3[43485] = 32'b00000000000000001011100101101101;
assign LUT_3[43486] = 32'b00000000000000000111000001110100;
assign LUT_3[43487] = 32'b00000000000000001101101101010001;
assign LUT_3[43488] = 32'b00000000000000000000001110110001;
assign LUT_3[43489] = 32'b00000000000000000110111010001110;
assign LUT_3[43490] = 32'b00000000000000000010010110010101;
assign LUT_3[43491] = 32'b00000000000000001001000001110010;
assign LUT_3[43492] = 32'b11111111111111111101011100100111;
assign LUT_3[43493] = 32'b00000000000000000100001000000100;
assign LUT_3[43494] = 32'b11111111111111111111100100001011;
assign LUT_3[43495] = 32'b00000000000000000110001111101000;
assign LUT_3[43496] = 32'b00000000000000000101100111110111;
assign LUT_3[43497] = 32'b00000000000000001100010011010100;
assign LUT_3[43498] = 32'b00000000000000000111101111011011;
assign LUT_3[43499] = 32'b00000000000000001110011010111000;
assign LUT_3[43500] = 32'b00000000000000000010110101101101;
assign LUT_3[43501] = 32'b00000000000000001001100001001010;
assign LUT_3[43502] = 32'b00000000000000000100111101010001;
assign LUT_3[43503] = 32'b00000000000000001011101000101110;
assign LUT_3[43504] = 32'b00000000000000000011100001110100;
assign LUT_3[43505] = 32'b00000000000000001010001101010001;
assign LUT_3[43506] = 32'b00000000000000000101101001011000;
assign LUT_3[43507] = 32'b00000000000000001100010100110101;
assign LUT_3[43508] = 32'b00000000000000000000101111101010;
assign LUT_3[43509] = 32'b00000000000000000111011011000111;
assign LUT_3[43510] = 32'b00000000000000000010110111001110;
assign LUT_3[43511] = 32'b00000000000000001001100010101011;
assign LUT_3[43512] = 32'b00000000000000001000111010111010;
assign LUT_3[43513] = 32'b00000000000000001111100110010111;
assign LUT_3[43514] = 32'b00000000000000001011000010011110;
assign LUT_3[43515] = 32'b00000000000000010001101101111011;
assign LUT_3[43516] = 32'b00000000000000000110001000110000;
assign LUT_3[43517] = 32'b00000000000000001100110100001101;
assign LUT_3[43518] = 32'b00000000000000001000010000010100;
assign LUT_3[43519] = 32'b00000000000000001110111011110001;
assign LUT_3[43520] = 32'b00000000000000000100000010010011;
assign LUT_3[43521] = 32'b00000000000000001010101101110000;
assign LUT_3[43522] = 32'b00000000000000000110001001110111;
assign LUT_3[43523] = 32'b00000000000000001100110101010100;
assign LUT_3[43524] = 32'b00000000000000000001010000001001;
assign LUT_3[43525] = 32'b00000000000000000111111011100110;
assign LUT_3[43526] = 32'b00000000000000000011010111101101;
assign LUT_3[43527] = 32'b00000000000000001010000011001010;
assign LUT_3[43528] = 32'b00000000000000001001011011011001;
assign LUT_3[43529] = 32'b00000000000000010000000110110110;
assign LUT_3[43530] = 32'b00000000000000001011100010111101;
assign LUT_3[43531] = 32'b00000000000000010010001110011010;
assign LUT_3[43532] = 32'b00000000000000000110101001001111;
assign LUT_3[43533] = 32'b00000000000000001101010100101100;
assign LUT_3[43534] = 32'b00000000000000001000110000110011;
assign LUT_3[43535] = 32'b00000000000000001111011100010000;
assign LUT_3[43536] = 32'b00000000000000000111010101010110;
assign LUT_3[43537] = 32'b00000000000000001110000000110011;
assign LUT_3[43538] = 32'b00000000000000001001011100111010;
assign LUT_3[43539] = 32'b00000000000000010000001000010111;
assign LUT_3[43540] = 32'b00000000000000000100100011001100;
assign LUT_3[43541] = 32'b00000000000000001011001110101001;
assign LUT_3[43542] = 32'b00000000000000000110101010110000;
assign LUT_3[43543] = 32'b00000000000000001101010110001101;
assign LUT_3[43544] = 32'b00000000000000001100101110011100;
assign LUT_3[43545] = 32'b00000000000000010011011001111001;
assign LUT_3[43546] = 32'b00000000000000001110110110000000;
assign LUT_3[43547] = 32'b00000000000000010101100001011101;
assign LUT_3[43548] = 32'b00000000000000001001111100010010;
assign LUT_3[43549] = 32'b00000000000000010000100111101111;
assign LUT_3[43550] = 32'b00000000000000001100000011110110;
assign LUT_3[43551] = 32'b00000000000000010010101111010011;
assign LUT_3[43552] = 32'b00000000000000000101010000110011;
assign LUT_3[43553] = 32'b00000000000000001011111100010000;
assign LUT_3[43554] = 32'b00000000000000000111011000010111;
assign LUT_3[43555] = 32'b00000000000000001110000011110100;
assign LUT_3[43556] = 32'b00000000000000000010011110101001;
assign LUT_3[43557] = 32'b00000000000000001001001010000110;
assign LUT_3[43558] = 32'b00000000000000000100100110001101;
assign LUT_3[43559] = 32'b00000000000000001011010001101010;
assign LUT_3[43560] = 32'b00000000000000001010101001111001;
assign LUT_3[43561] = 32'b00000000000000010001010101010110;
assign LUT_3[43562] = 32'b00000000000000001100110001011101;
assign LUT_3[43563] = 32'b00000000000000010011011100111010;
assign LUT_3[43564] = 32'b00000000000000000111110111101111;
assign LUT_3[43565] = 32'b00000000000000001110100011001100;
assign LUT_3[43566] = 32'b00000000000000001001111111010011;
assign LUT_3[43567] = 32'b00000000000000010000101010110000;
assign LUT_3[43568] = 32'b00000000000000001000100011110110;
assign LUT_3[43569] = 32'b00000000000000001111001111010011;
assign LUT_3[43570] = 32'b00000000000000001010101011011010;
assign LUT_3[43571] = 32'b00000000000000010001010110110111;
assign LUT_3[43572] = 32'b00000000000000000101110001101100;
assign LUT_3[43573] = 32'b00000000000000001100011101001001;
assign LUT_3[43574] = 32'b00000000000000000111111001010000;
assign LUT_3[43575] = 32'b00000000000000001110100100101101;
assign LUT_3[43576] = 32'b00000000000000001101111100111100;
assign LUT_3[43577] = 32'b00000000000000010100101000011001;
assign LUT_3[43578] = 32'b00000000000000010000000100100000;
assign LUT_3[43579] = 32'b00000000000000010110101111111101;
assign LUT_3[43580] = 32'b00000000000000001011001010110010;
assign LUT_3[43581] = 32'b00000000000000010001110110001111;
assign LUT_3[43582] = 32'b00000000000000001101010010010110;
assign LUT_3[43583] = 32'b00000000000000010011111101110011;
assign LUT_3[43584] = 32'b00000000000000000011111010111110;
assign LUT_3[43585] = 32'b00000000000000001010100110011011;
assign LUT_3[43586] = 32'b00000000000000000110000010100010;
assign LUT_3[43587] = 32'b00000000000000001100101101111111;
assign LUT_3[43588] = 32'b00000000000000000001001000110100;
assign LUT_3[43589] = 32'b00000000000000000111110100010001;
assign LUT_3[43590] = 32'b00000000000000000011010000011000;
assign LUT_3[43591] = 32'b00000000000000001001111011110101;
assign LUT_3[43592] = 32'b00000000000000001001010100000100;
assign LUT_3[43593] = 32'b00000000000000001111111111100001;
assign LUT_3[43594] = 32'b00000000000000001011011011101000;
assign LUT_3[43595] = 32'b00000000000000010010000111000101;
assign LUT_3[43596] = 32'b00000000000000000110100001111010;
assign LUT_3[43597] = 32'b00000000000000001101001101010111;
assign LUT_3[43598] = 32'b00000000000000001000101001011110;
assign LUT_3[43599] = 32'b00000000000000001111010100111011;
assign LUT_3[43600] = 32'b00000000000000000111001110000001;
assign LUT_3[43601] = 32'b00000000000000001101111001011110;
assign LUT_3[43602] = 32'b00000000000000001001010101100101;
assign LUT_3[43603] = 32'b00000000000000010000000001000010;
assign LUT_3[43604] = 32'b00000000000000000100011011110111;
assign LUT_3[43605] = 32'b00000000000000001011000111010100;
assign LUT_3[43606] = 32'b00000000000000000110100011011011;
assign LUT_3[43607] = 32'b00000000000000001101001110111000;
assign LUT_3[43608] = 32'b00000000000000001100100111000111;
assign LUT_3[43609] = 32'b00000000000000010011010010100100;
assign LUT_3[43610] = 32'b00000000000000001110101110101011;
assign LUT_3[43611] = 32'b00000000000000010101011010001000;
assign LUT_3[43612] = 32'b00000000000000001001110100111101;
assign LUT_3[43613] = 32'b00000000000000010000100000011010;
assign LUT_3[43614] = 32'b00000000000000001011111100100001;
assign LUT_3[43615] = 32'b00000000000000010010100111111110;
assign LUT_3[43616] = 32'b00000000000000000101001001011110;
assign LUT_3[43617] = 32'b00000000000000001011110100111011;
assign LUT_3[43618] = 32'b00000000000000000111010001000010;
assign LUT_3[43619] = 32'b00000000000000001101111100011111;
assign LUT_3[43620] = 32'b00000000000000000010010111010100;
assign LUT_3[43621] = 32'b00000000000000001001000010110001;
assign LUT_3[43622] = 32'b00000000000000000100011110111000;
assign LUT_3[43623] = 32'b00000000000000001011001010010101;
assign LUT_3[43624] = 32'b00000000000000001010100010100100;
assign LUT_3[43625] = 32'b00000000000000010001001110000001;
assign LUT_3[43626] = 32'b00000000000000001100101010001000;
assign LUT_3[43627] = 32'b00000000000000010011010101100101;
assign LUT_3[43628] = 32'b00000000000000000111110000011010;
assign LUT_3[43629] = 32'b00000000000000001110011011110111;
assign LUT_3[43630] = 32'b00000000000000001001110111111110;
assign LUT_3[43631] = 32'b00000000000000010000100011011011;
assign LUT_3[43632] = 32'b00000000000000001000011100100001;
assign LUT_3[43633] = 32'b00000000000000001111000111111110;
assign LUT_3[43634] = 32'b00000000000000001010100100000101;
assign LUT_3[43635] = 32'b00000000000000010001001111100010;
assign LUT_3[43636] = 32'b00000000000000000101101010010111;
assign LUT_3[43637] = 32'b00000000000000001100010101110100;
assign LUT_3[43638] = 32'b00000000000000000111110001111011;
assign LUT_3[43639] = 32'b00000000000000001110011101011000;
assign LUT_3[43640] = 32'b00000000000000001101110101100111;
assign LUT_3[43641] = 32'b00000000000000010100100001000100;
assign LUT_3[43642] = 32'b00000000000000001111111101001011;
assign LUT_3[43643] = 32'b00000000000000010110101000101000;
assign LUT_3[43644] = 32'b00000000000000001011000011011101;
assign LUT_3[43645] = 32'b00000000000000010001101110111010;
assign LUT_3[43646] = 32'b00000000000000001101001011000001;
assign LUT_3[43647] = 32'b00000000000000010011110110011110;
assign LUT_3[43648] = 32'b00000000000000000110001101010001;
assign LUT_3[43649] = 32'b00000000000000001100111000101110;
assign LUT_3[43650] = 32'b00000000000000001000010100110101;
assign LUT_3[43651] = 32'b00000000000000001111000000010010;
assign LUT_3[43652] = 32'b00000000000000000011011011000111;
assign LUT_3[43653] = 32'b00000000000000001010000110100100;
assign LUT_3[43654] = 32'b00000000000000000101100010101011;
assign LUT_3[43655] = 32'b00000000000000001100001110001000;
assign LUT_3[43656] = 32'b00000000000000001011100110010111;
assign LUT_3[43657] = 32'b00000000000000010010010001110100;
assign LUT_3[43658] = 32'b00000000000000001101101101111011;
assign LUT_3[43659] = 32'b00000000000000010100011001011000;
assign LUT_3[43660] = 32'b00000000000000001000110100001101;
assign LUT_3[43661] = 32'b00000000000000001111011111101010;
assign LUT_3[43662] = 32'b00000000000000001010111011110001;
assign LUT_3[43663] = 32'b00000000000000010001100111001110;
assign LUT_3[43664] = 32'b00000000000000001001100000010100;
assign LUT_3[43665] = 32'b00000000000000010000001011110001;
assign LUT_3[43666] = 32'b00000000000000001011100111111000;
assign LUT_3[43667] = 32'b00000000000000010010010011010101;
assign LUT_3[43668] = 32'b00000000000000000110101110001010;
assign LUT_3[43669] = 32'b00000000000000001101011001100111;
assign LUT_3[43670] = 32'b00000000000000001000110101101110;
assign LUT_3[43671] = 32'b00000000000000001111100001001011;
assign LUT_3[43672] = 32'b00000000000000001110111001011010;
assign LUT_3[43673] = 32'b00000000000000010101100100110111;
assign LUT_3[43674] = 32'b00000000000000010001000000111110;
assign LUT_3[43675] = 32'b00000000000000010111101100011011;
assign LUT_3[43676] = 32'b00000000000000001100000111010000;
assign LUT_3[43677] = 32'b00000000000000010010110010101101;
assign LUT_3[43678] = 32'b00000000000000001110001110110100;
assign LUT_3[43679] = 32'b00000000000000010100111010010001;
assign LUT_3[43680] = 32'b00000000000000000111011011110001;
assign LUT_3[43681] = 32'b00000000000000001110000111001110;
assign LUT_3[43682] = 32'b00000000000000001001100011010101;
assign LUT_3[43683] = 32'b00000000000000010000001110110010;
assign LUT_3[43684] = 32'b00000000000000000100101001100111;
assign LUT_3[43685] = 32'b00000000000000001011010101000100;
assign LUT_3[43686] = 32'b00000000000000000110110001001011;
assign LUT_3[43687] = 32'b00000000000000001101011100101000;
assign LUT_3[43688] = 32'b00000000000000001100110100110111;
assign LUT_3[43689] = 32'b00000000000000010011100000010100;
assign LUT_3[43690] = 32'b00000000000000001110111100011011;
assign LUT_3[43691] = 32'b00000000000000010101100111111000;
assign LUT_3[43692] = 32'b00000000000000001010000010101101;
assign LUT_3[43693] = 32'b00000000000000010000101110001010;
assign LUT_3[43694] = 32'b00000000000000001100001010010001;
assign LUT_3[43695] = 32'b00000000000000010010110101101110;
assign LUT_3[43696] = 32'b00000000000000001010101110110100;
assign LUT_3[43697] = 32'b00000000000000010001011010010001;
assign LUT_3[43698] = 32'b00000000000000001100110110011000;
assign LUT_3[43699] = 32'b00000000000000010011100001110101;
assign LUT_3[43700] = 32'b00000000000000000111111100101010;
assign LUT_3[43701] = 32'b00000000000000001110101000000111;
assign LUT_3[43702] = 32'b00000000000000001010000100001110;
assign LUT_3[43703] = 32'b00000000000000010000101111101011;
assign LUT_3[43704] = 32'b00000000000000010000000111111010;
assign LUT_3[43705] = 32'b00000000000000010110110011010111;
assign LUT_3[43706] = 32'b00000000000000010010001111011110;
assign LUT_3[43707] = 32'b00000000000000011000111010111011;
assign LUT_3[43708] = 32'b00000000000000001101010101110000;
assign LUT_3[43709] = 32'b00000000000000010100000001001101;
assign LUT_3[43710] = 32'b00000000000000001111011101010100;
assign LUT_3[43711] = 32'b00000000000000010110001000110001;
assign LUT_3[43712] = 32'b00000000000000000110000101111100;
assign LUT_3[43713] = 32'b00000000000000001100110001011001;
assign LUT_3[43714] = 32'b00000000000000001000001101100000;
assign LUT_3[43715] = 32'b00000000000000001110111000111101;
assign LUT_3[43716] = 32'b00000000000000000011010011110010;
assign LUT_3[43717] = 32'b00000000000000001001111111001111;
assign LUT_3[43718] = 32'b00000000000000000101011011010110;
assign LUT_3[43719] = 32'b00000000000000001100000110110011;
assign LUT_3[43720] = 32'b00000000000000001011011111000010;
assign LUT_3[43721] = 32'b00000000000000010010001010011111;
assign LUT_3[43722] = 32'b00000000000000001101100110100110;
assign LUT_3[43723] = 32'b00000000000000010100010010000011;
assign LUT_3[43724] = 32'b00000000000000001000101100111000;
assign LUT_3[43725] = 32'b00000000000000001111011000010101;
assign LUT_3[43726] = 32'b00000000000000001010110100011100;
assign LUT_3[43727] = 32'b00000000000000010001011111111001;
assign LUT_3[43728] = 32'b00000000000000001001011000111111;
assign LUT_3[43729] = 32'b00000000000000010000000100011100;
assign LUT_3[43730] = 32'b00000000000000001011100000100011;
assign LUT_3[43731] = 32'b00000000000000010010001100000000;
assign LUT_3[43732] = 32'b00000000000000000110100110110101;
assign LUT_3[43733] = 32'b00000000000000001101010010010010;
assign LUT_3[43734] = 32'b00000000000000001000101110011001;
assign LUT_3[43735] = 32'b00000000000000001111011001110110;
assign LUT_3[43736] = 32'b00000000000000001110110010000101;
assign LUT_3[43737] = 32'b00000000000000010101011101100010;
assign LUT_3[43738] = 32'b00000000000000010000111001101001;
assign LUT_3[43739] = 32'b00000000000000010111100101000110;
assign LUT_3[43740] = 32'b00000000000000001011111111111011;
assign LUT_3[43741] = 32'b00000000000000010010101011011000;
assign LUT_3[43742] = 32'b00000000000000001110000111011111;
assign LUT_3[43743] = 32'b00000000000000010100110010111100;
assign LUT_3[43744] = 32'b00000000000000000111010100011100;
assign LUT_3[43745] = 32'b00000000000000001101111111111001;
assign LUT_3[43746] = 32'b00000000000000001001011100000000;
assign LUT_3[43747] = 32'b00000000000000010000000111011101;
assign LUT_3[43748] = 32'b00000000000000000100100010010010;
assign LUT_3[43749] = 32'b00000000000000001011001101101111;
assign LUT_3[43750] = 32'b00000000000000000110101001110110;
assign LUT_3[43751] = 32'b00000000000000001101010101010011;
assign LUT_3[43752] = 32'b00000000000000001100101101100010;
assign LUT_3[43753] = 32'b00000000000000010011011000111111;
assign LUT_3[43754] = 32'b00000000000000001110110101000110;
assign LUT_3[43755] = 32'b00000000000000010101100000100011;
assign LUT_3[43756] = 32'b00000000000000001001111011011000;
assign LUT_3[43757] = 32'b00000000000000010000100110110101;
assign LUT_3[43758] = 32'b00000000000000001100000010111100;
assign LUT_3[43759] = 32'b00000000000000010010101110011001;
assign LUT_3[43760] = 32'b00000000000000001010100111011111;
assign LUT_3[43761] = 32'b00000000000000010001010010111100;
assign LUT_3[43762] = 32'b00000000000000001100101111000011;
assign LUT_3[43763] = 32'b00000000000000010011011010100000;
assign LUT_3[43764] = 32'b00000000000000000111110101010101;
assign LUT_3[43765] = 32'b00000000000000001110100000110010;
assign LUT_3[43766] = 32'b00000000000000001001111100111001;
assign LUT_3[43767] = 32'b00000000000000010000101000010110;
assign LUT_3[43768] = 32'b00000000000000010000000000100101;
assign LUT_3[43769] = 32'b00000000000000010110101100000010;
assign LUT_3[43770] = 32'b00000000000000010010001000001001;
assign LUT_3[43771] = 32'b00000000000000011000110011100110;
assign LUT_3[43772] = 32'b00000000000000001101001110011011;
assign LUT_3[43773] = 32'b00000000000000010011111001111000;
assign LUT_3[43774] = 32'b00000000000000001111010101111111;
assign LUT_3[43775] = 32'b00000000000000010110000001011100;
assign LUT_3[43776] = 32'b00000000000000000000010001110100;
assign LUT_3[43777] = 32'b00000000000000000110111101010001;
assign LUT_3[43778] = 32'b00000000000000000010011001011000;
assign LUT_3[43779] = 32'b00000000000000001001000100110101;
assign LUT_3[43780] = 32'b11111111111111111101011111101010;
assign LUT_3[43781] = 32'b00000000000000000100001011000111;
assign LUT_3[43782] = 32'b11111111111111111111100111001110;
assign LUT_3[43783] = 32'b00000000000000000110010010101011;
assign LUT_3[43784] = 32'b00000000000000000101101010111010;
assign LUT_3[43785] = 32'b00000000000000001100010110010111;
assign LUT_3[43786] = 32'b00000000000000000111110010011110;
assign LUT_3[43787] = 32'b00000000000000001110011101111011;
assign LUT_3[43788] = 32'b00000000000000000010111000110000;
assign LUT_3[43789] = 32'b00000000000000001001100100001101;
assign LUT_3[43790] = 32'b00000000000000000101000000010100;
assign LUT_3[43791] = 32'b00000000000000001011101011110001;
assign LUT_3[43792] = 32'b00000000000000000011100100110111;
assign LUT_3[43793] = 32'b00000000000000001010010000010100;
assign LUT_3[43794] = 32'b00000000000000000101101100011011;
assign LUT_3[43795] = 32'b00000000000000001100010111111000;
assign LUT_3[43796] = 32'b00000000000000000000110010101101;
assign LUT_3[43797] = 32'b00000000000000000111011110001010;
assign LUT_3[43798] = 32'b00000000000000000010111010010001;
assign LUT_3[43799] = 32'b00000000000000001001100101101110;
assign LUT_3[43800] = 32'b00000000000000001000111101111101;
assign LUT_3[43801] = 32'b00000000000000001111101001011010;
assign LUT_3[43802] = 32'b00000000000000001011000101100001;
assign LUT_3[43803] = 32'b00000000000000010001110000111110;
assign LUT_3[43804] = 32'b00000000000000000110001011110011;
assign LUT_3[43805] = 32'b00000000000000001100110111010000;
assign LUT_3[43806] = 32'b00000000000000001000010011010111;
assign LUT_3[43807] = 32'b00000000000000001110111110110100;
assign LUT_3[43808] = 32'b00000000000000000001100000010100;
assign LUT_3[43809] = 32'b00000000000000001000001011110001;
assign LUT_3[43810] = 32'b00000000000000000011100111111000;
assign LUT_3[43811] = 32'b00000000000000001010010011010101;
assign LUT_3[43812] = 32'b11111111111111111110101110001010;
assign LUT_3[43813] = 32'b00000000000000000101011001100111;
assign LUT_3[43814] = 32'b00000000000000000000110101101110;
assign LUT_3[43815] = 32'b00000000000000000111100001001011;
assign LUT_3[43816] = 32'b00000000000000000110111001011010;
assign LUT_3[43817] = 32'b00000000000000001101100100110111;
assign LUT_3[43818] = 32'b00000000000000001001000000111110;
assign LUT_3[43819] = 32'b00000000000000001111101100011011;
assign LUT_3[43820] = 32'b00000000000000000100000111010000;
assign LUT_3[43821] = 32'b00000000000000001010110010101101;
assign LUT_3[43822] = 32'b00000000000000000110001110110100;
assign LUT_3[43823] = 32'b00000000000000001100111010010001;
assign LUT_3[43824] = 32'b00000000000000000100110011010111;
assign LUT_3[43825] = 32'b00000000000000001011011110110100;
assign LUT_3[43826] = 32'b00000000000000000110111010111011;
assign LUT_3[43827] = 32'b00000000000000001101100110011000;
assign LUT_3[43828] = 32'b00000000000000000010000001001101;
assign LUT_3[43829] = 32'b00000000000000001000101100101010;
assign LUT_3[43830] = 32'b00000000000000000100001000110001;
assign LUT_3[43831] = 32'b00000000000000001010110100001110;
assign LUT_3[43832] = 32'b00000000000000001010001100011101;
assign LUT_3[43833] = 32'b00000000000000010000110111111010;
assign LUT_3[43834] = 32'b00000000000000001100010100000001;
assign LUT_3[43835] = 32'b00000000000000010010111111011110;
assign LUT_3[43836] = 32'b00000000000000000111011010010011;
assign LUT_3[43837] = 32'b00000000000000001110000101110000;
assign LUT_3[43838] = 32'b00000000000000001001100001110111;
assign LUT_3[43839] = 32'b00000000000000010000001101010100;
assign LUT_3[43840] = 32'b00000000000000000000001010011111;
assign LUT_3[43841] = 32'b00000000000000000110110101111100;
assign LUT_3[43842] = 32'b00000000000000000010010010000011;
assign LUT_3[43843] = 32'b00000000000000001000111101100000;
assign LUT_3[43844] = 32'b11111111111111111101011000010101;
assign LUT_3[43845] = 32'b00000000000000000100000011110010;
assign LUT_3[43846] = 32'b11111111111111111111011111111001;
assign LUT_3[43847] = 32'b00000000000000000110001011010110;
assign LUT_3[43848] = 32'b00000000000000000101100011100101;
assign LUT_3[43849] = 32'b00000000000000001100001111000010;
assign LUT_3[43850] = 32'b00000000000000000111101011001001;
assign LUT_3[43851] = 32'b00000000000000001110010110100110;
assign LUT_3[43852] = 32'b00000000000000000010110001011011;
assign LUT_3[43853] = 32'b00000000000000001001011100111000;
assign LUT_3[43854] = 32'b00000000000000000100111000111111;
assign LUT_3[43855] = 32'b00000000000000001011100100011100;
assign LUT_3[43856] = 32'b00000000000000000011011101100010;
assign LUT_3[43857] = 32'b00000000000000001010001000111111;
assign LUT_3[43858] = 32'b00000000000000000101100101000110;
assign LUT_3[43859] = 32'b00000000000000001100010000100011;
assign LUT_3[43860] = 32'b00000000000000000000101011011000;
assign LUT_3[43861] = 32'b00000000000000000111010110110101;
assign LUT_3[43862] = 32'b00000000000000000010110010111100;
assign LUT_3[43863] = 32'b00000000000000001001011110011001;
assign LUT_3[43864] = 32'b00000000000000001000110110101000;
assign LUT_3[43865] = 32'b00000000000000001111100010000101;
assign LUT_3[43866] = 32'b00000000000000001010111110001100;
assign LUT_3[43867] = 32'b00000000000000010001101001101001;
assign LUT_3[43868] = 32'b00000000000000000110000100011110;
assign LUT_3[43869] = 32'b00000000000000001100101111111011;
assign LUT_3[43870] = 32'b00000000000000001000001100000010;
assign LUT_3[43871] = 32'b00000000000000001110110111011111;
assign LUT_3[43872] = 32'b00000000000000000001011000111111;
assign LUT_3[43873] = 32'b00000000000000001000000100011100;
assign LUT_3[43874] = 32'b00000000000000000011100000100011;
assign LUT_3[43875] = 32'b00000000000000001010001100000000;
assign LUT_3[43876] = 32'b11111111111111111110100110110101;
assign LUT_3[43877] = 32'b00000000000000000101010010010010;
assign LUT_3[43878] = 32'b00000000000000000000101110011001;
assign LUT_3[43879] = 32'b00000000000000000111011001110110;
assign LUT_3[43880] = 32'b00000000000000000110110010000101;
assign LUT_3[43881] = 32'b00000000000000001101011101100010;
assign LUT_3[43882] = 32'b00000000000000001000111001101001;
assign LUT_3[43883] = 32'b00000000000000001111100101000110;
assign LUT_3[43884] = 32'b00000000000000000011111111111011;
assign LUT_3[43885] = 32'b00000000000000001010101011011000;
assign LUT_3[43886] = 32'b00000000000000000110000111011111;
assign LUT_3[43887] = 32'b00000000000000001100110010111100;
assign LUT_3[43888] = 32'b00000000000000000100101100000010;
assign LUT_3[43889] = 32'b00000000000000001011010111011111;
assign LUT_3[43890] = 32'b00000000000000000110110011100110;
assign LUT_3[43891] = 32'b00000000000000001101011111000011;
assign LUT_3[43892] = 32'b00000000000000000001111001111000;
assign LUT_3[43893] = 32'b00000000000000001000100101010101;
assign LUT_3[43894] = 32'b00000000000000000100000001011100;
assign LUT_3[43895] = 32'b00000000000000001010101100111001;
assign LUT_3[43896] = 32'b00000000000000001010000101001000;
assign LUT_3[43897] = 32'b00000000000000010000110000100101;
assign LUT_3[43898] = 32'b00000000000000001100001100101100;
assign LUT_3[43899] = 32'b00000000000000010010111000001001;
assign LUT_3[43900] = 32'b00000000000000000111010010111110;
assign LUT_3[43901] = 32'b00000000000000001101111110011011;
assign LUT_3[43902] = 32'b00000000000000001001011010100010;
assign LUT_3[43903] = 32'b00000000000000010000000101111111;
assign LUT_3[43904] = 32'b00000000000000000010011100110010;
assign LUT_3[43905] = 32'b00000000000000001001001000001111;
assign LUT_3[43906] = 32'b00000000000000000100100100010110;
assign LUT_3[43907] = 32'b00000000000000001011001111110011;
assign LUT_3[43908] = 32'b11111111111111111111101010101000;
assign LUT_3[43909] = 32'b00000000000000000110010110000101;
assign LUT_3[43910] = 32'b00000000000000000001110010001100;
assign LUT_3[43911] = 32'b00000000000000001000011101101001;
assign LUT_3[43912] = 32'b00000000000000000111110101111000;
assign LUT_3[43913] = 32'b00000000000000001110100001010101;
assign LUT_3[43914] = 32'b00000000000000001001111101011100;
assign LUT_3[43915] = 32'b00000000000000010000101000111001;
assign LUT_3[43916] = 32'b00000000000000000101000011101110;
assign LUT_3[43917] = 32'b00000000000000001011101111001011;
assign LUT_3[43918] = 32'b00000000000000000111001011010010;
assign LUT_3[43919] = 32'b00000000000000001101110110101111;
assign LUT_3[43920] = 32'b00000000000000000101101111110101;
assign LUT_3[43921] = 32'b00000000000000001100011011010010;
assign LUT_3[43922] = 32'b00000000000000000111110111011001;
assign LUT_3[43923] = 32'b00000000000000001110100010110110;
assign LUT_3[43924] = 32'b00000000000000000010111101101011;
assign LUT_3[43925] = 32'b00000000000000001001101001001000;
assign LUT_3[43926] = 32'b00000000000000000101000101001111;
assign LUT_3[43927] = 32'b00000000000000001011110000101100;
assign LUT_3[43928] = 32'b00000000000000001011001000111011;
assign LUT_3[43929] = 32'b00000000000000010001110100011000;
assign LUT_3[43930] = 32'b00000000000000001101010000011111;
assign LUT_3[43931] = 32'b00000000000000010011111011111100;
assign LUT_3[43932] = 32'b00000000000000001000010110110001;
assign LUT_3[43933] = 32'b00000000000000001111000010001110;
assign LUT_3[43934] = 32'b00000000000000001010011110010101;
assign LUT_3[43935] = 32'b00000000000000010001001001110010;
assign LUT_3[43936] = 32'b00000000000000000011101011010010;
assign LUT_3[43937] = 32'b00000000000000001010010110101111;
assign LUT_3[43938] = 32'b00000000000000000101110010110110;
assign LUT_3[43939] = 32'b00000000000000001100011110010011;
assign LUT_3[43940] = 32'b00000000000000000000111001001000;
assign LUT_3[43941] = 32'b00000000000000000111100100100101;
assign LUT_3[43942] = 32'b00000000000000000011000000101100;
assign LUT_3[43943] = 32'b00000000000000001001101100001001;
assign LUT_3[43944] = 32'b00000000000000001001000100011000;
assign LUT_3[43945] = 32'b00000000000000001111101111110101;
assign LUT_3[43946] = 32'b00000000000000001011001011111100;
assign LUT_3[43947] = 32'b00000000000000010001110111011001;
assign LUT_3[43948] = 32'b00000000000000000110010010001110;
assign LUT_3[43949] = 32'b00000000000000001100111101101011;
assign LUT_3[43950] = 32'b00000000000000001000011001110010;
assign LUT_3[43951] = 32'b00000000000000001111000101001111;
assign LUT_3[43952] = 32'b00000000000000000110111110010101;
assign LUT_3[43953] = 32'b00000000000000001101101001110010;
assign LUT_3[43954] = 32'b00000000000000001001000101111001;
assign LUT_3[43955] = 32'b00000000000000001111110001010110;
assign LUT_3[43956] = 32'b00000000000000000100001100001011;
assign LUT_3[43957] = 32'b00000000000000001010110111101000;
assign LUT_3[43958] = 32'b00000000000000000110010011101111;
assign LUT_3[43959] = 32'b00000000000000001100111111001100;
assign LUT_3[43960] = 32'b00000000000000001100010111011011;
assign LUT_3[43961] = 32'b00000000000000010011000010111000;
assign LUT_3[43962] = 32'b00000000000000001110011110111111;
assign LUT_3[43963] = 32'b00000000000000010101001010011100;
assign LUT_3[43964] = 32'b00000000000000001001100101010001;
assign LUT_3[43965] = 32'b00000000000000010000010000101110;
assign LUT_3[43966] = 32'b00000000000000001011101100110101;
assign LUT_3[43967] = 32'b00000000000000010010011000010010;
assign LUT_3[43968] = 32'b00000000000000000010010101011101;
assign LUT_3[43969] = 32'b00000000000000001001000000111010;
assign LUT_3[43970] = 32'b00000000000000000100011101000001;
assign LUT_3[43971] = 32'b00000000000000001011001000011110;
assign LUT_3[43972] = 32'b11111111111111111111100011010011;
assign LUT_3[43973] = 32'b00000000000000000110001110110000;
assign LUT_3[43974] = 32'b00000000000000000001101010110111;
assign LUT_3[43975] = 32'b00000000000000001000010110010100;
assign LUT_3[43976] = 32'b00000000000000000111101110100011;
assign LUT_3[43977] = 32'b00000000000000001110011010000000;
assign LUT_3[43978] = 32'b00000000000000001001110110000111;
assign LUT_3[43979] = 32'b00000000000000010000100001100100;
assign LUT_3[43980] = 32'b00000000000000000100111100011001;
assign LUT_3[43981] = 32'b00000000000000001011100111110110;
assign LUT_3[43982] = 32'b00000000000000000111000011111101;
assign LUT_3[43983] = 32'b00000000000000001101101111011010;
assign LUT_3[43984] = 32'b00000000000000000101101000100000;
assign LUT_3[43985] = 32'b00000000000000001100010011111101;
assign LUT_3[43986] = 32'b00000000000000000111110000000100;
assign LUT_3[43987] = 32'b00000000000000001110011011100001;
assign LUT_3[43988] = 32'b00000000000000000010110110010110;
assign LUT_3[43989] = 32'b00000000000000001001100001110011;
assign LUT_3[43990] = 32'b00000000000000000100111101111010;
assign LUT_3[43991] = 32'b00000000000000001011101001010111;
assign LUT_3[43992] = 32'b00000000000000001011000001100110;
assign LUT_3[43993] = 32'b00000000000000010001101101000011;
assign LUT_3[43994] = 32'b00000000000000001101001001001010;
assign LUT_3[43995] = 32'b00000000000000010011110100100111;
assign LUT_3[43996] = 32'b00000000000000001000001111011100;
assign LUT_3[43997] = 32'b00000000000000001110111010111001;
assign LUT_3[43998] = 32'b00000000000000001010010111000000;
assign LUT_3[43999] = 32'b00000000000000010001000010011101;
assign LUT_3[44000] = 32'b00000000000000000011100011111101;
assign LUT_3[44001] = 32'b00000000000000001010001111011010;
assign LUT_3[44002] = 32'b00000000000000000101101011100001;
assign LUT_3[44003] = 32'b00000000000000001100010110111110;
assign LUT_3[44004] = 32'b00000000000000000000110001110011;
assign LUT_3[44005] = 32'b00000000000000000111011101010000;
assign LUT_3[44006] = 32'b00000000000000000010111001010111;
assign LUT_3[44007] = 32'b00000000000000001001100100110100;
assign LUT_3[44008] = 32'b00000000000000001000111101000011;
assign LUT_3[44009] = 32'b00000000000000001111101000100000;
assign LUT_3[44010] = 32'b00000000000000001011000100100111;
assign LUT_3[44011] = 32'b00000000000000010001110000000100;
assign LUT_3[44012] = 32'b00000000000000000110001010111001;
assign LUT_3[44013] = 32'b00000000000000001100110110010110;
assign LUT_3[44014] = 32'b00000000000000001000010010011101;
assign LUT_3[44015] = 32'b00000000000000001110111101111010;
assign LUT_3[44016] = 32'b00000000000000000110110111000000;
assign LUT_3[44017] = 32'b00000000000000001101100010011101;
assign LUT_3[44018] = 32'b00000000000000001000111110100100;
assign LUT_3[44019] = 32'b00000000000000001111101010000001;
assign LUT_3[44020] = 32'b00000000000000000100000100110110;
assign LUT_3[44021] = 32'b00000000000000001010110000010011;
assign LUT_3[44022] = 32'b00000000000000000110001100011010;
assign LUT_3[44023] = 32'b00000000000000001100110111110111;
assign LUT_3[44024] = 32'b00000000000000001100010000000110;
assign LUT_3[44025] = 32'b00000000000000010010111011100011;
assign LUT_3[44026] = 32'b00000000000000001110010111101010;
assign LUT_3[44027] = 32'b00000000000000010101000011000111;
assign LUT_3[44028] = 32'b00000000000000001001011101111100;
assign LUT_3[44029] = 32'b00000000000000010000001001011001;
assign LUT_3[44030] = 32'b00000000000000001011100101100000;
assign LUT_3[44031] = 32'b00000000000000010010010000111101;
assign LUT_3[44032] = 32'b00000000000000000111010010000100;
assign LUT_3[44033] = 32'b00000000000000001101111101100001;
assign LUT_3[44034] = 32'b00000000000000001001011001101000;
assign LUT_3[44035] = 32'b00000000000000010000000101000101;
assign LUT_3[44036] = 32'b00000000000000000100011111111010;
assign LUT_3[44037] = 32'b00000000000000001011001011010111;
assign LUT_3[44038] = 32'b00000000000000000110100111011110;
assign LUT_3[44039] = 32'b00000000000000001101010010111011;
assign LUT_3[44040] = 32'b00000000000000001100101011001010;
assign LUT_3[44041] = 32'b00000000000000010011010110100111;
assign LUT_3[44042] = 32'b00000000000000001110110010101110;
assign LUT_3[44043] = 32'b00000000000000010101011110001011;
assign LUT_3[44044] = 32'b00000000000000001001111001000000;
assign LUT_3[44045] = 32'b00000000000000010000100100011101;
assign LUT_3[44046] = 32'b00000000000000001100000000100100;
assign LUT_3[44047] = 32'b00000000000000010010101100000001;
assign LUT_3[44048] = 32'b00000000000000001010100101000111;
assign LUT_3[44049] = 32'b00000000000000010001010000100100;
assign LUT_3[44050] = 32'b00000000000000001100101100101011;
assign LUT_3[44051] = 32'b00000000000000010011011000001000;
assign LUT_3[44052] = 32'b00000000000000000111110010111101;
assign LUT_3[44053] = 32'b00000000000000001110011110011010;
assign LUT_3[44054] = 32'b00000000000000001001111010100001;
assign LUT_3[44055] = 32'b00000000000000010000100101111110;
assign LUT_3[44056] = 32'b00000000000000001111111110001101;
assign LUT_3[44057] = 32'b00000000000000010110101001101010;
assign LUT_3[44058] = 32'b00000000000000010010000101110001;
assign LUT_3[44059] = 32'b00000000000000011000110001001110;
assign LUT_3[44060] = 32'b00000000000000001101001100000011;
assign LUT_3[44061] = 32'b00000000000000010011110111100000;
assign LUT_3[44062] = 32'b00000000000000001111010011100111;
assign LUT_3[44063] = 32'b00000000000000010101111111000100;
assign LUT_3[44064] = 32'b00000000000000001000100000100100;
assign LUT_3[44065] = 32'b00000000000000001111001100000001;
assign LUT_3[44066] = 32'b00000000000000001010101000001000;
assign LUT_3[44067] = 32'b00000000000000010001010011100101;
assign LUT_3[44068] = 32'b00000000000000000101101110011010;
assign LUT_3[44069] = 32'b00000000000000001100011001110111;
assign LUT_3[44070] = 32'b00000000000000000111110101111110;
assign LUT_3[44071] = 32'b00000000000000001110100001011011;
assign LUT_3[44072] = 32'b00000000000000001101111001101010;
assign LUT_3[44073] = 32'b00000000000000010100100101000111;
assign LUT_3[44074] = 32'b00000000000000010000000001001110;
assign LUT_3[44075] = 32'b00000000000000010110101100101011;
assign LUT_3[44076] = 32'b00000000000000001011000111100000;
assign LUT_3[44077] = 32'b00000000000000010001110010111101;
assign LUT_3[44078] = 32'b00000000000000001101001111000100;
assign LUT_3[44079] = 32'b00000000000000010011111010100001;
assign LUT_3[44080] = 32'b00000000000000001011110011100111;
assign LUT_3[44081] = 32'b00000000000000010010011111000100;
assign LUT_3[44082] = 32'b00000000000000001101111011001011;
assign LUT_3[44083] = 32'b00000000000000010100100110101000;
assign LUT_3[44084] = 32'b00000000000000001001000001011101;
assign LUT_3[44085] = 32'b00000000000000001111101100111010;
assign LUT_3[44086] = 32'b00000000000000001011001001000001;
assign LUT_3[44087] = 32'b00000000000000010001110100011110;
assign LUT_3[44088] = 32'b00000000000000010001001100101101;
assign LUT_3[44089] = 32'b00000000000000010111111000001010;
assign LUT_3[44090] = 32'b00000000000000010011010100010001;
assign LUT_3[44091] = 32'b00000000000000011001111111101110;
assign LUT_3[44092] = 32'b00000000000000001110011010100011;
assign LUT_3[44093] = 32'b00000000000000010101000110000000;
assign LUT_3[44094] = 32'b00000000000000010000100010000111;
assign LUT_3[44095] = 32'b00000000000000010111001101100100;
assign LUT_3[44096] = 32'b00000000000000000111001010101111;
assign LUT_3[44097] = 32'b00000000000000001101110110001100;
assign LUT_3[44098] = 32'b00000000000000001001010010010011;
assign LUT_3[44099] = 32'b00000000000000001111111101110000;
assign LUT_3[44100] = 32'b00000000000000000100011000100101;
assign LUT_3[44101] = 32'b00000000000000001011000100000010;
assign LUT_3[44102] = 32'b00000000000000000110100000001001;
assign LUT_3[44103] = 32'b00000000000000001101001011100110;
assign LUT_3[44104] = 32'b00000000000000001100100011110101;
assign LUT_3[44105] = 32'b00000000000000010011001111010010;
assign LUT_3[44106] = 32'b00000000000000001110101011011001;
assign LUT_3[44107] = 32'b00000000000000010101010110110110;
assign LUT_3[44108] = 32'b00000000000000001001110001101011;
assign LUT_3[44109] = 32'b00000000000000010000011101001000;
assign LUT_3[44110] = 32'b00000000000000001011111001001111;
assign LUT_3[44111] = 32'b00000000000000010010100100101100;
assign LUT_3[44112] = 32'b00000000000000001010011101110010;
assign LUT_3[44113] = 32'b00000000000000010001001001001111;
assign LUT_3[44114] = 32'b00000000000000001100100101010110;
assign LUT_3[44115] = 32'b00000000000000010011010000110011;
assign LUT_3[44116] = 32'b00000000000000000111101011101000;
assign LUT_3[44117] = 32'b00000000000000001110010111000101;
assign LUT_3[44118] = 32'b00000000000000001001110011001100;
assign LUT_3[44119] = 32'b00000000000000010000011110101001;
assign LUT_3[44120] = 32'b00000000000000001111110110111000;
assign LUT_3[44121] = 32'b00000000000000010110100010010101;
assign LUT_3[44122] = 32'b00000000000000010001111110011100;
assign LUT_3[44123] = 32'b00000000000000011000101001111001;
assign LUT_3[44124] = 32'b00000000000000001101000100101110;
assign LUT_3[44125] = 32'b00000000000000010011110000001011;
assign LUT_3[44126] = 32'b00000000000000001111001100010010;
assign LUT_3[44127] = 32'b00000000000000010101110111101111;
assign LUT_3[44128] = 32'b00000000000000001000011001001111;
assign LUT_3[44129] = 32'b00000000000000001111000100101100;
assign LUT_3[44130] = 32'b00000000000000001010100000110011;
assign LUT_3[44131] = 32'b00000000000000010001001100010000;
assign LUT_3[44132] = 32'b00000000000000000101100111000101;
assign LUT_3[44133] = 32'b00000000000000001100010010100010;
assign LUT_3[44134] = 32'b00000000000000000111101110101001;
assign LUT_3[44135] = 32'b00000000000000001110011010000110;
assign LUT_3[44136] = 32'b00000000000000001101110010010101;
assign LUT_3[44137] = 32'b00000000000000010100011101110010;
assign LUT_3[44138] = 32'b00000000000000001111111001111001;
assign LUT_3[44139] = 32'b00000000000000010110100101010110;
assign LUT_3[44140] = 32'b00000000000000001011000000001011;
assign LUT_3[44141] = 32'b00000000000000010001101011101000;
assign LUT_3[44142] = 32'b00000000000000001101000111101111;
assign LUT_3[44143] = 32'b00000000000000010011110011001100;
assign LUT_3[44144] = 32'b00000000000000001011101100010010;
assign LUT_3[44145] = 32'b00000000000000010010010111101111;
assign LUT_3[44146] = 32'b00000000000000001101110011110110;
assign LUT_3[44147] = 32'b00000000000000010100011111010011;
assign LUT_3[44148] = 32'b00000000000000001000111010001000;
assign LUT_3[44149] = 32'b00000000000000001111100101100101;
assign LUT_3[44150] = 32'b00000000000000001011000001101100;
assign LUT_3[44151] = 32'b00000000000000010001101101001001;
assign LUT_3[44152] = 32'b00000000000000010001000101011000;
assign LUT_3[44153] = 32'b00000000000000010111110000110101;
assign LUT_3[44154] = 32'b00000000000000010011001100111100;
assign LUT_3[44155] = 32'b00000000000000011001111000011001;
assign LUT_3[44156] = 32'b00000000000000001110010011001110;
assign LUT_3[44157] = 32'b00000000000000010100111110101011;
assign LUT_3[44158] = 32'b00000000000000010000011010110010;
assign LUT_3[44159] = 32'b00000000000000010111000110001111;
assign LUT_3[44160] = 32'b00000000000000001001011101000010;
assign LUT_3[44161] = 32'b00000000000000010000001000011111;
assign LUT_3[44162] = 32'b00000000000000001011100100100110;
assign LUT_3[44163] = 32'b00000000000000010010010000000011;
assign LUT_3[44164] = 32'b00000000000000000110101010111000;
assign LUT_3[44165] = 32'b00000000000000001101010110010101;
assign LUT_3[44166] = 32'b00000000000000001000110010011100;
assign LUT_3[44167] = 32'b00000000000000001111011101111001;
assign LUT_3[44168] = 32'b00000000000000001110110110001000;
assign LUT_3[44169] = 32'b00000000000000010101100001100101;
assign LUT_3[44170] = 32'b00000000000000010000111101101100;
assign LUT_3[44171] = 32'b00000000000000010111101001001001;
assign LUT_3[44172] = 32'b00000000000000001100000011111110;
assign LUT_3[44173] = 32'b00000000000000010010101111011011;
assign LUT_3[44174] = 32'b00000000000000001110001011100010;
assign LUT_3[44175] = 32'b00000000000000010100110110111111;
assign LUT_3[44176] = 32'b00000000000000001100110000000101;
assign LUT_3[44177] = 32'b00000000000000010011011011100010;
assign LUT_3[44178] = 32'b00000000000000001110110111101001;
assign LUT_3[44179] = 32'b00000000000000010101100011000110;
assign LUT_3[44180] = 32'b00000000000000001001111101111011;
assign LUT_3[44181] = 32'b00000000000000010000101001011000;
assign LUT_3[44182] = 32'b00000000000000001100000101011111;
assign LUT_3[44183] = 32'b00000000000000010010110000111100;
assign LUT_3[44184] = 32'b00000000000000010010001001001011;
assign LUT_3[44185] = 32'b00000000000000011000110100101000;
assign LUT_3[44186] = 32'b00000000000000010100010000101111;
assign LUT_3[44187] = 32'b00000000000000011010111100001100;
assign LUT_3[44188] = 32'b00000000000000001111010111000001;
assign LUT_3[44189] = 32'b00000000000000010110000010011110;
assign LUT_3[44190] = 32'b00000000000000010001011110100101;
assign LUT_3[44191] = 32'b00000000000000011000001010000010;
assign LUT_3[44192] = 32'b00000000000000001010101011100010;
assign LUT_3[44193] = 32'b00000000000000010001010110111111;
assign LUT_3[44194] = 32'b00000000000000001100110011000110;
assign LUT_3[44195] = 32'b00000000000000010011011110100011;
assign LUT_3[44196] = 32'b00000000000000000111111001011000;
assign LUT_3[44197] = 32'b00000000000000001110100100110101;
assign LUT_3[44198] = 32'b00000000000000001010000000111100;
assign LUT_3[44199] = 32'b00000000000000010000101100011001;
assign LUT_3[44200] = 32'b00000000000000010000000100101000;
assign LUT_3[44201] = 32'b00000000000000010110110000000101;
assign LUT_3[44202] = 32'b00000000000000010010001100001100;
assign LUT_3[44203] = 32'b00000000000000011000110111101001;
assign LUT_3[44204] = 32'b00000000000000001101010010011110;
assign LUT_3[44205] = 32'b00000000000000010011111101111011;
assign LUT_3[44206] = 32'b00000000000000001111011010000010;
assign LUT_3[44207] = 32'b00000000000000010110000101011111;
assign LUT_3[44208] = 32'b00000000000000001101111110100101;
assign LUT_3[44209] = 32'b00000000000000010100101010000010;
assign LUT_3[44210] = 32'b00000000000000010000000110001001;
assign LUT_3[44211] = 32'b00000000000000010110110001100110;
assign LUT_3[44212] = 32'b00000000000000001011001100011011;
assign LUT_3[44213] = 32'b00000000000000010001110111111000;
assign LUT_3[44214] = 32'b00000000000000001101010011111111;
assign LUT_3[44215] = 32'b00000000000000010011111111011100;
assign LUT_3[44216] = 32'b00000000000000010011010111101011;
assign LUT_3[44217] = 32'b00000000000000011010000011001000;
assign LUT_3[44218] = 32'b00000000000000010101011111001111;
assign LUT_3[44219] = 32'b00000000000000011100001010101100;
assign LUT_3[44220] = 32'b00000000000000010000100101100001;
assign LUT_3[44221] = 32'b00000000000000010111010000111110;
assign LUT_3[44222] = 32'b00000000000000010010101101000101;
assign LUT_3[44223] = 32'b00000000000000011001011000100010;
assign LUT_3[44224] = 32'b00000000000000001001010101101101;
assign LUT_3[44225] = 32'b00000000000000010000000001001010;
assign LUT_3[44226] = 32'b00000000000000001011011101010001;
assign LUT_3[44227] = 32'b00000000000000010010001000101110;
assign LUT_3[44228] = 32'b00000000000000000110100011100011;
assign LUT_3[44229] = 32'b00000000000000001101001111000000;
assign LUT_3[44230] = 32'b00000000000000001000101011000111;
assign LUT_3[44231] = 32'b00000000000000001111010110100100;
assign LUT_3[44232] = 32'b00000000000000001110101110110011;
assign LUT_3[44233] = 32'b00000000000000010101011010010000;
assign LUT_3[44234] = 32'b00000000000000010000110110010111;
assign LUT_3[44235] = 32'b00000000000000010111100001110100;
assign LUT_3[44236] = 32'b00000000000000001011111100101001;
assign LUT_3[44237] = 32'b00000000000000010010101000000110;
assign LUT_3[44238] = 32'b00000000000000001110000100001101;
assign LUT_3[44239] = 32'b00000000000000010100101111101010;
assign LUT_3[44240] = 32'b00000000000000001100101000110000;
assign LUT_3[44241] = 32'b00000000000000010011010100001101;
assign LUT_3[44242] = 32'b00000000000000001110110000010100;
assign LUT_3[44243] = 32'b00000000000000010101011011110001;
assign LUT_3[44244] = 32'b00000000000000001001110110100110;
assign LUT_3[44245] = 32'b00000000000000010000100010000011;
assign LUT_3[44246] = 32'b00000000000000001011111110001010;
assign LUT_3[44247] = 32'b00000000000000010010101001100111;
assign LUT_3[44248] = 32'b00000000000000010010000001110110;
assign LUT_3[44249] = 32'b00000000000000011000101101010011;
assign LUT_3[44250] = 32'b00000000000000010100001001011010;
assign LUT_3[44251] = 32'b00000000000000011010110100110111;
assign LUT_3[44252] = 32'b00000000000000001111001111101100;
assign LUT_3[44253] = 32'b00000000000000010101111011001001;
assign LUT_3[44254] = 32'b00000000000000010001010111010000;
assign LUT_3[44255] = 32'b00000000000000011000000010101101;
assign LUT_3[44256] = 32'b00000000000000001010100100001101;
assign LUT_3[44257] = 32'b00000000000000010001001111101010;
assign LUT_3[44258] = 32'b00000000000000001100101011110001;
assign LUT_3[44259] = 32'b00000000000000010011010111001110;
assign LUT_3[44260] = 32'b00000000000000000111110010000011;
assign LUT_3[44261] = 32'b00000000000000001110011101100000;
assign LUT_3[44262] = 32'b00000000000000001001111001100111;
assign LUT_3[44263] = 32'b00000000000000010000100101000100;
assign LUT_3[44264] = 32'b00000000000000001111111101010011;
assign LUT_3[44265] = 32'b00000000000000010110101000110000;
assign LUT_3[44266] = 32'b00000000000000010010000100110111;
assign LUT_3[44267] = 32'b00000000000000011000110000010100;
assign LUT_3[44268] = 32'b00000000000000001101001011001001;
assign LUT_3[44269] = 32'b00000000000000010011110110100110;
assign LUT_3[44270] = 32'b00000000000000001111010010101101;
assign LUT_3[44271] = 32'b00000000000000010101111110001010;
assign LUT_3[44272] = 32'b00000000000000001101110111010000;
assign LUT_3[44273] = 32'b00000000000000010100100010101101;
assign LUT_3[44274] = 32'b00000000000000001111111110110100;
assign LUT_3[44275] = 32'b00000000000000010110101010010001;
assign LUT_3[44276] = 32'b00000000000000001011000101000110;
assign LUT_3[44277] = 32'b00000000000000010001110000100011;
assign LUT_3[44278] = 32'b00000000000000001101001100101010;
assign LUT_3[44279] = 32'b00000000000000010011111000000111;
assign LUT_3[44280] = 32'b00000000000000010011010000010110;
assign LUT_3[44281] = 32'b00000000000000011001111011110011;
assign LUT_3[44282] = 32'b00000000000000010101010111111010;
assign LUT_3[44283] = 32'b00000000000000011100000011010111;
assign LUT_3[44284] = 32'b00000000000000010000011110001100;
assign LUT_3[44285] = 32'b00000000000000010111001001101001;
assign LUT_3[44286] = 32'b00000000000000010010100101110000;
assign LUT_3[44287] = 32'b00000000000000011001010001001101;
assign LUT_3[44288] = 32'b00000000000000000011100001100101;
assign LUT_3[44289] = 32'b00000000000000001010001101000010;
assign LUT_3[44290] = 32'b00000000000000000101101001001001;
assign LUT_3[44291] = 32'b00000000000000001100010100100110;
assign LUT_3[44292] = 32'b00000000000000000000101111011011;
assign LUT_3[44293] = 32'b00000000000000000111011010111000;
assign LUT_3[44294] = 32'b00000000000000000010110110111111;
assign LUT_3[44295] = 32'b00000000000000001001100010011100;
assign LUT_3[44296] = 32'b00000000000000001000111010101011;
assign LUT_3[44297] = 32'b00000000000000001111100110001000;
assign LUT_3[44298] = 32'b00000000000000001011000010001111;
assign LUT_3[44299] = 32'b00000000000000010001101101101100;
assign LUT_3[44300] = 32'b00000000000000000110001000100001;
assign LUT_3[44301] = 32'b00000000000000001100110011111110;
assign LUT_3[44302] = 32'b00000000000000001000010000000101;
assign LUT_3[44303] = 32'b00000000000000001110111011100010;
assign LUT_3[44304] = 32'b00000000000000000110110100101000;
assign LUT_3[44305] = 32'b00000000000000001101100000000101;
assign LUT_3[44306] = 32'b00000000000000001000111100001100;
assign LUT_3[44307] = 32'b00000000000000001111100111101001;
assign LUT_3[44308] = 32'b00000000000000000100000010011110;
assign LUT_3[44309] = 32'b00000000000000001010101101111011;
assign LUT_3[44310] = 32'b00000000000000000110001010000010;
assign LUT_3[44311] = 32'b00000000000000001100110101011111;
assign LUT_3[44312] = 32'b00000000000000001100001101101110;
assign LUT_3[44313] = 32'b00000000000000010010111001001011;
assign LUT_3[44314] = 32'b00000000000000001110010101010010;
assign LUT_3[44315] = 32'b00000000000000010101000000101111;
assign LUT_3[44316] = 32'b00000000000000001001011011100100;
assign LUT_3[44317] = 32'b00000000000000010000000111000001;
assign LUT_3[44318] = 32'b00000000000000001011100011001000;
assign LUT_3[44319] = 32'b00000000000000010010001110100101;
assign LUT_3[44320] = 32'b00000000000000000100110000000101;
assign LUT_3[44321] = 32'b00000000000000001011011011100010;
assign LUT_3[44322] = 32'b00000000000000000110110111101001;
assign LUT_3[44323] = 32'b00000000000000001101100011000110;
assign LUT_3[44324] = 32'b00000000000000000001111101111011;
assign LUT_3[44325] = 32'b00000000000000001000101001011000;
assign LUT_3[44326] = 32'b00000000000000000100000101011111;
assign LUT_3[44327] = 32'b00000000000000001010110000111100;
assign LUT_3[44328] = 32'b00000000000000001010001001001011;
assign LUT_3[44329] = 32'b00000000000000010000110100101000;
assign LUT_3[44330] = 32'b00000000000000001100010000101111;
assign LUT_3[44331] = 32'b00000000000000010010111100001100;
assign LUT_3[44332] = 32'b00000000000000000111010111000001;
assign LUT_3[44333] = 32'b00000000000000001110000010011110;
assign LUT_3[44334] = 32'b00000000000000001001011110100101;
assign LUT_3[44335] = 32'b00000000000000010000001010000010;
assign LUT_3[44336] = 32'b00000000000000001000000011001000;
assign LUT_3[44337] = 32'b00000000000000001110101110100101;
assign LUT_3[44338] = 32'b00000000000000001010001010101100;
assign LUT_3[44339] = 32'b00000000000000010000110110001001;
assign LUT_3[44340] = 32'b00000000000000000101010000111110;
assign LUT_3[44341] = 32'b00000000000000001011111100011011;
assign LUT_3[44342] = 32'b00000000000000000111011000100010;
assign LUT_3[44343] = 32'b00000000000000001110000011111111;
assign LUT_3[44344] = 32'b00000000000000001101011100001110;
assign LUT_3[44345] = 32'b00000000000000010100000111101011;
assign LUT_3[44346] = 32'b00000000000000001111100011110010;
assign LUT_3[44347] = 32'b00000000000000010110001111001111;
assign LUT_3[44348] = 32'b00000000000000001010101010000100;
assign LUT_3[44349] = 32'b00000000000000010001010101100001;
assign LUT_3[44350] = 32'b00000000000000001100110001101000;
assign LUT_3[44351] = 32'b00000000000000010011011101000101;
assign LUT_3[44352] = 32'b00000000000000000011011010010000;
assign LUT_3[44353] = 32'b00000000000000001010000101101101;
assign LUT_3[44354] = 32'b00000000000000000101100001110100;
assign LUT_3[44355] = 32'b00000000000000001100001101010001;
assign LUT_3[44356] = 32'b00000000000000000000101000000110;
assign LUT_3[44357] = 32'b00000000000000000111010011100011;
assign LUT_3[44358] = 32'b00000000000000000010101111101010;
assign LUT_3[44359] = 32'b00000000000000001001011011000111;
assign LUT_3[44360] = 32'b00000000000000001000110011010110;
assign LUT_3[44361] = 32'b00000000000000001111011110110011;
assign LUT_3[44362] = 32'b00000000000000001010111010111010;
assign LUT_3[44363] = 32'b00000000000000010001100110010111;
assign LUT_3[44364] = 32'b00000000000000000110000001001100;
assign LUT_3[44365] = 32'b00000000000000001100101100101001;
assign LUT_3[44366] = 32'b00000000000000001000001000110000;
assign LUT_3[44367] = 32'b00000000000000001110110100001101;
assign LUT_3[44368] = 32'b00000000000000000110101101010011;
assign LUT_3[44369] = 32'b00000000000000001101011000110000;
assign LUT_3[44370] = 32'b00000000000000001000110100110111;
assign LUT_3[44371] = 32'b00000000000000001111100000010100;
assign LUT_3[44372] = 32'b00000000000000000011111011001001;
assign LUT_3[44373] = 32'b00000000000000001010100110100110;
assign LUT_3[44374] = 32'b00000000000000000110000010101101;
assign LUT_3[44375] = 32'b00000000000000001100101110001010;
assign LUT_3[44376] = 32'b00000000000000001100000110011001;
assign LUT_3[44377] = 32'b00000000000000010010110001110110;
assign LUT_3[44378] = 32'b00000000000000001110001101111101;
assign LUT_3[44379] = 32'b00000000000000010100111001011010;
assign LUT_3[44380] = 32'b00000000000000001001010100001111;
assign LUT_3[44381] = 32'b00000000000000001111111111101100;
assign LUT_3[44382] = 32'b00000000000000001011011011110011;
assign LUT_3[44383] = 32'b00000000000000010010000111010000;
assign LUT_3[44384] = 32'b00000000000000000100101000110000;
assign LUT_3[44385] = 32'b00000000000000001011010100001101;
assign LUT_3[44386] = 32'b00000000000000000110110000010100;
assign LUT_3[44387] = 32'b00000000000000001101011011110001;
assign LUT_3[44388] = 32'b00000000000000000001110110100110;
assign LUT_3[44389] = 32'b00000000000000001000100010000011;
assign LUT_3[44390] = 32'b00000000000000000011111110001010;
assign LUT_3[44391] = 32'b00000000000000001010101001100111;
assign LUT_3[44392] = 32'b00000000000000001010000001110110;
assign LUT_3[44393] = 32'b00000000000000010000101101010011;
assign LUT_3[44394] = 32'b00000000000000001100001001011010;
assign LUT_3[44395] = 32'b00000000000000010010110100110111;
assign LUT_3[44396] = 32'b00000000000000000111001111101100;
assign LUT_3[44397] = 32'b00000000000000001101111011001001;
assign LUT_3[44398] = 32'b00000000000000001001010111010000;
assign LUT_3[44399] = 32'b00000000000000010000000010101101;
assign LUT_3[44400] = 32'b00000000000000000111111011110011;
assign LUT_3[44401] = 32'b00000000000000001110100111010000;
assign LUT_3[44402] = 32'b00000000000000001010000011010111;
assign LUT_3[44403] = 32'b00000000000000010000101110110100;
assign LUT_3[44404] = 32'b00000000000000000101001001101001;
assign LUT_3[44405] = 32'b00000000000000001011110101000110;
assign LUT_3[44406] = 32'b00000000000000000111010001001101;
assign LUT_3[44407] = 32'b00000000000000001101111100101010;
assign LUT_3[44408] = 32'b00000000000000001101010100111001;
assign LUT_3[44409] = 32'b00000000000000010100000000010110;
assign LUT_3[44410] = 32'b00000000000000001111011100011101;
assign LUT_3[44411] = 32'b00000000000000010110000111111010;
assign LUT_3[44412] = 32'b00000000000000001010100010101111;
assign LUT_3[44413] = 32'b00000000000000010001001110001100;
assign LUT_3[44414] = 32'b00000000000000001100101010010011;
assign LUT_3[44415] = 32'b00000000000000010011010101110000;
assign LUT_3[44416] = 32'b00000000000000000101101100100011;
assign LUT_3[44417] = 32'b00000000000000001100011000000000;
assign LUT_3[44418] = 32'b00000000000000000111110100000111;
assign LUT_3[44419] = 32'b00000000000000001110011111100100;
assign LUT_3[44420] = 32'b00000000000000000010111010011001;
assign LUT_3[44421] = 32'b00000000000000001001100101110110;
assign LUT_3[44422] = 32'b00000000000000000101000001111101;
assign LUT_3[44423] = 32'b00000000000000001011101101011010;
assign LUT_3[44424] = 32'b00000000000000001011000101101001;
assign LUT_3[44425] = 32'b00000000000000010001110001000110;
assign LUT_3[44426] = 32'b00000000000000001101001101001101;
assign LUT_3[44427] = 32'b00000000000000010011111000101010;
assign LUT_3[44428] = 32'b00000000000000001000010011011111;
assign LUT_3[44429] = 32'b00000000000000001110111110111100;
assign LUT_3[44430] = 32'b00000000000000001010011011000011;
assign LUT_3[44431] = 32'b00000000000000010001000110100000;
assign LUT_3[44432] = 32'b00000000000000001000111111100110;
assign LUT_3[44433] = 32'b00000000000000001111101011000011;
assign LUT_3[44434] = 32'b00000000000000001011000111001010;
assign LUT_3[44435] = 32'b00000000000000010001110010100111;
assign LUT_3[44436] = 32'b00000000000000000110001101011100;
assign LUT_3[44437] = 32'b00000000000000001100111000111001;
assign LUT_3[44438] = 32'b00000000000000001000010101000000;
assign LUT_3[44439] = 32'b00000000000000001111000000011101;
assign LUT_3[44440] = 32'b00000000000000001110011000101100;
assign LUT_3[44441] = 32'b00000000000000010101000100001001;
assign LUT_3[44442] = 32'b00000000000000010000100000010000;
assign LUT_3[44443] = 32'b00000000000000010111001011101101;
assign LUT_3[44444] = 32'b00000000000000001011100110100010;
assign LUT_3[44445] = 32'b00000000000000010010010001111111;
assign LUT_3[44446] = 32'b00000000000000001101101110000110;
assign LUT_3[44447] = 32'b00000000000000010100011001100011;
assign LUT_3[44448] = 32'b00000000000000000110111011000011;
assign LUT_3[44449] = 32'b00000000000000001101100110100000;
assign LUT_3[44450] = 32'b00000000000000001001000010100111;
assign LUT_3[44451] = 32'b00000000000000001111101110000100;
assign LUT_3[44452] = 32'b00000000000000000100001000111001;
assign LUT_3[44453] = 32'b00000000000000001010110100010110;
assign LUT_3[44454] = 32'b00000000000000000110010000011101;
assign LUT_3[44455] = 32'b00000000000000001100111011111010;
assign LUT_3[44456] = 32'b00000000000000001100010100001001;
assign LUT_3[44457] = 32'b00000000000000010010111111100110;
assign LUT_3[44458] = 32'b00000000000000001110011011101101;
assign LUT_3[44459] = 32'b00000000000000010101000111001010;
assign LUT_3[44460] = 32'b00000000000000001001100001111111;
assign LUT_3[44461] = 32'b00000000000000010000001101011100;
assign LUT_3[44462] = 32'b00000000000000001011101001100011;
assign LUT_3[44463] = 32'b00000000000000010010010101000000;
assign LUT_3[44464] = 32'b00000000000000001010001110000110;
assign LUT_3[44465] = 32'b00000000000000010000111001100011;
assign LUT_3[44466] = 32'b00000000000000001100010101101010;
assign LUT_3[44467] = 32'b00000000000000010011000001000111;
assign LUT_3[44468] = 32'b00000000000000000111011011111100;
assign LUT_3[44469] = 32'b00000000000000001110000111011001;
assign LUT_3[44470] = 32'b00000000000000001001100011100000;
assign LUT_3[44471] = 32'b00000000000000010000001110111101;
assign LUT_3[44472] = 32'b00000000000000001111100111001100;
assign LUT_3[44473] = 32'b00000000000000010110010010101001;
assign LUT_3[44474] = 32'b00000000000000010001101110110000;
assign LUT_3[44475] = 32'b00000000000000011000011010001101;
assign LUT_3[44476] = 32'b00000000000000001100110101000010;
assign LUT_3[44477] = 32'b00000000000000010011100000011111;
assign LUT_3[44478] = 32'b00000000000000001110111100100110;
assign LUT_3[44479] = 32'b00000000000000010101101000000011;
assign LUT_3[44480] = 32'b00000000000000000101100101001110;
assign LUT_3[44481] = 32'b00000000000000001100010000101011;
assign LUT_3[44482] = 32'b00000000000000000111101100110010;
assign LUT_3[44483] = 32'b00000000000000001110011000001111;
assign LUT_3[44484] = 32'b00000000000000000010110011000100;
assign LUT_3[44485] = 32'b00000000000000001001011110100001;
assign LUT_3[44486] = 32'b00000000000000000100111010101000;
assign LUT_3[44487] = 32'b00000000000000001011100110000101;
assign LUT_3[44488] = 32'b00000000000000001010111110010100;
assign LUT_3[44489] = 32'b00000000000000010001101001110001;
assign LUT_3[44490] = 32'b00000000000000001101000101111000;
assign LUT_3[44491] = 32'b00000000000000010011110001010101;
assign LUT_3[44492] = 32'b00000000000000001000001100001010;
assign LUT_3[44493] = 32'b00000000000000001110110111100111;
assign LUT_3[44494] = 32'b00000000000000001010010011101110;
assign LUT_3[44495] = 32'b00000000000000010000111111001011;
assign LUT_3[44496] = 32'b00000000000000001000111000010001;
assign LUT_3[44497] = 32'b00000000000000001111100011101110;
assign LUT_3[44498] = 32'b00000000000000001010111111110101;
assign LUT_3[44499] = 32'b00000000000000010001101011010010;
assign LUT_3[44500] = 32'b00000000000000000110000110000111;
assign LUT_3[44501] = 32'b00000000000000001100110001100100;
assign LUT_3[44502] = 32'b00000000000000001000001101101011;
assign LUT_3[44503] = 32'b00000000000000001110111001001000;
assign LUT_3[44504] = 32'b00000000000000001110010001010111;
assign LUT_3[44505] = 32'b00000000000000010100111100110100;
assign LUT_3[44506] = 32'b00000000000000010000011000111011;
assign LUT_3[44507] = 32'b00000000000000010111000100011000;
assign LUT_3[44508] = 32'b00000000000000001011011111001101;
assign LUT_3[44509] = 32'b00000000000000010010001010101010;
assign LUT_3[44510] = 32'b00000000000000001101100110110001;
assign LUT_3[44511] = 32'b00000000000000010100010010001110;
assign LUT_3[44512] = 32'b00000000000000000110110011101110;
assign LUT_3[44513] = 32'b00000000000000001101011111001011;
assign LUT_3[44514] = 32'b00000000000000001000111011010010;
assign LUT_3[44515] = 32'b00000000000000001111100110101111;
assign LUT_3[44516] = 32'b00000000000000000100000001100100;
assign LUT_3[44517] = 32'b00000000000000001010101101000001;
assign LUT_3[44518] = 32'b00000000000000000110001001001000;
assign LUT_3[44519] = 32'b00000000000000001100110100100101;
assign LUT_3[44520] = 32'b00000000000000001100001100110100;
assign LUT_3[44521] = 32'b00000000000000010010111000010001;
assign LUT_3[44522] = 32'b00000000000000001110010100011000;
assign LUT_3[44523] = 32'b00000000000000010100111111110101;
assign LUT_3[44524] = 32'b00000000000000001001011010101010;
assign LUT_3[44525] = 32'b00000000000000010000000110000111;
assign LUT_3[44526] = 32'b00000000000000001011100010001110;
assign LUT_3[44527] = 32'b00000000000000010010001101101011;
assign LUT_3[44528] = 32'b00000000000000001010000110110001;
assign LUT_3[44529] = 32'b00000000000000010000110010001110;
assign LUT_3[44530] = 32'b00000000000000001100001110010101;
assign LUT_3[44531] = 32'b00000000000000010010111001110010;
assign LUT_3[44532] = 32'b00000000000000000111010100100111;
assign LUT_3[44533] = 32'b00000000000000001110000000000100;
assign LUT_3[44534] = 32'b00000000000000001001011100001011;
assign LUT_3[44535] = 32'b00000000000000010000000111101000;
assign LUT_3[44536] = 32'b00000000000000001111011111110111;
assign LUT_3[44537] = 32'b00000000000000010110001011010100;
assign LUT_3[44538] = 32'b00000000000000010001100111011011;
assign LUT_3[44539] = 32'b00000000000000011000010010111000;
assign LUT_3[44540] = 32'b00000000000000001100101101101101;
assign LUT_3[44541] = 32'b00000000000000010011011001001010;
assign LUT_3[44542] = 32'b00000000000000001110110101010001;
assign LUT_3[44543] = 32'b00000000000000010101100000101110;
assign LUT_3[44544] = 32'b00000000000000001010100111010000;
assign LUT_3[44545] = 32'b00000000000000010001010010101101;
assign LUT_3[44546] = 32'b00000000000000001100101110110100;
assign LUT_3[44547] = 32'b00000000000000010011011010010001;
assign LUT_3[44548] = 32'b00000000000000000111110101000110;
assign LUT_3[44549] = 32'b00000000000000001110100000100011;
assign LUT_3[44550] = 32'b00000000000000001001111100101010;
assign LUT_3[44551] = 32'b00000000000000010000101000000111;
assign LUT_3[44552] = 32'b00000000000000010000000000010110;
assign LUT_3[44553] = 32'b00000000000000010110101011110011;
assign LUT_3[44554] = 32'b00000000000000010010000111111010;
assign LUT_3[44555] = 32'b00000000000000011000110011010111;
assign LUT_3[44556] = 32'b00000000000000001101001110001100;
assign LUT_3[44557] = 32'b00000000000000010011111001101001;
assign LUT_3[44558] = 32'b00000000000000001111010101110000;
assign LUT_3[44559] = 32'b00000000000000010110000001001101;
assign LUT_3[44560] = 32'b00000000000000001101111010010011;
assign LUT_3[44561] = 32'b00000000000000010100100101110000;
assign LUT_3[44562] = 32'b00000000000000010000000001110111;
assign LUT_3[44563] = 32'b00000000000000010110101101010100;
assign LUT_3[44564] = 32'b00000000000000001011001000001001;
assign LUT_3[44565] = 32'b00000000000000010001110011100110;
assign LUT_3[44566] = 32'b00000000000000001101001111101101;
assign LUT_3[44567] = 32'b00000000000000010011111011001010;
assign LUT_3[44568] = 32'b00000000000000010011010011011001;
assign LUT_3[44569] = 32'b00000000000000011001111110110110;
assign LUT_3[44570] = 32'b00000000000000010101011010111101;
assign LUT_3[44571] = 32'b00000000000000011100000110011010;
assign LUT_3[44572] = 32'b00000000000000010000100001001111;
assign LUT_3[44573] = 32'b00000000000000010111001100101100;
assign LUT_3[44574] = 32'b00000000000000010010101000110011;
assign LUT_3[44575] = 32'b00000000000000011001010100010000;
assign LUT_3[44576] = 32'b00000000000000001011110101110000;
assign LUT_3[44577] = 32'b00000000000000010010100001001101;
assign LUT_3[44578] = 32'b00000000000000001101111101010100;
assign LUT_3[44579] = 32'b00000000000000010100101000110001;
assign LUT_3[44580] = 32'b00000000000000001001000011100110;
assign LUT_3[44581] = 32'b00000000000000001111101111000011;
assign LUT_3[44582] = 32'b00000000000000001011001011001010;
assign LUT_3[44583] = 32'b00000000000000010001110110100111;
assign LUT_3[44584] = 32'b00000000000000010001001110110110;
assign LUT_3[44585] = 32'b00000000000000010111111010010011;
assign LUT_3[44586] = 32'b00000000000000010011010110011010;
assign LUT_3[44587] = 32'b00000000000000011010000001110111;
assign LUT_3[44588] = 32'b00000000000000001110011100101100;
assign LUT_3[44589] = 32'b00000000000000010101001000001001;
assign LUT_3[44590] = 32'b00000000000000010000100100010000;
assign LUT_3[44591] = 32'b00000000000000010111001111101101;
assign LUT_3[44592] = 32'b00000000000000001111001000110011;
assign LUT_3[44593] = 32'b00000000000000010101110100010000;
assign LUT_3[44594] = 32'b00000000000000010001010000010111;
assign LUT_3[44595] = 32'b00000000000000010111111011110100;
assign LUT_3[44596] = 32'b00000000000000001100010110101001;
assign LUT_3[44597] = 32'b00000000000000010011000010000110;
assign LUT_3[44598] = 32'b00000000000000001110011110001101;
assign LUT_3[44599] = 32'b00000000000000010101001001101010;
assign LUT_3[44600] = 32'b00000000000000010100100001111001;
assign LUT_3[44601] = 32'b00000000000000011011001101010110;
assign LUT_3[44602] = 32'b00000000000000010110101001011101;
assign LUT_3[44603] = 32'b00000000000000011101010100111010;
assign LUT_3[44604] = 32'b00000000000000010001101111101111;
assign LUT_3[44605] = 32'b00000000000000011000011011001100;
assign LUT_3[44606] = 32'b00000000000000010011110111010011;
assign LUT_3[44607] = 32'b00000000000000011010100010110000;
assign LUT_3[44608] = 32'b00000000000000001010011111111011;
assign LUT_3[44609] = 32'b00000000000000010001001011011000;
assign LUT_3[44610] = 32'b00000000000000001100100111011111;
assign LUT_3[44611] = 32'b00000000000000010011010010111100;
assign LUT_3[44612] = 32'b00000000000000000111101101110001;
assign LUT_3[44613] = 32'b00000000000000001110011001001110;
assign LUT_3[44614] = 32'b00000000000000001001110101010101;
assign LUT_3[44615] = 32'b00000000000000010000100000110010;
assign LUT_3[44616] = 32'b00000000000000001111111001000001;
assign LUT_3[44617] = 32'b00000000000000010110100100011110;
assign LUT_3[44618] = 32'b00000000000000010010000000100101;
assign LUT_3[44619] = 32'b00000000000000011000101100000010;
assign LUT_3[44620] = 32'b00000000000000001101000110110111;
assign LUT_3[44621] = 32'b00000000000000010011110010010100;
assign LUT_3[44622] = 32'b00000000000000001111001110011011;
assign LUT_3[44623] = 32'b00000000000000010101111001111000;
assign LUT_3[44624] = 32'b00000000000000001101110010111110;
assign LUT_3[44625] = 32'b00000000000000010100011110011011;
assign LUT_3[44626] = 32'b00000000000000001111111010100010;
assign LUT_3[44627] = 32'b00000000000000010110100101111111;
assign LUT_3[44628] = 32'b00000000000000001011000000110100;
assign LUT_3[44629] = 32'b00000000000000010001101100010001;
assign LUT_3[44630] = 32'b00000000000000001101001000011000;
assign LUT_3[44631] = 32'b00000000000000010011110011110101;
assign LUT_3[44632] = 32'b00000000000000010011001100000100;
assign LUT_3[44633] = 32'b00000000000000011001110111100001;
assign LUT_3[44634] = 32'b00000000000000010101010011101000;
assign LUT_3[44635] = 32'b00000000000000011011111111000101;
assign LUT_3[44636] = 32'b00000000000000010000011001111010;
assign LUT_3[44637] = 32'b00000000000000010111000101010111;
assign LUT_3[44638] = 32'b00000000000000010010100001011110;
assign LUT_3[44639] = 32'b00000000000000011001001100111011;
assign LUT_3[44640] = 32'b00000000000000001011101110011011;
assign LUT_3[44641] = 32'b00000000000000010010011001111000;
assign LUT_3[44642] = 32'b00000000000000001101110101111111;
assign LUT_3[44643] = 32'b00000000000000010100100001011100;
assign LUT_3[44644] = 32'b00000000000000001000111100010001;
assign LUT_3[44645] = 32'b00000000000000001111100111101110;
assign LUT_3[44646] = 32'b00000000000000001011000011110101;
assign LUT_3[44647] = 32'b00000000000000010001101111010010;
assign LUT_3[44648] = 32'b00000000000000010001000111100001;
assign LUT_3[44649] = 32'b00000000000000010111110010111110;
assign LUT_3[44650] = 32'b00000000000000010011001111000101;
assign LUT_3[44651] = 32'b00000000000000011001111010100010;
assign LUT_3[44652] = 32'b00000000000000001110010101010111;
assign LUT_3[44653] = 32'b00000000000000010101000000110100;
assign LUT_3[44654] = 32'b00000000000000010000011100111011;
assign LUT_3[44655] = 32'b00000000000000010111001000011000;
assign LUT_3[44656] = 32'b00000000000000001111000001011110;
assign LUT_3[44657] = 32'b00000000000000010101101100111011;
assign LUT_3[44658] = 32'b00000000000000010001001001000010;
assign LUT_3[44659] = 32'b00000000000000010111110100011111;
assign LUT_3[44660] = 32'b00000000000000001100001111010100;
assign LUT_3[44661] = 32'b00000000000000010010111010110001;
assign LUT_3[44662] = 32'b00000000000000001110010110111000;
assign LUT_3[44663] = 32'b00000000000000010101000010010101;
assign LUT_3[44664] = 32'b00000000000000010100011010100100;
assign LUT_3[44665] = 32'b00000000000000011011000110000001;
assign LUT_3[44666] = 32'b00000000000000010110100010001000;
assign LUT_3[44667] = 32'b00000000000000011101001101100101;
assign LUT_3[44668] = 32'b00000000000000010001101000011010;
assign LUT_3[44669] = 32'b00000000000000011000010011110111;
assign LUT_3[44670] = 32'b00000000000000010011101111111110;
assign LUT_3[44671] = 32'b00000000000000011010011011011011;
assign LUT_3[44672] = 32'b00000000000000001100110010001110;
assign LUT_3[44673] = 32'b00000000000000010011011101101011;
assign LUT_3[44674] = 32'b00000000000000001110111001110010;
assign LUT_3[44675] = 32'b00000000000000010101100101001111;
assign LUT_3[44676] = 32'b00000000000000001010000000000100;
assign LUT_3[44677] = 32'b00000000000000010000101011100001;
assign LUT_3[44678] = 32'b00000000000000001100000111101000;
assign LUT_3[44679] = 32'b00000000000000010010110011000101;
assign LUT_3[44680] = 32'b00000000000000010010001011010100;
assign LUT_3[44681] = 32'b00000000000000011000110110110001;
assign LUT_3[44682] = 32'b00000000000000010100010010111000;
assign LUT_3[44683] = 32'b00000000000000011010111110010101;
assign LUT_3[44684] = 32'b00000000000000001111011001001010;
assign LUT_3[44685] = 32'b00000000000000010110000100100111;
assign LUT_3[44686] = 32'b00000000000000010001100000101110;
assign LUT_3[44687] = 32'b00000000000000011000001100001011;
assign LUT_3[44688] = 32'b00000000000000010000000101010001;
assign LUT_3[44689] = 32'b00000000000000010110110000101110;
assign LUT_3[44690] = 32'b00000000000000010010001100110101;
assign LUT_3[44691] = 32'b00000000000000011000111000010010;
assign LUT_3[44692] = 32'b00000000000000001101010011000111;
assign LUT_3[44693] = 32'b00000000000000010011111110100100;
assign LUT_3[44694] = 32'b00000000000000001111011010101011;
assign LUT_3[44695] = 32'b00000000000000010110000110001000;
assign LUT_3[44696] = 32'b00000000000000010101011110010111;
assign LUT_3[44697] = 32'b00000000000000011100001001110100;
assign LUT_3[44698] = 32'b00000000000000010111100101111011;
assign LUT_3[44699] = 32'b00000000000000011110010001011000;
assign LUT_3[44700] = 32'b00000000000000010010101100001101;
assign LUT_3[44701] = 32'b00000000000000011001010111101010;
assign LUT_3[44702] = 32'b00000000000000010100110011110001;
assign LUT_3[44703] = 32'b00000000000000011011011111001110;
assign LUT_3[44704] = 32'b00000000000000001110000000101110;
assign LUT_3[44705] = 32'b00000000000000010100101100001011;
assign LUT_3[44706] = 32'b00000000000000010000001000010010;
assign LUT_3[44707] = 32'b00000000000000010110110011101111;
assign LUT_3[44708] = 32'b00000000000000001011001110100100;
assign LUT_3[44709] = 32'b00000000000000010001111010000001;
assign LUT_3[44710] = 32'b00000000000000001101010110001000;
assign LUT_3[44711] = 32'b00000000000000010100000001100101;
assign LUT_3[44712] = 32'b00000000000000010011011001110100;
assign LUT_3[44713] = 32'b00000000000000011010000101010001;
assign LUT_3[44714] = 32'b00000000000000010101100001011000;
assign LUT_3[44715] = 32'b00000000000000011100001100110101;
assign LUT_3[44716] = 32'b00000000000000010000100111101010;
assign LUT_3[44717] = 32'b00000000000000010111010011000111;
assign LUT_3[44718] = 32'b00000000000000010010101111001110;
assign LUT_3[44719] = 32'b00000000000000011001011010101011;
assign LUT_3[44720] = 32'b00000000000000010001010011110001;
assign LUT_3[44721] = 32'b00000000000000010111111111001110;
assign LUT_3[44722] = 32'b00000000000000010011011011010101;
assign LUT_3[44723] = 32'b00000000000000011010000110110010;
assign LUT_3[44724] = 32'b00000000000000001110100001100111;
assign LUT_3[44725] = 32'b00000000000000010101001101000100;
assign LUT_3[44726] = 32'b00000000000000010000101001001011;
assign LUT_3[44727] = 32'b00000000000000010111010100101000;
assign LUT_3[44728] = 32'b00000000000000010110101100110111;
assign LUT_3[44729] = 32'b00000000000000011101011000010100;
assign LUT_3[44730] = 32'b00000000000000011000110100011011;
assign LUT_3[44731] = 32'b00000000000000011111011111111000;
assign LUT_3[44732] = 32'b00000000000000010011111010101101;
assign LUT_3[44733] = 32'b00000000000000011010100110001010;
assign LUT_3[44734] = 32'b00000000000000010110000010010001;
assign LUT_3[44735] = 32'b00000000000000011100101101101110;
assign LUT_3[44736] = 32'b00000000000000001100101010111001;
assign LUT_3[44737] = 32'b00000000000000010011010110010110;
assign LUT_3[44738] = 32'b00000000000000001110110010011101;
assign LUT_3[44739] = 32'b00000000000000010101011101111010;
assign LUT_3[44740] = 32'b00000000000000001001111000101111;
assign LUT_3[44741] = 32'b00000000000000010000100100001100;
assign LUT_3[44742] = 32'b00000000000000001100000000010011;
assign LUT_3[44743] = 32'b00000000000000010010101011110000;
assign LUT_3[44744] = 32'b00000000000000010010000011111111;
assign LUT_3[44745] = 32'b00000000000000011000101111011100;
assign LUT_3[44746] = 32'b00000000000000010100001011100011;
assign LUT_3[44747] = 32'b00000000000000011010110111000000;
assign LUT_3[44748] = 32'b00000000000000001111010001110101;
assign LUT_3[44749] = 32'b00000000000000010101111101010010;
assign LUT_3[44750] = 32'b00000000000000010001011001011001;
assign LUT_3[44751] = 32'b00000000000000011000000100110110;
assign LUT_3[44752] = 32'b00000000000000001111111101111100;
assign LUT_3[44753] = 32'b00000000000000010110101001011001;
assign LUT_3[44754] = 32'b00000000000000010010000101100000;
assign LUT_3[44755] = 32'b00000000000000011000110000111101;
assign LUT_3[44756] = 32'b00000000000000001101001011110010;
assign LUT_3[44757] = 32'b00000000000000010011110111001111;
assign LUT_3[44758] = 32'b00000000000000001111010011010110;
assign LUT_3[44759] = 32'b00000000000000010101111110110011;
assign LUT_3[44760] = 32'b00000000000000010101010111000010;
assign LUT_3[44761] = 32'b00000000000000011100000010011111;
assign LUT_3[44762] = 32'b00000000000000010111011110100110;
assign LUT_3[44763] = 32'b00000000000000011110001010000011;
assign LUT_3[44764] = 32'b00000000000000010010100100111000;
assign LUT_3[44765] = 32'b00000000000000011001010000010101;
assign LUT_3[44766] = 32'b00000000000000010100101100011100;
assign LUT_3[44767] = 32'b00000000000000011011010111111001;
assign LUT_3[44768] = 32'b00000000000000001101111001011001;
assign LUT_3[44769] = 32'b00000000000000010100100100110110;
assign LUT_3[44770] = 32'b00000000000000010000000000111101;
assign LUT_3[44771] = 32'b00000000000000010110101100011010;
assign LUT_3[44772] = 32'b00000000000000001011000111001111;
assign LUT_3[44773] = 32'b00000000000000010001110010101100;
assign LUT_3[44774] = 32'b00000000000000001101001110110011;
assign LUT_3[44775] = 32'b00000000000000010011111010010000;
assign LUT_3[44776] = 32'b00000000000000010011010010011111;
assign LUT_3[44777] = 32'b00000000000000011001111101111100;
assign LUT_3[44778] = 32'b00000000000000010101011010000011;
assign LUT_3[44779] = 32'b00000000000000011100000101100000;
assign LUT_3[44780] = 32'b00000000000000010000100000010101;
assign LUT_3[44781] = 32'b00000000000000010111001011110010;
assign LUT_3[44782] = 32'b00000000000000010010100111111001;
assign LUT_3[44783] = 32'b00000000000000011001010011010110;
assign LUT_3[44784] = 32'b00000000000000010001001100011100;
assign LUT_3[44785] = 32'b00000000000000010111110111111001;
assign LUT_3[44786] = 32'b00000000000000010011010100000000;
assign LUT_3[44787] = 32'b00000000000000011001111111011101;
assign LUT_3[44788] = 32'b00000000000000001110011010010010;
assign LUT_3[44789] = 32'b00000000000000010101000101101111;
assign LUT_3[44790] = 32'b00000000000000010000100001110110;
assign LUT_3[44791] = 32'b00000000000000010111001101010011;
assign LUT_3[44792] = 32'b00000000000000010110100101100010;
assign LUT_3[44793] = 32'b00000000000000011101010000111111;
assign LUT_3[44794] = 32'b00000000000000011000101101000110;
assign LUT_3[44795] = 32'b00000000000000011111011000100011;
assign LUT_3[44796] = 32'b00000000000000010011110011011000;
assign LUT_3[44797] = 32'b00000000000000011010011110110101;
assign LUT_3[44798] = 32'b00000000000000010101111010111100;
assign LUT_3[44799] = 32'b00000000000000011100100110011001;
assign LUT_3[44800] = 32'b00000000000000000110110110110001;
assign LUT_3[44801] = 32'b00000000000000001101100010001110;
assign LUT_3[44802] = 32'b00000000000000001000111110010101;
assign LUT_3[44803] = 32'b00000000000000001111101001110010;
assign LUT_3[44804] = 32'b00000000000000000100000100100111;
assign LUT_3[44805] = 32'b00000000000000001010110000000100;
assign LUT_3[44806] = 32'b00000000000000000110001100001011;
assign LUT_3[44807] = 32'b00000000000000001100110111101000;
assign LUT_3[44808] = 32'b00000000000000001100001111110111;
assign LUT_3[44809] = 32'b00000000000000010010111011010100;
assign LUT_3[44810] = 32'b00000000000000001110010111011011;
assign LUT_3[44811] = 32'b00000000000000010101000010111000;
assign LUT_3[44812] = 32'b00000000000000001001011101101101;
assign LUT_3[44813] = 32'b00000000000000010000001001001010;
assign LUT_3[44814] = 32'b00000000000000001011100101010001;
assign LUT_3[44815] = 32'b00000000000000010010010000101110;
assign LUT_3[44816] = 32'b00000000000000001010001001110100;
assign LUT_3[44817] = 32'b00000000000000010000110101010001;
assign LUT_3[44818] = 32'b00000000000000001100010001011000;
assign LUT_3[44819] = 32'b00000000000000010010111100110101;
assign LUT_3[44820] = 32'b00000000000000000111010111101010;
assign LUT_3[44821] = 32'b00000000000000001110000011000111;
assign LUT_3[44822] = 32'b00000000000000001001011111001110;
assign LUT_3[44823] = 32'b00000000000000010000001010101011;
assign LUT_3[44824] = 32'b00000000000000001111100010111010;
assign LUT_3[44825] = 32'b00000000000000010110001110010111;
assign LUT_3[44826] = 32'b00000000000000010001101010011110;
assign LUT_3[44827] = 32'b00000000000000011000010101111011;
assign LUT_3[44828] = 32'b00000000000000001100110000110000;
assign LUT_3[44829] = 32'b00000000000000010011011100001101;
assign LUT_3[44830] = 32'b00000000000000001110111000010100;
assign LUT_3[44831] = 32'b00000000000000010101100011110001;
assign LUT_3[44832] = 32'b00000000000000001000000101010001;
assign LUT_3[44833] = 32'b00000000000000001110110000101110;
assign LUT_3[44834] = 32'b00000000000000001010001100110101;
assign LUT_3[44835] = 32'b00000000000000010000111000010010;
assign LUT_3[44836] = 32'b00000000000000000101010011000111;
assign LUT_3[44837] = 32'b00000000000000001011111110100100;
assign LUT_3[44838] = 32'b00000000000000000111011010101011;
assign LUT_3[44839] = 32'b00000000000000001110000110001000;
assign LUT_3[44840] = 32'b00000000000000001101011110010111;
assign LUT_3[44841] = 32'b00000000000000010100001001110100;
assign LUT_3[44842] = 32'b00000000000000001111100101111011;
assign LUT_3[44843] = 32'b00000000000000010110010001011000;
assign LUT_3[44844] = 32'b00000000000000001010101100001101;
assign LUT_3[44845] = 32'b00000000000000010001010111101010;
assign LUT_3[44846] = 32'b00000000000000001100110011110001;
assign LUT_3[44847] = 32'b00000000000000010011011111001110;
assign LUT_3[44848] = 32'b00000000000000001011011000010100;
assign LUT_3[44849] = 32'b00000000000000010010000011110001;
assign LUT_3[44850] = 32'b00000000000000001101011111111000;
assign LUT_3[44851] = 32'b00000000000000010100001011010101;
assign LUT_3[44852] = 32'b00000000000000001000100110001010;
assign LUT_3[44853] = 32'b00000000000000001111010001100111;
assign LUT_3[44854] = 32'b00000000000000001010101101101110;
assign LUT_3[44855] = 32'b00000000000000010001011001001011;
assign LUT_3[44856] = 32'b00000000000000010000110001011010;
assign LUT_3[44857] = 32'b00000000000000010111011100110111;
assign LUT_3[44858] = 32'b00000000000000010010111000111110;
assign LUT_3[44859] = 32'b00000000000000011001100100011011;
assign LUT_3[44860] = 32'b00000000000000001101111111010000;
assign LUT_3[44861] = 32'b00000000000000010100101010101101;
assign LUT_3[44862] = 32'b00000000000000010000000110110100;
assign LUT_3[44863] = 32'b00000000000000010110110010010001;
assign LUT_3[44864] = 32'b00000000000000000110101111011100;
assign LUT_3[44865] = 32'b00000000000000001101011010111001;
assign LUT_3[44866] = 32'b00000000000000001000110111000000;
assign LUT_3[44867] = 32'b00000000000000001111100010011101;
assign LUT_3[44868] = 32'b00000000000000000011111101010010;
assign LUT_3[44869] = 32'b00000000000000001010101000101111;
assign LUT_3[44870] = 32'b00000000000000000110000100110110;
assign LUT_3[44871] = 32'b00000000000000001100110000010011;
assign LUT_3[44872] = 32'b00000000000000001100001000100010;
assign LUT_3[44873] = 32'b00000000000000010010110011111111;
assign LUT_3[44874] = 32'b00000000000000001110010000000110;
assign LUT_3[44875] = 32'b00000000000000010100111011100011;
assign LUT_3[44876] = 32'b00000000000000001001010110011000;
assign LUT_3[44877] = 32'b00000000000000010000000001110101;
assign LUT_3[44878] = 32'b00000000000000001011011101111100;
assign LUT_3[44879] = 32'b00000000000000010010001001011001;
assign LUT_3[44880] = 32'b00000000000000001010000010011111;
assign LUT_3[44881] = 32'b00000000000000010000101101111100;
assign LUT_3[44882] = 32'b00000000000000001100001010000011;
assign LUT_3[44883] = 32'b00000000000000010010110101100000;
assign LUT_3[44884] = 32'b00000000000000000111010000010101;
assign LUT_3[44885] = 32'b00000000000000001101111011110010;
assign LUT_3[44886] = 32'b00000000000000001001010111111001;
assign LUT_3[44887] = 32'b00000000000000010000000011010110;
assign LUT_3[44888] = 32'b00000000000000001111011011100101;
assign LUT_3[44889] = 32'b00000000000000010110000111000010;
assign LUT_3[44890] = 32'b00000000000000010001100011001001;
assign LUT_3[44891] = 32'b00000000000000011000001110100110;
assign LUT_3[44892] = 32'b00000000000000001100101001011011;
assign LUT_3[44893] = 32'b00000000000000010011010100111000;
assign LUT_3[44894] = 32'b00000000000000001110110000111111;
assign LUT_3[44895] = 32'b00000000000000010101011100011100;
assign LUT_3[44896] = 32'b00000000000000000111111101111100;
assign LUT_3[44897] = 32'b00000000000000001110101001011001;
assign LUT_3[44898] = 32'b00000000000000001010000101100000;
assign LUT_3[44899] = 32'b00000000000000010000110000111101;
assign LUT_3[44900] = 32'b00000000000000000101001011110010;
assign LUT_3[44901] = 32'b00000000000000001011110111001111;
assign LUT_3[44902] = 32'b00000000000000000111010011010110;
assign LUT_3[44903] = 32'b00000000000000001101111110110011;
assign LUT_3[44904] = 32'b00000000000000001101010111000010;
assign LUT_3[44905] = 32'b00000000000000010100000010011111;
assign LUT_3[44906] = 32'b00000000000000001111011110100110;
assign LUT_3[44907] = 32'b00000000000000010110001010000011;
assign LUT_3[44908] = 32'b00000000000000001010100100111000;
assign LUT_3[44909] = 32'b00000000000000010001010000010101;
assign LUT_3[44910] = 32'b00000000000000001100101100011100;
assign LUT_3[44911] = 32'b00000000000000010011010111111001;
assign LUT_3[44912] = 32'b00000000000000001011010000111111;
assign LUT_3[44913] = 32'b00000000000000010001111100011100;
assign LUT_3[44914] = 32'b00000000000000001101011000100011;
assign LUT_3[44915] = 32'b00000000000000010100000100000000;
assign LUT_3[44916] = 32'b00000000000000001000011110110101;
assign LUT_3[44917] = 32'b00000000000000001111001010010010;
assign LUT_3[44918] = 32'b00000000000000001010100110011001;
assign LUT_3[44919] = 32'b00000000000000010001010001110110;
assign LUT_3[44920] = 32'b00000000000000010000101010000101;
assign LUT_3[44921] = 32'b00000000000000010111010101100010;
assign LUT_3[44922] = 32'b00000000000000010010110001101001;
assign LUT_3[44923] = 32'b00000000000000011001011101000110;
assign LUT_3[44924] = 32'b00000000000000001101110111111011;
assign LUT_3[44925] = 32'b00000000000000010100100011011000;
assign LUT_3[44926] = 32'b00000000000000001111111111011111;
assign LUT_3[44927] = 32'b00000000000000010110101010111100;
assign LUT_3[44928] = 32'b00000000000000001001000001101111;
assign LUT_3[44929] = 32'b00000000000000001111101101001100;
assign LUT_3[44930] = 32'b00000000000000001011001001010011;
assign LUT_3[44931] = 32'b00000000000000010001110100110000;
assign LUT_3[44932] = 32'b00000000000000000110001111100101;
assign LUT_3[44933] = 32'b00000000000000001100111011000010;
assign LUT_3[44934] = 32'b00000000000000001000010111001001;
assign LUT_3[44935] = 32'b00000000000000001111000010100110;
assign LUT_3[44936] = 32'b00000000000000001110011010110101;
assign LUT_3[44937] = 32'b00000000000000010101000110010010;
assign LUT_3[44938] = 32'b00000000000000010000100010011001;
assign LUT_3[44939] = 32'b00000000000000010111001101110110;
assign LUT_3[44940] = 32'b00000000000000001011101000101011;
assign LUT_3[44941] = 32'b00000000000000010010010100001000;
assign LUT_3[44942] = 32'b00000000000000001101110000001111;
assign LUT_3[44943] = 32'b00000000000000010100011011101100;
assign LUT_3[44944] = 32'b00000000000000001100010100110010;
assign LUT_3[44945] = 32'b00000000000000010011000000001111;
assign LUT_3[44946] = 32'b00000000000000001110011100010110;
assign LUT_3[44947] = 32'b00000000000000010101000111110011;
assign LUT_3[44948] = 32'b00000000000000001001100010101000;
assign LUT_3[44949] = 32'b00000000000000010000001110000101;
assign LUT_3[44950] = 32'b00000000000000001011101010001100;
assign LUT_3[44951] = 32'b00000000000000010010010101101001;
assign LUT_3[44952] = 32'b00000000000000010001101101111000;
assign LUT_3[44953] = 32'b00000000000000011000011001010101;
assign LUT_3[44954] = 32'b00000000000000010011110101011100;
assign LUT_3[44955] = 32'b00000000000000011010100000111001;
assign LUT_3[44956] = 32'b00000000000000001110111011101110;
assign LUT_3[44957] = 32'b00000000000000010101100111001011;
assign LUT_3[44958] = 32'b00000000000000010001000011010010;
assign LUT_3[44959] = 32'b00000000000000010111101110101111;
assign LUT_3[44960] = 32'b00000000000000001010010000001111;
assign LUT_3[44961] = 32'b00000000000000010000111011101100;
assign LUT_3[44962] = 32'b00000000000000001100010111110011;
assign LUT_3[44963] = 32'b00000000000000010011000011010000;
assign LUT_3[44964] = 32'b00000000000000000111011110000101;
assign LUT_3[44965] = 32'b00000000000000001110001001100010;
assign LUT_3[44966] = 32'b00000000000000001001100101101001;
assign LUT_3[44967] = 32'b00000000000000010000010001000110;
assign LUT_3[44968] = 32'b00000000000000001111101001010101;
assign LUT_3[44969] = 32'b00000000000000010110010100110010;
assign LUT_3[44970] = 32'b00000000000000010001110000111001;
assign LUT_3[44971] = 32'b00000000000000011000011100010110;
assign LUT_3[44972] = 32'b00000000000000001100110111001011;
assign LUT_3[44973] = 32'b00000000000000010011100010101000;
assign LUT_3[44974] = 32'b00000000000000001110111110101111;
assign LUT_3[44975] = 32'b00000000000000010101101010001100;
assign LUT_3[44976] = 32'b00000000000000001101100011010010;
assign LUT_3[44977] = 32'b00000000000000010100001110101111;
assign LUT_3[44978] = 32'b00000000000000001111101010110110;
assign LUT_3[44979] = 32'b00000000000000010110010110010011;
assign LUT_3[44980] = 32'b00000000000000001010110001001000;
assign LUT_3[44981] = 32'b00000000000000010001011100100101;
assign LUT_3[44982] = 32'b00000000000000001100111000101100;
assign LUT_3[44983] = 32'b00000000000000010011100100001001;
assign LUT_3[44984] = 32'b00000000000000010010111100011000;
assign LUT_3[44985] = 32'b00000000000000011001100111110101;
assign LUT_3[44986] = 32'b00000000000000010101000011111100;
assign LUT_3[44987] = 32'b00000000000000011011101111011001;
assign LUT_3[44988] = 32'b00000000000000010000001010001110;
assign LUT_3[44989] = 32'b00000000000000010110110101101011;
assign LUT_3[44990] = 32'b00000000000000010010010001110010;
assign LUT_3[44991] = 32'b00000000000000011000111101001111;
assign LUT_3[44992] = 32'b00000000000000001000111010011010;
assign LUT_3[44993] = 32'b00000000000000001111100101110111;
assign LUT_3[44994] = 32'b00000000000000001011000001111110;
assign LUT_3[44995] = 32'b00000000000000010001101101011011;
assign LUT_3[44996] = 32'b00000000000000000110001000010000;
assign LUT_3[44997] = 32'b00000000000000001100110011101101;
assign LUT_3[44998] = 32'b00000000000000001000001111110100;
assign LUT_3[44999] = 32'b00000000000000001110111011010001;
assign LUT_3[45000] = 32'b00000000000000001110010011100000;
assign LUT_3[45001] = 32'b00000000000000010100111110111101;
assign LUT_3[45002] = 32'b00000000000000010000011011000100;
assign LUT_3[45003] = 32'b00000000000000010111000110100001;
assign LUT_3[45004] = 32'b00000000000000001011100001010110;
assign LUT_3[45005] = 32'b00000000000000010010001100110011;
assign LUT_3[45006] = 32'b00000000000000001101101000111010;
assign LUT_3[45007] = 32'b00000000000000010100010100010111;
assign LUT_3[45008] = 32'b00000000000000001100001101011101;
assign LUT_3[45009] = 32'b00000000000000010010111000111010;
assign LUT_3[45010] = 32'b00000000000000001110010101000001;
assign LUT_3[45011] = 32'b00000000000000010101000000011110;
assign LUT_3[45012] = 32'b00000000000000001001011011010011;
assign LUT_3[45013] = 32'b00000000000000010000000110110000;
assign LUT_3[45014] = 32'b00000000000000001011100010110111;
assign LUT_3[45015] = 32'b00000000000000010010001110010100;
assign LUT_3[45016] = 32'b00000000000000010001100110100011;
assign LUT_3[45017] = 32'b00000000000000011000010010000000;
assign LUT_3[45018] = 32'b00000000000000010011101110000111;
assign LUT_3[45019] = 32'b00000000000000011010011001100100;
assign LUT_3[45020] = 32'b00000000000000001110110100011001;
assign LUT_3[45021] = 32'b00000000000000010101011111110110;
assign LUT_3[45022] = 32'b00000000000000010000111011111101;
assign LUT_3[45023] = 32'b00000000000000010111100111011010;
assign LUT_3[45024] = 32'b00000000000000001010001000111010;
assign LUT_3[45025] = 32'b00000000000000010000110100010111;
assign LUT_3[45026] = 32'b00000000000000001100010000011110;
assign LUT_3[45027] = 32'b00000000000000010010111011111011;
assign LUT_3[45028] = 32'b00000000000000000111010110110000;
assign LUT_3[45029] = 32'b00000000000000001110000010001101;
assign LUT_3[45030] = 32'b00000000000000001001011110010100;
assign LUT_3[45031] = 32'b00000000000000010000001001110001;
assign LUT_3[45032] = 32'b00000000000000001111100010000000;
assign LUT_3[45033] = 32'b00000000000000010110001101011101;
assign LUT_3[45034] = 32'b00000000000000010001101001100100;
assign LUT_3[45035] = 32'b00000000000000011000010101000001;
assign LUT_3[45036] = 32'b00000000000000001100101111110110;
assign LUT_3[45037] = 32'b00000000000000010011011011010011;
assign LUT_3[45038] = 32'b00000000000000001110110111011010;
assign LUT_3[45039] = 32'b00000000000000010101100010110111;
assign LUT_3[45040] = 32'b00000000000000001101011011111101;
assign LUT_3[45041] = 32'b00000000000000010100000111011010;
assign LUT_3[45042] = 32'b00000000000000001111100011100001;
assign LUT_3[45043] = 32'b00000000000000010110001110111110;
assign LUT_3[45044] = 32'b00000000000000001010101001110011;
assign LUT_3[45045] = 32'b00000000000000010001010101010000;
assign LUT_3[45046] = 32'b00000000000000001100110001010111;
assign LUT_3[45047] = 32'b00000000000000010011011100110100;
assign LUT_3[45048] = 32'b00000000000000010010110101000011;
assign LUT_3[45049] = 32'b00000000000000011001100000100000;
assign LUT_3[45050] = 32'b00000000000000010100111100100111;
assign LUT_3[45051] = 32'b00000000000000011011101000000100;
assign LUT_3[45052] = 32'b00000000000000010000000010111001;
assign LUT_3[45053] = 32'b00000000000000010110101110010110;
assign LUT_3[45054] = 32'b00000000000000010010001010011101;
assign LUT_3[45055] = 32'b00000000000000011000110101111010;
assign LUT_3[45056] = 32'b00000000000000000011001000010100;
assign LUT_3[45057] = 32'b00000000000000001001110011110001;
assign LUT_3[45058] = 32'b00000000000000000101001111111000;
assign LUT_3[45059] = 32'b00000000000000001011111011010101;
assign LUT_3[45060] = 32'b00000000000000000000010110001010;
assign LUT_3[45061] = 32'b00000000000000000111000001100111;
assign LUT_3[45062] = 32'b00000000000000000010011101101110;
assign LUT_3[45063] = 32'b00000000000000001001001001001011;
assign LUT_3[45064] = 32'b00000000000000001000100001011010;
assign LUT_3[45065] = 32'b00000000000000001111001100110111;
assign LUT_3[45066] = 32'b00000000000000001010101000111110;
assign LUT_3[45067] = 32'b00000000000000010001010100011011;
assign LUT_3[45068] = 32'b00000000000000000101101111010000;
assign LUT_3[45069] = 32'b00000000000000001100011010101101;
assign LUT_3[45070] = 32'b00000000000000000111110110110100;
assign LUT_3[45071] = 32'b00000000000000001110100010010001;
assign LUT_3[45072] = 32'b00000000000000000110011011010111;
assign LUT_3[45073] = 32'b00000000000000001101000110110100;
assign LUT_3[45074] = 32'b00000000000000001000100010111011;
assign LUT_3[45075] = 32'b00000000000000001111001110011000;
assign LUT_3[45076] = 32'b00000000000000000011101001001101;
assign LUT_3[45077] = 32'b00000000000000001010010100101010;
assign LUT_3[45078] = 32'b00000000000000000101110000110001;
assign LUT_3[45079] = 32'b00000000000000001100011100001110;
assign LUT_3[45080] = 32'b00000000000000001011110100011101;
assign LUT_3[45081] = 32'b00000000000000010010011111111010;
assign LUT_3[45082] = 32'b00000000000000001101111100000001;
assign LUT_3[45083] = 32'b00000000000000010100100111011110;
assign LUT_3[45084] = 32'b00000000000000001001000010010011;
assign LUT_3[45085] = 32'b00000000000000001111101101110000;
assign LUT_3[45086] = 32'b00000000000000001011001001110111;
assign LUT_3[45087] = 32'b00000000000000010001110101010100;
assign LUT_3[45088] = 32'b00000000000000000100010110110100;
assign LUT_3[45089] = 32'b00000000000000001011000010010001;
assign LUT_3[45090] = 32'b00000000000000000110011110011000;
assign LUT_3[45091] = 32'b00000000000000001101001001110101;
assign LUT_3[45092] = 32'b00000000000000000001100100101010;
assign LUT_3[45093] = 32'b00000000000000001000010000000111;
assign LUT_3[45094] = 32'b00000000000000000011101100001110;
assign LUT_3[45095] = 32'b00000000000000001010010111101011;
assign LUT_3[45096] = 32'b00000000000000001001101111111010;
assign LUT_3[45097] = 32'b00000000000000010000011011010111;
assign LUT_3[45098] = 32'b00000000000000001011110111011110;
assign LUT_3[45099] = 32'b00000000000000010010100010111011;
assign LUT_3[45100] = 32'b00000000000000000110111101110000;
assign LUT_3[45101] = 32'b00000000000000001101101001001101;
assign LUT_3[45102] = 32'b00000000000000001001000101010100;
assign LUT_3[45103] = 32'b00000000000000001111110000110001;
assign LUT_3[45104] = 32'b00000000000000000111101001110111;
assign LUT_3[45105] = 32'b00000000000000001110010101010100;
assign LUT_3[45106] = 32'b00000000000000001001110001011011;
assign LUT_3[45107] = 32'b00000000000000010000011100111000;
assign LUT_3[45108] = 32'b00000000000000000100110111101101;
assign LUT_3[45109] = 32'b00000000000000001011100011001010;
assign LUT_3[45110] = 32'b00000000000000000110111111010001;
assign LUT_3[45111] = 32'b00000000000000001101101010101110;
assign LUT_3[45112] = 32'b00000000000000001101000010111101;
assign LUT_3[45113] = 32'b00000000000000010011101110011010;
assign LUT_3[45114] = 32'b00000000000000001111001010100001;
assign LUT_3[45115] = 32'b00000000000000010101110101111110;
assign LUT_3[45116] = 32'b00000000000000001010010000110011;
assign LUT_3[45117] = 32'b00000000000000010000111100010000;
assign LUT_3[45118] = 32'b00000000000000001100011000010111;
assign LUT_3[45119] = 32'b00000000000000010011000011110100;
assign LUT_3[45120] = 32'b00000000000000000011000000111111;
assign LUT_3[45121] = 32'b00000000000000001001101100011100;
assign LUT_3[45122] = 32'b00000000000000000101001000100011;
assign LUT_3[45123] = 32'b00000000000000001011110100000000;
assign LUT_3[45124] = 32'b00000000000000000000001110110101;
assign LUT_3[45125] = 32'b00000000000000000110111010010010;
assign LUT_3[45126] = 32'b00000000000000000010010110011001;
assign LUT_3[45127] = 32'b00000000000000001001000001110110;
assign LUT_3[45128] = 32'b00000000000000001000011010000101;
assign LUT_3[45129] = 32'b00000000000000001111000101100010;
assign LUT_3[45130] = 32'b00000000000000001010100001101001;
assign LUT_3[45131] = 32'b00000000000000010001001101000110;
assign LUT_3[45132] = 32'b00000000000000000101100111111011;
assign LUT_3[45133] = 32'b00000000000000001100010011011000;
assign LUT_3[45134] = 32'b00000000000000000111101111011111;
assign LUT_3[45135] = 32'b00000000000000001110011010111100;
assign LUT_3[45136] = 32'b00000000000000000110010100000010;
assign LUT_3[45137] = 32'b00000000000000001100111111011111;
assign LUT_3[45138] = 32'b00000000000000001000011011100110;
assign LUT_3[45139] = 32'b00000000000000001111000111000011;
assign LUT_3[45140] = 32'b00000000000000000011100001111000;
assign LUT_3[45141] = 32'b00000000000000001010001101010101;
assign LUT_3[45142] = 32'b00000000000000000101101001011100;
assign LUT_3[45143] = 32'b00000000000000001100010100111001;
assign LUT_3[45144] = 32'b00000000000000001011101101001000;
assign LUT_3[45145] = 32'b00000000000000010010011000100101;
assign LUT_3[45146] = 32'b00000000000000001101110100101100;
assign LUT_3[45147] = 32'b00000000000000010100100000001001;
assign LUT_3[45148] = 32'b00000000000000001000111010111110;
assign LUT_3[45149] = 32'b00000000000000001111100110011011;
assign LUT_3[45150] = 32'b00000000000000001011000010100010;
assign LUT_3[45151] = 32'b00000000000000010001101101111111;
assign LUT_3[45152] = 32'b00000000000000000100001111011111;
assign LUT_3[45153] = 32'b00000000000000001010111010111100;
assign LUT_3[45154] = 32'b00000000000000000110010111000011;
assign LUT_3[45155] = 32'b00000000000000001101000010100000;
assign LUT_3[45156] = 32'b00000000000000000001011101010101;
assign LUT_3[45157] = 32'b00000000000000001000001000110010;
assign LUT_3[45158] = 32'b00000000000000000011100100111001;
assign LUT_3[45159] = 32'b00000000000000001010010000010110;
assign LUT_3[45160] = 32'b00000000000000001001101000100101;
assign LUT_3[45161] = 32'b00000000000000010000010100000010;
assign LUT_3[45162] = 32'b00000000000000001011110000001001;
assign LUT_3[45163] = 32'b00000000000000010010011011100110;
assign LUT_3[45164] = 32'b00000000000000000110110110011011;
assign LUT_3[45165] = 32'b00000000000000001101100001111000;
assign LUT_3[45166] = 32'b00000000000000001000111101111111;
assign LUT_3[45167] = 32'b00000000000000001111101001011100;
assign LUT_3[45168] = 32'b00000000000000000111100010100010;
assign LUT_3[45169] = 32'b00000000000000001110001101111111;
assign LUT_3[45170] = 32'b00000000000000001001101010000110;
assign LUT_3[45171] = 32'b00000000000000010000010101100011;
assign LUT_3[45172] = 32'b00000000000000000100110000011000;
assign LUT_3[45173] = 32'b00000000000000001011011011110101;
assign LUT_3[45174] = 32'b00000000000000000110110111111100;
assign LUT_3[45175] = 32'b00000000000000001101100011011001;
assign LUT_3[45176] = 32'b00000000000000001100111011101000;
assign LUT_3[45177] = 32'b00000000000000010011100111000101;
assign LUT_3[45178] = 32'b00000000000000001111000011001100;
assign LUT_3[45179] = 32'b00000000000000010101101110101001;
assign LUT_3[45180] = 32'b00000000000000001010001001011110;
assign LUT_3[45181] = 32'b00000000000000010000110100111011;
assign LUT_3[45182] = 32'b00000000000000001100010001000010;
assign LUT_3[45183] = 32'b00000000000000010010111100011111;
assign LUT_3[45184] = 32'b00000000000000000101010011010010;
assign LUT_3[45185] = 32'b00000000000000001011111110101111;
assign LUT_3[45186] = 32'b00000000000000000111011010110110;
assign LUT_3[45187] = 32'b00000000000000001110000110010011;
assign LUT_3[45188] = 32'b00000000000000000010100001001000;
assign LUT_3[45189] = 32'b00000000000000001001001100100101;
assign LUT_3[45190] = 32'b00000000000000000100101000101100;
assign LUT_3[45191] = 32'b00000000000000001011010100001001;
assign LUT_3[45192] = 32'b00000000000000001010101100011000;
assign LUT_3[45193] = 32'b00000000000000010001010111110101;
assign LUT_3[45194] = 32'b00000000000000001100110011111100;
assign LUT_3[45195] = 32'b00000000000000010011011111011001;
assign LUT_3[45196] = 32'b00000000000000000111111010001110;
assign LUT_3[45197] = 32'b00000000000000001110100101101011;
assign LUT_3[45198] = 32'b00000000000000001010000001110010;
assign LUT_3[45199] = 32'b00000000000000010000101101001111;
assign LUT_3[45200] = 32'b00000000000000001000100110010101;
assign LUT_3[45201] = 32'b00000000000000001111010001110010;
assign LUT_3[45202] = 32'b00000000000000001010101101111001;
assign LUT_3[45203] = 32'b00000000000000010001011001010110;
assign LUT_3[45204] = 32'b00000000000000000101110100001011;
assign LUT_3[45205] = 32'b00000000000000001100011111101000;
assign LUT_3[45206] = 32'b00000000000000000111111011101111;
assign LUT_3[45207] = 32'b00000000000000001110100111001100;
assign LUT_3[45208] = 32'b00000000000000001101111111011011;
assign LUT_3[45209] = 32'b00000000000000010100101010111000;
assign LUT_3[45210] = 32'b00000000000000010000000110111111;
assign LUT_3[45211] = 32'b00000000000000010110110010011100;
assign LUT_3[45212] = 32'b00000000000000001011001101010001;
assign LUT_3[45213] = 32'b00000000000000010001111000101110;
assign LUT_3[45214] = 32'b00000000000000001101010100110101;
assign LUT_3[45215] = 32'b00000000000000010100000000010010;
assign LUT_3[45216] = 32'b00000000000000000110100001110010;
assign LUT_3[45217] = 32'b00000000000000001101001101001111;
assign LUT_3[45218] = 32'b00000000000000001000101001010110;
assign LUT_3[45219] = 32'b00000000000000001111010100110011;
assign LUT_3[45220] = 32'b00000000000000000011101111101000;
assign LUT_3[45221] = 32'b00000000000000001010011011000101;
assign LUT_3[45222] = 32'b00000000000000000101110111001100;
assign LUT_3[45223] = 32'b00000000000000001100100010101001;
assign LUT_3[45224] = 32'b00000000000000001011111010111000;
assign LUT_3[45225] = 32'b00000000000000010010100110010101;
assign LUT_3[45226] = 32'b00000000000000001110000010011100;
assign LUT_3[45227] = 32'b00000000000000010100101101111001;
assign LUT_3[45228] = 32'b00000000000000001001001000101110;
assign LUT_3[45229] = 32'b00000000000000001111110100001011;
assign LUT_3[45230] = 32'b00000000000000001011010000010010;
assign LUT_3[45231] = 32'b00000000000000010001111011101111;
assign LUT_3[45232] = 32'b00000000000000001001110100110101;
assign LUT_3[45233] = 32'b00000000000000010000100000010010;
assign LUT_3[45234] = 32'b00000000000000001011111100011001;
assign LUT_3[45235] = 32'b00000000000000010010100111110110;
assign LUT_3[45236] = 32'b00000000000000000111000010101011;
assign LUT_3[45237] = 32'b00000000000000001101101110001000;
assign LUT_3[45238] = 32'b00000000000000001001001010001111;
assign LUT_3[45239] = 32'b00000000000000001111110101101100;
assign LUT_3[45240] = 32'b00000000000000001111001101111011;
assign LUT_3[45241] = 32'b00000000000000010101111001011000;
assign LUT_3[45242] = 32'b00000000000000010001010101011111;
assign LUT_3[45243] = 32'b00000000000000011000000000111100;
assign LUT_3[45244] = 32'b00000000000000001100011011110001;
assign LUT_3[45245] = 32'b00000000000000010011000111001110;
assign LUT_3[45246] = 32'b00000000000000001110100011010101;
assign LUT_3[45247] = 32'b00000000000000010101001110110010;
assign LUT_3[45248] = 32'b00000000000000000101001011111101;
assign LUT_3[45249] = 32'b00000000000000001011110111011010;
assign LUT_3[45250] = 32'b00000000000000000111010011100001;
assign LUT_3[45251] = 32'b00000000000000001101111110111110;
assign LUT_3[45252] = 32'b00000000000000000010011001110011;
assign LUT_3[45253] = 32'b00000000000000001001000101010000;
assign LUT_3[45254] = 32'b00000000000000000100100001010111;
assign LUT_3[45255] = 32'b00000000000000001011001100110100;
assign LUT_3[45256] = 32'b00000000000000001010100101000011;
assign LUT_3[45257] = 32'b00000000000000010001010000100000;
assign LUT_3[45258] = 32'b00000000000000001100101100100111;
assign LUT_3[45259] = 32'b00000000000000010011011000000100;
assign LUT_3[45260] = 32'b00000000000000000111110010111001;
assign LUT_3[45261] = 32'b00000000000000001110011110010110;
assign LUT_3[45262] = 32'b00000000000000001001111010011101;
assign LUT_3[45263] = 32'b00000000000000010000100101111010;
assign LUT_3[45264] = 32'b00000000000000001000011111000000;
assign LUT_3[45265] = 32'b00000000000000001111001010011101;
assign LUT_3[45266] = 32'b00000000000000001010100110100100;
assign LUT_3[45267] = 32'b00000000000000010001010010000001;
assign LUT_3[45268] = 32'b00000000000000000101101100110110;
assign LUT_3[45269] = 32'b00000000000000001100011000010011;
assign LUT_3[45270] = 32'b00000000000000000111110100011010;
assign LUT_3[45271] = 32'b00000000000000001110011111110111;
assign LUT_3[45272] = 32'b00000000000000001101111000000110;
assign LUT_3[45273] = 32'b00000000000000010100100011100011;
assign LUT_3[45274] = 32'b00000000000000001111111111101010;
assign LUT_3[45275] = 32'b00000000000000010110101011000111;
assign LUT_3[45276] = 32'b00000000000000001011000101111100;
assign LUT_3[45277] = 32'b00000000000000010001110001011001;
assign LUT_3[45278] = 32'b00000000000000001101001101100000;
assign LUT_3[45279] = 32'b00000000000000010011111000111101;
assign LUT_3[45280] = 32'b00000000000000000110011010011101;
assign LUT_3[45281] = 32'b00000000000000001101000101111010;
assign LUT_3[45282] = 32'b00000000000000001000100010000001;
assign LUT_3[45283] = 32'b00000000000000001111001101011110;
assign LUT_3[45284] = 32'b00000000000000000011101000010011;
assign LUT_3[45285] = 32'b00000000000000001010010011110000;
assign LUT_3[45286] = 32'b00000000000000000101101111110111;
assign LUT_3[45287] = 32'b00000000000000001100011011010100;
assign LUT_3[45288] = 32'b00000000000000001011110011100011;
assign LUT_3[45289] = 32'b00000000000000010010011111000000;
assign LUT_3[45290] = 32'b00000000000000001101111011000111;
assign LUT_3[45291] = 32'b00000000000000010100100110100100;
assign LUT_3[45292] = 32'b00000000000000001001000001011001;
assign LUT_3[45293] = 32'b00000000000000001111101100110110;
assign LUT_3[45294] = 32'b00000000000000001011001000111101;
assign LUT_3[45295] = 32'b00000000000000010001110100011010;
assign LUT_3[45296] = 32'b00000000000000001001101101100000;
assign LUT_3[45297] = 32'b00000000000000010000011000111101;
assign LUT_3[45298] = 32'b00000000000000001011110101000100;
assign LUT_3[45299] = 32'b00000000000000010010100000100001;
assign LUT_3[45300] = 32'b00000000000000000110111011010110;
assign LUT_3[45301] = 32'b00000000000000001101100110110011;
assign LUT_3[45302] = 32'b00000000000000001001000010111010;
assign LUT_3[45303] = 32'b00000000000000001111101110010111;
assign LUT_3[45304] = 32'b00000000000000001111000110100110;
assign LUT_3[45305] = 32'b00000000000000010101110010000011;
assign LUT_3[45306] = 32'b00000000000000010001001110001010;
assign LUT_3[45307] = 32'b00000000000000010111111001100111;
assign LUT_3[45308] = 32'b00000000000000001100010100011100;
assign LUT_3[45309] = 32'b00000000000000010010111111111001;
assign LUT_3[45310] = 32'b00000000000000001110011100000000;
assign LUT_3[45311] = 32'b00000000000000010101000111011101;
assign LUT_3[45312] = 32'b11111111111111111111010111110101;
assign LUT_3[45313] = 32'b00000000000000000110000011010010;
assign LUT_3[45314] = 32'b00000000000000000001011111011001;
assign LUT_3[45315] = 32'b00000000000000001000001010110110;
assign LUT_3[45316] = 32'b11111111111111111100100101101011;
assign LUT_3[45317] = 32'b00000000000000000011010001001000;
assign LUT_3[45318] = 32'b11111111111111111110101101001111;
assign LUT_3[45319] = 32'b00000000000000000101011000101100;
assign LUT_3[45320] = 32'b00000000000000000100110000111011;
assign LUT_3[45321] = 32'b00000000000000001011011100011000;
assign LUT_3[45322] = 32'b00000000000000000110111000011111;
assign LUT_3[45323] = 32'b00000000000000001101100011111100;
assign LUT_3[45324] = 32'b00000000000000000001111110110001;
assign LUT_3[45325] = 32'b00000000000000001000101010001110;
assign LUT_3[45326] = 32'b00000000000000000100000110010101;
assign LUT_3[45327] = 32'b00000000000000001010110001110010;
assign LUT_3[45328] = 32'b00000000000000000010101010111000;
assign LUT_3[45329] = 32'b00000000000000001001010110010101;
assign LUT_3[45330] = 32'b00000000000000000100110010011100;
assign LUT_3[45331] = 32'b00000000000000001011011101111001;
assign LUT_3[45332] = 32'b11111111111111111111111000101110;
assign LUT_3[45333] = 32'b00000000000000000110100100001011;
assign LUT_3[45334] = 32'b00000000000000000010000000010010;
assign LUT_3[45335] = 32'b00000000000000001000101011101111;
assign LUT_3[45336] = 32'b00000000000000001000000011111110;
assign LUT_3[45337] = 32'b00000000000000001110101111011011;
assign LUT_3[45338] = 32'b00000000000000001010001011100010;
assign LUT_3[45339] = 32'b00000000000000010000110110111111;
assign LUT_3[45340] = 32'b00000000000000000101010001110100;
assign LUT_3[45341] = 32'b00000000000000001011111101010001;
assign LUT_3[45342] = 32'b00000000000000000111011001011000;
assign LUT_3[45343] = 32'b00000000000000001110000100110101;
assign LUT_3[45344] = 32'b00000000000000000000100110010101;
assign LUT_3[45345] = 32'b00000000000000000111010001110010;
assign LUT_3[45346] = 32'b00000000000000000010101101111001;
assign LUT_3[45347] = 32'b00000000000000001001011001010110;
assign LUT_3[45348] = 32'b11111111111111111101110100001011;
assign LUT_3[45349] = 32'b00000000000000000100011111101000;
assign LUT_3[45350] = 32'b11111111111111111111111011101111;
assign LUT_3[45351] = 32'b00000000000000000110100111001100;
assign LUT_3[45352] = 32'b00000000000000000101111111011011;
assign LUT_3[45353] = 32'b00000000000000001100101010111000;
assign LUT_3[45354] = 32'b00000000000000001000000110111111;
assign LUT_3[45355] = 32'b00000000000000001110110010011100;
assign LUT_3[45356] = 32'b00000000000000000011001101010001;
assign LUT_3[45357] = 32'b00000000000000001001111000101110;
assign LUT_3[45358] = 32'b00000000000000000101010100110101;
assign LUT_3[45359] = 32'b00000000000000001100000000010010;
assign LUT_3[45360] = 32'b00000000000000000011111001011000;
assign LUT_3[45361] = 32'b00000000000000001010100100110101;
assign LUT_3[45362] = 32'b00000000000000000110000000111100;
assign LUT_3[45363] = 32'b00000000000000001100101100011001;
assign LUT_3[45364] = 32'b00000000000000000001000111001110;
assign LUT_3[45365] = 32'b00000000000000000111110010101011;
assign LUT_3[45366] = 32'b00000000000000000011001110110010;
assign LUT_3[45367] = 32'b00000000000000001001111010001111;
assign LUT_3[45368] = 32'b00000000000000001001010010011110;
assign LUT_3[45369] = 32'b00000000000000001111111101111011;
assign LUT_3[45370] = 32'b00000000000000001011011010000010;
assign LUT_3[45371] = 32'b00000000000000010010000101011111;
assign LUT_3[45372] = 32'b00000000000000000110100000010100;
assign LUT_3[45373] = 32'b00000000000000001101001011110001;
assign LUT_3[45374] = 32'b00000000000000001000100111111000;
assign LUT_3[45375] = 32'b00000000000000001111010011010101;
assign LUT_3[45376] = 32'b11111111111111111111010000100000;
assign LUT_3[45377] = 32'b00000000000000000101111011111101;
assign LUT_3[45378] = 32'b00000000000000000001011000000100;
assign LUT_3[45379] = 32'b00000000000000001000000011100001;
assign LUT_3[45380] = 32'b11111111111111111100011110010110;
assign LUT_3[45381] = 32'b00000000000000000011001001110011;
assign LUT_3[45382] = 32'b11111111111111111110100101111010;
assign LUT_3[45383] = 32'b00000000000000000101010001010111;
assign LUT_3[45384] = 32'b00000000000000000100101001100110;
assign LUT_3[45385] = 32'b00000000000000001011010101000011;
assign LUT_3[45386] = 32'b00000000000000000110110001001010;
assign LUT_3[45387] = 32'b00000000000000001101011100100111;
assign LUT_3[45388] = 32'b00000000000000000001110111011100;
assign LUT_3[45389] = 32'b00000000000000001000100010111001;
assign LUT_3[45390] = 32'b00000000000000000011111111000000;
assign LUT_3[45391] = 32'b00000000000000001010101010011101;
assign LUT_3[45392] = 32'b00000000000000000010100011100011;
assign LUT_3[45393] = 32'b00000000000000001001001111000000;
assign LUT_3[45394] = 32'b00000000000000000100101011000111;
assign LUT_3[45395] = 32'b00000000000000001011010110100100;
assign LUT_3[45396] = 32'b11111111111111111111110001011001;
assign LUT_3[45397] = 32'b00000000000000000110011100110110;
assign LUT_3[45398] = 32'b00000000000000000001111000111101;
assign LUT_3[45399] = 32'b00000000000000001000100100011010;
assign LUT_3[45400] = 32'b00000000000000000111111100101001;
assign LUT_3[45401] = 32'b00000000000000001110101000000110;
assign LUT_3[45402] = 32'b00000000000000001010000100001101;
assign LUT_3[45403] = 32'b00000000000000010000101111101010;
assign LUT_3[45404] = 32'b00000000000000000101001010011111;
assign LUT_3[45405] = 32'b00000000000000001011110101111100;
assign LUT_3[45406] = 32'b00000000000000000111010010000011;
assign LUT_3[45407] = 32'b00000000000000001101111101100000;
assign LUT_3[45408] = 32'b00000000000000000000011111000000;
assign LUT_3[45409] = 32'b00000000000000000111001010011101;
assign LUT_3[45410] = 32'b00000000000000000010100110100100;
assign LUT_3[45411] = 32'b00000000000000001001010010000001;
assign LUT_3[45412] = 32'b11111111111111111101101100110110;
assign LUT_3[45413] = 32'b00000000000000000100011000010011;
assign LUT_3[45414] = 32'b11111111111111111111110100011010;
assign LUT_3[45415] = 32'b00000000000000000110011111110111;
assign LUT_3[45416] = 32'b00000000000000000101111000000110;
assign LUT_3[45417] = 32'b00000000000000001100100011100011;
assign LUT_3[45418] = 32'b00000000000000000111111111101010;
assign LUT_3[45419] = 32'b00000000000000001110101011000111;
assign LUT_3[45420] = 32'b00000000000000000011000101111100;
assign LUT_3[45421] = 32'b00000000000000001001110001011001;
assign LUT_3[45422] = 32'b00000000000000000101001101100000;
assign LUT_3[45423] = 32'b00000000000000001011111000111101;
assign LUT_3[45424] = 32'b00000000000000000011110010000011;
assign LUT_3[45425] = 32'b00000000000000001010011101100000;
assign LUT_3[45426] = 32'b00000000000000000101111001100111;
assign LUT_3[45427] = 32'b00000000000000001100100101000100;
assign LUT_3[45428] = 32'b00000000000000000000111111111001;
assign LUT_3[45429] = 32'b00000000000000000111101011010110;
assign LUT_3[45430] = 32'b00000000000000000011000111011101;
assign LUT_3[45431] = 32'b00000000000000001001110010111010;
assign LUT_3[45432] = 32'b00000000000000001001001011001001;
assign LUT_3[45433] = 32'b00000000000000001111110110100110;
assign LUT_3[45434] = 32'b00000000000000001011010010101101;
assign LUT_3[45435] = 32'b00000000000000010001111110001010;
assign LUT_3[45436] = 32'b00000000000000000110011000111111;
assign LUT_3[45437] = 32'b00000000000000001101000100011100;
assign LUT_3[45438] = 32'b00000000000000001000100000100011;
assign LUT_3[45439] = 32'b00000000000000001111001100000000;
assign LUT_3[45440] = 32'b00000000000000000001100010110011;
assign LUT_3[45441] = 32'b00000000000000001000001110010000;
assign LUT_3[45442] = 32'b00000000000000000011101010010111;
assign LUT_3[45443] = 32'b00000000000000001010010101110100;
assign LUT_3[45444] = 32'b11111111111111111110110000101001;
assign LUT_3[45445] = 32'b00000000000000000101011100000110;
assign LUT_3[45446] = 32'b00000000000000000000111000001101;
assign LUT_3[45447] = 32'b00000000000000000111100011101010;
assign LUT_3[45448] = 32'b00000000000000000110111011111001;
assign LUT_3[45449] = 32'b00000000000000001101100111010110;
assign LUT_3[45450] = 32'b00000000000000001001000011011101;
assign LUT_3[45451] = 32'b00000000000000001111101110111010;
assign LUT_3[45452] = 32'b00000000000000000100001001101111;
assign LUT_3[45453] = 32'b00000000000000001010110101001100;
assign LUT_3[45454] = 32'b00000000000000000110010001010011;
assign LUT_3[45455] = 32'b00000000000000001100111100110000;
assign LUT_3[45456] = 32'b00000000000000000100110101110110;
assign LUT_3[45457] = 32'b00000000000000001011100001010011;
assign LUT_3[45458] = 32'b00000000000000000110111101011010;
assign LUT_3[45459] = 32'b00000000000000001101101000110111;
assign LUT_3[45460] = 32'b00000000000000000010000011101100;
assign LUT_3[45461] = 32'b00000000000000001000101111001001;
assign LUT_3[45462] = 32'b00000000000000000100001011010000;
assign LUT_3[45463] = 32'b00000000000000001010110110101101;
assign LUT_3[45464] = 32'b00000000000000001010001110111100;
assign LUT_3[45465] = 32'b00000000000000010000111010011001;
assign LUT_3[45466] = 32'b00000000000000001100010110100000;
assign LUT_3[45467] = 32'b00000000000000010011000001111101;
assign LUT_3[45468] = 32'b00000000000000000111011100110010;
assign LUT_3[45469] = 32'b00000000000000001110001000001111;
assign LUT_3[45470] = 32'b00000000000000001001100100010110;
assign LUT_3[45471] = 32'b00000000000000010000001111110011;
assign LUT_3[45472] = 32'b00000000000000000010110001010011;
assign LUT_3[45473] = 32'b00000000000000001001011100110000;
assign LUT_3[45474] = 32'b00000000000000000100111000110111;
assign LUT_3[45475] = 32'b00000000000000001011100100010100;
assign LUT_3[45476] = 32'b11111111111111111111111111001001;
assign LUT_3[45477] = 32'b00000000000000000110101010100110;
assign LUT_3[45478] = 32'b00000000000000000010000110101101;
assign LUT_3[45479] = 32'b00000000000000001000110010001010;
assign LUT_3[45480] = 32'b00000000000000001000001010011001;
assign LUT_3[45481] = 32'b00000000000000001110110101110110;
assign LUT_3[45482] = 32'b00000000000000001010010001111101;
assign LUT_3[45483] = 32'b00000000000000010000111101011010;
assign LUT_3[45484] = 32'b00000000000000000101011000001111;
assign LUT_3[45485] = 32'b00000000000000001100000011101100;
assign LUT_3[45486] = 32'b00000000000000000111011111110011;
assign LUT_3[45487] = 32'b00000000000000001110001011010000;
assign LUT_3[45488] = 32'b00000000000000000110000100010110;
assign LUT_3[45489] = 32'b00000000000000001100101111110011;
assign LUT_3[45490] = 32'b00000000000000001000001011111010;
assign LUT_3[45491] = 32'b00000000000000001110110111010111;
assign LUT_3[45492] = 32'b00000000000000000011010010001100;
assign LUT_3[45493] = 32'b00000000000000001001111101101001;
assign LUT_3[45494] = 32'b00000000000000000101011001110000;
assign LUT_3[45495] = 32'b00000000000000001100000101001101;
assign LUT_3[45496] = 32'b00000000000000001011011101011100;
assign LUT_3[45497] = 32'b00000000000000010010001000111001;
assign LUT_3[45498] = 32'b00000000000000001101100101000000;
assign LUT_3[45499] = 32'b00000000000000010100010000011101;
assign LUT_3[45500] = 32'b00000000000000001000101011010010;
assign LUT_3[45501] = 32'b00000000000000001111010110101111;
assign LUT_3[45502] = 32'b00000000000000001010110010110110;
assign LUT_3[45503] = 32'b00000000000000010001011110010011;
assign LUT_3[45504] = 32'b00000000000000000001011011011110;
assign LUT_3[45505] = 32'b00000000000000001000000110111011;
assign LUT_3[45506] = 32'b00000000000000000011100011000010;
assign LUT_3[45507] = 32'b00000000000000001010001110011111;
assign LUT_3[45508] = 32'b11111111111111111110101001010100;
assign LUT_3[45509] = 32'b00000000000000000101010100110001;
assign LUT_3[45510] = 32'b00000000000000000000110000111000;
assign LUT_3[45511] = 32'b00000000000000000111011100010101;
assign LUT_3[45512] = 32'b00000000000000000110110100100100;
assign LUT_3[45513] = 32'b00000000000000001101100000000001;
assign LUT_3[45514] = 32'b00000000000000001000111100001000;
assign LUT_3[45515] = 32'b00000000000000001111100111100101;
assign LUT_3[45516] = 32'b00000000000000000100000010011010;
assign LUT_3[45517] = 32'b00000000000000001010101101110111;
assign LUT_3[45518] = 32'b00000000000000000110001001111110;
assign LUT_3[45519] = 32'b00000000000000001100110101011011;
assign LUT_3[45520] = 32'b00000000000000000100101110100001;
assign LUT_3[45521] = 32'b00000000000000001011011001111110;
assign LUT_3[45522] = 32'b00000000000000000110110110000101;
assign LUT_3[45523] = 32'b00000000000000001101100001100010;
assign LUT_3[45524] = 32'b00000000000000000001111100010111;
assign LUT_3[45525] = 32'b00000000000000001000100111110100;
assign LUT_3[45526] = 32'b00000000000000000100000011111011;
assign LUT_3[45527] = 32'b00000000000000001010101111011000;
assign LUT_3[45528] = 32'b00000000000000001010000111100111;
assign LUT_3[45529] = 32'b00000000000000010000110011000100;
assign LUT_3[45530] = 32'b00000000000000001100001111001011;
assign LUT_3[45531] = 32'b00000000000000010010111010101000;
assign LUT_3[45532] = 32'b00000000000000000111010101011101;
assign LUT_3[45533] = 32'b00000000000000001110000000111010;
assign LUT_3[45534] = 32'b00000000000000001001011101000001;
assign LUT_3[45535] = 32'b00000000000000010000001000011110;
assign LUT_3[45536] = 32'b00000000000000000010101001111110;
assign LUT_3[45537] = 32'b00000000000000001001010101011011;
assign LUT_3[45538] = 32'b00000000000000000100110001100010;
assign LUT_3[45539] = 32'b00000000000000001011011100111111;
assign LUT_3[45540] = 32'b11111111111111111111110111110100;
assign LUT_3[45541] = 32'b00000000000000000110100011010001;
assign LUT_3[45542] = 32'b00000000000000000001111111011000;
assign LUT_3[45543] = 32'b00000000000000001000101010110101;
assign LUT_3[45544] = 32'b00000000000000001000000011000100;
assign LUT_3[45545] = 32'b00000000000000001110101110100001;
assign LUT_3[45546] = 32'b00000000000000001010001010101000;
assign LUT_3[45547] = 32'b00000000000000010000110110000101;
assign LUT_3[45548] = 32'b00000000000000000101010000111010;
assign LUT_3[45549] = 32'b00000000000000001011111100010111;
assign LUT_3[45550] = 32'b00000000000000000111011000011110;
assign LUT_3[45551] = 32'b00000000000000001110000011111011;
assign LUT_3[45552] = 32'b00000000000000000101111101000001;
assign LUT_3[45553] = 32'b00000000000000001100101000011110;
assign LUT_3[45554] = 32'b00000000000000001000000100100101;
assign LUT_3[45555] = 32'b00000000000000001110110000000010;
assign LUT_3[45556] = 32'b00000000000000000011001010110111;
assign LUT_3[45557] = 32'b00000000000000001001110110010100;
assign LUT_3[45558] = 32'b00000000000000000101010010011011;
assign LUT_3[45559] = 32'b00000000000000001011111101111000;
assign LUT_3[45560] = 32'b00000000000000001011010110000111;
assign LUT_3[45561] = 32'b00000000000000010010000001100100;
assign LUT_3[45562] = 32'b00000000000000001101011101101011;
assign LUT_3[45563] = 32'b00000000000000010100001001001000;
assign LUT_3[45564] = 32'b00000000000000001000100011111101;
assign LUT_3[45565] = 32'b00000000000000001111001111011010;
assign LUT_3[45566] = 32'b00000000000000001010101011100001;
assign LUT_3[45567] = 32'b00000000000000010001010110111110;
assign LUT_3[45568] = 32'b00000000000000000110011101100000;
assign LUT_3[45569] = 32'b00000000000000001101001000111101;
assign LUT_3[45570] = 32'b00000000000000001000100101000100;
assign LUT_3[45571] = 32'b00000000000000001111010000100001;
assign LUT_3[45572] = 32'b00000000000000000011101011010110;
assign LUT_3[45573] = 32'b00000000000000001010010110110011;
assign LUT_3[45574] = 32'b00000000000000000101110010111010;
assign LUT_3[45575] = 32'b00000000000000001100011110010111;
assign LUT_3[45576] = 32'b00000000000000001011110110100110;
assign LUT_3[45577] = 32'b00000000000000010010100010000011;
assign LUT_3[45578] = 32'b00000000000000001101111110001010;
assign LUT_3[45579] = 32'b00000000000000010100101001100111;
assign LUT_3[45580] = 32'b00000000000000001001000100011100;
assign LUT_3[45581] = 32'b00000000000000001111101111111001;
assign LUT_3[45582] = 32'b00000000000000001011001100000000;
assign LUT_3[45583] = 32'b00000000000000010001110111011101;
assign LUT_3[45584] = 32'b00000000000000001001110000100011;
assign LUT_3[45585] = 32'b00000000000000010000011100000000;
assign LUT_3[45586] = 32'b00000000000000001011111000000111;
assign LUT_3[45587] = 32'b00000000000000010010100011100100;
assign LUT_3[45588] = 32'b00000000000000000110111110011001;
assign LUT_3[45589] = 32'b00000000000000001101101001110110;
assign LUT_3[45590] = 32'b00000000000000001001000101111101;
assign LUT_3[45591] = 32'b00000000000000001111110001011010;
assign LUT_3[45592] = 32'b00000000000000001111001001101001;
assign LUT_3[45593] = 32'b00000000000000010101110101000110;
assign LUT_3[45594] = 32'b00000000000000010001010001001101;
assign LUT_3[45595] = 32'b00000000000000010111111100101010;
assign LUT_3[45596] = 32'b00000000000000001100010111011111;
assign LUT_3[45597] = 32'b00000000000000010011000010111100;
assign LUT_3[45598] = 32'b00000000000000001110011111000011;
assign LUT_3[45599] = 32'b00000000000000010101001010100000;
assign LUT_3[45600] = 32'b00000000000000000111101100000000;
assign LUT_3[45601] = 32'b00000000000000001110010111011101;
assign LUT_3[45602] = 32'b00000000000000001001110011100100;
assign LUT_3[45603] = 32'b00000000000000010000011111000001;
assign LUT_3[45604] = 32'b00000000000000000100111001110110;
assign LUT_3[45605] = 32'b00000000000000001011100101010011;
assign LUT_3[45606] = 32'b00000000000000000111000001011010;
assign LUT_3[45607] = 32'b00000000000000001101101100110111;
assign LUT_3[45608] = 32'b00000000000000001101000101000110;
assign LUT_3[45609] = 32'b00000000000000010011110000100011;
assign LUT_3[45610] = 32'b00000000000000001111001100101010;
assign LUT_3[45611] = 32'b00000000000000010101111000000111;
assign LUT_3[45612] = 32'b00000000000000001010010010111100;
assign LUT_3[45613] = 32'b00000000000000010000111110011001;
assign LUT_3[45614] = 32'b00000000000000001100011010100000;
assign LUT_3[45615] = 32'b00000000000000010011000101111101;
assign LUT_3[45616] = 32'b00000000000000001010111111000011;
assign LUT_3[45617] = 32'b00000000000000010001101010100000;
assign LUT_3[45618] = 32'b00000000000000001101000110100111;
assign LUT_3[45619] = 32'b00000000000000010011110010000100;
assign LUT_3[45620] = 32'b00000000000000001000001100111001;
assign LUT_3[45621] = 32'b00000000000000001110111000010110;
assign LUT_3[45622] = 32'b00000000000000001010010100011101;
assign LUT_3[45623] = 32'b00000000000000010000111111111010;
assign LUT_3[45624] = 32'b00000000000000010000011000001001;
assign LUT_3[45625] = 32'b00000000000000010111000011100110;
assign LUT_3[45626] = 32'b00000000000000010010011111101101;
assign LUT_3[45627] = 32'b00000000000000011001001011001010;
assign LUT_3[45628] = 32'b00000000000000001101100101111111;
assign LUT_3[45629] = 32'b00000000000000010100010001011100;
assign LUT_3[45630] = 32'b00000000000000001111101101100011;
assign LUT_3[45631] = 32'b00000000000000010110011001000000;
assign LUT_3[45632] = 32'b00000000000000000110010110001011;
assign LUT_3[45633] = 32'b00000000000000001101000001101000;
assign LUT_3[45634] = 32'b00000000000000001000011101101111;
assign LUT_3[45635] = 32'b00000000000000001111001001001100;
assign LUT_3[45636] = 32'b00000000000000000011100100000001;
assign LUT_3[45637] = 32'b00000000000000001010001111011110;
assign LUT_3[45638] = 32'b00000000000000000101101011100101;
assign LUT_3[45639] = 32'b00000000000000001100010111000010;
assign LUT_3[45640] = 32'b00000000000000001011101111010001;
assign LUT_3[45641] = 32'b00000000000000010010011010101110;
assign LUT_3[45642] = 32'b00000000000000001101110110110101;
assign LUT_3[45643] = 32'b00000000000000010100100010010010;
assign LUT_3[45644] = 32'b00000000000000001000111101000111;
assign LUT_3[45645] = 32'b00000000000000001111101000100100;
assign LUT_3[45646] = 32'b00000000000000001011000100101011;
assign LUT_3[45647] = 32'b00000000000000010001110000001000;
assign LUT_3[45648] = 32'b00000000000000001001101001001110;
assign LUT_3[45649] = 32'b00000000000000010000010100101011;
assign LUT_3[45650] = 32'b00000000000000001011110000110010;
assign LUT_3[45651] = 32'b00000000000000010010011100001111;
assign LUT_3[45652] = 32'b00000000000000000110110111000100;
assign LUT_3[45653] = 32'b00000000000000001101100010100001;
assign LUT_3[45654] = 32'b00000000000000001000111110101000;
assign LUT_3[45655] = 32'b00000000000000001111101010000101;
assign LUT_3[45656] = 32'b00000000000000001111000010010100;
assign LUT_3[45657] = 32'b00000000000000010101101101110001;
assign LUT_3[45658] = 32'b00000000000000010001001001111000;
assign LUT_3[45659] = 32'b00000000000000010111110101010101;
assign LUT_3[45660] = 32'b00000000000000001100010000001010;
assign LUT_3[45661] = 32'b00000000000000010010111011100111;
assign LUT_3[45662] = 32'b00000000000000001110010111101110;
assign LUT_3[45663] = 32'b00000000000000010101000011001011;
assign LUT_3[45664] = 32'b00000000000000000111100100101011;
assign LUT_3[45665] = 32'b00000000000000001110010000001000;
assign LUT_3[45666] = 32'b00000000000000001001101100001111;
assign LUT_3[45667] = 32'b00000000000000010000010111101100;
assign LUT_3[45668] = 32'b00000000000000000100110010100001;
assign LUT_3[45669] = 32'b00000000000000001011011101111110;
assign LUT_3[45670] = 32'b00000000000000000110111010000101;
assign LUT_3[45671] = 32'b00000000000000001101100101100010;
assign LUT_3[45672] = 32'b00000000000000001100111101110001;
assign LUT_3[45673] = 32'b00000000000000010011101001001110;
assign LUT_3[45674] = 32'b00000000000000001111000101010101;
assign LUT_3[45675] = 32'b00000000000000010101110000110010;
assign LUT_3[45676] = 32'b00000000000000001010001011100111;
assign LUT_3[45677] = 32'b00000000000000010000110111000100;
assign LUT_3[45678] = 32'b00000000000000001100010011001011;
assign LUT_3[45679] = 32'b00000000000000010010111110101000;
assign LUT_3[45680] = 32'b00000000000000001010110111101110;
assign LUT_3[45681] = 32'b00000000000000010001100011001011;
assign LUT_3[45682] = 32'b00000000000000001100111111010010;
assign LUT_3[45683] = 32'b00000000000000010011101010101111;
assign LUT_3[45684] = 32'b00000000000000001000000101100100;
assign LUT_3[45685] = 32'b00000000000000001110110001000001;
assign LUT_3[45686] = 32'b00000000000000001010001101001000;
assign LUT_3[45687] = 32'b00000000000000010000111000100101;
assign LUT_3[45688] = 32'b00000000000000010000010000110100;
assign LUT_3[45689] = 32'b00000000000000010110111100010001;
assign LUT_3[45690] = 32'b00000000000000010010011000011000;
assign LUT_3[45691] = 32'b00000000000000011001000011110101;
assign LUT_3[45692] = 32'b00000000000000001101011110101010;
assign LUT_3[45693] = 32'b00000000000000010100001010000111;
assign LUT_3[45694] = 32'b00000000000000001111100110001110;
assign LUT_3[45695] = 32'b00000000000000010110010001101011;
assign LUT_3[45696] = 32'b00000000000000001000101000011110;
assign LUT_3[45697] = 32'b00000000000000001111010011111011;
assign LUT_3[45698] = 32'b00000000000000001010110000000010;
assign LUT_3[45699] = 32'b00000000000000010001011011011111;
assign LUT_3[45700] = 32'b00000000000000000101110110010100;
assign LUT_3[45701] = 32'b00000000000000001100100001110001;
assign LUT_3[45702] = 32'b00000000000000000111111101111000;
assign LUT_3[45703] = 32'b00000000000000001110101001010101;
assign LUT_3[45704] = 32'b00000000000000001110000001100100;
assign LUT_3[45705] = 32'b00000000000000010100101101000001;
assign LUT_3[45706] = 32'b00000000000000010000001001001000;
assign LUT_3[45707] = 32'b00000000000000010110110100100101;
assign LUT_3[45708] = 32'b00000000000000001011001111011010;
assign LUT_3[45709] = 32'b00000000000000010001111010110111;
assign LUT_3[45710] = 32'b00000000000000001101010110111110;
assign LUT_3[45711] = 32'b00000000000000010100000010011011;
assign LUT_3[45712] = 32'b00000000000000001011111011100001;
assign LUT_3[45713] = 32'b00000000000000010010100110111110;
assign LUT_3[45714] = 32'b00000000000000001110000011000101;
assign LUT_3[45715] = 32'b00000000000000010100101110100010;
assign LUT_3[45716] = 32'b00000000000000001001001001010111;
assign LUT_3[45717] = 32'b00000000000000001111110100110100;
assign LUT_3[45718] = 32'b00000000000000001011010000111011;
assign LUT_3[45719] = 32'b00000000000000010001111100011000;
assign LUT_3[45720] = 32'b00000000000000010001010100100111;
assign LUT_3[45721] = 32'b00000000000000011000000000000100;
assign LUT_3[45722] = 32'b00000000000000010011011100001011;
assign LUT_3[45723] = 32'b00000000000000011010000111101000;
assign LUT_3[45724] = 32'b00000000000000001110100010011101;
assign LUT_3[45725] = 32'b00000000000000010101001101111010;
assign LUT_3[45726] = 32'b00000000000000010000101010000001;
assign LUT_3[45727] = 32'b00000000000000010111010101011110;
assign LUT_3[45728] = 32'b00000000000000001001110110111110;
assign LUT_3[45729] = 32'b00000000000000010000100010011011;
assign LUT_3[45730] = 32'b00000000000000001011111110100010;
assign LUT_3[45731] = 32'b00000000000000010010101001111111;
assign LUT_3[45732] = 32'b00000000000000000111000100110100;
assign LUT_3[45733] = 32'b00000000000000001101110000010001;
assign LUT_3[45734] = 32'b00000000000000001001001100011000;
assign LUT_3[45735] = 32'b00000000000000001111110111110101;
assign LUT_3[45736] = 32'b00000000000000001111010000000100;
assign LUT_3[45737] = 32'b00000000000000010101111011100001;
assign LUT_3[45738] = 32'b00000000000000010001010111101000;
assign LUT_3[45739] = 32'b00000000000000011000000011000101;
assign LUT_3[45740] = 32'b00000000000000001100011101111010;
assign LUT_3[45741] = 32'b00000000000000010011001001010111;
assign LUT_3[45742] = 32'b00000000000000001110100101011110;
assign LUT_3[45743] = 32'b00000000000000010101010000111011;
assign LUT_3[45744] = 32'b00000000000000001101001010000001;
assign LUT_3[45745] = 32'b00000000000000010011110101011110;
assign LUT_3[45746] = 32'b00000000000000001111010001100101;
assign LUT_3[45747] = 32'b00000000000000010101111101000010;
assign LUT_3[45748] = 32'b00000000000000001010010111110111;
assign LUT_3[45749] = 32'b00000000000000010001000011010100;
assign LUT_3[45750] = 32'b00000000000000001100011111011011;
assign LUT_3[45751] = 32'b00000000000000010011001010111000;
assign LUT_3[45752] = 32'b00000000000000010010100011000111;
assign LUT_3[45753] = 32'b00000000000000011001001110100100;
assign LUT_3[45754] = 32'b00000000000000010100101010101011;
assign LUT_3[45755] = 32'b00000000000000011011010110001000;
assign LUT_3[45756] = 32'b00000000000000001111110000111101;
assign LUT_3[45757] = 32'b00000000000000010110011100011010;
assign LUT_3[45758] = 32'b00000000000000010001111000100001;
assign LUT_3[45759] = 32'b00000000000000011000100011111110;
assign LUT_3[45760] = 32'b00000000000000001000100001001001;
assign LUT_3[45761] = 32'b00000000000000001111001100100110;
assign LUT_3[45762] = 32'b00000000000000001010101000101101;
assign LUT_3[45763] = 32'b00000000000000010001010100001010;
assign LUT_3[45764] = 32'b00000000000000000101101110111111;
assign LUT_3[45765] = 32'b00000000000000001100011010011100;
assign LUT_3[45766] = 32'b00000000000000000111110110100011;
assign LUT_3[45767] = 32'b00000000000000001110100010000000;
assign LUT_3[45768] = 32'b00000000000000001101111010001111;
assign LUT_3[45769] = 32'b00000000000000010100100101101100;
assign LUT_3[45770] = 32'b00000000000000010000000001110011;
assign LUT_3[45771] = 32'b00000000000000010110101101010000;
assign LUT_3[45772] = 32'b00000000000000001011001000000101;
assign LUT_3[45773] = 32'b00000000000000010001110011100010;
assign LUT_3[45774] = 32'b00000000000000001101001111101001;
assign LUT_3[45775] = 32'b00000000000000010011111011000110;
assign LUT_3[45776] = 32'b00000000000000001011110100001100;
assign LUT_3[45777] = 32'b00000000000000010010011111101001;
assign LUT_3[45778] = 32'b00000000000000001101111011110000;
assign LUT_3[45779] = 32'b00000000000000010100100111001101;
assign LUT_3[45780] = 32'b00000000000000001001000010000010;
assign LUT_3[45781] = 32'b00000000000000001111101101011111;
assign LUT_3[45782] = 32'b00000000000000001011001001100110;
assign LUT_3[45783] = 32'b00000000000000010001110101000011;
assign LUT_3[45784] = 32'b00000000000000010001001101010010;
assign LUT_3[45785] = 32'b00000000000000010111111000101111;
assign LUT_3[45786] = 32'b00000000000000010011010100110110;
assign LUT_3[45787] = 32'b00000000000000011010000000010011;
assign LUT_3[45788] = 32'b00000000000000001110011011001000;
assign LUT_3[45789] = 32'b00000000000000010101000110100101;
assign LUT_3[45790] = 32'b00000000000000010000100010101100;
assign LUT_3[45791] = 32'b00000000000000010111001110001001;
assign LUT_3[45792] = 32'b00000000000000001001101111101001;
assign LUT_3[45793] = 32'b00000000000000010000011011000110;
assign LUT_3[45794] = 32'b00000000000000001011110111001101;
assign LUT_3[45795] = 32'b00000000000000010010100010101010;
assign LUT_3[45796] = 32'b00000000000000000110111101011111;
assign LUT_3[45797] = 32'b00000000000000001101101000111100;
assign LUT_3[45798] = 32'b00000000000000001001000101000011;
assign LUT_3[45799] = 32'b00000000000000001111110000100000;
assign LUT_3[45800] = 32'b00000000000000001111001000101111;
assign LUT_3[45801] = 32'b00000000000000010101110100001100;
assign LUT_3[45802] = 32'b00000000000000010001010000010011;
assign LUT_3[45803] = 32'b00000000000000010111111011110000;
assign LUT_3[45804] = 32'b00000000000000001100010110100101;
assign LUT_3[45805] = 32'b00000000000000010011000010000010;
assign LUT_3[45806] = 32'b00000000000000001110011110001001;
assign LUT_3[45807] = 32'b00000000000000010101001001100110;
assign LUT_3[45808] = 32'b00000000000000001101000010101100;
assign LUT_3[45809] = 32'b00000000000000010011101110001001;
assign LUT_3[45810] = 32'b00000000000000001111001010010000;
assign LUT_3[45811] = 32'b00000000000000010101110101101101;
assign LUT_3[45812] = 32'b00000000000000001010010000100010;
assign LUT_3[45813] = 32'b00000000000000010000111011111111;
assign LUT_3[45814] = 32'b00000000000000001100011000000110;
assign LUT_3[45815] = 32'b00000000000000010011000011100011;
assign LUT_3[45816] = 32'b00000000000000010010011011110010;
assign LUT_3[45817] = 32'b00000000000000011001000111001111;
assign LUT_3[45818] = 32'b00000000000000010100100011010110;
assign LUT_3[45819] = 32'b00000000000000011011001110110011;
assign LUT_3[45820] = 32'b00000000000000001111101001101000;
assign LUT_3[45821] = 32'b00000000000000010110010101000101;
assign LUT_3[45822] = 32'b00000000000000010001110001001100;
assign LUT_3[45823] = 32'b00000000000000011000011100101001;
assign LUT_3[45824] = 32'b00000000000000000010101101000001;
assign LUT_3[45825] = 32'b00000000000000001001011000011110;
assign LUT_3[45826] = 32'b00000000000000000100110100100101;
assign LUT_3[45827] = 32'b00000000000000001011100000000010;
assign LUT_3[45828] = 32'b11111111111111111111111010110111;
assign LUT_3[45829] = 32'b00000000000000000110100110010100;
assign LUT_3[45830] = 32'b00000000000000000010000010011011;
assign LUT_3[45831] = 32'b00000000000000001000101101111000;
assign LUT_3[45832] = 32'b00000000000000001000000110000111;
assign LUT_3[45833] = 32'b00000000000000001110110001100100;
assign LUT_3[45834] = 32'b00000000000000001010001101101011;
assign LUT_3[45835] = 32'b00000000000000010000111001001000;
assign LUT_3[45836] = 32'b00000000000000000101010011111101;
assign LUT_3[45837] = 32'b00000000000000001011111111011010;
assign LUT_3[45838] = 32'b00000000000000000111011011100001;
assign LUT_3[45839] = 32'b00000000000000001110000110111110;
assign LUT_3[45840] = 32'b00000000000000000110000000000100;
assign LUT_3[45841] = 32'b00000000000000001100101011100001;
assign LUT_3[45842] = 32'b00000000000000001000000111101000;
assign LUT_3[45843] = 32'b00000000000000001110110011000101;
assign LUT_3[45844] = 32'b00000000000000000011001101111010;
assign LUT_3[45845] = 32'b00000000000000001001111001010111;
assign LUT_3[45846] = 32'b00000000000000000101010101011110;
assign LUT_3[45847] = 32'b00000000000000001100000000111011;
assign LUT_3[45848] = 32'b00000000000000001011011001001010;
assign LUT_3[45849] = 32'b00000000000000010010000100100111;
assign LUT_3[45850] = 32'b00000000000000001101100000101110;
assign LUT_3[45851] = 32'b00000000000000010100001100001011;
assign LUT_3[45852] = 32'b00000000000000001000100111000000;
assign LUT_3[45853] = 32'b00000000000000001111010010011101;
assign LUT_3[45854] = 32'b00000000000000001010101110100100;
assign LUT_3[45855] = 32'b00000000000000010001011010000001;
assign LUT_3[45856] = 32'b00000000000000000011111011100001;
assign LUT_3[45857] = 32'b00000000000000001010100110111110;
assign LUT_3[45858] = 32'b00000000000000000110000011000101;
assign LUT_3[45859] = 32'b00000000000000001100101110100010;
assign LUT_3[45860] = 32'b00000000000000000001001001010111;
assign LUT_3[45861] = 32'b00000000000000000111110100110100;
assign LUT_3[45862] = 32'b00000000000000000011010000111011;
assign LUT_3[45863] = 32'b00000000000000001001111100011000;
assign LUT_3[45864] = 32'b00000000000000001001010100100111;
assign LUT_3[45865] = 32'b00000000000000010000000000000100;
assign LUT_3[45866] = 32'b00000000000000001011011100001011;
assign LUT_3[45867] = 32'b00000000000000010010000111101000;
assign LUT_3[45868] = 32'b00000000000000000110100010011101;
assign LUT_3[45869] = 32'b00000000000000001101001101111010;
assign LUT_3[45870] = 32'b00000000000000001000101010000001;
assign LUT_3[45871] = 32'b00000000000000001111010101011110;
assign LUT_3[45872] = 32'b00000000000000000111001110100100;
assign LUT_3[45873] = 32'b00000000000000001101111010000001;
assign LUT_3[45874] = 32'b00000000000000001001010110001000;
assign LUT_3[45875] = 32'b00000000000000010000000001100101;
assign LUT_3[45876] = 32'b00000000000000000100011100011010;
assign LUT_3[45877] = 32'b00000000000000001011000111110111;
assign LUT_3[45878] = 32'b00000000000000000110100011111110;
assign LUT_3[45879] = 32'b00000000000000001101001111011011;
assign LUT_3[45880] = 32'b00000000000000001100100111101010;
assign LUT_3[45881] = 32'b00000000000000010011010011000111;
assign LUT_3[45882] = 32'b00000000000000001110101111001110;
assign LUT_3[45883] = 32'b00000000000000010101011010101011;
assign LUT_3[45884] = 32'b00000000000000001001110101100000;
assign LUT_3[45885] = 32'b00000000000000010000100000111101;
assign LUT_3[45886] = 32'b00000000000000001011111101000100;
assign LUT_3[45887] = 32'b00000000000000010010101000100001;
assign LUT_3[45888] = 32'b00000000000000000010100101101100;
assign LUT_3[45889] = 32'b00000000000000001001010001001001;
assign LUT_3[45890] = 32'b00000000000000000100101101010000;
assign LUT_3[45891] = 32'b00000000000000001011011000101101;
assign LUT_3[45892] = 32'b11111111111111111111110011100010;
assign LUT_3[45893] = 32'b00000000000000000110011110111111;
assign LUT_3[45894] = 32'b00000000000000000001111011000110;
assign LUT_3[45895] = 32'b00000000000000001000100110100011;
assign LUT_3[45896] = 32'b00000000000000000111111110110010;
assign LUT_3[45897] = 32'b00000000000000001110101010001111;
assign LUT_3[45898] = 32'b00000000000000001010000110010110;
assign LUT_3[45899] = 32'b00000000000000010000110001110011;
assign LUT_3[45900] = 32'b00000000000000000101001100101000;
assign LUT_3[45901] = 32'b00000000000000001011111000000101;
assign LUT_3[45902] = 32'b00000000000000000111010100001100;
assign LUT_3[45903] = 32'b00000000000000001101111111101001;
assign LUT_3[45904] = 32'b00000000000000000101111000101111;
assign LUT_3[45905] = 32'b00000000000000001100100100001100;
assign LUT_3[45906] = 32'b00000000000000001000000000010011;
assign LUT_3[45907] = 32'b00000000000000001110101011110000;
assign LUT_3[45908] = 32'b00000000000000000011000110100101;
assign LUT_3[45909] = 32'b00000000000000001001110010000010;
assign LUT_3[45910] = 32'b00000000000000000101001110001001;
assign LUT_3[45911] = 32'b00000000000000001011111001100110;
assign LUT_3[45912] = 32'b00000000000000001011010001110101;
assign LUT_3[45913] = 32'b00000000000000010001111101010010;
assign LUT_3[45914] = 32'b00000000000000001101011001011001;
assign LUT_3[45915] = 32'b00000000000000010100000100110110;
assign LUT_3[45916] = 32'b00000000000000001000011111101011;
assign LUT_3[45917] = 32'b00000000000000001111001011001000;
assign LUT_3[45918] = 32'b00000000000000001010100111001111;
assign LUT_3[45919] = 32'b00000000000000010001010010101100;
assign LUT_3[45920] = 32'b00000000000000000011110100001100;
assign LUT_3[45921] = 32'b00000000000000001010011111101001;
assign LUT_3[45922] = 32'b00000000000000000101111011110000;
assign LUT_3[45923] = 32'b00000000000000001100100111001101;
assign LUT_3[45924] = 32'b00000000000000000001000010000010;
assign LUT_3[45925] = 32'b00000000000000000111101101011111;
assign LUT_3[45926] = 32'b00000000000000000011001001100110;
assign LUT_3[45927] = 32'b00000000000000001001110101000011;
assign LUT_3[45928] = 32'b00000000000000001001001101010010;
assign LUT_3[45929] = 32'b00000000000000001111111000101111;
assign LUT_3[45930] = 32'b00000000000000001011010100110110;
assign LUT_3[45931] = 32'b00000000000000010010000000010011;
assign LUT_3[45932] = 32'b00000000000000000110011011001000;
assign LUT_3[45933] = 32'b00000000000000001101000110100101;
assign LUT_3[45934] = 32'b00000000000000001000100010101100;
assign LUT_3[45935] = 32'b00000000000000001111001110001001;
assign LUT_3[45936] = 32'b00000000000000000111000111001111;
assign LUT_3[45937] = 32'b00000000000000001101110010101100;
assign LUT_3[45938] = 32'b00000000000000001001001110110011;
assign LUT_3[45939] = 32'b00000000000000001111111010010000;
assign LUT_3[45940] = 32'b00000000000000000100010101000101;
assign LUT_3[45941] = 32'b00000000000000001011000000100010;
assign LUT_3[45942] = 32'b00000000000000000110011100101001;
assign LUT_3[45943] = 32'b00000000000000001101001000000110;
assign LUT_3[45944] = 32'b00000000000000001100100000010101;
assign LUT_3[45945] = 32'b00000000000000010011001011110010;
assign LUT_3[45946] = 32'b00000000000000001110100111111001;
assign LUT_3[45947] = 32'b00000000000000010101010011010110;
assign LUT_3[45948] = 32'b00000000000000001001101110001011;
assign LUT_3[45949] = 32'b00000000000000010000011001101000;
assign LUT_3[45950] = 32'b00000000000000001011110101101111;
assign LUT_3[45951] = 32'b00000000000000010010100001001100;
assign LUT_3[45952] = 32'b00000000000000000100110111111111;
assign LUT_3[45953] = 32'b00000000000000001011100011011100;
assign LUT_3[45954] = 32'b00000000000000000110111111100011;
assign LUT_3[45955] = 32'b00000000000000001101101011000000;
assign LUT_3[45956] = 32'b00000000000000000010000101110101;
assign LUT_3[45957] = 32'b00000000000000001000110001010010;
assign LUT_3[45958] = 32'b00000000000000000100001101011001;
assign LUT_3[45959] = 32'b00000000000000001010111000110110;
assign LUT_3[45960] = 32'b00000000000000001010010001000101;
assign LUT_3[45961] = 32'b00000000000000010000111100100010;
assign LUT_3[45962] = 32'b00000000000000001100011000101001;
assign LUT_3[45963] = 32'b00000000000000010011000100000110;
assign LUT_3[45964] = 32'b00000000000000000111011110111011;
assign LUT_3[45965] = 32'b00000000000000001110001010011000;
assign LUT_3[45966] = 32'b00000000000000001001100110011111;
assign LUT_3[45967] = 32'b00000000000000010000010001111100;
assign LUT_3[45968] = 32'b00000000000000001000001011000010;
assign LUT_3[45969] = 32'b00000000000000001110110110011111;
assign LUT_3[45970] = 32'b00000000000000001010010010100110;
assign LUT_3[45971] = 32'b00000000000000010000111110000011;
assign LUT_3[45972] = 32'b00000000000000000101011000111000;
assign LUT_3[45973] = 32'b00000000000000001100000100010101;
assign LUT_3[45974] = 32'b00000000000000000111100000011100;
assign LUT_3[45975] = 32'b00000000000000001110001011111001;
assign LUT_3[45976] = 32'b00000000000000001101100100001000;
assign LUT_3[45977] = 32'b00000000000000010100001111100101;
assign LUT_3[45978] = 32'b00000000000000001111101011101100;
assign LUT_3[45979] = 32'b00000000000000010110010111001001;
assign LUT_3[45980] = 32'b00000000000000001010110001111110;
assign LUT_3[45981] = 32'b00000000000000010001011101011011;
assign LUT_3[45982] = 32'b00000000000000001100111001100010;
assign LUT_3[45983] = 32'b00000000000000010011100100111111;
assign LUT_3[45984] = 32'b00000000000000000110000110011111;
assign LUT_3[45985] = 32'b00000000000000001100110001111100;
assign LUT_3[45986] = 32'b00000000000000001000001110000011;
assign LUT_3[45987] = 32'b00000000000000001110111001100000;
assign LUT_3[45988] = 32'b00000000000000000011010100010101;
assign LUT_3[45989] = 32'b00000000000000001001111111110010;
assign LUT_3[45990] = 32'b00000000000000000101011011111001;
assign LUT_3[45991] = 32'b00000000000000001100000111010110;
assign LUT_3[45992] = 32'b00000000000000001011011111100101;
assign LUT_3[45993] = 32'b00000000000000010010001011000010;
assign LUT_3[45994] = 32'b00000000000000001101100111001001;
assign LUT_3[45995] = 32'b00000000000000010100010010100110;
assign LUT_3[45996] = 32'b00000000000000001000101101011011;
assign LUT_3[45997] = 32'b00000000000000001111011000111000;
assign LUT_3[45998] = 32'b00000000000000001010110100111111;
assign LUT_3[45999] = 32'b00000000000000010001100000011100;
assign LUT_3[46000] = 32'b00000000000000001001011001100010;
assign LUT_3[46001] = 32'b00000000000000010000000100111111;
assign LUT_3[46002] = 32'b00000000000000001011100001000110;
assign LUT_3[46003] = 32'b00000000000000010010001100100011;
assign LUT_3[46004] = 32'b00000000000000000110100111011000;
assign LUT_3[46005] = 32'b00000000000000001101010010110101;
assign LUT_3[46006] = 32'b00000000000000001000101110111100;
assign LUT_3[46007] = 32'b00000000000000001111011010011001;
assign LUT_3[46008] = 32'b00000000000000001110110010101000;
assign LUT_3[46009] = 32'b00000000000000010101011110000101;
assign LUT_3[46010] = 32'b00000000000000010000111010001100;
assign LUT_3[46011] = 32'b00000000000000010111100101101001;
assign LUT_3[46012] = 32'b00000000000000001100000000011110;
assign LUT_3[46013] = 32'b00000000000000010010101011111011;
assign LUT_3[46014] = 32'b00000000000000001110001000000010;
assign LUT_3[46015] = 32'b00000000000000010100110011011111;
assign LUT_3[46016] = 32'b00000000000000000100110000101010;
assign LUT_3[46017] = 32'b00000000000000001011011100000111;
assign LUT_3[46018] = 32'b00000000000000000110111000001110;
assign LUT_3[46019] = 32'b00000000000000001101100011101011;
assign LUT_3[46020] = 32'b00000000000000000001111110100000;
assign LUT_3[46021] = 32'b00000000000000001000101001111101;
assign LUT_3[46022] = 32'b00000000000000000100000110000100;
assign LUT_3[46023] = 32'b00000000000000001010110001100001;
assign LUT_3[46024] = 32'b00000000000000001010001001110000;
assign LUT_3[46025] = 32'b00000000000000010000110101001101;
assign LUT_3[46026] = 32'b00000000000000001100010001010100;
assign LUT_3[46027] = 32'b00000000000000010010111100110001;
assign LUT_3[46028] = 32'b00000000000000000111010111100110;
assign LUT_3[46029] = 32'b00000000000000001110000011000011;
assign LUT_3[46030] = 32'b00000000000000001001011111001010;
assign LUT_3[46031] = 32'b00000000000000010000001010100111;
assign LUT_3[46032] = 32'b00000000000000001000000011101101;
assign LUT_3[46033] = 32'b00000000000000001110101111001010;
assign LUT_3[46034] = 32'b00000000000000001010001011010001;
assign LUT_3[46035] = 32'b00000000000000010000110110101110;
assign LUT_3[46036] = 32'b00000000000000000101010001100011;
assign LUT_3[46037] = 32'b00000000000000001011111101000000;
assign LUT_3[46038] = 32'b00000000000000000111011001000111;
assign LUT_3[46039] = 32'b00000000000000001110000100100100;
assign LUT_3[46040] = 32'b00000000000000001101011100110011;
assign LUT_3[46041] = 32'b00000000000000010100001000010000;
assign LUT_3[46042] = 32'b00000000000000001111100100010111;
assign LUT_3[46043] = 32'b00000000000000010110001111110100;
assign LUT_3[46044] = 32'b00000000000000001010101010101001;
assign LUT_3[46045] = 32'b00000000000000010001010110000110;
assign LUT_3[46046] = 32'b00000000000000001100110010001101;
assign LUT_3[46047] = 32'b00000000000000010011011101101010;
assign LUT_3[46048] = 32'b00000000000000000101111111001010;
assign LUT_3[46049] = 32'b00000000000000001100101010100111;
assign LUT_3[46050] = 32'b00000000000000001000000110101110;
assign LUT_3[46051] = 32'b00000000000000001110110010001011;
assign LUT_3[46052] = 32'b00000000000000000011001101000000;
assign LUT_3[46053] = 32'b00000000000000001001111000011101;
assign LUT_3[46054] = 32'b00000000000000000101010100100100;
assign LUT_3[46055] = 32'b00000000000000001100000000000001;
assign LUT_3[46056] = 32'b00000000000000001011011000010000;
assign LUT_3[46057] = 32'b00000000000000010010000011101101;
assign LUT_3[46058] = 32'b00000000000000001101011111110100;
assign LUT_3[46059] = 32'b00000000000000010100001011010001;
assign LUT_3[46060] = 32'b00000000000000001000100110000110;
assign LUT_3[46061] = 32'b00000000000000001111010001100011;
assign LUT_3[46062] = 32'b00000000000000001010101101101010;
assign LUT_3[46063] = 32'b00000000000000010001011001000111;
assign LUT_3[46064] = 32'b00000000000000001001010010001101;
assign LUT_3[46065] = 32'b00000000000000001111111101101010;
assign LUT_3[46066] = 32'b00000000000000001011011001110001;
assign LUT_3[46067] = 32'b00000000000000010010000101001110;
assign LUT_3[46068] = 32'b00000000000000000110100000000011;
assign LUT_3[46069] = 32'b00000000000000001101001011100000;
assign LUT_3[46070] = 32'b00000000000000001000100111100111;
assign LUT_3[46071] = 32'b00000000000000001111010011000100;
assign LUT_3[46072] = 32'b00000000000000001110101011010011;
assign LUT_3[46073] = 32'b00000000000000010101010110110000;
assign LUT_3[46074] = 32'b00000000000000010000110010110111;
assign LUT_3[46075] = 32'b00000000000000010111011110010100;
assign LUT_3[46076] = 32'b00000000000000001011111001001001;
assign LUT_3[46077] = 32'b00000000000000010010100100100110;
assign LUT_3[46078] = 32'b00000000000000001110000000101101;
assign LUT_3[46079] = 32'b00000000000000010100101100001010;
assign LUT_3[46080] = 32'b00000000000000001001101101010001;
assign LUT_3[46081] = 32'b00000000000000010000011000101110;
assign LUT_3[46082] = 32'b00000000000000001011110100110101;
assign LUT_3[46083] = 32'b00000000000000010010100000010010;
assign LUT_3[46084] = 32'b00000000000000000110111011000111;
assign LUT_3[46085] = 32'b00000000000000001101100110100100;
assign LUT_3[46086] = 32'b00000000000000001001000010101011;
assign LUT_3[46087] = 32'b00000000000000001111101110001000;
assign LUT_3[46088] = 32'b00000000000000001111000110010111;
assign LUT_3[46089] = 32'b00000000000000010101110001110100;
assign LUT_3[46090] = 32'b00000000000000010001001101111011;
assign LUT_3[46091] = 32'b00000000000000010111111001011000;
assign LUT_3[46092] = 32'b00000000000000001100010100001101;
assign LUT_3[46093] = 32'b00000000000000010010111111101010;
assign LUT_3[46094] = 32'b00000000000000001110011011110001;
assign LUT_3[46095] = 32'b00000000000000010101000111001110;
assign LUT_3[46096] = 32'b00000000000000001101000000010100;
assign LUT_3[46097] = 32'b00000000000000010011101011110001;
assign LUT_3[46098] = 32'b00000000000000001111000111111000;
assign LUT_3[46099] = 32'b00000000000000010101110011010101;
assign LUT_3[46100] = 32'b00000000000000001010001110001010;
assign LUT_3[46101] = 32'b00000000000000010000111001100111;
assign LUT_3[46102] = 32'b00000000000000001100010101101110;
assign LUT_3[46103] = 32'b00000000000000010011000001001011;
assign LUT_3[46104] = 32'b00000000000000010010011001011010;
assign LUT_3[46105] = 32'b00000000000000011001000100110111;
assign LUT_3[46106] = 32'b00000000000000010100100000111110;
assign LUT_3[46107] = 32'b00000000000000011011001100011011;
assign LUT_3[46108] = 32'b00000000000000001111100111010000;
assign LUT_3[46109] = 32'b00000000000000010110010010101101;
assign LUT_3[46110] = 32'b00000000000000010001101110110100;
assign LUT_3[46111] = 32'b00000000000000011000011010010001;
assign LUT_3[46112] = 32'b00000000000000001010111011110001;
assign LUT_3[46113] = 32'b00000000000000010001100111001110;
assign LUT_3[46114] = 32'b00000000000000001101000011010101;
assign LUT_3[46115] = 32'b00000000000000010011101110110010;
assign LUT_3[46116] = 32'b00000000000000001000001001100111;
assign LUT_3[46117] = 32'b00000000000000001110110101000100;
assign LUT_3[46118] = 32'b00000000000000001010010001001011;
assign LUT_3[46119] = 32'b00000000000000010000111100101000;
assign LUT_3[46120] = 32'b00000000000000010000010100110111;
assign LUT_3[46121] = 32'b00000000000000010111000000010100;
assign LUT_3[46122] = 32'b00000000000000010010011100011011;
assign LUT_3[46123] = 32'b00000000000000011001000111111000;
assign LUT_3[46124] = 32'b00000000000000001101100010101101;
assign LUT_3[46125] = 32'b00000000000000010100001110001010;
assign LUT_3[46126] = 32'b00000000000000001111101010010001;
assign LUT_3[46127] = 32'b00000000000000010110010101101110;
assign LUT_3[46128] = 32'b00000000000000001110001110110100;
assign LUT_3[46129] = 32'b00000000000000010100111010010001;
assign LUT_3[46130] = 32'b00000000000000010000010110011000;
assign LUT_3[46131] = 32'b00000000000000010111000001110101;
assign LUT_3[46132] = 32'b00000000000000001011011100101010;
assign LUT_3[46133] = 32'b00000000000000010010001000000111;
assign LUT_3[46134] = 32'b00000000000000001101100100001110;
assign LUT_3[46135] = 32'b00000000000000010100001111101011;
assign LUT_3[46136] = 32'b00000000000000010011100111111010;
assign LUT_3[46137] = 32'b00000000000000011010010011010111;
assign LUT_3[46138] = 32'b00000000000000010101101111011110;
assign LUT_3[46139] = 32'b00000000000000011100011010111011;
assign LUT_3[46140] = 32'b00000000000000010000110101110000;
assign LUT_3[46141] = 32'b00000000000000010111100001001101;
assign LUT_3[46142] = 32'b00000000000000010010111101010100;
assign LUT_3[46143] = 32'b00000000000000011001101000110001;
assign LUT_3[46144] = 32'b00000000000000001001100101111100;
assign LUT_3[46145] = 32'b00000000000000010000010001011001;
assign LUT_3[46146] = 32'b00000000000000001011101101100000;
assign LUT_3[46147] = 32'b00000000000000010010011000111101;
assign LUT_3[46148] = 32'b00000000000000000110110011110010;
assign LUT_3[46149] = 32'b00000000000000001101011111001111;
assign LUT_3[46150] = 32'b00000000000000001000111011010110;
assign LUT_3[46151] = 32'b00000000000000001111100110110011;
assign LUT_3[46152] = 32'b00000000000000001110111111000010;
assign LUT_3[46153] = 32'b00000000000000010101101010011111;
assign LUT_3[46154] = 32'b00000000000000010001000110100110;
assign LUT_3[46155] = 32'b00000000000000010111110010000011;
assign LUT_3[46156] = 32'b00000000000000001100001100111000;
assign LUT_3[46157] = 32'b00000000000000010010111000010101;
assign LUT_3[46158] = 32'b00000000000000001110010100011100;
assign LUT_3[46159] = 32'b00000000000000010100111111111001;
assign LUT_3[46160] = 32'b00000000000000001100111000111111;
assign LUT_3[46161] = 32'b00000000000000010011100100011100;
assign LUT_3[46162] = 32'b00000000000000001111000000100011;
assign LUT_3[46163] = 32'b00000000000000010101101100000000;
assign LUT_3[46164] = 32'b00000000000000001010000110110101;
assign LUT_3[46165] = 32'b00000000000000010000110010010010;
assign LUT_3[46166] = 32'b00000000000000001100001110011001;
assign LUT_3[46167] = 32'b00000000000000010010111001110110;
assign LUT_3[46168] = 32'b00000000000000010010010010000101;
assign LUT_3[46169] = 32'b00000000000000011000111101100010;
assign LUT_3[46170] = 32'b00000000000000010100011001101001;
assign LUT_3[46171] = 32'b00000000000000011011000101000110;
assign LUT_3[46172] = 32'b00000000000000001111011111111011;
assign LUT_3[46173] = 32'b00000000000000010110001011011000;
assign LUT_3[46174] = 32'b00000000000000010001100111011111;
assign LUT_3[46175] = 32'b00000000000000011000010010111100;
assign LUT_3[46176] = 32'b00000000000000001010110100011100;
assign LUT_3[46177] = 32'b00000000000000010001011111111001;
assign LUT_3[46178] = 32'b00000000000000001100111100000000;
assign LUT_3[46179] = 32'b00000000000000010011100111011101;
assign LUT_3[46180] = 32'b00000000000000001000000010010010;
assign LUT_3[46181] = 32'b00000000000000001110101101101111;
assign LUT_3[46182] = 32'b00000000000000001010001001110110;
assign LUT_3[46183] = 32'b00000000000000010000110101010011;
assign LUT_3[46184] = 32'b00000000000000010000001101100010;
assign LUT_3[46185] = 32'b00000000000000010110111000111111;
assign LUT_3[46186] = 32'b00000000000000010010010101000110;
assign LUT_3[46187] = 32'b00000000000000011001000000100011;
assign LUT_3[46188] = 32'b00000000000000001101011011011000;
assign LUT_3[46189] = 32'b00000000000000010100000110110101;
assign LUT_3[46190] = 32'b00000000000000001111100010111100;
assign LUT_3[46191] = 32'b00000000000000010110001110011001;
assign LUT_3[46192] = 32'b00000000000000001110000111011111;
assign LUT_3[46193] = 32'b00000000000000010100110010111100;
assign LUT_3[46194] = 32'b00000000000000010000001111000011;
assign LUT_3[46195] = 32'b00000000000000010110111010100000;
assign LUT_3[46196] = 32'b00000000000000001011010101010101;
assign LUT_3[46197] = 32'b00000000000000010010000000110010;
assign LUT_3[46198] = 32'b00000000000000001101011100111001;
assign LUT_3[46199] = 32'b00000000000000010100001000010110;
assign LUT_3[46200] = 32'b00000000000000010011100000100101;
assign LUT_3[46201] = 32'b00000000000000011010001100000010;
assign LUT_3[46202] = 32'b00000000000000010101101000001001;
assign LUT_3[46203] = 32'b00000000000000011100010011100110;
assign LUT_3[46204] = 32'b00000000000000010000101110011011;
assign LUT_3[46205] = 32'b00000000000000010111011001111000;
assign LUT_3[46206] = 32'b00000000000000010010110101111111;
assign LUT_3[46207] = 32'b00000000000000011001100001011100;
assign LUT_3[46208] = 32'b00000000000000001011111000001111;
assign LUT_3[46209] = 32'b00000000000000010010100011101100;
assign LUT_3[46210] = 32'b00000000000000001101111111110011;
assign LUT_3[46211] = 32'b00000000000000010100101011010000;
assign LUT_3[46212] = 32'b00000000000000001001000110000101;
assign LUT_3[46213] = 32'b00000000000000001111110001100010;
assign LUT_3[46214] = 32'b00000000000000001011001101101001;
assign LUT_3[46215] = 32'b00000000000000010001111001000110;
assign LUT_3[46216] = 32'b00000000000000010001010001010101;
assign LUT_3[46217] = 32'b00000000000000010111111100110010;
assign LUT_3[46218] = 32'b00000000000000010011011000111001;
assign LUT_3[46219] = 32'b00000000000000011010000100010110;
assign LUT_3[46220] = 32'b00000000000000001110011111001011;
assign LUT_3[46221] = 32'b00000000000000010101001010101000;
assign LUT_3[46222] = 32'b00000000000000010000100110101111;
assign LUT_3[46223] = 32'b00000000000000010111010010001100;
assign LUT_3[46224] = 32'b00000000000000001111001011010010;
assign LUT_3[46225] = 32'b00000000000000010101110110101111;
assign LUT_3[46226] = 32'b00000000000000010001010010110110;
assign LUT_3[46227] = 32'b00000000000000010111111110010011;
assign LUT_3[46228] = 32'b00000000000000001100011001001000;
assign LUT_3[46229] = 32'b00000000000000010011000100100101;
assign LUT_3[46230] = 32'b00000000000000001110100000101100;
assign LUT_3[46231] = 32'b00000000000000010101001100001001;
assign LUT_3[46232] = 32'b00000000000000010100100100011000;
assign LUT_3[46233] = 32'b00000000000000011011001111110101;
assign LUT_3[46234] = 32'b00000000000000010110101011111100;
assign LUT_3[46235] = 32'b00000000000000011101010111011001;
assign LUT_3[46236] = 32'b00000000000000010001110010001110;
assign LUT_3[46237] = 32'b00000000000000011000011101101011;
assign LUT_3[46238] = 32'b00000000000000010011111001110010;
assign LUT_3[46239] = 32'b00000000000000011010100101001111;
assign LUT_3[46240] = 32'b00000000000000001101000110101111;
assign LUT_3[46241] = 32'b00000000000000010011110010001100;
assign LUT_3[46242] = 32'b00000000000000001111001110010011;
assign LUT_3[46243] = 32'b00000000000000010101111001110000;
assign LUT_3[46244] = 32'b00000000000000001010010100100101;
assign LUT_3[46245] = 32'b00000000000000010001000000000010;
assign LUT_3[46246] = 32'b00000000000000001100011100001001;
assign LUT_3[46247] = 32'b00000000000000010011000111100110;
assign LUT_3[46248] = 32'b00000000000000010010011111110101;
assign LUT_3[46249] = 32'b00000000000000011001001011010010;
assign LUT_3[46250] = 32'b00000000000000010100100111011001;
assign LUT_3[46251] = 32'b00000000000000011011010010110110;
assign LUT_3[46252] = 32'b00000000000000001111101101101011;
assign LUT_3[46253] = 32'b00000000000000010110011001001000;
assign LUT_3[46254] = 32'b00000000000000010001110101001111;
assign LUT_3[46255] = 32'b00000000000000011000100000101100;
assign LUT_3[46256] = 32'b00000000000000010000011001110010;
assign LUT_3[46257] = 32'b00000000000000010111000101001111;
assign LUT_3[46258] = 32'b00000000000000010010100001010110;
assign LUT_3[46259] = 32'b00000000000000011001001100110011;
assign LUT_3[46260] = 32'b00000000000000001101100111101000;
assign LUT_3[46261] = 32'b00000000000000010100010011000101;
assign LUT_3[46262] = 32'b00000000000000001111101111001100;
assign LUT_3[46263] = 32'b00000000000000010110011010101001;
assign LUT_3[46264] = 32'b00000000000000010101110010111000;
assign LUT_3[46265] = 32'b00000000000000011100011110010101;
assign LUT_3[46266] = 32'b00000000000000010111111010011100;
assign LUT_3[46267] = 32'b00000000000000011110100101111001;
assign LUT_3[46268] = 32'b00000000000000010011000000101110;
assign LUT_3[46269] = 32'b00000000000000011001101100001011;
assign LUT_3[46270] = 32'b00000000000000010101001000010010;
assign LUT_3[46271] = 32'b00000000000000011011110011101111;
assign LUT_3[46272] = 32'b00000000000000001011110000111010;
assign LUT_3[46273] = 32'b00000000000000010010011100010111;
assign LUT_3[46274] = 32'b00000000000000001101111000011110;
assign LUT_3[46275] = 32'b00000000000000010100100011111011;
assign LUT_3[46276] = 32'b00000000000000001000111110110000;
assign LUT_3[46277] = 32'b00000000000000001111101010001101;
assign LUT_3[46278] = 32'b00000000000000001011000110010100;
assign LUT_3[46279] = 32'b00000000000000010001110001110001;
assign LUT_3[46280] = 32'b00000000000000010001001010000000;
assign LUT_3[46281] = 32'b00000000000000010111110101011101;
assign LUT_3[46282] = 32'b00000000000000010011010001100100;
assign LUT_3[46283] = 32'b00000000000000011001111101000001;
assign LUT_3[46284] = 32'b00000000000000001110010111110110;
assign LUT_3[46285] = 32'b00000000000000010101000011010011;
assign LUT_3[46286] = 32'b00000000000000010000011111011010;
assign LUT_3[46287] = 32'b00000000000000010111001010110111;
assign LUT_3[46288] = 32'b00000000000000001111000011111101;
assign LUT_3[46289] = 32'b00000000000000010101101111011010;
assign LUT_3[46290] = 32'b00000000000000010001001011100001;
assign LUT_3[46291] = 32'b00000000000000010111110110111110;
assign LUT_3[46292] = 32'b00000000000000001100010001110011;
assign LUT_3[46293] = 32'b00000000000000010010111101010000;
assign LUT_3[46294] = 32'b00000000000000001110011001010111;
assign LUT_3[46295] = 32'b00000000000000010101000100110100;
assign LUT_3[46296] = 32'b00000000000000010100011101000011;
assign LUT_3[46297] = 32'b00000000000000011011001000100000;
assign LUT_3[46298] = 32'b00000000000000010110100100100111;
assign LUT_3[46299] = 32'b00000000000000011101010000000100;
assign LUT_3[46300] = 32'b00000000000000010001101010111001;
assign LUT_3[46301] = 32'b00000000000000011000010110010110;
assign LUT_3[46302] = 32'b00000000000000010011110010011101;
assign LUT_3[46303] = 32'b00000000000000011010011101111010;
assign LUT_3[46304] = 32'b00000000000000001100111111011010;
assign LUT_3[46305] = 32'b00000000000000010011101010110111;
assign LUT_3[46306] = 32'b00000000000000001111000110111110;
assign LUT_3[46307] = 32'b00000000000000010101110010011011;
assign LUT_3[46308] = 32'b00000000000000001010001101010000;
assign LUT_3[46309] = 32'b00000000000000010000111000101101;
assign LUT_3[46310] = 32'b00000000000000001100010100110100;
assign LUT_3[46311] = 32'b00000000000000010011000000010001;
assign LUT_3[46312] = 32'b00000000000000010010011000100000;
assign LUT_3[46313] = 32'b00000000000000011001000011111101;
assign LUT_3[46314] = 32'b00000000000000010100100000000100;
assign LUT_3[46315] = 32'b00000000000000011011001011100001;
assign LUT_3[46316] = 32'b00000000000000001111100110010110;
assign LUT_3[46317] = 32'b00000000000000010110010001110011;
assign LUT_3[46318] = 32'b00000000000000010001101101111010;
assign LUT_3[46319] = 32'b00000000000000011000011001010111;
assign LUT_3[46320] = 32'b00000000000000010000010010011101;
assign LUT_3[46321] = 32'b00000000000000010110111101111010;
assign LUT_3[46322] = 32'b00000000000000010010011010000001;
assign LUT_3[46323] = 32'b00000000000000011001000101011110;
assign LUT_3[46324] = 32'b00000000000000001101100000010011;
assign LUT_3[46325] = 32'b00000000000000010100001011110000;
assign LUT_3[46326] = 32'b00000000000000001111100111110111;
assign LUT_3[46327] = 32'b00000000000000010110010011010100;
assign LUT_3[46328] = 32'b00000000000000010101101011100011;
assign LUT_3[46329] = 32'b00000000000000011100010111000000;
assign LUT_3[46330] = 32'b00000000000000010111110011000111;
assign LUT_3[46331] = 32'b00000000000000011110011110100100;
assign LUT_3[46332] = 32'b00000000000000010010111001011001;
assign LUT_3[46333] = 32'b00000000000000011001100100110110;
assign LUT_3[46334] = 32'b00000000000000010101000000111101;
assign LUT_3[46335] = 32'b00000000000000011011101100011010;
assign LUT_3[46336] = 32'b00000000000000000101111100110010;
assign LUT_3[46337] = 32'b00000000000000001100101000001111;
assign LUT_3[46338] = 32'b00000000000000001000000100010110;
assign LUT_3[46339] = 32'b00000000000000001110101111110011;
assign LUT_3[46340] = 32'b00000000000000000011001010101000;
assign LUT_3[46341] = 32'b00000000000000001001110110000101;
assign LUT_3[46342] = 32'b00000000000000000101010010001100;
assign LUT_3[46343] = 32'b00000000000000001011111101101001;
assign LUT_3[46344] = 32'b00000000000000001011010101111000;
assign LUT_3[46345] = 32'b00000000000000010010000001010101;
assign LUT_3[46346] = 32'b00000000000000001101011101011100;
assign LUT_3[46347] = 32'b00000000000000010100001000111001;
assign LUT_3[46348] = 32'b00000000000000001000100011101110;
assign LUT_3[46349] = 32'b00000000000000001111001111001011;
assign LUT_3[46350] = 32'b00000000000000001010101011010010;
assign LUT_3[46351] = 32'b00000000000000010001010110101111;
assign LUT_3[46352] = 32'b00000000000000001001001111110101;
assign LUT_3[46353] = 32'b00000000000000001111111011010010;
assign LUT_3[46354] = 32'b00000000000000001011010111011001;
assign LUT_3[46355] = 32'b00000000000000010010000010110110;
assign LUT_3[46356] = 32'b00000000000000000110011101101011;
assign LUT_3[46357] = 32'b00000000000000001101001001001000;
assign LUT_3[46358] = 32'b00000000000000001000100101001111;
assign LUT_3[46359] = 32'b00000000000000001111010000101100;
assign LUT_3[46360] = 32'b00000000000000001110101000111011;
assign LUT_3[46361] = 32'b00000000000000010101010100011000;
assign LUT_3[46362] = 32'b00000000000000010000110000011111;
assign LUT_3[46363] = 32'b00000000000000010111011011111100;
assign LUT_3[46364] = 32'b00000000000000001011110110110001;
assign LUT_3[46365] = 32'b00000000000000010010100010001110;
assign LUT_3[46366] = 32'b00000000000000001101111110010101;
assign LUT_3[46367] = 32'b00000000000000010100101001110010;
assign LUT_3[46368] = 32'b00000000000000000111001011010010;
assign LUT_3[46369] = 32'b00000000000000001101110110101111;
assign LUT_3[46370] = 32'b00000000000000001001010010110110;
assign LUT_3[46371] = 32'b00000000000000001111111110010011;
assign LUT_3[46372] = 32'b00000000000000000100011001001000;
assign LUT_3[46373] = 32'b00000000000000001011000100100101;
assign LUT_3[46374] = 32'b00000000000000000110100000101100;
assign LUT_3[46375] = 32'b00000000000000001101001100001001;
assign LUT_3[46376] = 32'b00000000000000001100100100011000;
assign LUT_3[46377] = 32'b00000000000000010011001111110101;
assign LUT_3[46378] = 32'b00000000000000001110101011111100;
assign LUT_3[46379] = 32'b00000000000000010101010111011001;
assign LUT_3[46380] = 32'b00000000000000001001110010001110;
assign LUT_3[46381] = 32'b00000000000000010000011101101011;
assign LUT_3[46382] = 32'b00000000000000001011111001110010;
assign LUT_3[46383] = 32'b00000000000000010010100101001111;
assign LUT_3[46384] = 32'b00000000000000001010011110010101;
assign LUT_3[46385] = 32'b00000000000000010001001001110010;
assign LUT_3[46386] = 32'b00000000000000001100100101111001;
assign LUT_3[46387] = 32'b00000000000000010011010001010110;
assign LUT_3[46388] = 32'b00000000000000000111101100001011;
assign LUT_3[46389] = 32'b00000000000000001110010111101000;
assign LUT_3[46390] = 32'b00000000000000001001110011101111;
assign LUT_3[46391] = 32'b00000000000000010000011111001100;
assign LUT_3[46392] = 32'b00000000000000001111110111011011;
assign LUT_3[46393] = 32'b00000000000000010110100010111000;
assign LUT_3[46394] = 32'b00000000000000010001111110111111;
assign LUT_3[46395] = 32'b00000000000000011000101010011100;
assign LUT_3[46396] = 32'b00000000000000001101000101010001;
assign LUT_3[46397] = 32'b00000000000000010011110000101110;
assign LUT_3[46398] = 32'b00000000000000001111001100110101;
assign LUT_3[46399] = 32'b00000000000000010101111000010010;
assign LUT_3[46400] = 32'b00000000000000000101110101011101;
assign LUT_3[46401] = 32'b00000000000000001100100000111010;
assign LUT_3[46402] = 32'b00000000000000000111111101000001;
assign LUT_3[46403] = 32'b00000000000000001110101000011110;
assign LUT_3[46404] = 32'b00000000000000000011000011010011;
assign LUT_3[46405] = 32'b00000000000000001001101110110000;
assign LUT_3[46406] = 32'b00000000000000000101001010110111;
assign LUT_3[46407] = 32'b00000000000000001011110110010100;
assign LUT_3[46408] = 32'b00000000000000001011001110100011;
assign LUT_3[46409] = 32'b00000000000000010001111010000000;
assign LUT_3[46410] = 32'b00000000000000001101010110000111;
assign LUT_3[46411] = 32'b00000000000000010100000001100100;
assign LUT_3[46412] = 32'b00000000000000001000011100011001;
assign LUT_3[46413] = 32'b00000000000000001111000111110110;
assign LUT_3[46414] = 32'b00000000000000001010100011111101;
assign LUT_3[46415] = 32'b00000000000000010001001111011010;
assign LUT_3[46416] = 32'b00000000000000001001001000100000;
assign LUT_3[46417] = 32'b00000000000000001111110011111101;
assign LUT_3[46418] = 32'b00000000000000001011010000000100;
assign LUT_3[46419] = 32'b00000000000000010001111011100001;
assign LUT_3[46420] = 32'b00000000000000000110010110010110;
assign LUT_3[46421] = 32'b00000000000000001101000001110011;
assign LUT_3[46422] = 32'b00000000000000001000011101111010;
assign LUT_3[46423] = 32'b00000000000000001111001001010111;
assign LUT_3[46424] = 32'b00000000000000001110100001100110;
assign LUT_3[46425] = 32'b00000000000000010101001101000011;
assign LUT_3[46426] = 32'b00000000000000010000101001001010;
assign LUT_3[46427] = 32'b00000000000000010111010100100111;
assign LUT_3[46428] = 32'b00000000000000001011101111011100;
assign LUT_3[46429] = 32'b00000000000000010010011010111001;
assign LUT_3[46430] = 32'b00000000000000001101110111000000;
assign LUT_3[46431] = 32'b00000000000000010100100010011101;
assign LUT_3[46432] = 32'b00000000000000000111000011111101;
assign LUT_3[46433] = 32'b00000000000000001101101111011010;
assign LUT_3[46434] = 32'b00000000000000001001001011100001;
assign LUT_3[46435] = 32'b00000000000000001111110110111110;
assign LUT_3[46436] = 32'b00000000000000000100010001110011;
assign LUT_3[46437] = 32'b00000000000000001010111101010000;
assign LUT_3[46438] = 32'b00000000000000000110011001010111;
assign LUT_3[46439] = 32'b00000000000000001101000100110100;
assign LUT_3[46440] = 32'b00000000000000001100011101000011;
assign LUT_3[46441] = 32'b00000000000000010011001000100000;
assign LUT_3[46442] = 32'b00000000000000001110100100100111;
assign LUT_3[46443] = 32'b00000000000000010101010000000100;
assign LUT_3[46444] = 32'b00000000000000001001101010111001;
assign LUT_3[46445] = 32'b00000000000000010000010110010110;
assign LUT_3[46446] = 32'b00000000000000001011110010011101;
assign LUT_3[46447] = 32'b00000000000000010010011101111010;
assign LUT_3[46448] = 32'b00000000000000001010010111000000;
assign LUT_3[46449] = 32'b00000000000000010001000010011101;
assign LUT_3[46450] = 32'b00000000000000001100011110100100;
assign LUT_3[46451] = 32'b00000000000000010011001010000001;
assign LUT_3[46452] = 32'b00000000000000000111100100110110;
assign LUT_3[46453] = 32'b00000000000000001110010000010011;
assign LUT_3[46454] = 32'b00000000000000001001101100011010;
assign LUT_3[46455] = 32'b00000000000000010000010111110111;
assign LUT_3[46456] = 32'b00000000000000001111110000000110;
assign LUT_3[46457] = 32'b00000000000000010110011011100011;
assign LUT_3[46458] = 32'b00000000000000010001110111101010;
assign LUT_3[46459] = 32'b00000000000000011000100011000111;
assign LUT_3[46460] = 32'b00000000000000001100111101111100;
assign LUT_3[46461] = 32'b00000000000000010011101001011001;
assign LUT_3[46462] = 32'b00000000000000001111000101100000;
assign LUT_3[46463] = 32'b00000000000000010101110000111101;
assign LUT_3[46464] = 32'b00000000000000001000000111110000;
assign LUT_3[46465] = 32'b00000000000000001110110011001101;
assign LUT_3[46466] = 32'b00000000000000001010001111010100;
assign LUT_3[46467] = 32'b00000000000000010000111010110001;
assign LUT_3[46468] = 32'b00000000000000000101010101100110;
assign LUT_3[46469] = 32'b00000000000000001100000001000011;
assign LUT_3[46470] = 32'b00000000000000000111011101001010;
assign LUT_3[46471] = 32'b00000000000000001110001000100111;
assign LUT_3[46472] = 32'b00000000000000001101100000110110;
assign LUT_3[46473] = 32'b00000000000000010100001100010011;
assign LUT_3[46474] = 32'b00000000000000001111101000011010;
assign LUT_3[46475] = 32'b00000000000000010110010011110111;
assign LUT_3[46476] = 32'b00000000000000001010101110101100;
assign LUT_3[46477] = 32'b00000000000000010001011010001001;
assign LUT_3[46478] = 32'b00000000000000001100110110010000;
assign LUT_3[46479] = 32'b00000000000000010011100001101101;
assign LUT_3[46480] = 32'b00000000000000001011011010110011;
assign LUT_3[46481] = 32'b00000000000000010010000110010000;
assign LUT_3[46482] = 32'b00000000000000001101100010010111;
assign LUT_3[46483] = 32'b00000000000000010100001101110100;
assign LUT_3[46484] = 32'b00000000000000001000101000101001;
assign LUT_3[46485] = 32'b00000000000000001111010100000110;
assign LUT_3[46486] = 32'b00000000000000001010110000001101;
assign LUT_3[46487] = 32'b00000000000000010001011011101010;
assign LUT_3[46488] = 32'b00000000000000010000110011111001;
assign LUT_3[46489] = 32'b00000000000000010111011111010110;
assign LUT_3[46490] = 32'b00000000000000010010111011011101;
assign LUT_3[46491] = 32'b00000000000000011001100110111010;
assign LUT_3[46492] = 32'b00000000000000001110000001101111;
assign LUT_3[46493] = 32'b00000000000000010100101101001100;
assign LUT_3[46494] = 32'b00000000000000010000001001010011;
assign LUT_3[46495] = 32'b00000000000000010110110100110000;
assign LUT_3[46496] = 32'b00000000000000001001010110010000;
assign LUT_3[46497] = 32'b00000000000000010000000001101101;
assign LUT_3[46498] = 32'b00000000000000001011011101110100;
assign LUT_3[46499] = 32'b00000000000000010010001001010001;
assign LUT_3[46500] = 32'b00000000000000000110100100000110;
assign LUT_3[46501] = 32'b00000000000000001101001111100011;
assign LUT_3[46502] = 32'b00000000000000001000101011101010;
assign LUT_3[46503] = 32'b00000000000000001111010111000111;
assign LUT_3[46504] = 32'b00000000000000001110101111010110;
assign LUT_3[46505] = 32'b00000000000000010101011010110011;
assign LUT_3[46506] = 32'b00000000000000010000110110111010;
assign LUT_3[46507] = 32'b00000000000000010111100010010111;
assign LUT_3[46508] = 32'b00000000000000001011111101001100;
assign LUT_3[46509] = 32'b00000000000000010010101000101001;
assign LUT_3[46510] = 32'b00000000000000001110000100110000;
assign LUT_3[46511] = 32'b00000000000000010100110000001101;
assign LUT_3[46512] = 32'b00000000000000001100101001010011;
assign LUT_3[46513] = 32'b00000000000000010011010100110000;
assign LUT_3[46514] = 32'b00000000000000001110110000110111;
assign LUT_3[46515] = 32'b00000000000000010101011100010100;
assign LUT_3[46516] = 32'b00000000000000001001110111001001;
assign LUT_3[46517] = 32'b00000000000000010000100010100110;
assign LUT_3[46518] = 32'b00000000000000001011111110101101;
assign LUT_3[46519] = 32'b00000000000000010010101010001010;
assign LUT_3[46520] = 32'b00000000000000010010000010011001;
assign LUT_3[46521] = 32'b00000000000000011000101101110110;
assign LUT_3[46522] = 32'b00000000000000010100001001111101;
assign LUT_3[46523] = 32'b00000000000000011010110101011010;
assign LUT_3[46524] = 32'b00000000000000001111010000001111;
assign LUT_3[46525] = 32'b00000000000000010101111011101100;
assign LUT_3[46526] = 32'b00000000000000010001010111110011;
assign LUT_3[46527] = 32'b00000000000000011000000011010000;
assign LUT_3[46528] = 32'b00000000000000001000000000011011;
assign LUT_3[46529] = 32'b00000000000000001110101011111000;
assign LUT_3[46530] = 32'b00000000000000001010000111111111;
assign LUT_3[46531] = 32'b00000000000000010000110011011100;
assign LUT_3[46532] = 32'b00000000000000000101001110010001;
assign LUT_3[46533] = 32'b00000000000000001011111001101110;
assign LUT_3[46534] = 32'b00000000000000000111010101110101;
assign LUT_3[46535] = 32'b00000000000000001110000001010010;
assign LUT_3[46536] = 32'b00000000000000001101011001100001;
assign LUT_3[46537] = 32'b00000000000000010100000100111110;
assign LUT_3[46538] = 32'b00000000000000001111100001000101;
assign LUT_3[46539] = 32'b00000000000000010110001100100010;
assign LUT_3[46540] = 32'b00000000000000001010100111010111;
assign LUT_3[46541] = 32'b00000000000000010001010010110100;
assign LUT_3[46542] = 32'b00000000000000001100101110111011;
assign LUT_3[46543] = 32'b00000000000000010011011010011000;
assign LUT_3[46544] = 32'b00000000000000001011010011011110;
assign LUT_3[46545] = 32'b00000000000000010001111110111011;
assign LUT_3[46546] = 32'b00000000000000001101011011000010;
assign LUT_3[46547] = 32'b00000000000000010100000110011111;
assign LUT_3[46548] = 32'b00000000000000001000100001010100;
assign LUT_3[46549] = 32'b00000000000000001111001100110001;
assign LUT_3[46550] = 32'b00000000000000001010101000111000;
assign LUT_3[46551] = 32'b00000000000000010001010100010101;
assign LUT_3[46552] = 32'b00000000000000010000101100100100;
assign LUT_3[46553] = 32'b00000000000000010111011000000001;
assign LUT_3[46554] = 32'b00000000000000010010110100001000;
assign LUT_3[46555] = 32'b00000000000000011001011111100101;
assign LUT_3[46556] = 32'b00000000000000001101111010011010;
assign LUT_3[46557] = 32'b00000000000000010100100101110111;
assign LUT_3[46558] = 32'b00000000000000010000000001111110;
assign LUT_3[46559] = 32'b00000000000000010110101101011011;
assign LUT_3[46560] = 32'b00000000000000001001001110111011;
assign LUT_3[46561] = 32'b00000000000000001111111010011000;
assign LUT_3[46562] = 32'b00000000000000001011010110011111;
assign LUT_3[46563] = 32'b00000000000000010010000001111100;
assign LUT_3[46564] = 32'b00000000000000000110011100110001;
assign LUT_3[46565] = 32'b00000000000000001101001000001110;
assign LUT_3[46566] = 32'b00000000000000001000100100010101;
assign LUT_3[46567] = 32'b00000000000000001111001111110010;
assign LUT_3[46568] = 32'b00000000000000001110101000000001;
assign LUT_3[46569] = 32'b00000000000000010101010011011110;
assign LUT_3[46570] = 32'b00000000000000010000101111100101;
assign LUT_3[46571] = 32'b00000000000000010111011011000010;
assign LUT_3[46572] = 32'b00000000000000001011110101110111;
assign LUT_3[46573] = 32'b00000000000000010010100001010100;
assign LUT_3[46574] = 32'b00000000000000001101111101011011;
assign LUT_3[46575] = 32'b00000000000000010100101000111000;
assign LUT_3[46576] = 32'b00000000000000001100100001111110;
assign LUT_3[46577] = 32'b00000000000000010011001101011011;
assign LUT_3[46578] = 32'b00000000000000001110101001100010;
assign LUT_3[46579] = 32'b00000000000000010101010100111111;
assign LUT_3[46580] = 32'b00000000000000001001101111110100;
assign LUT_3[46581] = 32'b00000000000000010000011011010001;
assign LUT_3[46582] = 32'b00000000000000001011110111011000;
assign LUT_3[46583] = 32'b00000000000000010010100010110101;
assign LUT_3[46584] = 32'b00000000000000010001111011000100;
assign LUT_3[46585] = 32'b00000000000000011000100110100001;
assign LUT_3[46586] = 32'b00000000000000010100000010101000;
assign LUT_3[46587] = 32'b00000000000000011010101110000101;
assign LUT_3[46588] = 32'b00000000000000001111001000111010;
assign LUT_3[46589] = 32'b00000000000000010101110100010111;
assign LUT_3[46590] = 32'b00000000000000010001010000011110;
assign LUT_3[46591] = 32'b00000000000000010111111011111011;
assign LUT_3[46592] = 32'b00000000000000001101000010011101;
assign LUT_3[46593] = 32'b00000000000000010011101101111010;
assign LUT_3[46594] = 32'b00000000000000001111001010000001;
assign LUT_3[46595] = 32'b00000000000000010101110101011110;
assign LUT_3[46596] = 32'b00000000000000001010010000010011;
assign LUT_3[46597] = 32'b00000000000000010000111011110000;
assign LUT_3[46598] = 32'b00000000000000001100010111110111;
assign LUT_3[46599] = 32'b00000000000000010011000011010100;
assign LUT_3[46600] = 32'b00000000000000010010011011100011;
assign LUT_3[46601] = 32'b00000000000000011001000111000000;
assign LUT_3[46602] = 32'b00000000000000010100100011000111;
assign LUT_3[46603] = 32'b00000000000000011011001110100100;
assign LUT_3[46604] = 32'b00000000000000001111101001011001;
assign LUT_3[46605] = 32'b00000000000000010110010100110110;
assign LUT_3[46606] = 32'b00000000000000010001110000111101;
assign LUT_3[46607] = 32'b00000000000000011000011100011010;
assign LUT_3[46608] = 32'b00000000000000010000010101100000;
assign LUT_3[46609] = 32'b00000000000000010111000000111101;
assign LUT_3[46610] = 32'b00000000000000010010011101000100;
assign LUT_3[46611] = 32'b00000000000000011001001000100001;
assign LUT_3[46612] = 32'b00000000000000001101100011010110;
assign LUT_3[46613] = 32'b00000000000000010100001110110011;
assign LUT_3[46614] = 32'b00000000000000001111101010111010;
assign LUT_3[46615] = 32'b00000000000000010110010110010111;
assign LUT_3[46616] = 32'b00000000000000010101101110100110;
assign LUT_3[46617] = 32'b00000000000000011100011010000011;
assign LUT_3[46618] = 32'b00000000000000010111110110001010;
assign LUT_3[46619] = 32'b00000000000000011110100001100111;
assign LUT_3[46620] = 32'b00000000000000010010111100011100;
assign LUT_3[46621] = 32'b00000000000000011001100111111001;
assign LUT_3[46622] = 32'b00000000000000010101000100000000;
assign LUT_3[46623] = 32'b00000000000000011011101111011101;
assign LUT_3[46624] = 32'b00000000000000001110010000111101;
assign LUT_3[46625] = 32'b00000000000000010100111100011010;
assign LUT_3[46626] = 32'b00000000000000010000011000100001;
assign LUT_3[46627] = 32'b00000000000000010111000011111110;
assign LUT_3[46628] = 32'b00000000000000001011011110110011;
assign LUT_3[46629] = 32'b00000000000000010010001010010000;
assign LUT_3[46630] = 32'b00000000000000001101100110010111;
assign LUT_3[46631] = 32'b00000000000000010100010001110100;
assign LUT_3[46632] = 32'b00000000000000010011101010000011;
assign LUT_3[46633] = 32'b00000000000000011010010101100000;
assign LUT_3[46634] = 32'b00000000000000010101110001100111;
assign LUT_3[46635] = 32'b00000000000000011100011101000100;
assign LUT_3[46636] = 32'b00000000000000010000110111111001;
assign LUT_3[46637] = 32'b00000000000000010111100011010110;
assign LUT_3[46638] = 32'b00000000000000010010111111011101;
assign LUT_3[46639] = 32'b00000000000000011001101010111010;
assign LUT_3[46640] = 32'b00000000000000010001100100000000;
assign LUT_3[46641] = 32'b00000000000000011000001111011101;
assign LUT_3[46642] = 32'b00000000000000010011101011100100;
assign LUT_3[46643] = 32'b00000000000000011010010111000001;
assign LUT_3[46644] = 32'b00000000000000001110110001110110;
assign LUT_3[46645] = 32'b00000000000000010101011101010011;
assign LUT_3[46646] = 32'b00000000000000010000111001011010;
assign LUT_3[46647] = 32'b00000000000000010111100100110111;
assign LUT_3[46648] = 32'b00000000000000010110111101000110;
assign LUT_3[46649] = 32'b00000000000000011101101000100011;
assign LUT_3[46650] = 32'b00000000000000011001000100101010;
assign LUT_3[46651] = 32'b00000000000000011111110000000111;
assign LUT_3[46652] = 32'b00000000000000010100001010111100;
assign LUT_3[46653] = 32'b00000000000000011010110110011001;
assign LUT_3[46654] = 32'b00000000000000010110010010100000;
assign LUT_3[46655] = 32'b00000000000000011100111101111101;
assign LUT_3[46656] = 32'b00000000000000001100111011001000;
assign LUT_3[46657] = 32'b00000000000000010011100110100101;
assign LUT_3[46658] = 32'b00000000000000001111000010101100;
assign LUT_3[46659] = 32'b00000000000000010101101110001001;
assign LUT_3[46660] = 32'b00000000000000001010001000111110;
assign LUT_3[46661] = 32'b00000000000000010000110100011011;
assign LUT_3[46662] = 32'b00000000000000001100010000100010;
assign LUT_3[46663] = 32'b00000000000000010010111011111111;
assign LUT_3[46664] = 32'b00000000000000010010010100001110;
assign LUT_3[46665] = 32'b00000000000000011000111111101011;
assign LUT_3[46666] = 32'b00000000000000010100011011110010;
assign LUT_3[46667] = 32'b00000000000000011011000111001111;
assign LUT_3[46668] = 32'b00000000000000001111100010000100;
assign LUT_3[46669] = 32'b00000000000000010110001101100001;
assign LUT_3[46670] = 32'b00000000000000010001101001101000;
assign LUT_3[46671] = 32'b00000000000000011000010101000101;
assign LUT_3[46672] = 32'b00000000000000010000001110001011;
assign LUT_3[46673] = 32'b00000000000000010110111001101000;
assign LUT_3[46674] = 32'b00000000000000010010010101101111;
assign LUT_3[46675] = 32'b00000000000000011001000001001100;
assign LUT_3[46676] = 32'b00000000000000001101011100000001;
assign LUT_3[46677] = 32'b00000000000000010100000111011110;
assign LUT_3[46678] = 32'b00000000000000001111100011100101;
assign LUT_3[46679] = 32'b00000000000000010110001111000010;
assign LUT_3[46680] = 32'b00000000000000010101100111010001;
assign LUT_3[46681] = 32'b00000000000000011100010010101110;
assign LUT_3[46682] = 32'b00000000000000010111101110110101;
assign LUT_3[46683] = 32'b00000000000000011110011010010010;
assign LUT_3[46684] = 32'b00000000000000010010110101000111;
assign LUT_3[46685] = 32'b00000000000000011001100000100100;
assign LUT_3[46686] = 32'b00000000000000010100111100101011;
assign LUT_3[46687] = 32'b00000000000000011011101000001000;
assign LUT_3[46688] = 32'b00000000000000001110001001101000;
assign LUT_3[46689] = 32'b00000000000000010100110101000101;
assign LUT_3[46690] = 32'b00000000000000010000010001001100;
assign LUT_3[46691] = 32'b00000000000000010110111100101001;
assign LUT_3[46692] = 32'b00000000000000001011010111011110;
assign LUT_3[46693] = 32'b00000000000000010010000010111011;
assign LUT_3[46694] = 32'b00000000000000001101011111000010;
assign LUT_3[46695] = 32'b00000000000000010100001010011111;
assign LUT_3[46696] = 32'b00000000000000010011100010101110;
assign LUT_3[46697] = 32'b00000000000000011010001110001011;
assign LUT_3[46698] = 32'b00000000000000010101101010010010;
assign LUT_3[46699] = 32'b00000000000000011100010101101111;
assign LUT_3[46700] = 32'b00000000000000010000110000100100;
assign LUT_3[46701] = 32'b00000000000000010111011100000001;
assign LUT_3[46702] = 32'b00000000000000010010111000001000;
assign LUT_3[46703] = 32'b00000000000000011001100011100101;
assign LUT_3[46704] = 32'b00000000000000010001011100101011;
assign LUT_3[46705] = 32'b00000000000000011000001000001000;
assign LUT_3[46706] = 32'b00000000000000010011100100001111;
assign LUT_3[46707] = 32'b00000000000000011010001111101100;
assign LUT_3[46708] = 32'b00000000000000001110101010100001;
assign LUT_3[46709] = 32'b00000000000000010101010101111110;
assign LUT_3[46710] = 32'b00000000000000010000110010000101;
assign LUT_3[46711] = 32'b00000000000000010111011101100010;
assign LUT_3[46712] = 32'b00000000000000010110110101110001;
assign LUT_3[46713] = 32'b00000000000000011101100001001110;
assign LUT_3[46714] = 32'b00000000000000011000111101010101;
assign LUT_3[46715] = 32'b00000000000000011111101000110010;
assign LUT_3[46716] = 32'b00000000000000010100000011100111;
assign LUT_3[46717] = 32'b00000000000000011010101111000100;
assign LUT_3[46718] = 32'b00000000000000010110001011001011;
assign LUT_3[46719] = 32'b00000000000000011100110110101000;
assign LUT_3[46720] = 32'b00000000000000001111001101011011;
assign LUT_3[46721] = 32'b00000000000000010101111000111000;
assign LUT_3[46722] = 32'b00000000000000010001010100111111;
assign LUT_3[46723] = 32'b00000000000000011000000000011100;
assign LUT_3[46724] = 32'b00000000000000001100011011010001;
assign LUT_3[46725] = 32'b00000000000000010011000110101110;
assign LUT_3[46726] = 32'b00000000000000001110100010110101;
assign LUT_3[46727] = 32'b00000000000000010101001110010010;
assign LUT_3[46728] = 32'b00000000000000010100100110100001;
assign LUT_3[46729] = 32'b00000000000000011011010001111110;
assign LUT_3[46730] = 32'b00000000000000010110101110000101;
assign LUT_3[46731] = 32'b00000000000000011101011001100010;
assign LUT_3[46732] = 32'b00000000000000010001110100010111;
assign LUT_3[46733] = 32'b00000000000000011000011111110100;
assign LUT_3[46734] = 32'b00000000000000010011111011111011;
assign LUT_3[46735] = 32'b00000000000000011010100111011000;
assign LUT_3[46736] = 32'b00000000000000010010100000011110;
assign LUT_3[46737] = 32'b00000000000000011001001011111011;
assign LUT_3[46738] = 32'b00000000000000010100101000000010;
assign LUT_3[46739] = 32'b00000000000000011011010011011111;
assign LUT_3[46740] = 32'b00000000000000001111101110010100;
assign LUT_3[46741] = 32'b00000000000000010110011001110001;
assign LUT_3[46742] = 32'b00000000000000010001110101111000;
assign LUT_3[46743] = 32'b00000000000000011000100001010101;
assign LUT_3[46744] = 32'b00000000000000010111111001100100;
assign LUT_3[46745] = 32'b00000000000000011110100101000001;
assign LUT_3[46746] = 32'b00000000000000011010000001001000;
assign LUT_3[46747] = 32'b00000000000000100000101100100101;
assign LUT_3[46748] = 32'b00000000000000010101000111011010;
assign LUT_3[46749] = 32'b00000000000000011011110010110111;
assign LUT_3[46750] = 32'b00000000000000010111001110111110;
assign LUT_3[46751] = 32'b00000000000000011101111010011011;
assign LUT_3[46752] = 32'b00000000000000010000011011111011;
assign LUT_3[46753] = 32'b00000000000000010111000111011000;
assign LUT_3[46754] = 32'b00000000000000010010100011011111;
assign LUT_3[46755] = 32'b00000000000000011001001110111100;
assign LUT_3[46756] = 32'b00000000000000001101101001110001;
assign LUT_3[46757] = 32'b00000000000000010100010101001110;
assign LUT_3[46758] = 32'b00000000000000001111110001010101;
assign LUT_3[46759] = 32'b00000000000000010110011100110010;
assign LUT_3[46760] = 32'b00000000000000010101110101000001;
assign LUT_3[46761] = 32'b00000000000000011100100000011110;
assign LUT_3[46762] = 32'b00000000000000010111111100100101;
assign LUT_3[46763] = 32'b00000000000000011110101000000010;
assign LUT_3[46764] = 32'b00000000000000010011000010110111;
assign LUT_3[46765] = 32'b00000000000000011001101110010100;
assign LUT_3[46766] = 32'b00000000000000010101001010011011;
assign LUT_3[46767] = 32'b00000000000000011011110101111000;
assign LUT_3[46768] = 32'b00000000000000010011101110111110;
assign LUT_3[46769] = 32'b00000000000000011010011010011011;
assign LUT_3[46770] = 32'b00000000000000010101110110100010;
assign LUT_3[46771] = 32'b00000000000000011100100001111111;
assign LUT_3[46772] = 32'b00000000000000010000111100110100;
assign LUT_3[46773] = 32'b00000000000000010111101000010001;
assign LUT_3[46774] = 32'b00000000000000010011000100011000;
assign LUT_3[46775] = 32'b00000000000000011001101111110101;
assign LUT_3[46776] = 32'b00000000000000011001001000000100;
assign LUT_3[46777] = 32'b00000000000000011111110011100001;
assign LUT_3[46778] = 32'b00000000000000011011001111101000;
assign LUT_3[46779] = 32'b00000000000000100001111011000101;
assign LUT_3[46780] = 32'b00000000000000010110010101111010;
assign LUT_3[46781] = 32'b00000000000000011101000001010111;
assign LUT_3[46782] = 32'b00000000000000011000011101011110;
assign LUT_3[46783] = 32'b00000000000000011111001000111011;
assign LUT_3[46784] = 32'b00000000000000001111000110000110;
assign LUT_3[46785] = 32'b00000000000000010101110001100011;
assign LUT_3[46786] = 32'b00000000000000010001001101101010;
assign LUT_3[46787] = 32'b00000000000000010111111001000111;
assign LUT_3[46788] = 32'b00000000000000001100010011111100;
assign LUT_3[46789] = 32'b00000000000000010010111111011001;
assign LUT_3[46790] = 32'b00000000000000001110011011100000;
assign LUT_3[46791] = 32'b00000000000000010101000110111101;
assign LUT_3[46792] = 32'b00000000000000010100011111001100;
assign LUT_3[46793] = 32'b00000000000000011011001010101001;
assign LUT_3[46794] = 32'b00000000000000010110100110110000;
assign LUT_3[46795] = 32'b00000000000000011101010010001101;
assign LUT_3[46796] = 32'b00000000000000010001101101000010;
assign LUT_3[46797] = 32'b00000000000000011000011000011111;
assign LUT_3[46798] = 32'b00000000000000010011110100100110;
assign LUT_3[46799] = 32'b00000000000000011010100000000011;
assign LUT_3[46800] = 32'b00000000000000010010011001001001;
assign LUT_3[46801] = 32'b00000000000000011001000100100110;
assign LUT_3[46802] = 32'b00000000000000010100100000101101;
assign LUT_3[46803] = 32'b00000000000000011011001100001010;
assign LUT_3[46804] = 32'b00000000000000001111100110111111;
assign LUT_3[46805] = 32'b00000000000000010110010010011100;
assign LUT_3[46806] = 32'b00000000000000010001101110100011;
assign LUT_3[46807] = 32'b00000000000000011000011010000000;
assign LUT_3[46808] = 32'b00000000000000010111110010001111;
assign LUT_3[46809] = 32'b00000000000000011110011101101100;
assign LUT_3[46810] = 32'b00000000000000011001111001110011;
assign LUT_3[46811] = 32'b00000000000000100000100101010000;
assign LUT_3[46812] = 32'b00000000000000010101000000000101;
assign LUT_3[46813] = 32'b00000000000000011011101011100010;
assign LUT_3[46814] = 32'b00000000000000010111000111101001;
assign LUT_3[46815] = 32'b00000000000000011101110011000110;
assign LUT_3[46816] = 32'b00000000000000010000010100100110;
assign LUT_3[46817] = 32'b00000000000000010111000000000011;
assign LUT_3[46818] = 32'b00000000000000010010011100001010;
assign LUT_3[46819] = 32'b00000000000000011001000111100111;
assign LUT_3[46820] = 32'b00000000000000001101100010011100;
assign LUT_3[46821] = 32'b00000000000000010100001101111001;
assign LUT_3[46822] = 32'b00000000000000001111101010000000;
assign LUT_3[46823] = 32'b00000000000000010110010101011101;
assign LUT_3[46824] = 32'b00000000000000010101101101101100;
assign LUT_3[46825] = 32'b00000000000000011100011001001001;
assign LUT_3[46826] = 32'b00000000000000010111110101010000;
assign LUT_3[46827] = 32'b00000000000000011110100000101101;
assign LUT_3[46828] = 32'b00000000000000010010111011100010;
assign LUT_3[46829] = 32'b00000000000000011001100110111111;
assign LUT_3[46830] = 32'b00000000000000010101000011000110;
assign LUT_3[46831] = 32'b00000000000000011011101110100011;
assign LUT_3[46832] = 32'b00000000000000010011100111101001;
assign LUT_3[46833] = 32'b00000000000000011010010011000110;
assign LUT_3[46834] = 32'b00000000000000010101101111001101;
assign LUT_3[46835] = 32'b00000000000000011100011010101010;
assign LUT_3[46836] = 32'b00000000000000010000110101011111;
assign LUT_3[46837] = 32'b00000000000000010111100000111100;
assign LUT_3[46838] = 32'b00000000000000010010111101000011;
assign LUT_3[46839] = 32'b00000000000000011001101000100000;
assign LUT_3[46840] = 32'b00000000000000011001000000101111;
assign LUT_3[46841] = 32'b00000000000000011111101100001100;
assign LUT_3[46842] = 32'b00000000000000011011001000010011;
assign LUT_3[46843] = 32'b00000000000000100001110011110000;
assign LUT_3[46844] = 32'b00000000000000010110001110100101;
assign LUT_3[46845] = 32'b00000000000000011100111010000010;
assign LUT_3[46846] = 32'b00000000000000011000010110001001;
assign LUT_3[46847] = 32'b00000000000000011111000001100110;
assign LUT_3[46848] = 32'b00000000000000001001010001111110;
assign LUT_3[46849] = 32'b00000000000000001111111101011011;
assign LUT_3[46850] = 32'b00000000000000001011011001100010;
assign LUT_3[46851] = 32'b00000000000000010010000100111111;
assign LUT_3[46852] = 32'b00000000000000000110011111110100;
assign LUT_3[46853] = 32'b00000000000000001101001011010001;
assign LUT_3[46854] = 32'b00000000000000001000100111011000;
assign LUT_3[46855] = 32'b00000000000000001111010010110101;
assign LUT_3[46856] = 32'b00000000000000001110101011000100;
assign LUT_3[46857] = 32'b00000000000000010101010110100001;
assign LUT_3[46858] = 32'b00000000000000010000110010101000;
assign LUT_3[46859] = 32'b00000000000000010111011110000101;
assign LUT_3[46860] = 32'b00000000000000001011111000111010;
assign LUT_3[46861] = 32'b00000000000000010010100100010111;
assign LUT_3[46862] = 32'b00000000000000001110000000011110;
assign LUT_3[46863] = 32'b00000000000000010100101011111011;
assign LUT_3[46864] = 32'b00000000000000001100100101000001;
assign LUT_3[46865] = 32'b00000000000000010011010000011110;
assign LUT_3[46866] = 32'b00000000000000001110101100100101;
assign LUT_3[46867] = 32'b00000000000000010101011000000010;
assign LUT_3[46868] = 32'b00000000000000001001110010110111;
assign LUT_3[46869] = 32'b00000000000000010000011110010100;
assign LUT_3[46870] = 32'b00000000000000001011111010011011;
assign LUT_3[46871] = 32'b00000000000000010010100101111000;
assign LUT_3[46872] = 32'b00000000000000010001111110000111;
assign LUT_3[46873] = 32'b00000000000000011000101001100100;
assign LUT_3[46874] = 32'b00000000000000010100000101101011;
assign LUT_3[46875] = 32'b00000000000000011010110001001000;
assign LUT_3[46876] = 32'b00000000000000001111001011111101;
assign LUT_3[46877] = 32'b00000000000000010101110111011010;
assign LUT_3[46878] = 32'b00000000000000010001010011100001;
assign LUT_3[46879] = 32'b00000000000000010111111110111110;
assign LUT_3[46880] = 32'b00000000000000001010100000011110;
assign LUT_3[46881] = 32'b00000000000000010001001011111011;
assign LUT_3[46882] = 32'b00000000000000001100101000000010;
assign LUT_3[46883] = 32'b00000000000000010011010011011111;
assign LUT_3[46884] = 32'b00000000000000000111101110010100;
assign LUT_3[46885] = 32'b00000000000000001110011001110001;
assign LUT_3[46886] = 32'b00000000000000001001110101111000;
assign LUT_3[46887] = 32'b00000000000000010000100001010101;
assign LUT_3[46888] = 32'b00000000000000001111111001100100;
assign LUT_3[46889] = 32'b00000000000000010110100101000001;
assign LUT_3[46890] = 32'b00000000000000010010000001001000;
assign LUT_3[46891] = 32'b00000000000000011000101100100101;
assign LUT_3[46892] = 32'b00000000000000001101000111011010;
assign LUT_3[46893] = 32'b00000000000000010011110010110111;
assign LUT_3[46894] = 32'b00000000000000001111001110111110;
assign LUT_3[46895] = 32'b00000000000000010101111010011011;
assign LUT_3[46896] = 32'b00000000000000001101110011100001;
assign LUT_3[46897] = 32'b00000000000000010100011110111110;
assign LUT_3[46898] = 32'b00000000000000001111111011000101;
assign LUT_3[46899] = 32'b00000000000000010110100110100010;
assign LUT_3[46900] = 32'b00000000000000001011000001010111;
assign LUT_3[46901] = 32'b00000000000000010001101100110100;
assign LUT_3[46902] = 32'b00000000000000001101001000111011;
assign LUT_3[46903] = 32'b00000000000000010011110100011000;
assign LUT_3[46904] = 32'b00000000000000010011001100100111;
assign LUT_3[46905] = 32'b00000000000000011001111000000100;
assign LUT_3[46906] = 32'b00000000000000010101010100001011;
assign LUT_3[46907] = 32'b00000000000000011011111111101000;
assign LUT_3[46908] = 32'b00000000000000010000011010011101;
assign LUT_3[46909] = 32'b00000000000000010111000101111010;
assign LUT_3[46910] = 32'b00000000000000010010100010000001;
assign LUT_3[46911] = 32'b00000000000000011001001101011110;
assign LUT_3[46912] = 32'b00000000000000001001001010101001;
assign LUT_3[46913] = 32'b00000000000000001111110110000110;
assign LUT_3[46914] = 32'b00000000000000001011010010001101;
assign LUT_3[46915] = 32'b00000000000000010001111101101010;
assign LUT_3[46916] = 32'b00000000000000000110011000011111;
assign LUT_3[46917] = 32'b00000000000000001101000011111100;
assign LUT_3[46918] = 32'b00000000000000001000100000000011;
assign LUT_3[46919] = 32'b00000000000000001111001011100000;
assign LUT_3[46920] = 32'b00000000000000001110100011101111;
assign LUT_3[46921] = 32'b00000000000000010101001111001100;
assign LUT_3[46922] = 32'b00000000000000010000101011010011;
assign LUT_3[46923] = 32'b00000000000000010111010110110000;
assign LUT_3[46924] = 32'b00000000000000001011110001100101;
assign LUT_3[46925] = 32'b00000000000000010010011101000010;
assign LUT_3[46926] = 32'b00000000000000001101111001001001;
assign LUT_3[46927] = 32'b00000000000000010100100100100110;
assign LUT_3[46928] = 32'b00000000000000001100011101101100;
assign LUT_3[46929] = 32'b00000000000000010011001001001001;
assign LUT_3[46930] = 32'b00000000000000001110100101010000;
assign LUT_3[46931] = 32'b00000000000000010101010000101101;
assign LUT_3[46932] = 32'b00000000000000001001101011100010;
assign LUT_3[46933] = 32'b00000000000000010000010110111111;
assign LUT_3[46934] = 32'b00000000000000001011110011000110;
assign LUT_3[46935] = 32'b00000000000000010010011110100011;
assign LUT_3[46936] = 32'b00000000000000010001110110110010;
assign LUT_3[46937] = 32'b00000000000000011000100010001111;
assign LUT_3[46938] = 32'b00000000000000010011111110010110;
assign LUT_3[46939] = 32'b00000000000000011010101001110011;
assign LUT_3[46940] = 32'b00000000000000001111000100101000;
assign LUT_3[46941] = 32'b00000000000000010101110000000101;
assign LUT_3[46942] = 32'b00000000000000010001001100001100;
assign LUT_3[46943] = 32'b00000000000000010111110111101001;
assign LUT_3[46944] = 32'b00000000000000001010011001001001;
assign LUT_3[46945] = 32'b00000000000000010001000100100110;
assign LUT_3[46946] = 32'b00000000000000001100100000101101;
assign LUT_3[46947] = 32'b00000000000000010011001100001010;
assign LUT_3[46948] = 32'b00000000000000000111100110111111;
assign LUT_3[46949] = 32'b00000000000000001110010010011100;
assign LUT_3[46950] = 32'b00000000000000001001101110100011;
assign LUT_3[46951] = 32'b00000000000000010000011010000000;
assign LUT_3[46952] = 32'b00000000000000001111110010001111;
assign LUT_3[46953] = 32'b00000000000000010110011101101100;
assign LUT_3[46954] = 32'b00000000000000010001111001110011;
assign LUT_3[46955] = 32'b00000000000000011000100101010000;
assign LUT_3[46956] = 32'b00000000000000001101000000000101;
assign LUT_3[46957] = 32'b00000000000000010011101011100010;
assign LUT_3[46958] = 32'b00000000000000001111000111101001;
assign LUT_3[46959] = 32'b00000000000000010101110011000110;
assign LUT_3[46960] = 32'b00000000000000001101101100001100;
assign LUT_3[46961] = 32'b00000000000000010100010111101001;
assign LUT_3[46962] = 32'b00000000000000001111110011110000;
assign LUT_3[46963] = 32'b00000000000000010110011111001101;
assign LUT_3[46964] = 32'b00000000000000001010111010000010;
assign LUT_3[46965] = 32'b00000000000000010001100101011111;
assign LUT_3[46966] = 32'b00000000000000001101000001100110;
assign LUT_3[46967] = 32'b00000000000000010011101101000011;
assign LUT_3[46968] = 32'b00000000000000010011000101010010;
assign LUT_3[46969] = 32'b00000000000000011001110000101111;
assign LUT_3[46970] = 32'b00000000000000010101001100110110;
assign LUT_3[46971] = 32'b00000000000000011011111000010011;
assign LUT_3[46972] = 32'b00000000000000010000010011001000;
assign LUT_3[46973] = 32'b00000000000000010110111110100101;
assign LUT_3[46974] = 32'b00000000000000010010011010101100;
assign LUT_3[46975] = 32'b00000000000000011001000110001001;
assign LUT_3[46976] = 32'b00000000000000001011011100111100;
assign LUT_3[46977] = 32'b00000000000000010010001000011001;
assign LUT_3[46978] = 32'b00000000000000001101100100100000;
assign LUT_3[46979] = 32'b00000000000000010100001111111101;
assign LUT_3[46980] = 32'b00000000000000001000101010110010;
assign LUT_3[46981] = 32'b00000000000000001111010110001111;
assign LUT_3[46982] = 32'b00000000000000001010110010010110;
assign LUT_3[46983] = 32'b00000000000000010001011101110011;
assign LUT_3[46984] = 32'b00000000000000010000110110000010;
assign LUT_3[46985] = 32'b00000000000000010111100001011111;
assign LUT_3[46986] = 32'b00000000000000010010111101100110;
assign LUT_3[46987] = 32'b00000000000000011001101001000011;
assign LUT_3[46988] = 32'b00000000000000001110000011111000;
assign LUT_3[46989] = 32'b00000000000000010100101111010101;
assign LUT_3[46990] = 32'b00000000000000010000001011011100;
assign LUT_3[46991] = 32'b00000000000000010110110110111001;
assign LUT_3[46992] = 32'b00000000000000001110101111111111;
assign LUT_3[46993] = 32'b00000000000000010101011011011100;
assign LUT_3[46994] = 32'b00000000000000010000110111100011;
assign LUT_3[46995] = 32'b00000000000000010111100011000000;
assign LUT_3[46996] = 32'b00000000000000001011111101110101;
assign LUT_3[46997] = 32'b00000000000000010010101001010010;
assign LUT_3[46998] = 32'b00000000000000001110000101011001;
assign LUT_3[46999] = 32'b00000000000000010100110000110110;
assign LUT_3[47000] = 32'b00000000000000010100001001000101;
assign LUT_3[47001] = 32'b00000000000000011010110100100010;
assign LUT_3[47002] = 32'b00000000000000010110010000101001;
assign LUT_3[47003] = 32'b00000000000000011100111100000110;
assign LUT_3[47004] = 32'b00000000000000010001010110111011;
assign LUT_3[47005] = 32'b00000000000000011000000010011000;
assign LUT_3[47006] = 32'b00000000000000010011011110011111;
assign LUT_3[47007] = 32'b00000000000000011010001001111100;
assign LUT_3[47008] = 32'b00000000000000001100101011011100;
assign LUT_3[47009] = 32'b00000000000000010011010110111001;
assign LUT_3[47010] = 32'b00000000000000001110110011000000;
assign LUT_3[47011] = 32'b00000000000000010101011110011101;
assign LUT_3[47012] = 32'b00000000000000001001111001010010;
assign LUT_3[47013] = 32'b00000000000000010000100100101111;
assign LUT_3[47014] = 32'b00000000000000001100000000110110;
assign LUT_3[47015] = 32'b00000000000000010010101100010011;
assign LUT_3[47016] = 32'b00000000000000010010000100100010;
assign LUT_3[47017] = 32'b00000000000000011000101111111111;
assign LUT_3[47018] = 32'b00000000000000010100001100000110;
assign LUT_3[47019] = 32'b00000000000000011010110111100011;
assign LUT_3[47020] = 32'b00000000000000001111010010011000;
assign LUT_3[47021] = 32'b00000000000000010101111101110101;
assign LUT_3[47022] = 32'b00000000000000010001011001111100;
assign LUT_3[47023] = 32'b00000000000000011000000101011001;
assign LUT_3[47024] = 32'b00000000000000001111111110011111;
assign LUT_3[47025] = 32'b00000000000000010110101001111100;
assign LUT_3[47026] = 32'b00000000000000010010000110000011;
assign LUT_3[47027] = 32'b00000000000000011000110001100000;
assign LUT_3[47028] = 32'b00000000000000001101001100010101;
assign LUT_3[47029] = 32'b00000000000000010011110111110010;
assign LUT_3[47030] = 32'b00000000000000001111010011111001;
assign LUT_3[47031] = 32'b00000000000000010101111111010110;
assign LUT_3[47032] = 32'b00000000000000010101010111100101;
assign LUT_3[47033] = 32'b00000000000000011100000011000010;
assign LUT_3[47034] = 32'b00000000000000010111011111001001;
assign LUT_3[47035] = 32'b00000000000000011110001010100110;
assign LUT_3[47036] = 32'b00000000000000010010100101011011;
assign LUT_3[47037] = 32'b00000000000000011001010000111000;
assign LUT_3[47038] = 32'b00000000000000010100101100111111;
assign LUT_3[47039] = 32'b00000000000000011011011000011100;
assign LUT_3[47040] = 32'b00000000000000001011010101100111;
assign LUT_3[47041] = 32'b00000000000000010010000001000100;
assign LUT_3[47042] = 32'b00000000000000001101011101001011;
assign LUT_3[47043] = 32'b00000000000000010100001000101000;
assign LUT_3[47044] = 32'b00000000000000001000100011011101;
assign LUT_3[47045] = 32'b00000000000000001111001110111010;
assign LUT_3[47046] = 32'b00000000000000001010101011000001;
assign LUT_3[47047] = 32'b00000000000000010001010110011110;
assign LUT_3[47048] = 32'b00000000000000010000101110101101;
assign LUT_3[47049] = 32'b00000000000000010111011010001010;
assign LUT_3[47050] = 32'b00000000000000010010110110010001;
assign LUT_3[47051] = 32'b00000000000000011001100001101110;
assign LUT_3[47052] = 32'b00000000000000001101111100100011;
assign LUT_3[47053] = 32'b00000000000000010100101000000000;
assign LUT_3[47054] = 32'b00000000000000010000000100000111;
assign LUT_3[47055] = 32'b00000000000000010110101111100100;
assign LUT_3[47056] = 32'b00000000000000001110101000101010;
assign LUT_3[47057] = 32'b00000000000000010101010100000111;
assign LUT_3[47058] = 32'b00000000000000010000110000001110;
assign LUT_3[47059] = 32'b00000000000000010111011011101011;
assign LUT_3[47060] = 32'b00000000000000001011110110100000;
assign LUT_3[47061] = 32'b00000000000000010010100001111101;
assign LUT_3[47062] = 32'b00000000000000001101111110000100;
assign LUT_3[47063] = 32'b00000000000000010100101001100001;
assign LUT_3[47064] = 32'b00000000000000010100000001110000;
assign LUT_3[47065] = 32'b00000000000000011010101101001101;
assign LUT_3[47066] = 32'b00000000000000010110001001010100;
assign LUT_3[47067] = 32'b00000000000000011100110100110001;
assign LUT_3[47068] = 32'b00000000000000010001001111100110;
assign LUT_3[47069] = 32'b00000000000000010111111011000011;
assign LUT_3[47070] = 32'b00000000000000010011010111001010;
assign LUT_3[47071] = 32'b00000000000000011010000010100111;
assign LUT_3[47072] = 32'b00000000000000001100100100000111;
assign LUT_3[47073] = 32'b00000000000000010011001111100100;
assign LUT_3[47074] = 32'b00000000000000001110101011101011;
assign LUT_3[47075] = 32'b00000000000000010101010111001000;
assign LUT_3[47076] = 32'b00000000000000001001110001111101;
assign LUT_3[47077] = 32'b00000000000000010000011101011010;
assign LUT_3[47078] = 32'b00000000000000001011111001100001;
assign LUT_3[47079] = 32'b00000000000000010010100100111110;
assign LUT_3[47080] = 32'b00000000000000010001111101001101;
assign LUT_3[47081] = 32'b00000000000000011000101000101010;
assign LUT_3[47082] = 32'b00000000000000010100000100110001;
assign LUT_3[47083] = 32'b00000000000000011010110000001110;
assign LUT_3[47084] = 32'b00000000000000001111001011000011;
assign LUT_3[47085] = 32'b00000000000000010101110110100000;
assign LUT_3[47086] = 32'b00000000000000010001010010100111;
assign LUT_3[47087] = 32'b00000000000000010111111110000100;
assign LUT_3[47088] = 32'b00000000000000001111110111001010;
assign LUT_3[47089] = 32'b00000000000000010110100010100111;
assign LUT_3[47090] = 32'b00000000000000010001111110101110;
assign LUT_3[47091] = 32'b00000000000000011000101010001011;
assign LUT_3[47092] = 32'b00000000000000001101000101000000;
assign LUT_3[47093] = 32'b00000000000000010011110000011101;
assign LUT_3[47094] = 32'b00000000000000001111001100100100;
assign LUT_3[47095] = 32'b00000000000000010101111000000001;
assign LUT_3[47096] = 32'b00000000000000010101010000010000;
assign LUT_3[47097] = 32'b00000000000000011011111011101101;
assign LUT_3[47098] = 32'b00000000000000010111010111110100;
assign LUT_3[47099] = 32'b00000000000000011110000011010001;
assign LUT_3[47100] = 32'b00000000000000010010011110000110;
assign LUT_3[47101] = 32'b00000000000000011001001001100011;
assign LUT_3[47102] = 32'b00000000000000010100100101101010;
assign LUT_3[47103] = 32'b00000000000000011011010001000111;
assign LUT_3[47104] = 32'b00000000000000000100111110100010;
assign LUT_3[47105] = 32'b00000000000000001011101001111111;
assign LUT_3[47106] = 32'b00000000000000000111000110000110;
assign LUT_3[47107] = 32'b00000000000000001101110001100011;
assign LUT_3[47108] = 32'b00000000000000000010001100011000;
assign LUT_3[47109] = 32'b00000000000000001000110111110101;
assign LUT_3[47110] = 32'b00000000000000000100010011111100;
assign LUT_3[47111] = 32'b00000000000000001010111111011001;
assign LUT_3[47112] = 32'b00000000000000001010010111101000;
assign LUT_3[47113] = 32'b00000000000000010001000011000101;
assign LUT_3[47114] = 32'b00000000000000001100011111001100;
assign LUT_3[47115] = 32'b00000000000000010011001010101001;
assign LUT_3[47116] = 32'b00000000000000000111100101011110;
assign LUT_3[47117] = 32'b00000000000000001110010000111011;
assign LUT_3[47118] = 32'b00000000000000001001101101000010;
assign LUT_3[47119] = 32'b00000000000000010000011000011111;
assign LUT_3[47120] = 32'b00000000000000001000010001100101;
assign LUT_3[47121] = 32'b00000000000000001110111101000010;
assign LUT_3[47122] = 32'b00000000000000001010011001001001;
assign LUT_3[47123] = 32'b00000000000000010001000100100110;
assign LUT_3[47124] = 32'b00000000000000000101011111011011;
assign LUT_3[47125] = 32'b00000000000000001100001010111000;
assign LUT_3[47126] = 32'b00000000000000000111100110111111;
assign LUT_3[47127] = 32'b00000000000000001110010010011100;
assign LUT_3[47128] = 32'b00000000000000001101101010101011;
assign LUT_3[47129] = 32'b00000000000000010100010110001000;
assign LUT_3[47130] = 32'b00000000000000001111110010001111;
assign LUT_3[47131] = 32'b00000000000000010110011101101100;
assign LUT_3[47132] = 32'b00000000000000001010111000100001;
assign LUT_3[47133] = 32'b00000000000000010001100011111110;
assign LUT_3[47134] = 32'b00000000000000001101000000000101;
assign LUT_3[47135] = 32'b00000000000000010011101011100010;
assign LUT_3[47136] = 32'b00000000000000000110001101000010;
assign LUT_3[47137] = 32'b00000000000000001100111000011111;
assign LUT_3[47138] = 32'b00000000000000001000010100100110;
assign LUT_3[47139] = 32'b00000000000000001111000000000011;
assign LUT_3[47140] = 32'b00000000000000000011011010111000;
assign LUT_3[47141] = 32'b00000000000000001010000110010101;
assign LUT_3[47142] = 32'b00000000000000000101100010011100;
assign LUT_3[47143] = 32'b00000000000000001100001101111001;
assign LUT_3[47144] = 32'b00000000000000001011100110001000;
assign LUT_3[47145] = 32'b00000000000000010010010001100101;
assign LUT_3[47146] = 32'b00000000000000001101101101101100;
assign LUT_3[47147] = 32'b00000000000000010100011001001001;
assign LUT_3[47148] = 32'b00000000000000001000110011111110;
assign LUT_3[47149] = 32'b00000000000000001111011111011011;
assign LUT_3[47150] = 32'b00000000000000001010111011100010;
assign LUT_3[47151] = 32'b00000000000000010001100110111111;
assign LUT_3[47152] = 32'b00000000000000001001100000000101;
assign LUT_3[47153] = 32'b00000000000000010000001011100010;
assign LUT_3[47154] = 32'b00000000000000001011100111101001;
assign LUT_3[47155] = 32'b00000000000000010010010011000110;
assign LUT_3[47156] = 32'b00000000000000000110101101111011;
assign LUT_3[47157] = 32'b00000000000000001101011001011000;
assign LUT_3[47158] = 32'b00000000000000001000110101011111;
assign LUT_3[47159] = 32'b00000000000000001111100000111100;
assign LUT_3[47160] = 32'b00000000000000001110111001001011;
assign LUT_3[47161] = 32'b00000000000000010101100100101000;
assign LUT_3[47162] = 32'b00000000000000010001000000101111;
assign LUT_3[47163] = 32'b00000000000000010111101100001100;
assign LUT_3[47164] = 32'b00000000000000001100000111000001;
assign LUT_3[47165] = 32'b00000000000000010010110010011110;
assign LUT_3[47166] = 32'b00000000000000001110001110100101;
assign LUT_3[47167] = 32'b00000000000000010100111010000010;
assign LUT_3[47168] = 32'b00000000000000000100110111001101;
assign LUT_3[47169] = 32'b00000000000000001011100010101010;
assign LUT_3[47170] = 32'b00000000000000000110111110110001;
assign LUT_3[47171] = 32'b00000000000000001101101010001110;
assign LUT_3[47172] = 32'b00000000000000000010000101000011;
assign LUT_3[47173] = 32'b00000000000000001000110000100000;
assign LUT_3[47174] = 32'b00000000000000000100001100100111;
assign LUT_3[47175] = 32'b00000000000000001010111000000100;
assign LUT_3[47176] = 32'b00000000000000001010010000010011;
assign LUT_3[47177] = 32'b00000000000000010000111011110000;
assign LUT_3[47178] = 32'b00000000000000001100010111110111;
assign LUT_3[47179] = 32'b00000000000000010011000011010100;
assign LUT_3[47180] = 32'b00000000000000000111011110001001;
assign LUT_3[47181] = 32'b00000000000000001110001001100110;
assign LUT_3[47182] = 32'b00000000000000001001100101101101;
assign LUT_3[47183] = 32'b00000000000000010000010001001010;
assign LUT_3[47184] = 32'b00000000000000001000001010010000;
assign LUT_3[47185] = 32'b00000000000000001110110101101101;
assign LUT_3[47186] = 32'b00000000000000001010010001110100;
assign LUT_3[47187] = 32'b00000000000000010000111101010001;
assign LUT_3[47188] = 32'b00000000000000000101011000000110;
assign LUT_3[47189] = 32'b00000000000000001100000011100011;
assign LUT_3[47190] = 32'b00000000000000000111011111101010;
assign LUT_3[47191] = 32'b00000000000000001110001011000111;
assign LUT_3[47192] = 32'b00000000000000001101100011010110;
assign LUT_3[47193] = 32'b00000000000000010100001110110011;
assign LUT_3[47194] = 32'b00000000000000001111101010111010;
assign LUT_3[47195] = 32'b00000000000000010110010110010111;
assign LUT_3[47196] = 32'b00000000000000001010110001001100;
assign LUT_3[47197] = 32'b00000000000000010001011100101001;
assign LUT_3[47198] = 32'b00000000000000001100111000110000;
assign LUT_3[47199] = 32'b00000000000000010011100100001101;
assign LUT_3[47200] = 32'b00000000000000000110000101101101;
assign LUT_3[47201] = 32'b00000000000000001100110001001010;
assign LUT_3[47202] = 32'b00000000000000001000001101010001;
assign LUT_3[47203] = 32'b00000000000000001110111000101110;
assign LUT_3[47204] = 32'b00000000000000000011010011100011;
assign LUT_3[47205] = 32'b00000000000000001001111111000000;
assign LUT_3[47206] = 32'b00000000000000000101011011000111;
assign LUT_3[47207] = 32'b00000000000000001100000110100100;
assign LUT_3[47208] = 32'b00000000000000001011011110110011;
assign LUT_3[47209] = 32'b00000000000000010010001010010000;
assign LUT_3[47210] = 32'b00000000000000001101100110010111;
assign LUT_3[47211] = 32'b00000000000000010100010001110100;
assign LUT_3[47212] = 32'b00000000000000001000101100101001;
assign LUT_3[47213] = 32'b00000000000000001111011000000110;
assign LUT_3[47214] = 32'b00000000000000001010110100001101;
assign LUT_3[47215] = 32'b00000000000000010001011111101010;
assign LUT_3[47216] = 32'b00000000000000001001011000110000;
assign LUT_3[47217] = 32'b00000000000000010000000100001101;
assign LUT_3[47218] = 32'b00000000000000001011100000010100;
assign LUT_3[47219] = 32'b00000000000000010010001011110001;
assign LUT_3[47220] = 32'b00000000000000000110100110100110;
assign LUT_3[47221] = 32'b00000000000000001101010010000011;
assign LUT_3[47222] = 32'b00000000000000001000101110001010;
assign LUT_3[47223] = 32'b00000000000000001111011001100111;
assign LUT_3[47224] = 32'b00000000000000001110110001110110;
assign LUT_3[47225] = 32'b00000000000000010101011101010011;
assign LUT_3[47226] = 32'b00000000000000010000111001011010;
assign LUT_3[47227] = 32'b00000000000000010111100100110111;
assign LUT_3[47228] = 32'b00000000000000001011111111101100;
assign LUT_3[47229] = 32'b00000000000000010010101011001001;
assign LUT_3[47230] = 32'b00000000000000001110000111010000;
assign LUT_3[47231] = 32'b00000000000000010100110010101101;
assign LUT_3[47232] = 32'b00000000000000000111001001100000;
assign LUT_3[47233] = 32'b00000000000000001101110100111101;
assign LUT_3[47234] = 32'b00000000000000001001010001000100;
assign LUT_3[47235] = 32'b00000000000000001111111100100001;
assign LUT_3[47236] = 32'b00000000000000000100010111010110;
assign LUT_3[47237] = 32'b00000000000000001011000010110011;
assign LUT_3[47238] = 32'b00000000000000000110011110111010;
assign LUT_3[47239] = 32'b00000000000000001101001010010111;
assign LUT_3[47240] = 32'b00000000000000001100100010100110;
assign LUT_3[47241] = 32'b00000000000000010011001110000011;
assign LUT_3[47242] = 32'b00000000000000001110101010001010;
assign LUT_3[47243] = 32'b00000000000000010101010101100111;
assign LUT_3[47244] = 32'b00000000000000001001110000011100;
assign LUT_3[47245] = 32'b00000000000000010000011011111001;
assign LUT_3[47246] = 32'b00000000000000001011111000000000;
assign LUT_3[47247] = 32'b00000000000000010010100011011101;
assign LUT_3[47248] = 32'b00000000000000001010011100100011;
assign LUT_3[47249] = 32'b00000000000000010001001000000000;
assign LUT_3[47250] = 32'b00000000000000001100100100000111;
assign LUT_3[47251] = 32'b00000000000000010011001111100100;
assign LUT_3[47252] = 32'b00000000000000000111101010011001;
assign LUT_3[47253] = 32'b00000000000000001110010101110110;
assign LUT_3[47254] = 32'b00000000000000001001110001111101;
assign LUT_3[47255] = 32'b00000000000000010000011101011010;
assign LUT_3[47256] = 32'b00000000000000001111110101101001;
assign LUT_3[47257] = 32'b00000000000000010110100001000110;
assign LUT_3[47258] = 32'b00000000000000010001111101001101;
assign LUT_3[47259] = 32'b00000000000000011000101000101010;
assign LUT_3[47260] = 32'b00000000000000001101000011011111;
assign LUT_3[47261] = 32'b00000000000000010011101110111100;
assign LUT_3[47262] = 32'b00000000000000001111001011000011;
assign LUT_3[47263] = 32'b00000000000000010101110110100000;
assign LUT_3[47264] = 32'b00000000000000001000011000000000;
assign LUT_3[47265] = 32'b00000000000000001111000011011101;
assign LUT_3[47266] = 32'b00000000000000001010011111100100;
assign LUT_3[47267] = 32'b00000000000000010001001011000001;
assign LUT_3[47268] = 32'b00000000000000000101100101110110;
assign LUT_3[47269] = 32'b00000000000000001100010001010011;
assign LUT_3[47270] = 32'b00000000000000000111101101011010;
assign LUT_3[47271] = 32'b00000000000000001110011000110111;
assign LUT_3[47272] = 32'b00000000000000001101110001000110;
assign LUT_3[47273] = 32'b00000000000000010100011100100011;
assign LUT_3[47274] = 32'b00000000000000001111111000101010;
assign LUT_3[47275] = 32'b00000000000000010110100100000111;
assign LUT_3[47276] = 32'b00000000000000001010111110111100;
assign LUT_3[47277] = 32'b00000000000000010001101010011001;
assign LUT_3[47278] = 32'b00000000000000001101000110100000;
assign LUT_3[47279] = 32'b00000000000000010011110001111101;
assign LUT_3[47280] = 32'b00000000000000001011101011000011;
assign LUT_3[47281] = 32'b00000000000000010010010110100000;
assign LUT_3[47282] = 32'b00000000000000001101110010100111;
assign LUT_3[47283] = 32'b00000000000000010100011110000100;
assign LUT_3[47284] = 32'b00000000000000001000111000111001;
assign LUT_3[47285] = 32'b00000000000000001111100100010110;
assign LUT_3[47286] = 32'b00000000000000001011000000011101;
assign LUT_3[47287] = 32'b00000000000000010001101011111010;
assign LUT_3[47288] = 32'b00000000000000010001000100001001;
assign LUT_3[47289] = 32'b00000000000000010111101111100110;
assign LUT_3[47290] = 32'b00000000000000010011001011101101;
assign LUT_3[47291] = 32'b00000000000000011001110111001010;
assign LUT_3[47292] = 32'b00000000000000001110010001111111;
assign LUT_3[47293] = 32'b00000000000000010100111101011100;
assign LUT_3[47294] = 32'b00000000000000010000011001100011;
assign LUT_3[47295] = 32'b00000000000000010111000101000000;
assign LUT_3[47296] = 32'b00000000000000000111000010001011;
assign LUT_3[47297] = 32'b00000000000000001101101101101000;
assign LUT_3[47298] = 32'b00000000000000001001001001101111;
assign LUT_3[47299] = 32'b00000000000000001111110101001100;
assign LUT_3[47300] = 32'b00000000000000000100010000000001;
assign LUT_3[47301] = 32'b00000000000000001010111011011110;
assign LUT_3[47302] = 32'b00000000000000000110010111100101;
assign LUT_3[47303] = 32'b00000000000000001101000011000010;
assign LUT_3[47304] = 32'b00000000000000001100011011010001;
assign LUT_3[47305] = 32'b00000000000000010011000110101110;
assign LUT_3[47306] = 32'b00000000000000001110100010110101;
assign LUT_3[47307] = 32'b00000000000000010101001110010010;
assign LUT_3[47308] = 32'b00000000000000001001101001000111;
assign LUT_3[47309] = 32'b00000000000000010000010100100100;
assign LUT_3[47310] = 32'b00000000000000001011110000101011;
assign LUT_3[47311] = 32'b00000000000000010010011100001000;
assign LUT_3[47312] = 32'b00000000000000001010010101001110;
assign LUT_3[47313] = 32'b00000000000000010001000000101011;
assign LUT_3[47314] = 32'b00000000000000001100011100110010;
assign LUT_3[47315] = 32'b00000000000000010011001000001111;
assign LUT_3[47316] = 32'b00000000000000000111100011000100;
assign LUT_3[47317] = 32'b00000000000000001110001110100001;
assign LUT_3[47318] = 32'b00000000000000001001101010101000;
assign LUT_3[47319] = 32'b00000000000000010000010110000101;
assign LUT_3[47320] = 32'b00000000000000001111101110010100;
assign LUT_3[47321] = 32'b00000000000000010110011001110001;
assign LUT_3[47322] = 32'b00000000000000010001110101111000;
assign LUT_3[47323] = 32'b00000000000000011000100001010101;
assign LUT_3[47324] = 32'b00000000000000001100111100001010;
assign LUT_3[47325] = 32'b00000000000000010011100111100111;
assign LUT_3[47326] = 32'b00000000000000001111000011101110;
assign LUT_3[47327] = 32'b00000000000000010101101111001011;
assign LUT_3[47328] = 32'b00000000000000001000010000101011;
assign LUT_3[47329] = 32'b00000000000000001110111100001000;
assign LUT_3[47330] = 32'b00000000000000001010011000001111;
assign LUT_3[47331] = 32'b00000000000000010001000011101100;
assign LUT_3[47332] = 32'b00000000000000000101011110100001;
assign LUT_3[47333] = 32'b00000000000000001100001001111110;
assign LUT_3[47334] = 32'b00000000000000000111100110000101;
assign LUT_3[47335] = 32'b00000000000000001110010001100010;
assign LUT_3[47336] = 32'b00000000000000001101101001110001;
assign LUT_3[47337] = 32'b00000000000000010100010101001110;
assign LUT_3[47338] = 32'b00000000000000001111110001010101;
assign LUT_3[47339] = 32'b00000000000000010110011100110010;
assign LUT_3[47340] = 32'b00000000000000001010110111100111;
assign LUT_3[47341] = 32'b00000000000000010001100011000100;
assign LUT_3[47342] = 32'b00000000000000001100111111001011;
assign LUT_3[47343] = 32'b00000000000000010011101010101000;
assign LUT_3[47344] = 32'b00000000000000001011100011101110;
assign LUT_3[47345] = 32'b00000000000000010010001111001011;
assign LUT_3[47346] = 32'b00000000000000001101101011010010;
assign LUT_3[47347] = 32'b00000000000000010100010110101111;
assign LUT_3[47348] = 32'b00000000000000001000110001100100;
assign LUT_3[47349] = 32'b00000000000000001111011101000001;
assign LUT_3[47350] = 32'b00000000000000001010111001001000;
assign LUT_3[47351] = 32'b00000000000000010001100100100101;
assign LUT_3[47352] = 32'b00000000000000010000111100110100;
assign LUT_3[47353] = 32'b00000000000000010111101000010001;
assign LUT_3[47354] = 32'b00000000000000010011000100011000;
assign LUT_3[47355] = 32'b00000000000000011001101111110101;
assign LUT_3[47356] = 32'b00000000000000001110001010101010;
assign LUT_3[47357] = 32'b00000000000000010100110110000111;
assign LUT_3[47358] = 32'b00000000000000010000010010001110;
assign LUT_3[47359] = 32'b00000000000000010110111101101011;
assign LUT_3[47360] = 32'b00000000000000000001001110000011;
assign LUT_3[47361] = 32'b00000000000000000111111001100000;
assign LUT_3[47362] = 32'b00000000000000000011010101100111;
assign LUT_3[47363] = 32'b00000000000000001010000001000100;
assign LUT_3[47364] = 32'b11111111111111111110011011111001;
assign LUT_3[47365] = 32'b00000000000000000101000111010110;
assign LUT_3[47366] = 32'b00000000000000000000100011011101;
assign LUT_3[47367] = 32'b00000000000000000111001110111010;
assign LUT_3[47368] = 32'b00000000000000000110100111001001;
assign LUT_3[47369] = 32'b00000000000000001101010010100110;
assign LUT_3[47370] = 32'b00000000000000001000101110101101;
assign LUT_3[47371] = 32'b00000000000000001111011010001010;
assign LUT_3[47372] = 32'b00000000000000000011110100111111;
assign LUT_3[47373] = 32'b00000000000000001010100000011100;
assign LUT_3[47374] = 32'b00000000000000000101111100100011;
assign LUT_3[47375] = 32'b00000000000000001100101000000000;
assign LUT_3[47376] = 32'b00000000000000000100100001000110;
assign LUT_3[47377] = 32'b00000000000000001011001100100011;
assign LUT_3[47378] = 32'b00000000000000000110101000101010;
assign LUT_3[47379] = 32'b00000000000000001101010100000111;
assign LUT_3[47380] = 32'b00000000000000000001101110111100;
assign LUT_3[47381] = 32'b00000000000000001000011010011001;
assign LUT_3[47382] = 32'b00000000000000000011110110100000;
assign LUT_3[47383] = 32'b00000000000000001010100001111101;
assign LUT_3[47384] = 32'b00000000000000001001111010001100;
assign LUT_3[47385] = 32'b00000000000000010000100101101001;
assign LUT_3[47386] = 32'b00000000000000001100000001110000;
assign LUT_3[47387] = 32'b00000000000000010010101101001101;
assign LUT_3[47388] = 32'b00000000000000000111001000000010;
assign LUT_3[47389] = 32'b00000000000000001101110011011111;
assign LUT_3[47390] = 32'b00000000000000001001001111100110;
assign LUT_3[47391] = 32'b00000000000000001111111011000011;
assign LUT_3[47392] = 32'b00000000000000000010011100100011;
assign LUT_3[47393] = 32'b00000000000000001001001000000000;
assign LUT_3[47394] = 32'b00000000000000000100100100000111;
assign LUT_3[47395] = 32'b00000000000000001011001111100100;
assign LUT_3[47396] = 32'b11111111111111111111101010011001;
assign LUT_3[47397] = 32'b00000000000000000110010101110110;
assign LUT_3[47398] = 32'b00000000000000000001110001111101;
assign LUT_3[47399] = 32'b00000000000000001000011101011010;
assign LUT_3[47400] = 32'b00000000000000000111110101101001;
assign LUT_3[47401] = 32'b00000000000000001110100001000110;
assign LUT_3[47402] = 32'b00000000000000001001111101001101;
assign LUT_3[47403] = 32'b00000000000000010000101000101010;
assign LUT_3[47404] = 32'b00000000000000000101000011011111;
assign LUT_3[47405] = 32'b00000000000000001011101110111100;
assign LUT_3[47406] = 32'b00000000000000000111001011000011;
assign LUT_3[47407] = 32'b00000000000000001101110110100000;
assign LUT_3[47408] = 32'b00000000000000000101101111100110;
assign LUT_3[47409] = 32'b00000000000000001100011011000011;
assign LUT_3[47410] = 32'b00000000000000000111110111001010;
assign LUT_3[47411] = 32'b00000000000000001110100010100111;
assign LUT_3[47412] = 32'b00000000000000000010111101011100;
assign LUT_3[47413] = 32'b00000000000000001001101000111001;
assign LUT_3[47414] = 32'b00000000000000000101000101000000;
assign LUT_3[47415] = 32'b00000000000000001011110000011101;
assign LUT_3[47416] = 32'b00000000000000001011001000101100;
assign LUT_3[47417] = 32'b00000000000000010001110100001001;
assign LUT_3[47418] = 32'b00000000000000001101010000010000;
assign LUT_3[47419] = 32'b00000000000000010011111011101101;
assign LUT_3[47420] = 32'b00000000000000001000010110100010;
assign LUT_3[47421] = 32'b00000000000000001111000001111111;
assign LUT_3[47422] = 32'b00000000000000001010011110000110;
assign LUT_3[47423] = 32'b00000000000000010001001001100011;
assign LUT_3[47424] = 32'b00000000000000000001000110101110;
assign LUT_3[47425] = 32'b00000000000000000111110010001011;
assign LUT_3[47426] = 32'b00000000000000000011001110010010;
assign LUT_3[47427] = 32'b00000000000000001001111001101111;
assign LUT_3[47428] = 32'b11111111111111111110010100100100;
assign LUT_3[47429] = 32'b00000000000000000101000000000001;
assign LUT_3[47430] = 32'b00000000000000000000011100001000;
assign LUT_3[47431] = 32'b00000000000000000111000111100101;
assign LUT_3[47432] = 32'b00000000000000000110011111110100;
assign LUT_3[47433] = 32'b00000000000000001101001011010001;
assign LUT_3[47434] = 32'b00000000000000001000100111011000;
assign LUT_3[47435] = 32'b00000000000000001111010010110101;
assign LUT_3[47436] = 32'b00000000000000000011101101101010;
assign LUT_3[47437] = 32'b00000000000000001010011001000111;
assign LUT_3[47438] = 32'b00000000000000000101110101001110;
assign LUT_3[47439] = 32'b00000000000000001100100000101011;
assign LUT_3[47440] = 32'b00000000000000000100011001110001;
assign LUT_3[47441] = 32'b00000000000000001011000101001110;
assign LUT_3[47442] = 32'b00000000000000000110100001010101;
assign LUT_3[47443] = 32'b00000000000000001101001100110010;
assign LUT_3[47444] = 32'b00000000000000000001100111100111;
assign LUT_3[47445] = 32'b00000000000000001000010011000100;
assign LUT_3[47446] = 32'b00000000000000000011101111001011;
assign LUT_3[47447] = 32'b00000000000000001010011010101000;
assign LUT_3[47448] = 32'b00000000000000001001110010110111;
assign LUT_3[47449] = 32'b00000000000000010000011110010100;
assign LUT_3[47450] = 32'b00000000000000001011111010011011;
assign LUT_3[47451] = 32'b00000000000000010010100101111000;
assign LUT_3[47452] = 32'b00000000000000000111000000101101;
assign LUT_3[47453] = 32'b00000000000000001101101100001010;
assign LUT_3[47454] = 32'b00000000000000001001001000010001;
assign LUT_3[47455] = 32'b00000000000000001111110011101110;
assign LUT_3[47456] = 32'b00000000000000000010010101001110;
assign LUT_3[47457] = 32'b00000000000000001001000000101011;
assign LUT_3[47458] = 32'b00000000000000000100011100110010;
assign LUT_3[47459] = 32'b00000000000000001011001000001111;
assign LUT_3[47460] = 32'b11111111111111111111100011000100;
assign LUT_3[47461] = 32'b00000000000000000110001110100001;
assign LUT_3[47462] = 32'b00000000000000000001101010101000;
assign LUT_3[47463] = 32'b00000000000000001000010110000101;
assign LUT_3[47464] = 32'b00000000000000000111101110010100;
assign LUT_3[47465] = 32'b00000000000000001110011001110001;
assign LUT_3[47466] = 32'b00000000000000001001110101111000;
assign LUT_3[47467] = 32'b00000000000000010000100001010101;
assign LUT_3[47468] = 32'b00000000000000000100111100001010;
assign LUT_3[47469] = 32'b00000000000000001011100111100111;
assign LUT_3[47470] = 32'b00000000000000000111000011101110;
assign LUT_3[47471] = 32'b00000000000000001101101111001011;
assign LUT_3[47472] = 32'b00000000000000000101101000010001;
assign LUT_3[47473] = 32'b00000000000000001100010011101110;
assign LUT_3[47474] = 32'b00000000000000000111101111110101;
assign LUT_3[47475] = 32'b00000000000000001110011011010010;
assign LUT_3[47476] = 32'b00000000000000000010110110000111;
assign LUT_3[47477] = 32'b00000000000000001001100001100100;
assign LUT_3[47478] = 32'b00000000000000000100111101101011;
assign LUT_3[47479] = 32'b00000000000000001011101001001000;
assign LUT_3[47480] = 32'b00000000000000001011000001010111;
assign LUT_3[47481] = 32'b00000000000000010001101100110100;
assign LUT_3[47482] = 32'b00000000000000001101001000111011;
assign LUT_3[47483] = 32'b00000000000000010011110100011000;
assign LUT_3[47484] = 32'b00000000000000001000001111001101;
assign LUT_3[47485] = 32'b00000000000000001110111010101010;
assign LUT_3[47486] = 32'b00000000000000001010010110110001;
assign LUT_3[47487] = 32'b00000000000000010001000010001110;
assign LUT_3[47488] = 32'b00000000000000000011011001000001;
assign LUT_3[47489] = 32'b00000000000000001010000100011110;
assign LUT_3[47490] = 32'b00000000000000000101100000100101;
assign LUT_3[47491] = 32'b00000000000000001100001100000010;
assign LUT_3[47492] = 32'b00000000000000000000100110110111;
assign LUT_3[47493] = 32'b00000000000000000111010010010100;
assign LUT_3[47494] = 32'b00000000000000000010101110011011;
assign LUT_3[47495] = 32'b00000000000000001001011001111000;
assign LUT_3[47496] = 32'b00000000000000001000110010000111;
assign LUT_3[47497] = 32'b00000000000000001111011101100100;
assign LUT_3[47498] = 32'b00000000000000001010111001101011;
assign LUT_3[47499] = 32'b00000000000000010001100101001000;
assign LUT_3[47500] = 32'b00000000000000000101111111111101;
assign LUT_3[47501] = 32'b00000000000000001100101011011010;
assign LUT_3[47502] = 32'b00000000000000001000000111100001;
assign LUT_3[47503] = 32'b00000000000000001110110010111110;
assign LUT_3[47504] = 32'b00000000000000000110101100000100;
assign LUT_3[47505] = 32'b00000000000000001101010111100001;
assign LUT_3[47506] = 32'b00000000000000001000110011101000;
assign LUT_3[47507] = 32'b00000000000000001111011111000101;
assign LUT_3[47508] = 32'b00000000000000000011111001111010;
assign LUT_3[47509] = 32'b00000000000000001010100101010111;
assign LUT_3[47510] = 32'b00000000000000000110000001011110;
assign LUT_3[47511] = 32'b00000000000000001100101100111011;
assign LUT_3[47512] = 32'b00000000000000001100000101001010;
assign LUT_3[47513] = 32'b00000000000000010010110000100111;
assign LUT_3[47514] = 32'b00000000000000001110001100101110;
assign LUT_3[47515] = 32'b00000000000000010100111000001011;
assign LUT_3[47516] = 32'b00000000000000001001010011000000;
assign LUT_3[47517] = 32'b00000000000000001111111110011101;
assign LUT_3[47518] = 32'b00000000000000001011011010100100;
assign LUT_3[47519] = 32'b00000000000000010010000110000001;
assign LUT_3[47520] = 32'b00000000000000000100100111100001;
assign LUT_3[47521] = 32'b00000000000000001011010010111110;
assign LUT_3[47522] = 32'b00000000000000000110101111000101;
assign LUT_3[47523] = 32'b00000000000000001101011010100010;
assign LUT_3[47524] = 32'b00000000000000000001110101010111;
assign LUT_3[47525] = 32'b00000000000000001000100000110100;
assign LUT_3[47526] = 32'b00000000000000000011111100111011;
assign LUT_3[47527] = 32'b00000000000000001010101000011000;
assign LUT_3[47528] = 32'b00000000000000001010000000100111;
assign LUT_3[47529] = 32'b00000000000000010000101100000100;
assign LUT_3[47530] = 32'b00000000000000001100001000001011;
assign LUT_3[47531] = 32'b00000000000000010010110011101000;
assign LUT_3[47532] = 32'b00000000000000000111001110011101;
assign LUT_3[47533] = 32'b00000000000000001101111001111010;
assign LUT_3[47534] = 32'b00000000000000001001010110000001;
assign LUT_3[47535] = 32'b00000000000000010000000001011110;
assign LUT_3[47536] = 32'b00000000000000000111111010100100;
assign LUT_3[47537] = 32'b00000000000000001110100110000001;
assign LUT_3[47538] = 32'b00000000000000001010000010001000;
assign LUT_3[47539] = 32'b00000000000000010000101101100101;
assign LUT_3[47540] = 32'b00000000000000000101001000011010;
assign LUT_3[47541] = 32'b00000000000000001011110011110111;
assign LUT_3[47542] = 32'b00000000000000000111001111111110;
assign LUT_3[47543] = 32'b00000000000000001101111011011011;
assign LUT_3[47544] = 32'b00000000000000001101010011101010;
assign LUT_3[47545] = 32'b00000000000000010011111111000111;
assign LUT_3[47546] = 32'b00000000000000001111011011001110;
assign LUT_3[47547] = 32'b00000000000000010110000110101011;
assign LUT_3[47548] = 32'b00000000000000001010100001100000;
assign LUT_3[47549] = 32'b00000000000000010001001100111101;
assign LUT_3[47550] = 32'b00000000000000001100101001000100;
assign LUT_3[47551] = 32'b00000000000000010011010100100001;
assign LUT_3[47552] = 32'b00000000000000000011010001101100;
assign LUT_3[47553] = 32'b00000000000000001001111101001001;
assign LUT_3[47554] = 32'b00000000000000000101011001010000;
assign LUT_3[47555] = 32'b00000000000000001100000100101101;
assign LUT_3[47556] = 32'b00000000000000000000011111100010;
assign LUT_3[47557] = 32'b00000000000000000111001010111111;
assign LUT_3[47558] = 32'b00000000000000000010100111000110;
assign LUT_3[47559] = 32'b00000000000000001001010010100011;
assign LUT_3[47560] = 32'b00000000000000001000101010110010;
assign LUT_3[47561] = 32'b00000000000000001111010110001111;
assign LUT_3[47562] = 32'b00000000000000001010110010010110;
assign LUT_3[47563] = 32'b00000000000000010001011101110011;
assign LUT_3[47564] = 32'b00000000000000000101111000101000;
assign LUT_3[47565] = 32'b00000000000000001100100100000101;
assign LUT_3[47566] = 32'b00000000000000001000000000001100;
assign LUT_3[47567] = 32'b00000000000000001110101011101001;
assign LUT_3[47568] = 32'b00000000000000000110100100101111;
assign LUT_3[47569] = 32'b00000000000000001101010000001100;
assign LUT_3[47570] = 32'b00000000000000001000101100010011;
assign LUT_3[47571] = 32'b00000000000000001111010111110000;
assign LUT_3[47572] = 32'b00000000000000000011110010100101;
assign LUT_3[47573] = 32'b00000000000000001010011110000010;
assign LUT_3[47574] = 32'b00000000000000000101111010001001;
assign LUT_3[47575] = 32'b00000000000000001100100101100110;
assign LUT_3[47576] = 32'b00000000000000001011111101110101;
assign LUT_3[47577] = 32'b00000000000000010010101001010010;
assign LUT_3[47578] = 32'b00000000000000001110000101011001;
assign LUT_3[47579] = 32'b00000000000000010100110000110110;
assign LUT_3[47580] = 32'b00000000000000001001001011101011;
assign LUT_3[47581] = 32'b00000000000000001111110111001000;
assign LUT_3[47582] = 32'b00000000000000001011010011001111;
assign LUT_3[47583] = 32'b00000000000000010001111110101100;
assign LUT_3[47584] = 32'b00000000000000000100100000001100;
assign LUT_3[47585] = 32'b00000000000000001011001011101001;
assign LUT_3[47586] = 32'b00000000000000000110100111110000;
assign LUT_3[47587] = 32'b00000000000000001101010011001101;
assign LUT_3[47588] = 32'b00000000000000000001101110000010;
assign LUT_3[47589] = 32'b00000000000000001000011001011111;
assign LUT_3[47590] = 32'b00000000000000000011110101100110;
assign LUT_3[47591] = 32'b00000000000000001010100001000011;
assign LUT_3[47592] = 32'b00000000000000001001111001010010;
assign LUT_3[47593] = 32'b00000000000000010000100100101111;
assign LUT_3[47594] = 32'b00000000000000001100000000110110;
assign LUT_3[47595] = 32'b00000000000000010010101100010011;
assign LUT_3[47596] = 32'b00000000000000000111000111001000;
assign LUT_3[47597] = 32'b00000000000000001101110010100101;
assign LUT_3[47598] = 32'b00000000000000001001001110101100;
assign LUT_3[47599] = 32'b00000000000000001111111010001001;
assign LUT_3[47600] = 32'b00000000000000000111110011001111;
assign LUT_3[47601] = 32'b00000000000000001110011110101100;
assign LUT_3[47602] = 32'b00000000000000001001111010110011;
assign LUT_3[47603] = 32'b00000000000000010000100110010000;
assign LUT_3[47604] = 32'b00000000000000000101000001000101;
assign LUT_3[47605] = 32'b00000000000000001011101100100010;
assign LUT_3[47606] = 32'b00000000000000000111001000101001;
assign LUT_3[47607] = 32'b00000000000000001101110100000110;
assign LUT_3[47608] = 32'b00000000000000001101001100010101;
assign LUT_3[47609] = 32'b00000000000000010011110111110010;
assign LUT_3[47610] = 32'b00000000000000001111010011111001;
assign LUT_3[47611] = 32'b00000000000000010101111111010110;
assign LUT_3[47612] = 32'b00000000000000001010011010001011;
assign LUT_3[47613] = 32'b00000000000000010001000101101000;
assign LUT_3[47614] = 32'b00000000000000001100100001101111;
assign LUT_3[47615] = 32'b00000000000000010011001101001100;
assign LUT_3[47616] = 32'b00000000000000001000010011101110;
assign LUT_3[47617] = 32'b00000000000000001110111111001011;
assign LUT_3[47618] = 32'b00000000000000001010011011010010;
assign LUT_3[47619] = 32'b00000000000000010001000110101111;
assign LUT_3[47620] = 32'b00000000000000000101100001100100;
assign LUT_3[47621] = 32'b00000000000000001100001101000001;
assign LUT_3[47622] = 32'b00000000000000000111101001001000;
assign LUT_3[47623] = 32'b00000000000000001110010100100101;
assign LUT_3[47624] = 32'b00000000000000001101101100110100;
assign LUT_3[47625] = 32'b00000000000000010100011000010001;
assign LUT_3[47626] = 32'b00000000000000001111110100011000;
assign LUT_3[47627] = 32'b00000000000000010110011111110101;
assign LUT_3[47628] = 32'b00000000000000001010111010101010;
assign LUT_3[47629] = 32'b00000000000000010001100110000111;
assign LUT_3[47630] = 32'b00000000000000001101000010001110;
assign LUT_3[47631] = 32'b00000000000000010011101101101011;
assign LUT_3[47632] = 32'b00000000000000001011100110110001;
assign LUT_3[47633] = 32'b00000000000000010010010010001110;
assign LUT_3[47634] = 32'b00000000000000001101101110010101;
assign LUT_3[47635] = 32'b00000000000000010100011001110010;
assign LUT_3[47636] = 32'b00000000000000001000110100100111;
assign LUT_3[47637] = 32'b00000000000000001111100000000100;
assign LUT_3[47638] = 32'b00000000000000001010111100001011;
assign LUT_3[47639] = 32'b00000000000000010001100111101000;
assign LUT_3[47640] = 32'b00000000000000010000111111110111;
assign LUT_3[47641] = 32'b00000000000000010111101011010100;
assign LUT_3[47642] = 32'b00000000000000010011000111011011;
assign LUT_3[47643] = 32'b00000000000000011001110010111000;
assign LUT_3[47644] = 32'b00000000000000001110001101101101;
assign LUT_3[47645] = 32'b00000000000000010100111001001010;
assign LUT_3[47646] = 32'b00000000000000010000010101010001;
assign LUT_3[47647] = 32'b00000000000000010111000000101110;
assign LUT_3[47648] = 32'b00000000000000001001100010001110;
assign LUT_3[47649] = 32'b00000000000000010000001101101011;
assign LUT_3[47650] = 32'b00000000000000001011101001110010;
assign LUT_3[47651] = 32'b00000000000000010010010101001111;
assign LUT_3[47652] = 32'b00000000000000000110110000000100;
assign LUT_3[47653] = 32'b00000000000000001101011011100001;
assign LUT_3[47654] = 32'b00000000000000001000110111101000;
assign LUT_3[47655] = 32'b00000000000000001111100011000101;
assign LUT_3[47656] = 32'b00000000000000001110111011010100;
assign LUT_3[47657] = 32'b00000000000000010101100110110001;
assign LUT_3[47658] = 32'b00000000000000010001000010111000;
assign LUT_3[47659] = 32'b00000000000000010111101110010101;
assign LUT_3[47660] = 32'b00000000000000001100001001001010;
assign LUT_3[47661] = 32'b00000000000000010010110100100111;
assign LUT_3[47662] = 32'b00000000000000001110010000101110;
assign LUT_3[47663] = 32'b00000000000000010100111100001011;
assign LUT_3[47664] = 32'b00000000000000001100110101010001;
assign LUT_3[47665] = 32'b00000000000000010011100000101110;
assign LUT_3[47666] = 32'b00000000000000001110111100110101;
assign LUT_3[47667] = 32'b00000000000000010101101000010010;
assign LUT_3[47668] = 32'b00000000000000001010000011000111;
assign LUT_3[47669] = 32'b00000000000000010000101110100100;
assign LUT_3[47670] = 32'b00000000000000001100001010101011;
assign LUT_3[47671] = 32'b00000000000000010010110110001000;
assign LUT_3[47672] = 32'b00000000000000010010001110010111;
assign LUT_3[47673] = 32'b00000000000000011000111001110100;
assign LUT_3[47674] = 32'b00000000000000010100010101111011;
assign LUT_3[47675] = 32'b00000000000000011011000001011000;
assign LUT_3[47676] = 32'b00000000000000001111011100001101;
assign LUT_3[47677] = 32'b00000000000000010110000111101010;
assign LUT_3[47678] = 32'b00000000000000010001100011110001;
assign LUT_3[47679] = 32'b00000000000000011000001111001110;
assign LUT_3[47680] = 32'b00000000000000001000001100011001;
assign LUT_3[47681] = 32'b00000000000000001110110111110110;
assign LUT_3[47682] = 32'b00000000000000001010010011111101;
assign LUT_3[47683] = 32'b00000000000000010000111111011010;
assign LUT_3[47684] = 32'b00000000000000000101011010001111;
assign LUT_3[47685] = 32'b00000000000000001100000101101100;
assign LUT_3[47686] = 32'b00000000000000000111100001110011;
assign LUT_3[47687] = 32'b00000000000000001110001101010000;
assign LUT_3[47688] = 32'b00000000000000001101100101011111;
assign LUT_3[47689] = 32'b00000000000000010100010000111100;
assign LUT_3[47690] = 32'b00000000000000001111101101000011;
assign LUT_3[47691] = 32'b00000000000000010110011000100000;
assign LUT_3[47692] = 32'b00000000000000001010110011010101;
assign LUT_3[47693] = 32'b00000000000000010001011110110010;
assign LUT_3[47694] = 32'b00000000000000001100111010111001;
assign LUT_3[47695] = 32'b00000000000000010011100110010110;
assign LUT_3[47696] = 32'b00000000000000001011011111011100;
assign LUT_3[47697] = 32'b00000000000000010010001010111001;
assign LUT_3[47698] = 32'b00000000000000001101100111000000;
assign LUT_3[47699] = 32'b00000000000000010100010010011101;
assign LUT_3[47700] = 32'b00000000000000001000101101010010;
assign LUT_3[47701] = 32'b00000000000000001111011000101111;
assign LUT_3[47702] = 32'b00000000000000001010110100110110;
assign LUT_3[47703] = 32'b00000000000000010001100000010011;
assign LUT_3[47704] = 32'b00000000000000010000111000100010;
assign LUT_3[47705] = 32'b00000000000000010111100011111111;
assign LUT_3[47706] = 32'b00000000000000010011000000000110;
assign LUT_3[47707] = 32'b00000000000000011001101011100011;
assign LUT_3[47708] = 32'b00000000000000001110000110011000;
assign LUT_3[47709] = 32'b00000000000000010100110001110101;
assign LUT_3[47710] = 32'b00000000000000010000001101111100;
assign LUT_3[47711] = 32'b00000000000000010110111001011001;
assign LUT_3[47712] = 32'b00000000000000001001011010111001;
assign LUT_3[47713] = 32'b00000000000000010000000110010110;
assign LUT_3[47714] = 32'b00000000000000001011100010011101;
assign LUT_3[47715] = 32'b00000000000000010010001101111010;
assign LUT_3[47716] = 32'b00000000000000000110101000101111;
assign LUT_3[47717] = 32'b00000000000000001101010100001100;
assign LUT_3[47718] = 32'b00000000000000001000110000010011;
assign LUT_3[47719] = 32'b00000000000000001111011011110000;
assign LUT_3[47720] = 32'b00000000000000001110110011111111;
assign LUT_3[47721] = 32'b00000000000000010101011111011100;
assign LUT_3[47722] = 32'b00000000000000010000111011100011;
assign LUT_3[47723] = 32'b00000000000000010111100111000000;
assign LUT_3[47724] = 32'b00000000000000001100000001110101;
assign LUT_3[47725] = 32'b00000000000000010010101101010010;
assign LUT_3[47726] = 32'b00000000000000001110001001011001;
assign LUT_3[47727] = 32'b00000000000000010100110100110110;
assign LUT_3[47728] = 32'b00000000000000001100101101111100;
assign LUT_3[47729] = 32'b00000000000000010011011001011001;
assign LUT_3[47730] = 32'b00000000000000001110110101100000;
assign LUT_3[47731] = 32'b00000000000000010101100000111101;
assign LUT_3[47732] = 32'b00000000000000001001111011110010;
assign LUT_3[47733] = 32'b00000000000000010000100111001111;
assign LUT_3[47734] = 32'b00000000000000001100000011010110;
assign LUT_3[47735] = 32'b00000000000000010010101110110011;
assign LUT_3[47736] = 32'b00000000000000010010000111000010;
assign LUT_3[47737] = 32'b00000000000000011000110010011111;
assign LUT_3[47738] = 32'b00000000000000010100001110100110;
assign LUT_3[47739] = 32'b00000000000000011010111010000011;
assign LUT_3[47740] = 32'b00000000000000001111010100111000;
assign LUT_3[47741] = 32'b00000000000000010110000000010101;
assign LUT_3[47742] = 32'b00000000000000010001011100011100;
assign LUT_3[47743] = 32'b00000000000000011000000111111001;
assign LUT_3[47744] = 32'b00000000000000001010011110101100;
assign LUT_3[47745] = 32'b00000000000000010001001010001001;
assign LUT_3[47746] = 32'b00000000000000001100100110010000;
assign LUT_3[47747] = 32'b00000000000000010011010001101101;
assign LUT_3[47748] = 32'b00000000000000000111101100100010;
assign LUT_3[47749] = 32'b00000000000000001110010111111111;
assign LUT_3[47750] = 32'b00000000000000001001110100000110;
assign LUT_3[47751] = 32'b00000000000000010000011111100011;
assign LUT_3[47752] = 32'b00000000000000001111110111110010;
assign LUT_3[47753] = 32'b00000000000000010110100011001111;
assign LUT_3[47754] = 32'b00000000000000010001111111010110;
assign LUT_3[47755] = 32'b00000000000000011000101010110011;
assign LUT_3[47756] = 32'b00000000000000001101000101101000;
assign LUT_3[47757] = 32'b00000000000000010011110001000101;
assign LUT_3[47758] = 32'b00000000000000001111001101001100;
assign LUT_3[47759] = 32'b00000000000000010101111000101001;
assign LUT_3[47760] = 32'b00000000000000001101110001101111;
assign LUT_3[47761] = 32'b00000000000000010100011101001100;
assign LUT_3[47762] = 32'b00000000000000001111111001010011;
assign LUT_3[47763] = 32'b00000000000000010110100100110000;
assign LUT_3[47764] = 32'b00000000000000001010111111100101;
assign LUT_3[47765] = 32'b00000000000000010001101011000010;
assign LUT_3[47766] = 32'b00000000000000001101000111001001;
assign LUT_3[47767] = 32'b00000000000000010011110010100110;
assign LUT_3[47768] = 32'b00000000000000010011001010110101;
assign LUT_3[47769] = 32'b00000000000000011001110110010010;
assign LUT_3[47770] = 32'b00000000000000010101010010011001;
assign LUT_3[47771] = 32'b00000000000000011011111101110110;
assign LUT_3[47772] = 32'b00000000000000010000011000101011;
assign LUT_3[47773] = 32'b00000000000000010111000100001000;
assign LUT_3[47774] = 32'b00000000000000010010100000001111;
assign LUT_3[47775] = 32'b00000000000000011001001011101100;
assign LUT_3[47776] = 32'b00000000000000001011101101001100;
assign LUT_3[47777] = 32'b00000000000000010010011000101001;
assign LUT_3[47778] = 32'b00000000000000001101110100110000;
assign LUT_3[47779] = 32'b00000000000000010100100000001101;
assign LUT_3[47780] = 32'b00000000000000001000111011000010;
assign LUT_3[47781] = 32'b00000000000000001111100110011111;
assign LUT_3[47782] = 32'b00000000000000001011000010100110;
assign LUT_3[47783] = 32'b00000000000000010001101110000011;
assign LUT_3[47784] = 32'b00000000000000010001000110010010;
assign LUT_3[47785] = 32'b00000000000000010111110001101111;
assign LUT_3[47786] = 32'b00000000000000010011001101110110;
assign LUT_3[47787] = 32'b00000000000000011001111001010011;
assign LUT_3[47788] = 32'b00000000000000001110010100001000;
assign LUT_3[47789] = 32'b00000000000000010100111111100101;
assign LUT_3[47790] = 32'b00000000000000010000011011101100;
assign LUT_3[47791] = 32'b00000000000000010111000111001001;
assign LUT_3[47792] = 32'b00000000000000001111000000001111;
assign LUT_3[47793] = 32'b00000000000000010101101011101100;
assign LUT_3[47794] = 32'b00000000000000010001000111110011;
assign LUT_3[47795] = 32'b00000000000000010111110011010000;
assign LUT_3[47796] = 32'b00000000000000001100001110000101;
assign LUT_3[47797] = 32'b00000000000000010010111001100010;
assign LUT_3[47798] = 32'b00000000000000001110010101101001;
assign LUT_3[47799] = 32'b00000000000000010101000001000110;
assign LUT_3[47800] = 32'b00000000000000010100011001010101;
assign LUT_3[47801] = 32'b00000000000000011011000100110010;
assign LUT_3[47802] = 32'b00000000000000010110100000111001;
assign LUT_3[47803] = 32'b00000000000000011101001100010110;
assign LUT_3[47804] = 32'b00000000000000010001100111001011;
assign LUT_3[47805] = 32'b00000000000000011000010010101000;
assign LUT_3[47806] = 32'b00000000000000010011101110101111;
assign LUT_3[47807] = 32'b00000000000000011010011010001100;
assign LUT_3[47808] = 32'b00000000000000001010010111010111;
assign LUT_3[47809] = 32'b00000000000000010001000010110100;
assign LUT_3[47810] = 32'b00000000000000001100011110111011;
assign LUT_3[47811] = 32'b00000000000000010011001010011000;
assign LUT_3[47812] = 32'b00000000000000000111100101001101;
assign LUT_3[47813] = 32'b00000000000000001110010000101010;
assign LUT_3[47814] = 32'b00000000000000001001101100110001;
assign LUT_3[47815] = 32'b00000000000000010000011000001110;
assign LUT_3[47816] = 32'b00000000000000001111110000011101;
assign LUT_3[47817] = 32'b00000000000000010110011011111010;
assign LUT_3[47818] = 32'b00000000000000010001111000000001;
assign LUT_3[47819] = 32'b00000000000000011000100011011110;
assign LUT_3[47820] = 32'b00000000000000001100111110010011;
assign LUT_3[47821] = 32'b00000000000000010011101001110000;
assign LUT_3[47822] = 32'b00000000000000001111000101110111;
assign LUT_3[47823] = 32'b00000000000000010101110001010100;
assign LUT_3[47824] = 32'b00000000000000001101101010011010;
assign LUT_3[47825] = 32'b00000000000000010100010101110111;
assign LUT_3[47826] = 32'b00000000000000001111110001111110;
assign LUT_3[47827] = 32'b00000000000000010110011101011011;
assign LUT_3[47828] = 32'b00000000000000001010111000010000;
assign LUT_3[47829] = 32'b00000000000000010001100011101101;
assign LUT_3[47830] = 32'b00000000000000001100111111110100;
assign LUT_3[47831] = 32'b00000000000000010011101011010001;
assign LUT_3[47832] = 32'b00000000000000010011000011100000;
assign LUT_3[47833] = 32'b00000000000000011001101110111101;
assign LUT_3[47834] = 32'b00000000000000010101001011000100;
assign LUT_3[47835] = 32'b00000000000000011011110110100001;
assign LUT_3[47836] = 32'b00000000000000010000010001010110;
assign LUT_3[47837] = 32'b00000000000000010110111100110011;
assign LUT_3[47838] = 32'b00000000000000010010011000111010;
assign LUT_3[47839] = 32'b00000000000000011001000100010111;
assign LUT_3[47840] = 32'b00000000000000001011100101110111;
assign LUT_3[47841] = 32'b00000000000000010010010001010100;
assign LUT_3[47842] = 32'b00000000000000001101101101011011;
assign LUT_3[47843] = 32'b00000000000000010100011000111000;
assign LUT_3[47844] = 32'b00000000000000001000110011101101;
assign LUT_3[47845] = 32'b00000000000000001111011111001010;
assign LUT_3[47846] = 32'b00000000000000001010111011010001;
assign LUT_3[47847] = 32'b00000000000000010001100110101110;
assign LUT_3[47848] = 32'b00000000000000010000111110111101;
assign LUT_3[47849] = 32'b00000000000000010111101010011010;
assign LUT_3[47850] = 32'b00000000000000010011000110100001;
assign LUT_3[47851] = 32'b00000000000000011001110001111110;
assign LUT_3[47852] = 32'b00000000000000001110001100110011;
assign LUT_3[47853] = 32'b00000000000000010100111000010000;
assign LUT_3[47854] = 32'b00000000000000010000010100010111;
assign LUT_3[47855] = 32'b00000000000000010110111111110100;
assign LUT_3[47856] = 32'b00000000000000001110111000111010;
assign LUT_3[47857] = 32'b00000000000000010101100100010111;
assign LUT_3[47858] = 32'b00000000000000010001000000011110;
assign LUT_3[47859] = 32'b00000000000000010111101011111011;
assign LUT_3[47860] = 32'b00000000000000001100000110110000;
assign LUT_3[47861] = 32'b00000000000000010010110010001101;
assign LUT_3[47862] = 32'b00000000000000001110001110010100;
assign LUT_3[47863] = 32'b00000000000000010100111001110001;
assign LUT_3[47864] = 32'b00000000000000010100010010000000;
assign LUT_3[47865] = 32'b00000000000000011010111101011101;
assign LUT_3[47866] = 32'b00000000000000010110011001100100;
assign LUT_3[47867] = 32'b00000000000000011101000101000001;
assign LUT_3[47868] = 32'b00000000000000010001011111110110;
assign LUT_3[47869] = 32'b00000000000000011000001011010011;
assign LUT_3[47870] = 32'b00000000000000010011100111011010;
assign LUT_3[47871] = 32'b00000000000000011010010010110111;
assign LUT_3[47872] = 32'b00000000000000000100100011001111;
assign LUT_3[47873] = 32'b00000000000000001011001110101100;
assign LUT_3[47874] = 32'b00000000000000000110101010110011;
assign LUT_3[47875] = 32'b00000000000000001101010110010000;
assign LUT_3[47876] = 32'b00000000000000000001110001000101;
assign LUT_3[47877] = 32'b00000000000000001000011100100010;
assign LUT_3[47878] = 32'b00000000000000000011111000101001;
assign LUT_3[47879] = 32'b00000000000000001010100100000110;
assign LUT_3[47880] = 32'b00000000000000001001111100010101;
assign LUT_3[47881] = 32'b00000000000000010000100111110010;
assign LUT_3[47882] = 32'b00000000000000001100000011111001;
assign LUT_3[47883] = 32'b00000000000000010010101111010110;
assign LUT_3[47884] = 32'b00000000000000000111001010001011;
assign LUT_3[47885] = 32'b00000000000000001101110101101000;
assign LUT_3[47886] = 32'b00000000000000001001010001101111;
assign LUT_3[47887] = 32'b00000000000000001111111101001100;
assign LUT_3[47888] = 32'b00000000000000000111110110010010;
assign LUT_3[47889] = 32'b00000000000000001110100001101111;
assign LUT_3[47890] = 32'b00000000000000001001111101110110;
assign LUT_3[47891] = 32'b00000000000000010000101001010011;
assign LUT_3[47892] = 32'b00000000000000000101000100001000;
assign LUT_3[47893] = 32'b00000000000000001011101111100101;
assign LUT_3[47894] = 32'b00000000000000000111001011101100;
assign LUT_3[47895] = 32'b00000000000000001101110111001001;
assign LUT_3[47896] = 32'b00000000000000001101001111011000;
assign LUT_3[47897] = 32'b00000000000000010011111010110101;
assign LUT_3[47898] = 32'b00000000000000001111010110111100;
assign LUT_3[47899] = 32'b00000000000000010110000010011001;
assign LUT_3[47900] = 32'b00000000000000001010011101001110;
assign LUT_3[47901] = 32'b00000000000000010001001000101011;
assign LUT_3[47902] = 32'b00000000000000001100100100110010;
assign LUT_3[47903] = 32'b00000000000000010011010000001111;
assign LUT_3[47904] = 32'b00000000000000000101110001101111;
assign LUT_3[47905] = 32'b00000000000000001100011101001100;
assign LUT_3[47906] = 32'b00000000000000000111111001010011;
assign LUT_3[47907] = 32'b00000000000000001110100100110000;
assign LUT_3[47908] = 32'b00000000000000000010111111100101;
assign LUT_3[47909] = 32'b00000000000000001001101011000010;
assign LUT_3[47910] = 32'b00000000000000000101000111001001;
assign LUT_3[47911] = 32'b00000000000000001011110010100110;
assign LUT_3[47912] = 32'b00000000000000001011001010110101;
assign LUT_3[47913] = 32'b00000000000000010001110110010010;
assign LUT_3[47914] = 32'b00000000000000001101010010011001;
assign LUT_3[47915] = 32'b00000000000000010011111101110110;
assign LUT_3[47916] = 32'b00000000000000001000011000101011;
assign LUT_3[47917] = 32'b00000000000000001111000100001000;
assign LUT_3[47918] = 32'b00000000000000001010100000001111;
assign LUT_3[47919] = 32'b00000000000000010001001011101100;
assign LUT_3[47920] = 32'b00000000000000001001000100110010;
assign LUT_3[47921] = 32'b00000000000000001111110000001111;
assign LUT_3[47922] = 32'b00000000000000001011001100010110;
assign LUT_3[47923] = 32'b00000000000000010001110111110011;
assign LUT_3[47924] = 32'b00000000000000000110010010101000;
assign LUT_3[47925] = 32'b00000000000000001100111110000101;
assign LUT_3[47926] = 32'b00000000000000001000011010001100;
assign LUT_3[47927] = 32'b00000000000000001111000101101001;
assign LUT_3[47928] = 32'b00000000000000001110011101111000;
assign LUT_3[47929] = 32'b00000000000000010101001001010101;
assign LUT_3[47930] = 32'b00000000000000010000100101011100;
assign LUT_3[47931] = 32'b00000000000000010111010000111001;
assign LUT_3[47932] = 32'b00000000000000001011101011101110;
assign LUT_3[47933] = 32'b00000000000000010010010111001011;
assign LUT_3[47934] = 32'b00000000000000001101110011010010;
assign LUT_3[47935] = 32'b00000000000000010100011110101111;
assign LUT_3[47936] = 32'b00000000000000000100011011111010;
assign LUT_3[47937] = 32'b00000000000000001011000111010111;
assign LUT_3[47938] = 32'b00000000000000000110100011011110;
assign LUT_3[47939] = 32'b00000000000000001101001110111011;
assign LUT_3[47940] = 32'b00000000000000000001101001110000;
assign LUT_3[47941] = 32'b00000000000000001000010101001101;
assign LUT_3[47942] = 32'b00000000000000000011110001010100;
assign LUT_3[47943] = 32'b00000000000000001010011100110001;
assign LUT_3[47944] = 32'b00000000000000001001110101000000;
assign LUT_3[47945] = 32'b00000000000000010000100000011101;
assign LUT_3[47946] = 32'b00000000000000001011111100100100;
assign LUT_3[47947] = 32'b00000000000000010010101000000001;
assign LUT_3[47948] = 32'b00000000000000000111000010110110;
assign LUT_3[47949] = 32'b00000000000000001101101110010011;
assign LUT_3[47950] = 32'b00000000000000001001001010011010;
assign LUT_3[47951] = 32'b00000000000000001111110101110111;
assign LUT_3[47952] = 32'b00000000000000000111101110111101;
assign LUT_3[47953] = 32'b00000000000000001110011010011010;
assign LUT_3[47954] = 32'b00000000000000001001110110100001;
assign LUT_3[47955] = 32'b00000000000000010000100001111110;
assign LUT_3[47956] = 32'b00000000000000000100111100110011;
assign LUT_3[47957] = 32'b00000000000000001011101000010000;
assign LUT_3[47958] = 32'b00000000000000000111000100010111;
assign LUT_3[47959] = 32'b00000000000000001101101111110100;
assign LUT_3[47960] = 32'b00000000000000001101001000000011;
assign LUT_3[47961] = 32'b00000000000000010011110011100000;
assign LUT_3[47962] = 32'b00000000000000001111001111100111;
assign LUT_3[47963] = 32'b00000000000000010101111011000100;
assign LUT_3[47964] = 32'b00000000000000001010010101111001;
assign LUT_3[47965] = 32'b00000000000000010001000001010110;
assign LUT_3[47966] = 32'b00000000000000001100011101011101;
assign LUT_3[47967] = 32'b00000000000000010011001000111010;
assign LUT_3[47968] = 32'b00000000000000000101101010011010;
assign LUT_3[47969] = 32'b00000000000000001100010101110111;
assign LUT_3[47970] = 32'b00000000000000000111110001111110;
assign LUT_3[47971] = 32'b00000000000000001110011101011011;
assign LUT_3[47972] = 32'b00000000000000000010111000010000;
assign LUT_3[47973] = 32'b00000000000000001001100011101101;
assign LUT_3[47974] = 32'b00000000000000000100111111110100;
assign LUT_3[47975] = 32'b00000000000000001011101011010001;
assign LUT_3[47976] = 32'b00000000000000001011000011100000;
assign LUT_3[47977] = 32'b00000000000000010001101110111101;
assign LUT_3[47978] = 32'b00000000000000001101001011000100;
assign LUT_3[47979] = 32'b00000000000000010011110110100001;
assign LUT_3[47980] = 32'b00000000000000001000010001010110;
assign LUT_3[47981] = 32'b00000000000000001110111100110011;
assign LUT_3[47982] = 32'b00000000000000001010011000111010;
assign LUT_3[47983] = 32'b00000000000000010001000100010111;
assign LUT_3[47984] = 32'b00000000000000001000111101011101;
assign LUT_3[47985] = 32'b00000000000000001111101000111010;
assign LUT_3[47986] = 32'b00000000000000001011000101000001;
assign LUT_3[47987] = 32'b00000000000000010001110000011110;
assign LUT_3[47988] = 32'b00000000000000000110001011010011;
assign LUT_3[47989] = 32'b00000000000000001100110110110000;
assign LUT_3[47990] = 32'b00000000000000001000010010110111;
assign LUT_3[47991] = 32'b00000000000000001110111110010100;
assign LUT_3[47992] = 32'b00000000000000001110010110100011;
assign LUT_3[47993] = 32'b00000000000000010101000010000000;
assign LUT_3[47994] = 32'b00000000000000010000011110000111;
assign LUT_3[47995] = 32'b00000000000000010111001001100100;
assign LUT_3[47996] = 32'b00000000000000001011100100011001;
assign LUT_3[47997] = 32'b00000000000000010010001111110110;
assign LUT_3[47998] = 32'b00000000000000001101101011111101;
assign LUT_3[47999] = 32'b00000000000000010100010111011010;
assign LUT_3[48000] = 32'b00000000000000000110101110001101;
assign LUT_3[48001] = 32'b00000000000000001101011001101010;
assign LUT_3[48002] = 32'b00000000000000001000110101110001;
assign LUT_3[48003] = 32'b00000000000000001111100001001110;
assign LUT_3[48004] = 32'b00000000000000000011111100000011;
assign LUT_3[48005] = 32'b00000000000000001010100111100000;
assign LUT_3[48006] = 32'b00000000000000000110000011100111;
assign LUT_3[48007] = 32'b00000000000000001100101111000100;
assign LUT_3[48008] = 32'b00000000000000001100000111010011;
assign LUT_3[48009] = 32'b00000000000000010010110010110000;
assign LUT_3[48010] = 32'b00000000000000001110001110110111;
assign LUT_3[48011] = 32'b00000000000000010100111010010100;
assign LUT_3[48012] = 32'b00000000000000001001010101001001;
assign LUT_3[48013] = 32'b00000000000000010000000000100110;
assign LUT_3[48014] = 32'b00000000000000001011011100101101;
assign LUT_3[48015] = 32'b00000000000000010010001000001010;
assign LUT_3[48016] = 32'b00000000000000001010000001010000;
assign LUT_3[48017] = 32'b00000000000000010000101100101101;
assign LUT_3[48018] = 32'b00000000000000001100001000110100;
assign LUT_3[48019] = 32'b00000000000000010010110100010001;
assign LUT_3[48020] = 32'b00000000000000000111001111000110;
assign LUT_3[48021] = 32'b00000000000000001101111010100011;
assign LUT_3[48022] = 32'b00000000000000001001010110101010;
assign LUT_3[48023] = 32'b00000000000000010000000010000111;
assign LUT_3[48024] = 32'b00000000000000001111011010010110;
assign LUT_3[48025] = 32'b00000000000000010110000101110011;
assign LUT_3[48026] = 32'b00000000000000010001100001111010;
assign LUT_3[48027] = 32'b00000000000000011000001101010111;
assign LUT_3[48028] = 32'b00000000000000001100101000001100;
assign LUT_3[48029] = 32'b00000000000000010011010011101001;
assign LUT_3[48030] = 32'b00000000000000001110101111110000;
assign LUT_3[48031] = 32'b00000000000000010101011011001101;
assign LUT_3[48032] = 32'b00000000000000000111111100101101;
assign LUT_3[48033] = 32'b00000000000000001110101000001010;
assign LUT_3[48034] = 32'b00000000000000001010000100010001;
assign LUT_3[48035] = 32'b00000000000000010000101111101110;
assign LUT_3[48036] = 32'b00000000000000000101001010100011;
assign LUT_3[48037] = 32'b00000000000000001011110110000000;
assign LUT_3[48038] = 32'b00000000000000000111010010000111;
assign LUT_3[48039] = 32'b00000000000000001101111101100100;
assign LUT_3[48040] = 32'b00000000000000001101010101110011;
assign LUT_3[48041] = 32'b00000000000000010100000001010000;
assign LUT_3[48042] = 32'b00000000000000001111011101010111;
assign LUT_3[48043] = 32'b00000000000000010110001000110100;
assign LUT_3[48044] = 32'b00000000000000001010100011101001;
assign LUT_3[48045] = 32'b00000000000000010001001111000110;
assign LUT_3[48046] = 32'b00000000000000001100101011001101;
assign LUT_3[48047] = 32'b00000000000000010011010110101010;
assign LUT_3[48048] = 32'b00000000000000001011001111110000;
assign LUT_3[48049] = 32'b00000000000000010001111011001101;
assign LUT_3[48050] = 32'b00000000000000001101010111010100;
assign LUT_3[48051] = 32'b00000000000000010100000010110001;
assign LUT_3[48052] = 32'b00000000000000001000011101100110;
assign LUT_3[48053] = 32'b00000000000000001111001001000011;
assign LUT_3[48054] = 32'b00000000000000001010100101001010;
assign LUT_3[48055] = 32'b00000000000000010001010000100111;
assign LUT_3[48056] = 32'b00000000000000010000101000110110;
assign LUT_3[48057] = 32'b00000000000000010111010100010011;
assign LUT_3[48058] = 32'b00000000000000010010110000011010;
assign LUT_3[48059] = 32'b00000000000000011001011011110111;
assign LUT_3[48060] = 32'b00000000000000001101110110101100;
assign LUT_3[48061] = 32'b00000000000000010100100010001001;
assign LUT_3[48062] = 32'b00000000000000001111111110010000;
assign LUT_3[48063] = 32'b00000000000000010110101001101101;
assign LUT_3[48064] = 32'b00000000000000000110100110111000;
assign LUT_3[48065] = 32'b00000000000000001101010010010101;
assign LUT_3[48066] = 32'b00000000000000001000101110011100;
assign LUT_3[48067] = 32'b00000000000000001111011001111001;
assign LUT_3[48068] = 32'b00000000000000000011110100101110;
assign LUT_3[48069] = 32'b00000000000000001010100000001011;
assign LUT_3[48070] = 32'b00000000000000000101111100010010;
assign LUT_3[48071] = 32'b00000000000000001100100111101111;
assign LUT_3[48072] = 32'b00000000000000001011111111111110;
assign LUT_3[48073] = 32'b00000000000000010010101011011011;
assign LUT_3[48074] = 32'b00000000000000001110000111100010;
assign LUT_3[48075] = 32'b00000000000000010100110010111111;
assign LUT_3[48076] = 32'b00000000000000001001001101110100;
assign LUT_3[48077] = 32'b00000000000000001111111001010001;
assign LUT_3[48078] = 32'b00000000000000001011010101011000;
assign LUT_3[48079] = 32'b00000000000000010010000000110101;
assign LUT_3[48080] = 32'b00000000000000001001111001111011;
assign LUT_3[48081] = 32'b00000000000000010000100101011000;
assign LUT_3[48082] = 32'b00000000000000001100000001011111;
assign LUT_3[48083] = 32'b00000000000000010010101100111100;
assign LUT_3[48084] = 32'b00000000000000000111000111110001;
assign LUT_3[48085] = 32'b00000000000000001101110011001110;
assign LUT_3[48086] = 32'b00000000000000001001001111010101;
assign LUT_3[48087] = 32'b00000000000000001111111010110010;
assign LUT_3[48088] = 32'b00000000000000001111010011000001;
assign LUT_3[48089] = 32'b00000000000000010101111110011110;
assign LUT_3[48090] = 32'b00000000000000010001011010100101;
assign LUT_3[48091] = 32'b00000000000000011000000110000010;
assign LUT_3[48092] = 32'b00000000000000001100100000110111;
assign LUT_3[48093] = 32'b00000000000000010011001100010100;
assign LUT_3[48094] = 32'b00000000000000001110101000011011;
assign LUT_3[48095] = 32'b00000000000000010101010011111000;
assign LUT_3[48096] = 32'b00000000000000000111110101011000;
assign LUT_3[48097] = 32'b00000000000000001110100000110101;
assign LUT_3[48098] = 32'b00000000000000001001111100111100;
assign LUT_3[48099] = 32'b00000000000000010000101000011001;
assign LUT_3[48100] = 32'b00000000000000000101000011001110;
assign LUT_3[48101] = 32'b00000000000000001011101110101011;
assign LUT_3[48102] = 32'b00000000000000000111001010110010;
assign LUT_3[48103] = 32'b00000000000000001101110110001111;
assign LUT_3[48104] = 32'b00000000000000001101001110011110;
assign LUT_3[48105] = 32'b00000000000000010011111001111011;
assign LUT_3[48106] = 32'b00000000000000001111010110000010;
assign LUT_3[48107] = 32'b00000000000000010110000001011111;
assign LUT_3[48108] = 32'b00000000000000001010011100010100;
assign LUT_3[48109] = 32'b00000000000000010001000111110001;
assign LUT_3[48110] = 32'b00000000000000001100100011111000;
assign LUT_3[48111] = 32'b00000000000000010011001111010101;
assign LUT_3[48112] = 32'b00000000000000001011001000011011;
assign LUT_3[48113] = 32'b00000000000000010001110011111000;
assign LUT_3[48114] = 32'b00000000000000001101001111111111;
assign LUT_3[48115] = 32'b00000000000000010011111011011100;
assign LUT_3[48116] = 32'b00000000000000001000010110010001;
assign LUT_3[48117] = 32'b00000000000000001111000001101110;
assign LUT_3[48118] = 32'b00000000000000001010011101110101;
assign LUT_3[48119] = 32'b00000000000000010001001001010010;
assign LUT_3[48120] = 32'b00000000000000010000100001100001;
assign LUT_3[48121] = 32'b00000000000000010111001100111110;
assign LUT_3[48122] = 32'b00000000000000010010101001000101;
assign LUT_3[48123] = 32'b00000000000000011001010100100010;
assign LUT_3[48124] = 32'b00000000000000001101101111010111;
assign LUT_3[48125] = 32'b00000000000000010100011010110100;
assign LUT_3[48126] = 32'b00000000000000001111110110111011;
assign LUT_3[48127] = 32'b00000000000000010110100010011000;
assign LUT_3[48128] = 32'b00000000000000001011100011011111;
assign LUT_3[48129] = 32'b00000000000000010010001110111100;
assign LUT_3[48130] = 32'b00000000000000001101101011000011;
assign LUT_3[48131] = 32'b00000000000000010100010110100000;
assign LUT_3[48132] = 32'b00000000000000001000110001010101;
assign LUT_3[48133] = 32'b00000000000000001111011100110010;
assign LUT_3[48134] = 32'b00000000000000001010111000111001;
assign LUT_3[48135] = 32'b00000000000000010001100100010110;
assign LUT_3[48136] = 32'b00000000000000010000111100100101;
assign LUT_3[48137] = 32'b00000000000000010111101000000010;
assign LUT_3[48138] = 32'b00000000000000010011000100001001;
assign LUT_3[48139] = 32'b00000000000000011001101111100110;
assign LUT_3[48140] = 32'b00000000000000001110001010011011;
assign LUT_3[48141] = 32'b00000000000000010100110101111000;
assign LUT_3[48142] = 32'b00000000000000010000010001111111;
assign LUT_3[48143] = 32'b00000000000000010110111101011100;
assign LUT_3[48144] = 32'b00000000000000001110110110100010;
assign LUT_3[48145] = 32'b00000000000000010101100001111111;
assign LUT_3[48146] = 32'b00000000000000010000111110000110;
assign LUT_3[48147] = 32'b00000000000000010111101001100011;
assign LUT_3[48148] = 32'b00000000000000001100000100011000;
assign LUT_3[48149] = 32'b00000000000000010010101111110101;
assign LUT_3[48150] = 32'b00000000000000001110001011111100;
assign LUT_3[48151] = 32'b00000000000000010100110111011001;
assign LUT_3[48152] = 32'b00000000000000010100001111101000;
assign LUT_3[48153] = 32'b00000000000000011010111011000101;
assign LUT_3[48154] = 32'b00000000000000010110010111001100;
assign LUT_3[48155] = 32'b00000000000000011101000010101001;
assign LUT_3[48156] = 32'b00000000000000010001011101011110;
assign LUT_3[48157] = 32'b00000000000000011000001000111011;
assign LUT_3[48158] = 32'b00000000000000010011100101000010;
assign LUT_3[48159] = 32'b00000000000000011010010000011111;
assign LUT_3[48160] = 32'b00000000000000001100110001111111;
assign LUT_3[48161] = 32'b00000000000000010011011101011100;
assign LUT_3[48162] = 32'b00000000000000001110111001100011;
assign LUT_3[48163] = 32'b00000000000000010101100101000000;
assign LUT_3[48164] = 32'b00000000000000001001111111110101;
assign LUT_3[48165] = 32'b00000000000000010000101011010010;
assign LUT_3[48166] = 32'b00000000000000001100000111011001;
assign LUT_3[48167] = 32'b00000000000000010010110010110110;
assign LUT_3[48168] = 32'b00000000000000010010001011000101;
assign LUT_3[48169] = 32'b00000000000000011000110110100010;
assign LUT_3[48170] = 32'b00000000000000010100010010101001;
assign LUT_3[48171] = 32'b00000000000000011010111110000110;
assign LUT_3[48172] = 32'b00000000000000001111011000111011;
assign LUT_3[48173] = 32'b00000000000000010110000100011000;
assign LUT_3[48174] = 32'b00000000000000010001100000011111;
assign LUT_3[48175] = 32'b00000000000000011000001011111100;
assign LUT_3[48176] = 32'b00000000000000010000000101000010;
assign LUT_3[48177] = 32'b00000000000000010110110000011111;
assign LUT_3[48178] = 32'b00000000000000010010001100100110;
assign LUT_3[48179] = 32'b00000000000000011000111000000011;
assign LUT_3[48180] = 32'b00000000000000001101010010111000;
assign LUT_3[48181] = 32'b00000000000000010011111110010101;
assign LUT_3[48182] = 32'b00000000000000001111011010011100;
assign LUT_3[48183] = 32'b00000000000000010110000101111001;
assign LUT_3[48184] = 32'b00000000000000010101011110001000;
assign LUT_3[48185] = 32'b00000000000000011100001001100101;
assign LUT_3[48186] = 32'b00000000000000010111100101101100;
assign LUT_3[48187] = 32'b00000000000000011110010001001001;
assign LUT_3[48188] = 32'b00000000000000010010101011111110;
assign LUT_3[48189] = 32'b00000000000000011001010111011011;
assign LUT_3[48190] = 32'b00000000000000010100110011100010;
assign LUT_3[48191] = 32'b00000000000000011011011110111111;
assign LUT_3[48192] = 32'b00000000000000001011011100001010;
assign LUT_3[48193] = 32'b00000000000000010010000111100111;
assign LUT_3[48194] = 32'b00000000000000001101100011101110;
assign LUT_3[48195] = 32'b00000000000000010100001111001011;
assign LUT_3[48196] = 32'b00000000000000001000101010000000;
assign LUT_3[48197] = 32'b00000000000000001111010101011101;
assign LUT_3[48198] = 32'b00000000000000001010110001100100;
assign LUT_3[48199] = 32'b00000000000000010001011101000001;
assign LUT_3[48200] = 32'b00000000000000010000110101010000;
assign LUT_3[48201] = 32'b00000000000000010111100000101101;
assign LUT_3[48202] = 32'b00000000000000010010111100110100;
assign LUT_3[48203] = 32'b00000000000000011001101000010001;
assign LUT_3[48204] = 32'b00000000000000001110000011000110;
assign LUT_3[48205] = 32'b00000000000000010100101110100011;
assign LUT_3[48206] = 32'b00000000000000010000001010101010;
assign LUT_3[48207] = 32'b00000000000000010110110110000111;
assign LUT_3[48208] = 32'b00000000000000001110101111001101;
assign LUT_3[48209] = 32'b00000000000000010101011010101010;
assign LUT_3[48210] = 32'b00000000000000010000110110110001;
assign LUT_3[48211] = 32'b00000000000000010111100010001110;
assign LUT_3[48212] = 32'b00000000000000001011111101000011;
assign LUT_3[48213] = 32'b00000000000000010010101000100000;
assign LUT_3[48214] = 32'b00000000000000001110000100100111;
assign LUT_3[48215] = 32'b00000000000000010100110000000100;
assign LUT_3[48216] = 32'b00000000000000010100001000010011;
assign LUT_3[48217] = 32'b00000000000000011010110011110000;
assign LUT_3[48218] = 32'b00000000000000010110001111110111;
assign LUT_3[48219] = 32'b00000000000000011100111011010100;
assign LUT_3[48220] = 32'b00000000000000010001010110001001;
assign LUT_3[48221] = 32'b00000000000000011000000001100110;
assign LUT_3[48222] = 32'b00000000000000010011011101101101;
assign LUT_3[48223] = 32'b00000000000000011010001001001010;
assign LUT_3[48224] = 32'b00000000000000001100101010101010;
assign LUT_3[48225] = 32'b00000000000000010011010110000111;
assign LUT_3[48226] = 32'b00000000000000001110110010001110;
assign LUT_3[48227] = 32'b00000000000000010101011101101011;
assign LUT_3[48228] = 32'b00000000000000001001111000100000;
assign LUT_3[48229] = 32'b00000000000000010000100011111101;
assign LUT_3[48230] = 32'b00000000000000001100000000000100;
assign LUT_3[48231] = 32'b00000000000000010010101011100001;
assign LUT_3[48232] = 32'b00000000000000010010000011110000;
assign LUT_3[48233] = 32'b00000000000000011000101111001101;
assign LUT_3[48234] = 32'b00000000000000010100001011010100;
assign LUT_3[48235] = 32'b00000000000000011010110110110001;
assign LUT_3[48236] = 32'b00000000000000001111010001100110;
assign LUT_3[48237] = 32'b00000000000000010101111101000011;
assign LUT_3[48238] = 32'b00000000000000010001011001001010;
assign LUT_3[48239] = 32'b00000000000000011000000100100111;
assign LUT_3[48240] = 32'b00000000000000001111111101101101;
assign LUT_3[48241] = 32'b00000000000000010110101001001010;
assign LUT_3[48242] = 32'b00000000000000010010000101010001;
assign LUT_3[48243] = 32'b00000000000000011000110000101110;
assign LUT_3[48244] = 32'b00000000000000001101001011100011;
assign LUT_3[48245] = 32'b00000000000000010011110111000000;
assign LUT_3[48246] = 32'b00000000000000001111010011000111;
assign LUT_3[48247] = 32'b00000000000000010101111110100100;
assign LUT_3[48248] = 32'b00000000000000010101010110110011;
assign LUT_3[48249] = 32'b00000000000000011100000010010000;
assign LUT_3[48250] = 32'b00000000000000010111011110010111;
assign LUT_3[48251] = 32'b00000000000000011110001001110100;
assign LUT_3[48252] = 32'b00000000000000010010100100101001;
assign LUT_3[48253] = 32'b00000000000000011001010000000110;
assign LUT_3[48254] = 32'b00000000000000010100101100001101;
assign LUT_3[48255] = 32'b00000000000000011011010111101010;
assign LUT_3[48256] = 32'b00000000000000001101101110011101;
assign LUT_3[48257] = 32'b00000000000000010100011001111010;
assign LUT_3[48258] = 32'b00000000000000001111110110000001;
assign LUT_3[48259] = 32'b00000000000000010110100001011110;
assign LUT_3[48260] = 32'b00000000000000001010111100010011;
assign LUT_3[48261] = 32'b00000000000000010001100111110000;
assign LUT_3[48262] = 32'b00000000000000001101000011110111;
assign LUT_3[48263] = 32'b00000000000000010011101111010100;
assign LUT_3[48264] = 32'b00000000000000010011000111100011;
assign LUT_3[48265] = 32'b00000000000000011001110011000000;
assign LUT_3[48266] = 32'b00000000000000010101001111000111;
assign LUT_3[48267] = 32'b00000000000000011011111010100100;
assign LUT_3[48268] = 32'b00000000000000010000010101011001;
assign LUT_3[48269] = 32'b00000000000000010111000000110110;
assign LUT_3[48270] = 32'b00000000000000010010011100111101;
assign LUT_3[48271] = 32'b00000000000000011001001000011010;
assign LUT_3[48272] = 32'b00000000000000010001000001100000;
assign LUT_3[48273] = 32'b00000000000000010111101100111101;
assign LUT_3[48274] = 32'b00000000000000010011001001000100;
assign LUT_3[48275] = 32'b00000000000000011001110100100001;
assign LUT_3[48276] = 32'b00000000000000001110001111010110;
assign LUT_3[48277] = 32'b00000000000000010100111010110011;
assign LUT_3[48278] = 32'b00000000000000010000010110111010;
assign LUT_3[48279] = 32'b00000000000000010111000010010111;
assign LUT_3[48280] = 32'b00000000000000010110011010100110;
assign LUT_3[48281] = 32'b00000000000000011101000110000011;
assign LUT_3[48282] = 32'b00000000000000011000100010001010;
assign LUT_3[48283] = 32'b00000000000000011111001101100111;
assign LUT_3[48284] = 32'b00000000000000010011101000011100;
assign LUT_3[48285] = 32'b00000000000000011010010011111001;
assign LUT_3[48286] = 32'b00000000000000010101110000000000;
assign LUT_3[48287] = 32'b00000000000000011100011011011101;
assign LUT_3[48288] = 32'b00000000000000001110111100111101;
assign LUT_3[48289] = 32'b00000000000000010101101000011010;
assign LUT_3[48290] = 32'b00000000000000010001000100100001;
assign LUT_3[48291] = 32'b00000000000000010111101111111110;
assign LUT_3[48292] = 32'b00000000000000001100001010110011;
assign LUT_3[48293] = 32'b00000000000000010010110110010000;
assign LUT_3[48294] = 32'b00000000000000001110010010010111;
assign LUT_3[48295] = 32'b00000000000000010100111101110100;
assign LUT_3[48296] = 32'b00000000000000010100010110000011;
assign LUT_3[48297] = 32'b00000000000000011011000001100000;
assign LUT_3[48298] = 32'b00000000000000010110011101100111;
assign LUT_3[48299] = 32'b00000000000000011101001001000100;
assign LUT_3[48300] = 32'b00000000000000010001100011111001;
assign LUT_3[48301] = 32'b00000000000000011000001111010110;
assign LUT_3[48302] = 32'b00000000000000010011101011011101;
assign LUT_3[48303] = 32'b00000000000000011010010110111010;
assign LUT_3[48304] = 32'b00000000000000010010010000000000;
assign LUT_3[48305] = 32'b00000000000000011000111011011101;
assign LUT_3[48306] = 32'b00000000000000010100010111100100;
assign LUT_3[48307] = 32'b00000000000000011011000011000001;
assign LUT_3[48308] = 32'b00000000000000001111011101110110;
assign LUT_3[48309] = 32'b00000000000000010110001001010011;
assign LUT_3[48310] = 32'b00000000000000010001100101011010;
assign LUT_3[48311] = 32'b00000000000000011000010000110111;
assign LUT_3[48312] = 32'b00000000000000010111101001000110;
assign LUT_3[48313] = 32'b00000000000000011110010100100011;
assign LUT_3[48314] = 32'b00000000000000011001110000101010;
assign LUT_3[48315] = 32'b00000000000000100000011100000111;
assign LUT_3[48316] = 32'b00000000000000010100110110111100;
assign LUT_3[48317] = 32'b00000000000000011011100010011001;
assign LUT_3[48318] = 32'b00000000000000010110111110100000;
assign LUT_3[48319] = 32'b00000000000000011101101001111101;
assign LUT_3[48320] = 32'b00000000000000001101100111001000;
assign LUT_3[48321] = 32'b00000000000000010100010010100101;
assign LUT_3[48322] = 32'b00000000000000001111101110101100;
assign LUT_3[48323] = 32'b00000000000000010110011010001001;
assign LUT_3[48324] = 32'b00000000000000001010110100111110;
assign LUT_3[48325] = 32'b00000000000000010001100000011011;
assign LUT_3[48326] = 32'b00000000000000001100111100100010;
assign LUT_3[48327] = 32'b00000000000000010011100111111111;
assign LUT_3[48328] = 32'b00000000000000010011000000001110;
assign LUT_3[48329] = 32'b00000000000000011001101011101011;
assign LUT_3[48330] = 32'b00000000000000010101000111110010;
assign LUT_3[48331] = 32'b00000000000000011011110011001111;
assign LUT_3[48332] = 32'b00000000000000010000001110000100;
assign LUT_3[48333] = 32'b00000000000000010110111001100001;
assign LUT_3[48334] = 32'b00000000000000010010010101101000;
assign LUT_3[48335] = 32'b00000000000000011001000001000101;
assign LUT_3[48336] = 32'b00000000000000010000111010001011;
assign LUT_3[48337] = 32'b00000000000000010111100101101000;
assign LUT_3[48338] = 32'b00000000000000010011000001101111;
assign LUT_3[48339] = 32'b00000000000000011001101101001100;
assign LUT_3[48340] = 32'b00000000000000001110001000000001;
assign LUT_3[48341] = 32'b00000000000000010100110011011110;
assign LUT_3[48342] = 32'b00000000000000010000001111100101;
assign LUT_3[48343] = 32'b00000000000000010110111011000010;
assign LUT_3[48344] = 32'b00000000000000010110010011010001;
assign LUT_3[48345] = 32'b00000000000000011100111110101110;
assign LUT_3[48346] = 32'b00000000000000011000011010110101;
assign LUT_3[48347] = 32'b00000000000000011111000110010010;
assign LUT_3[48348] = 32'b00000000000000010011100001000111;
assign LUT_3[48349] = 32'b00000000000000011010001100100100;
assign LUT_3[48350] = 32'b00000000000000010101101000101011;
assign LUT_3[48351] = 32'b00000000000000011100010100001000;
assign LUT_3[48352] = 32'b00000000000000001110110101101000;
assign LUT_3[48353] = 32'b00000000000000010101100001000101;
assign LUT_3[48354] = 32'b00000000000000010000111101001100;
assign LUT_3[48355] = 32'b00000000000000010111101000101001;
assign LUT_3[48356] = 32'b00000000000000001100000011011110;
assign LUT_3[48357] = 32'b00000000000000010010101110111011;
assign LUT_3[48358] = 32'b00000000000000001110001011000010;
assign LUT_3[48359] = 32'b00000000000000010100110110011111;
assign LUT_3[48360] = 32'b00000000000000010100001110101110;
assign LUT_3[48361] = 32'b00000000000000011010111010001011;
assign LUT_3[48362] = 32'b00000000000000010110010110010010;
assign LUT_3[48363] = 32'b00000000000000011101000001101111;
assign LUT_3[48364] = 32'b00000000000000010001011100100100;
assign LUT_3[48365] = 32'b00000000000000011000001000000001;
assign LUT_3[48366] = 32'b00000000000000010011100100001000;
assign LUT_3[48367] = 32'b00000000000000011010001111100101;
assign LUT_3[48368] = 32'b00000000000000010010001000101011;
assign LUT_3[48369] = 32'b00000000000000011000110100001000;
assign LUT_3[48370] = 32'b00000000000000010100010000001111;
assign LUT_3[48371] = 32'b00000000000000011010111011101100;
assign LUT_3[48372] = 32'b00000000000000001111010110100001;
assign LUT_3[48373] = 32'b00000000000000010110000001111110;
assign LUT_3[48374] = 32'b00000000000000010001011110000101;
assign LUT_3[48375] = 32'b00000000000000011000001001100010;
assign LUT_3[48376] = 32'b00000000000000010111100001110001;
assign LUT_3[48377] = 32'b00000000000000011110001101001110;
assign LUT_3[48378] = 32'b00000000000000011001101001010101;
assign LUT_3[48379] = 32'b00000000000000100000010100110010;
assign LUT_3[48380] = 32'b00000000000000010100101111100111;
assign LUT_3[48381] = 32'b00000000000000011011011011000100;
assign LUT_3[48382] = 32'b00000000000000010110110111001011;
assign LUT_3[48383] = 32'b00000000000000011101100010101000;
assign LUT_3[48384] = 32'b00000000000000000111110011000000;
assign LUT_3[48385] = 32'b00000000000000001110011110011101;
assign LUT_3[48386] = 32'b00000000000000001001111010100100;
assign LUT_3[48387] = 32'b00000000000000010000100110000001;
assign LUT_3[48388] = 32'b00000000000000000101000000110110;
assign LUT_3[48389] = 32'b00000000000000001011101100010011;
assign LUT_3[48390] = 32'b00000000000000000111001000011010;
assign LUT_3[48391] = 32'b00000000000000001101110011110111;
assign LUT_3[48392] = 32'b00000000000000001101001100000110;
assign LUT_3[48393] = 32'b00000000000000010011110111100011;
assign LUT_3[48394] = 32'b00000000000000001111010011101010;
assign LUT_3[48395] = 32'b00000000000000010101111111000111;
assign LUT_3[48396] = 32'b00000000000000001010011001111100;
assign LUT_3[48397] = 32'b00000000000000010001000101011001;
assign LUT_3[48398] = 32'b00000000000000001100100001100000;
assign LUT_3[48399] = 32'b00000000000000010011001100111101;
assign LUT_3[48400] = 32'b00000000000000001011000110000011;
assign LUT_3[48401] = 32'b00000000000000010001110001100000;
assign LUT_3[48402] = 32'b00000000000000001101001101100111;
assign LUT_3[48403] = 32'b00000000000000010011111001000100;
assign LUT_3[48404] = 32'b00000000000000001000010011111001;
assign LUT_3[48405] = 32'b00000000000000001110111111010110;
assign LUT_3[48406] = 32'b00000000000000001010011011011101;
assign LUT_3[48407] = 32'b00000000000000010001000110111010;
assign LUT_3[48408] = 32'b00000000000000010000011111001001;
assign LUT_3[48409] = 32'b00000000000000010111001010100110;
assign LUT_3[48410] = 32'b00000000000000010010100110101101;
assign LUT_3[48411] = 32'b00000000000000011001010010001010;
assign LUT_3[48412] = 32'b00000000000000001101101100111111;
assign LUT_3[48413] = 32'b00000000000000010100011000011100;
assign LUT_3[48414] = 32'b00000000000000001111110100100011;
assign LUT_3[48415] = 32'b00000000000000010110100000000000;
assign LUT_3[48416] = 32'b00000000000000001001000001100000;
assign LUT_3[48417] = 32'b00000000000000001111101100111101;
assign LUT_3[48418] = 32'b00000000000000001011001001000100;
assign LUT_3[48419] = 32'b00000000000000010001110100100001;
assign LUT_3[48420] = 32'b00000000000000000110001111010110;
assign LUT_3[48421] = 32'b00000000000000001100111010110011;
assign LUT_3[48422] = 32'b00000000000000001000010110111010;
assign LUT_3[48423] = 32'b00000000000000001111000010010111;
assign LUT_3[48424] = 32'b00000000000000001110011010100110;
assign LUT_3[48425] = 32'b00000000000000010101000110000011;
assign LUT_3[48426] = 32'b00000000000000010000100010001010;
assign LUT_3[48427] = 32'b00000000000000010111001101100111;
assign LUT_3[48428] = 32'b00000000000000001011101000011100;
assign LUT_3[48429] = 32'b00000000000000010010010011111001;
assign LUT_3[48430] = 32'b00000000000000001101110000000000;
assign LUT_3[48431] = 32'b00000000000000010100011011011101;
assign LUT_3[48432] = 32'b00000000000000001100010100100011;
assign LUT_3[48433] = 32'b00000000000000010011000000000000;
assign LUT_3[48434] = 32'b00000000000000001110011100000111;
assign LUT_3[48435] = 32'b00000000000000010101000111100100;
assign LUT_3[48436] = 32'b00000000000000001001100010011001;
assign LUT_3[48437] = 32'b00000000000000010000001101110110;
assign LUT_3[48438] = 32'b00000000000000001011101001111101;
assign LUT_3[48439] = 32'b00000000000000010010010101011010;
assign LUT_3[48440] = 32'b00000000000000010001101101101001;
assign LUT_3[48441] = 32'b00000000000000011000011001000110;
assign LUT_3[48442] = 32'b00000000000000010011110101001101;
assign LUT_3[48443] = 32'b00000000000000011010100000101010;
assign LUT_3[48444] = 32'b00000000000000001110111011011111;
assign LUT_3[48445] = 32'b00000000000000010101100110111100;
assign LUT_3[48446] = 32'b00000000000000010001000011000011;
assign LUT_3[48447] = 32'b00000000000000010111101110100000;
assign LUT_3[48448] = 32'b00000000000000000111101011101011;
assign LUT_3[48449] = 32'b00000000000000001110010111001000;
assign LUT_3[48450] = 32'b00000000000000001001110011001111;
assign LUT_3[48451] = 32'b00000000000000010000011110101100;
assign LUT_3[48452] = 32'b00000000000000000100111001100001;
assign LUT_3[48453] = 32'b00000000000000001011100100111110;
assign LUT_3[48454] = 32'b00000000000000000111000001000101;
assign LUT_3[48455] = 32'b00000000000000001101101100100010;
assign LUT_3[48456] = 32'b00000000000000001101000100110001;
assign LUT_3[48457] = 32'b00000000000000010011110000001110;
assign LUT_3[48458] = 32'b00000000000000001111001100010101;
assign LUT_3[48459] = 32'b00000000000000010101110111110010;
assign LUT_3[48460] = 32'b00000000000000001010010010100111;
assign LUT_3[48461] = 32'b00000000000000010000111110000100;
assign LUT_3[48462] = 32'b00000000000000001100011010001011;
assign LUT_3[48463] = 32'b00000000000000010011000101101000;
assign LUT_3[48464] = 32'b00000000000000001010111110101110;
assign LUT_3[48465] = 32'b00000000000000010001101010001011;
assign LUT_3[48466] = 32'b00000000000000001101000110010010;
assign LUT_3[48467] = 32'b00000000000000010011110001101111;
assign LUT_3[48468] = 32'b00000000000000001000001100100100;
assign LUT_3[48469] = 32'b00000000000000001110111000000001;
assign LUT_3[48470] = 32'b00000000000000001010010100001000;
assign LUT_3[48471] = 32'b00000000000000010000111111100101;
assign LUT_3[48472] = 32'b00000000000000010000010111110100;
assign LUT_3[48473] = 32'b00000000000000010111000011010001;
assign LUT_3[48474] = 32'b00000000000000010010011111011000;
assign LUT_3[48475] = 32'b00000000000000011001001010110101;
assign LUT_3[48476] = 32'b00000000000000001101100101101010;
assign LUT_3[48477] = 32'b00000000000000010100010001000111;
assign LUT_3[48478] = 32'b00000000000000001111101101001110;
assign LUT_3[48479] = 32'b00000000000000010110011000101011;
assign LUT_3[48480] = 32'b00000000000000001000111010001011;
assign LUT_3[48481] = 32'b00000000000000001111100101101000;
assign LUT_3[48482] = 32'b00000000000000001011000001101111;
assign LUT_3[48483] = 32'b00000000000000010001101101001100;
assign LUT_3[48484] = 32'b00000000000000000110001000000001;
assign LUT_3[48485] = 32'b00000000000000001100110011011110;
assign LUT_3[48486] = 32'b00000000000000001000001111100101;
assign LUT_3[48487] = 32'b00000000000000001110111011000010;
assign LUT_3[48488] = 32'b00000000000000001110010011010001;
assign LUT_3[48489] = 32'b00000000000000010100111110101110;
assign LUT_3[48490] = 32'b00000000000000010000011010110101;
assign LUT_3[48491] = 32'b00000000000000010111000110010010;
assign LUT_3[48492] = 32'b00000000000000001011100001000111;
assign LUT_3[48493] = 32'b00000000000000010010001100100100;
assign LUT_3[48494] = 32'b00000000000000001101101000101011;
assign LUT_3[48495] = 32'b00000000000000010100010100001000;
assign LUT_3[48496] = 32'b00000000000000001100001101001110;
assign LUT_3[48497] = 32'b00000000000000010010111000101011;
assign LUT_3[48498] = 32'b00000000000000001110010100110010;
assign LUT_3[48499] = 32'b00000000000000010101000000001111;
assign LUT_3[48500] = 32'b00000000000000001001011011000100;
assign LUT_3[48501] = 32'b00000000000000010000000110100001;
assign LUT_3[48502] = 32'b00000000000000001011100010101000;
assign LUT_3[48503] = 32'b00000000000000010010001110000101;
assign LUT_3[48504] = 32'b00000000000000010001100110010100;
assign LUT_3[48505] = 32'b00000000000000011000010001110001;
assign LUT_3[48506] = 32'b00000000000000010011101101111000;
assign LUT_3[48507] = 32'b00000000000000011010011001010101;
assign LUT_3[48508] = 32'b00000000000000001110110100001010;
assign LUT_3[48509] = 32'b00000000000000010101011111100111;
assign LUT_3[48510] = 32'b00000000000000010000111011101110;
assign LUT_3[48511] = 32'b00000000000000010111100111001011;
assign LUT_3[48512] = 32'b00000000000000001001111101111110;
assign LUT_3[48513] = 32'b00000000000000010000101001011011;
assign LUT_3[48514] = 32'b00000000000000001100000101100010;
assign LUT_3[48515] = 32'b00000000000000010010110000111111;
assign LUT_3[48516] = 32'b00000000000000000111001011110100;
assign LUT_3[48517] = 32'b00000000000000001101110111010001;
assign LUT_3[48518] = 32'b00000000000000001001010011011000;
assign LUT_3[48519] = 32'b00000000000000001111111110110101;
assign LUT_3[48520] = 32'b00000000000000001111010111000100;
assign LUT_3[48521] = 32'b00000000000000010110000010100001;
assign LUT_3[48522] = 32'b00000000000000010001011110101000;
assign LUT_3[48523] = 32'b00000000000000011000001010000101;
assign LUT_3[48524] = 32'b00000000000000001100100100111010;
assign LUT_3[48525] = 32'b00000000000000010011010000010111;
assign LUT_3[48526] = 32'b00000000000000001110101100011110;
assign LUT_3[48527] = 32'b00000000000000010101010111111011;
assign LUT_3[48528] = 32'b00000000000000001101010001000001;
assign LUT_3[48529] = 32'b00000000000000010011111100011110;
assign LUT_3[48530] = 32'b00000000000000001111011000100101;
assign LUT_3[48531] = 32'b00000000000000010110000100000010;
assign LUT_3[48532] = 32'b00000000000000001010011110110111;
assign LUT_3[48533] = 32'b00000000000000010001001010010100;
assign LUT_3[48534] = 32'b00000000000000001100100110011011;
assign LUT_3[48535] = 32'b00000000000000010011010001111000;
assign LUT_3[48536] = 32'b00000000000000010010101010000111;
assign LUT_3[48537] = 32'b00000000000000011001010101100100;
assign LUT_3[48538] = 32'b00000000000000010100110001101011;
assign LUT_3[48539] = 32'b00000000000000011011011101001000;
assign LUT_3[48540] = 32'b00000000000000001111110111111101;
assign LUT_3[48541] = 32'b00000000000000010110100011011010;
assign LUT_3[48542] = 32'b00000000000000010001111111100001;
assign LUT_3[48543] = 32'b00000000000000011000101010111110;
assign LUT_3[48544] = 32'b00000000000000001011001100011110;
assign LUT_3[48545] = 32'b00000000000000010001110111111011;
assign LUT_3[48546] = 32'b00000000000000001101010100000010;
assign LUT_3[48547] = 32'b00000000000000010011111111011111;
assign LUT_3[48548] = 32'b00000000000000001000011010010100;
assign LUT_3[48549] = 32'b00000000000000001111000101110001;
assign LUT_3[48550] = 32'b00000000000000001010100001111000;
assign LUT_3[48551] = 32'b00000000000000010001001101010101;
assign LUT_3[48552] = 32'b00000000000000010000100101100100;
assign LUT_3[48553] = 32'b00000000000000010111010001000001;
assign LUT_3[48554] = 32'b00000000000000010010101101001000;
assign LUT_3[48555] = 32'b00000000000000011001011000100101;
assign LUT_3[48556] = 32'b00000000000000001101110011011010;
assign LUT_3[48557] = 32'b00000000000000010100011110110111;
assign LUT_3[48558] = 32'b00000000000000001111111010111110;
assign LUT_3[48559] = 32'b00000000000000010110100110011011;
assign LUT_3[48560] = 32'b00000000000000001110011111100001;
assign LUT_3[48561] = 32'b00000000000000010101001010111110;
assign LUT_3[48562] = 32'b00000000000000010000100111000101;
assign LUT_3[48563] = 32'b00000000000000010111010010100010;
assign LUT_3[48564] = 32'b00000000000000001011101101010111;
assign LUT_3[48565] = 32'b00000000000000010010011000110100;
assign LUT_3[48566] = 32'b00000000000000001101110100111011;
assign LUT_3[48567] = 32'b00000000000000010100100000011000;
assign LUT_3[48568] = 32'b00000000000000010011111000100111;
assign LUT_3[48569] = 32'b00000000000000011010100100000100;
assign LUT_3[48570] = 32'b00000000000000010110000000001011;
assign LUT_3[48571] = 32'b00000000000000011100101011101000;
assign LUT_3[48572] = 32'b00000000000000010001000110011101;
assign LUT_3[48573] = 32'b00000000000000010111110001111010;
assign LUT_3[48574] = 32'b00000000000000010011001110000001;
assign LUT_3[48575] = 32'b00000000000000011001111001011110;
assign LUT_3[48576] = 32'b00000000000000001001110110101001;
assign LUT_3[48577] = 32'b00000000000000010000100010000110;
assign LUT_3[48578] = 32'b00000000000000001011111110001101;
assign LUT_3[48579] = 32'b00000000000000010010101001101010;
assign LUT_3[48580] = 32'b00000000000000000111000100011111;
assign LUT_3[48581] = 32'b00000000000000001101101111111100;
assign LUT_3[48582] = 32'b00000000000000001001001100000011;
assign LUT_3[48583] = 32'b00000000000000001111110111100000;
assign LUT_3[48584] = 32'b00000000000000001111001111101111;
assign LUT_3[48585] = 32'b00000000000000010101111011001100;
assign LUT_3[48586] = 32'b00000000000000010001010111010011;
assign LUT_3[48587] = 32'b00000000000000011000000010110000;
assign LUT_3[48588] = 32'b00000000000000001100011101100101;
assign LUT_3[48589] = 32'b00000000000000010011001001000010;
assign LUT_3[48590] = 32'b00000000000000001110100101001001;
assign LUT_3[48591] = 32'b00000000000000010101010000100110;
assign LUT_3[48592] = 32'b00000000000000001101001001101100;
assign LUT_3[48593] = 32'b00000000000000010011110101001001;
assign LUT_3[48594] = 32'b00000000000000001111010001010000;
assign LUT_3[48595] = 32'b00000000000000010101111100101101;
assign LUT_3[48596] = 32'b00000000000000001010010111100010;
assign LUT_3[48597] = 32'b00000000000000010001000010111111;
assign LUT_3[48598] = 32'b00000000000000001100011111000110;
assign LUT_3[48599] = 32'b00000000000000010011001010100011;
assign LUT_3[48600] = 32'b00000000000000010010100010110010;
assign LUT_3[48601] = 32'b00000000000000011001001110001111;
assign LUT_3[48602] = 32'b00000000000000010100101010010110;
assign LUT_3[48603] = 32'b00000000000000011011010101110011;
assign LUT_3[48604] = 32'b00000000000000001111110000101000;
assign LUT_3[48605] = 32'b00000000000000010110011100000101;
assign LUT_3[48606] = 32'b00000000000000010001111000001100;
assign LUT_3[48607] = 32'b00000000000000011000100011101001;
assign LUT_3[48608] = 32'b00000000000000001011000101001001;
assign LUT_3[48609] = 32'b00000000000000010001110000100110;
assign LUT_3[48610] = 32'b00000000000000001101001100101101;
assign LUT_3[48611] = 32'b00000000000000010011111000001010;
assign LUT_3[48612] = 32'b00000000000000001000010010111111;
assign LUT_3[48613] = 32'b00000000000000001110111110011100;
assign LUT_3[48614] = 32'b00000000000000001010011010100011;
assign LUT_3[48615] = 32'b00000000000000010001000110000000;
assign LUT_3[48616] = 32'b00000000000000010000011110001111;
assign LUT_3[48617] = 32'b00000000000000010111001001101100;
assign LUT_3[48618] = 32'b00000000000000010010100101110011;
assign LUT_3[48619] = 32'b00000000000000011001010001010000;
assign LUT_3[48620] = 32'b00000000000000001101101100000101;
assign LUT_3[48621] = 32'b00000000000000010100010111100010;
assign LUT_3[48622] = 32'b00000000000000001111110011101001;
assign LUT_3[48623] = 32'b00000000000000010110011111000110;
assign LUT_3[48624] = 32'b00000000000000001110011000001100;
assign LUT_3[48625] = 32'b00000000000000010101000011101001;
assign LUT_3[48626] = 32'b00000000000000010000011111110000;
assign LUT_3[48627] = 32'b00000000000000010111001011001101;
assign LUT_3[48628] = 32'b00000000000000001011100110000010;
assign LUT_3[48629] = 32'b00000000000000010010010001011111;
assign LUT_3[48630] = 32'b00000000000000001101101101100110;
assign LUT_3[48631] = 32'b00000000000000010100011001000011;
assign LUT_3[48632] = 32'b00000000000000010011110001010010;
assign LUT_3[48633] = 32'b00000000000000011010011100101111;
assign LUT_3[48634] = 32'b00000000000000010101111000110110;
assign LUT_3[48635] = 32'b00000000000000011100100100010011;
assign LUT_3[48636] = 32'b00000000000000010000111111001000;
assign LUT_3[48637] = 32'b00000000000000010111101010100101;
assign LUT_3[48638] = 32'b00000000000000010011000110101100;
assign LUT_3[48639] = 32'b00000000000000011001110010001001;
assign LUT_3[48640] = 32'b00000000000000001110111000101011;
assign LUT_3[48641] = 32'b00000000000000010101100100001000;
assign LUT_3[48642] = 32'b00000000000000010001000000001111;
assign LUT_3[48643] = 32'b00000000000000010111101011101100;
assign LUT_3[48644] = 32'b00000000000000001100000110100001;
assign LUT_3[48645] = 32'b00000000000000010010110001111110;
assign LUT_3[48646] = 32'b00000000000000001110001110000101;
assign LUT_3[48647] = 32'b00000000000000010100111001100010;
assign LUT_3[48648] = 32'b00000000000000010100010001110001;
assign LUT_3[48649] = 32'b00000000000000011010111101001110;
assign LUT_3[48650] = 32'b00000000000000010110011001010101;
assign LUT_3[48651] = 32'b00000000000000011101000100110010;
assign LUT_3[48652] = 32'b00000000000000010001011111100111;
assign LUT_3[48653] = 32'b00000000000000011000001011000100;
assign LUT_3[48654] = 32'b00000000000000010011100111001011;
assign LUT_3[48655] = 32'b00000000000000011010010010101000;
assign LUT_3[48656] = 32'b00000000000000010010001011101110;
assign LUT_3[48657] = 32'b00000000000000011000110111001011;
assign LUT_3[48658] = 32'b00000000000000010100010011010010;
assign LUT_3[48659] = 32'b00000000000000011010111110101111;
assign LUT_3[48660] = 32'b00000000000000001111011001100100;
assign LUT_3[48661] = 32'b00000000000000010110000101000001;
assign LUT_3[48662] = 32'b00000000000000010001100001001000;
assign LUT_3[48663] = 32'b00000000000000011000001100100101;
assign LUT_3[48664] = 32'b00000000000000010111100100110100;
assign LUT_3[48665] = 32'b00000000000000011110010000010001;
assign LUT_3[48666] = 32'b00000000000000011001101100011000;
assign LUT_3[48667] = 32'b00000000000000100000010111110101;
assign LUT_3[48668] = 32'b00000000000000010100110010101010;
assign LUT_3[48669] = 32'b00000000000000011011011110000111;
assign LUT_3[48670] = 32'b00000000000000010110111010001110;
assign LUT_3[48671] = 32'b00000000000000011101100101101011;
assign LUT_3[48672] = 32'b00000000000000010000000111001011;
assign LUT_3[48673] = 32'b00000000000000010110110010101000;
assign LUT_3[48674] = 32'b00000000000000010010001110101111;
assign LUT_3[48675] = 32'b00000000000000011000111010001100;
assign LUT_3[48676] = 32'b00000000000000001101010101000001;
assign LUT_3[48677] = 32'b00000000000000010100000000011110;
assign LUT_3[48678] = 32'b00000000000000001111011100100101;
assign LUT_3[48679] = 32'b00000000000000010110001000000010;
assign LUT_3[48680] = 32'b00000000000000010101100000010001;
assign LUT_3[48681] = 32'b00000000000000011100001011101110;
assign LUT_3[48682] = 32'b00000000000000010111100111110101;
assign LUT_3[48683] = 32'b00000000000000011110010011010010;
assign LUT_3[48684] = 32'b00000000000000010010101110000111;
assign LUT_3[48685] = 32'b00000000000000011001011001100100;
assign LUT_3[48686] = 32'b00000000000000010100110101101011;
assign LUT_3[48687] = 32'b00000000000000011011100001001000;
assign LUT_3[48688] = 32'b00000000000000010011011010001110;
assign LUT_3[48689] = 32'b00000000000000011010000101101011;
assign LUT_3[48690] = 32'b00000000000000010101100001110010;
assign LUT_3[48691] = 32'b00000000000000011100001101001111;
assign LUT_3[48692] = 32'b00000000000000010000101000000100;
assign LUT_3[48693] = 32'b00000000000000010111010011100001;
assign LUT_3[48694] = 32'b00000000000000010010101111101000;
assign LUT_3[48695] = 32'b00000000000000011001011011000101;
assign LUT_3[48696] = 32'b00000000000000011000110011010100;
assign LUT_3[48697] = 32'b00000000000000011111011110110001;
assign LUT_3[48698] = 32'b00000000000000011010111010111000;
assign LUT_3[48699] = 32'b00000000000000100001100110010101;
assign LUT_3[48700] = 32'b00000000000000010110000001001010;
assign LUT_3[48701] = 32'b00000000000000011100101100100111;
assign LUT_3[48702] = 32'b00000000000000011000001000101110;
assign LUT_3[48703] = 32'b00000000000000011110110100001011;
assign LUT_3[48704] = 32'b00000000000000001110110001010110;
assign LUT_3[48705] = 32'b00000000000000010101011100110011;
assign LUT_3[48706] = 32'b00000000000000010000111000111010;
assign LUT_3[48707] = 32'b00000000000000010111100100010111;
assign LUT_3[48708] = 32'b00000000000000001011111111001100;
assign LUT_3[48709] = 32'b00000000000000010010101010101001;
assign LUT_3[48710] = 32'b00000000000000001110000110110000;
assign LUT_3[48711] = 32'b00000000000000010100110010001101;
assign LUT_3[48712] = 32'b00000000000000010100001010011100;
assign LUT_3[48713] = 32'b00000000000000011010110101111001;
assign LUT_3[48714] = 32'b00000000000000010110010010000000;
assign LUT_3[48715] = 32'b00000000000000011100111101011101;
assign LUT_3[48716] = 32'b00000000000000010001011000010010;
assign LUT_3[48717] = 32'b00000000000000011000000011101111;
assign LUT_3[48718] = 32'b00000000000000010011011111110110;
assign LUT_3[48719] = 32'b00000000000000011010001011010011;
assign LUT_3[48720] = 32'b00000000000000010010000100011001;
assign LUT_3[48721] = 32'b00000000000000011000101111110110;
assign LUT_3[48722] = 32'b00000000000000010100001011111101;
assign LUT_3[48723] = 32'b00000000000000011010110111011010;
assign LUT_3[48724] = 32'b00000000000000001111010010001111;
assign LUT_3[48725] = 32'b00000000000000010101111101101100;
assign LUT_3[48726] = 32'b00000000000000010001011001110011;
assign LUT_3[48727] = 32'b00000000000000011000000101010000;
assign LUT_3[48728] = 32'b00000000000000010111011101011111;
assign LUT_3[48729] = 32'b00000000000000011110001000111100;
assign LUT_3[48730] = 32'b00000000000000011001100101000011;
assign LUT_3[48731] = 32'b00000000000000100000010000100000;
assign LUT_3[48732] = 32'b00000000000000010100101011010101;
assign LUT_3[48733] = 32'b00000000000000011011010110110010;
assign LUT_3[48734] = 32'b00000000000000010110110010111001;
assign LUT_3[48735] = 32'b00000000000000011101011110010110;
assign LUT_3[48736] = 32'b00000000000000001111111111110110;
assign LUT_3[48737] = 32'b00000000000000010110101011010011;
assign LUT_3[48738] = 32'b00000000000000010010000111011010;
assign LUT_3[48739] = 32'b00000000000000011000110010110111;
assign LUT_3[48740] = 32'b00000000000000001101001101101100;
assign LUT_3[48741] = 32'b00000000000000010011111001001001;
assign LUT_3[48742] = 32'b00000000000000001111010101010000;
assign LUT_3[48743] = 32'b00000000000000010110000000101101;
assign LUT_3[48744] = 32'b00000000000000010101011000111100;
assign LUT_3[48745] = 32'b00000000000000011100000100011001;
assign LUT_3[48746] = 32'b00000000000000010111100000100000;
assign LUT_3[48747] = 32'b00000000000000011110001011111101;
assign LUT_3[48748] = 32'b00000000000000010010100110110010;
assign LUT_3[48749] = 32'b00000000000000011001010010001111;
assign LUT_3[48750] = 32'b00000000000000010100101110010110;
assign LUT_3[48751] = 32'b00000000000000011011011001110011;
assign LUT_3[48752] = 32'b00000000000000010011010010111001;
assign LUT_3[48753] = 32'b00000000000000011001111110010110;
assign LUT_3[48754] = 32'b00000000000000010101011010011101;
assign LUT_3[48755] = 32'b00000000000000011100000101111010;
assign LUT_3[48756] = 32'b00000000000000010000100000101111;
assign LUT_3[48757] = 32'b00000000000000010111001100001100;
assign LUT_3[48758] = 32'b00000000000000010010101000010011;
assign LUT_3[48759] = 32'b00000000000000011001010011110000;
assign LUT_3[48760] = 32'b00000000000000011000101011111111;
assign LUT_3[48761] = 32'b00000000000000011111010111011100;
assign LUT_3[48762] = 32'b00000000000000011010110011100011;
assign LUT_3[48763] = 32'b00000000000000100001011111000000;
assign LUT_3[48764] = 32'b00000000000000010101111001110101;
assign LUT_3[48765] = 32'b00000000000000011100100101010010;
assign LUT_3[48766] = 32'b00000000000000011000000001011001;
assign LUT_3[48767] = 32'b00000000000000011110101100110110;
assign LUT_3[48768] = 32'b00000000000000010001000011101001;
assign LUT_3[48769] = 32'b00000000000000010111101111000110;
assign LUT_3[48770] = 32'b00000000000000010011001011001101;
assign LUT_3[48771] = 32'b00000000000000011001110110101010;
assign LUT_3[48772] = 32'b00000000000000001110010001011111;
assign LUT_3[48773] = 32'b00000000000000010100111100111100;
assign LUT_3[48774] = 32'b00000000000000010000011001000011;
assign LUT_3[48775] = 32'b00000000000000010111000100100000;
assign LUT_3[48776] = 32'b00000000000000010110011100101111;
assign LUT_3[48777] = 32'b00000000000000011101001000001100;
assign LUT_3[48778] = 32'b00000000000000011000100100010011;
assign LUT_3[48779] = 32'b00000000000000011111001111110000;
assign LUT_3[48780] = 32'b00000000000000010011101010100101;
assign LUT_3[48781] = 32'b00000000000000011010010110000010;
assign LUT_3[48782] = 32'b00000000000000010101110010001001;
assign LUT_3[48783] = 32'b00000000000000011100011101100110;
assign LUT_3[48784] = 32'b00000000000000010100010110101100;
assign LUT_3[48785] = 32'b00000000000000011011000010001001;
assign LUT_3[48786] = 32'b00000000000000010110011110010000;
assign LUT_3[48787] = 32'b00000000000000011101001001101101;
assign LUT_3[48788] = 32'b00000000000000010001100100100010;
assign LUT_3[48789] = 32'b00000000000000011000001111111111;
assign LUT_3[48790] = 32'b00000000000000010011101100000110;
assign LUT_3[48791] = 32'b00000000000000011010010111100011;
assign LUT_3[48792] = 32'b00000000000000011001101111110010;
assign LUT_3[48793] = 32'b00000000000000100000011011001111;
assign LUT_3[48794] = 32'b00000000000000011011110111010110;
assign LUT_3[48795] = 32'b00000000000000100010100010110011;
assign LUT_3[48796] = 32'b00000000000000010110111101101000;
assign LUT_3[48797] = 32'b00000000000000011101101001000101;
assign LUT_3[48798] = 32'b00000000000000011001000101001100;
assign LUT_3[48799] = 32'b00000000000000011111110000101001;
assign LUT_3[48800] = 32'b00000000000000010010010010001001;
assign LUT_3[48801] = 32'b00000000000000011000111101100110;
assign LUT_3[48802] = 32'b00000000000000010100011001101101;
assign LUT_3[48803] = 32'b00000000000000011011000101001010;
assign LUT_3[48804] = 32'b00000000000000001111011111111111;
assign LUT_3[48805] = 32'b00000000000000010110001011011100;
assign LUT_3[48806] = 32'b00000000000000010001100111100011;
assign LUT_3[48807] = 32'b00000000000000011000010011000000;
assign LUT_3[48808] = 32'b00000000000000010111101011001111;
assign LUT_3[48809] = 32'b00000000000000011110010110101100;
assign LUT_3[48810] = 32'b00000000000000011001110010110011;
assign LUT_3[48811] = 32'b00000000000000100000011110010000;
assign LUT_3[48812] = 32'b00000000000000010100111001000101;
assign LUT_3[48813] = 32'b00000000000000011011100100100010;
assign LUT_3[48814] = 32'b00000000000000010111000000101001;
assign LUT_3[48815] = 32'b00000000000000011101101100000110;
assign LUT_3[48816] = 32'b00000000000000010101100101001100;
assign LUT_3[48817] = 32'b00000000000000011100010000101001;
assign LUT_3[48818] = 32'b00000000000000010111101100110000;
assign LUT_3[48819] = 32'b00000000000000011110011000001101;
assign LUT_3[48820] = 32'b00000000000000010010110011000010;
assign LUT_3[48821] = 32'b00000000000000011001011110011111;
assign LUT_3[48822] = 32'b00000000000000010100111010100110;
assign LUT_3[48823] = 32'b00000000000000011011100110000011;
assign LUT_3[48824] = 32'b00000000000000011010111110010010;
assign LUT_3[48825] = 32'b00000000000000100001101001101111;
assign LUT_3[48826] = 32'b00000000000000011101000101110110;
assign LUT_3[48827] = 32'b00000000000000100011110001010011;
assign LUT_3[48828] = 32'b00000000000000011000001100001000;
assign LUT_3[48829] = 32'b00000000000000011110110111100101;
assign LUT_3[48830] = 32'b00000000000000011010010011101100;
assign LUT_3[48831] = 32'b00000000000000100000111111001001;
assign LUT_3[48832] = 32'b00000000000000010000111100010100;
assign LUT_3[48833] = 32'b00000000000000010111100111110001;
assign LUT_3[48834] = 32'b00000000000000010011000011111000;
assign LUT_3[48835] = 32'b00000000000000011001101111010101;
assign LUT_3[48836] = 32'b00000000000000001110001010001010;
assign LUT_3[48837] = 32'b00000000000000010100110101100111;
assign LUT_3[48838] = 32'b00000000000000010000010001101110;
assign LUT_3[48839] = 32'b00000000000000010110111101001011;
assign LUT_3[48840] = 32'b00000000000000010110010101011010;
assign LUT_3[48841] = 32'b00000000000000011101000000110111;
assign LUT_3[48842] = 32'b00000000000000011000011100111110;
assign LUT_3[48843] = 32'b00000000000000011111001000011011;
assign LUT_3[48844] = 32'b00000000000000010011100011010000;
assign LUT_3[48845] = 32'b00000000000000011010001110101101;
assign LUT_3[48846] = 32'b00000000000000010101101010110100;
assign LUT_3[48847] = 32'b00000000000000011100010110010001;
assign LUT_3[48848] = 32'b00000000000000010100001111010111;
assign LUT_3[48849] = 32'b00000000000000011010111010110100;
assign LUT_3[48850] = 32'b00000000000000010110010110111011;
assign LUT_3[48851] = 32'b00000000000000011101000010011000;
assign LUT_3[48852] = 32'b00000000000000010001011101001101;
assign LUT_3[48853] = 32'b00000000000000011000001000101010;
assign LUT_3[48854] = 32'b00000000000000010011100100110001;
assign LUT_3[48855] = 32'b00000000000000011010010000001110;
assign LUT_3[48856] = 32'b00000000000000011001101000011101;
assign LUT_3[48857] = 32'b00000000000000100000010011111010;
assign LUT_3[48858] = 32'b00000000000000011011110000000001;
assign LUT_3[48859] = 32'b00000000000000100010011011011110;
assign LUT_3[48860] = 32'b00000000000000010110110110010011;
assign LUT_3[48861] = 32'b00000000000000011101100001110000;
assign LUT_3[48862] = 32'b00000000000000011000111101110111;
assign LUT_3[48863] = 32'b00000000000000011111101001010100;
assign LUT_3[48864] = 32'b00000000000000010010001010110100;
assign LUT_3[48865] = 32'b00000000000000011000110110010001;
assign LUT_3[48866] = 32'b00000000000000010100010010011000;
assign LUT_3[48867] = 32'b00000000000000011010111101110101;
assign LUT_3[48868] = 32'b00000000000000001111011000101010;
assign LUT_3[48869] = 32'b00000000000000010110000100000111;
assign LUT_3[48870] = 32'b00000000000000010001100000001110;
assign LUT_3[48871] = 32'b00000000000000011000001011101011;
assign LUT_3[48872] = 32'b00000000000000010111100011111010;
assign LUT_3[48873] = 32'b00000000000000011110001111010111;
assign LUT_3[48874] = 32'b00000000000000011001101011011110;
assign LUT_3[48875] = 32'b00000000000000100000010110111011;
assign LUT_3[48876] = 32'b00000000000000010100110001110000;
assign LUT_3[48877] = 32'b00000000000000011011011101001101;
assign LUT_3[48878] = 32'b00000000000000010110111001010100;
assign LUT_3[48879] = 32'b00000000000000011101100100110001;
assign LUT_3[48880] = 32'b00000000000000010101011101110111;
assign LUT_3[48881] = 32'b00000000000000011100001001010100;
assign LUT_3[48882] = 32'b00000000000000010111100101011011;
assign LUT_3[48883] = 32'b00000000000000011110010000111000;
assign LUT_3[48884] = 32'b00000000000000010010101011101101;
assign LUT_3[48885] = 32'b00000000000000011001010111001010;
assign LUT_3[48886] = 32'b00000000000000010100110011010001;
assign LUT_3[48887] = 32'b00000000000000011011011110101110;
assign LUT_3[48888] = 32'b00000000000000011010110110111101;
assign LUT_3[48889] = 32'b00000000000000100001100010011010;
assign LUT_3[48890] = 32'b00000000000000011100111110100001;
assign LUT_3[48891] = 32'b00000000000000100011101001111110;
assign LUT_3[48892] = 32'b00000000000000011000000100110011;
assign LUT_3[48893] = 32'b00000000000000011110110000010000;
assign LUT_3[48894] = 32'b00000000000000011010001100010111;
assign LUT_3[48895] = 32'b00000000000000100000110111110100;
assign LUT_3[48896] = 32'b00000000000000001011001000001100;
assign LUT_3[48897] = 32'b00000000000000010001110011101001;
assign LUT_3[48898] = 32'b00000000000000001101001111110000;
assign LUT_3[48899] = 32'b00000000000000010011111011001101;
assign LUT_3[48900] = 32'b00000000000000001000010110000010;
assign LUT_3[48901] = 32'b00000000000000001111000001011111;
assign LUT_3[48902] = 32'b00000000000000001010011101100110;
assign LUT_3[48903] = 32'b00000000000000010001001001000011;
assign LUT_3[48904] = 32'b00000000000000010000100001010010;
assign LUT_3[48905] = 32'b00000000000000010111001100101111;
assign LUT_3[48906] = 32'b00000000000000010010101000110110;
assign LUT_3[48907] = 32'b00000000000000011001010100010011;
assign LUT_3[48908] = 32'b00000000000000001101101111001000;
assign LUT_3[48909] = 32'b00000000000000010100011010100101;
assign LUT_3[48910] = 32'b00000000000000001111110110101100;
assign LUT_3[48911] = 32'b00000000000000010110100010001001;
assign LUT_3[48912] = 32'b00000000000000001110011011001111;
assign LUT_3[48913] = 32'b00000000000000010101000110101100;
assign LUT_3[48914] = 32'b00000000000000010000100010110011;
assign LUT_3[48915] = 32'b00000000000000010111001110010000;
assign LUT_3[48916] = 32'b00000000000000001011101001000101;
assign LUT_3[48917] = 32'b00000000000000010010010100100010;
assign LUT_3[48918] = 32'b00000000000000001101110000101001;
assign LUT_3[48919] = 32'b00000000000000010100011100000110;
assign LUT_3[48920] = 32'b00000000000000010011110100010101;
assign LUT_3[48921] = 32'b00000000000000011010011111110010;
assign LUT_3[48922] = 32'b00000000000000010101111011111001;
assign LUT_3[48923] = 32'b00000000000000011100100111010110;
assign LUT_3[48924] = 32'b00000000000000010001000010001011;
assign LUT_3[48925] = 32'b00000000000000010111101101101000;
assign LUT_3[48926] = 32'b00000000000000010011001001101111;
assign LUT_3[48927] = 32'b00000000000000011001110101001100;
assign LUT_3[48928] = 32'b00000000000000001100010110101100;
assign LUT_3[48929] = 32'b00000000000000010011000010001001;
assign LUT_3[48930] = 32'b00000000000000001110011110010000;
assign LUT_3[48931] = 32'b00000000000000010101001001101101;
assign LUT_3[48932] = 32'b00000000000000001001100100100010;
assign LUT_3[48933] = 32'b00000000000000010000001111111111;
assign LUT_3[48934] = 32'b00000000000000001011101100000110;
assign LUT_3[48935] = 32'b00000000000000010010010111100011;
assign LUT_3[48936] = 32'b00000000000000010001101111110010;
assign LUT_3[48937] = 32'b00000000000000011000011011001111;
assign LUT_3[48938] = 32'b00000000000000010011110111010110;
assign LUT_3[48939] = 32'b00000000000000011010100010110011;
assign LUT_3[48940] = 32'b00000000000000001110111101101000;
assign LUT_3[48941] = 32'b00000000000000010101101001000101;
assign LUT_3[48942] = 32'b00000000000000010001000101001100;
assign LUT_3[48943] = 32'b00000000000000010111110000101001;
assign LUT_3[48944] = 32'b00000000000000001111101001101111;
assign LUT_3[48945] = 32'b00000000000000010110010101001100;
assign LUT_3[48946] = 32'b00000000000000010001110001010011;
assign LUT_3[48947] = 32'b00000000000000011000011100110000;
assign LUT_3[48948] = 32'b00000000000000001100110111100101;
assign LUT_3[48949] = 32'b00000000000000010011100011000010;
assign LUT_3[48950] = 32'b00000000000000001110111111001001;
assign LUT_3[48951] = 32'b00000000000000010101101010100110;
assign LUT_3[48952] = 32'b00000000000000010101000010110101;
assign LUT_3[48953] = 32'b00000000000000011011101110010010;
assign LUT_3[48954] = 32'b00000000000000010111001010011001;
assign LUT_3[48955] = 32'b00000000000000011101110101110110;
assign LUT_3[48956] = 32'b00000000000000010010010000101011;
assign LUT_3[48957] = 32'b00000000000000011000111100001000;
assign LUT_3[48958] = 32'b00000000000000010100011000001111;
assign LUT_3[48959] = 32'b00000000000000011011000011101100;
assign LUT_3[48960] = 32'b00000000000000001011000000110111;
assign LUT_3[48961] = 32'b00000000000000010001101100010100;
assign LUT_3[48962] = 32'b00000000000000001101001000011011;
assign LUT_3[48963] = 32'b00000000000000010011110011111000;
assign LUT_3[48964] = 32'b00000000000000001000001110101101;
assign LUT_3[48965] = 32'b00000000000000001110111010001010;
assign LUT_3[48966] = 32'b00000000000000001010010110010001;
assign LUT_3[48967] = 32'b00000000000000010001000001101110;
assign LUT_3[48968] = 32'b00000000000000010000011001111101;
assign LUT_3[48969] = 32'b00000000000000010111000101011010;
assign LUT_3[48970] = 32'b00000000000000010010100001100001;
assign LUT_3[48971] = 32'b00000000000000011001001100111110;
assign LUT_3[48972] = 32'b00000000000000001101100111110011;
assign LUT_3[48973] = 32'b00000000000000010100010011010000;
assign LUT_3[48974] = 32'b00000000000000001111101111010111;
assign LUT_3[48975] = 32'b00000000000000010110011010110100;
assign LUT_3[48976] = 32'b00000000000000001110010011111010;
assign LUT_3[48977] = 32'b00000000000000010100111111010111;
assign LUT_3[48978] = 32'b00000000000000010000011011011110;
assign LUT_3[48979] = 32'b00000000000000010111000110111011;
assign LUT_3[48980] = 32'b00000000000000001011100001110000;
assign LUT_3[48981] = 32'b00000000000000010010001101001101;
assign LUT_3[48982] = 32'b00000000000000001101101001010100;
assign LUT_3[48983] = 32'b00000000000000010100010100110001;
assign LUT_3[48984] = 32'b00000000000000010011101101000000;
assign LUT_3[48985] = 32'b00000000000000011010011000011101;
assign LUT_3[48986] = 32'b00000000000000010101110100100100;
assign LUT_3[48987] = 32'b00000000000000011100100000000001;
assign LUT_3[48988] = 32'b00000000000000010000111010110110;
assign LUT_3[48989] = 32'b00000000000000010111100110010011;
assign LUT_3[48990] = 32'b00000000000000010011000010011010;
assign LUT_3[48991] = 32'b00000000000000011001101101110111;
assign LUT_3[48992] = 32'b00000000000000001100001111010111;
assign LUT_3[48993] = 32'b00000000000000010010111010110100;
assign LUT_3[48994] = 32'b00000000000000001110010110111011;
assign LUT_3[48995] = 32'b00000000000000010101000010011000;
assign LUT_3[48996] = 32'b00000000000000001001011101001101;
assign LUT_3[48997] = 32'b00000000000000010000001000101010;
assign LUT_3[48998] = 32'b00000000000000001011100100110001;
assign LUT_3[48999] = 32'b00000000000000010010010000001110;
assign LUT_3[49000] = 32'b00000000000000010001101000011101;
assign LUT_3[49001] = 32'b00000000000000011000010011111010;
assign LUT_3[49002] = 32'b00000000000000010011110000000001;
assign LUT_3[49003] = 32'b00000000000000011010011011011110;
assign LUT_3[49004] = 32'b00000000000000001110110110010011;
assign LUT_3[49005] = 32'b00000000000000010101100001110000;
assign LUT_3[49006] = 32'b00000000000000010000111101110111;
assign LUT_3[49007] = 32'b00000000000000010111101001010100;
assign LUT_3[49008] = 32'b00000000000000001111100010011010;
assign LUT_3[49009] = 32'b00000000000000010110001101110111;
assign LUT_3[49010] = 32'b00000000000000010001101001111110;
assign LUT_3[49011] = 32'b00000000000000011000010101011011;
assign LUT_3[49012] = 32'b00000000000000001100110000010000;
assign LUT_3[49013] = 32'b00000000000000010011011011101101;
assign LUT_3[49014] = 32'b00000000000000001110110111110100;
assign LUT_3[49015] = 32'b00000000000000010101100011010001;
assign LUT_3[49016] = 32'b00000000000000010100111011100000;
assign LUT_3[49017] = 32'b00000000000000011011100110111101;
assign LUT_3[49018] = 32'b00000000000000010111000011000100;
assign LUT_3[49019] = 32'b00000000000000011101101110100001;
assign LUT_3[49020] = 32'b00000000000000010010001001010110;
assign LUT_3[49021] = 32'b00000000000000011000110100110011;
assign LUT_3[49022] = 32'b00000000000000010100010000111010;
assign LUT_3[49023] = 32'b00000000000000011010111100010111;
assign LUT_3[49024] = 32'b00000000000000001101010011001010;
assign LUT_3[49025] = 32'b00000000000000010011111110100111;
assign LUT_3[49026] = 32'b00000000000000001111011010101110;
assign LUT_3[49027] = 32'b00000000000000010110000110001011;
assign LUT_3[49028] = 32'b00000000000000001010100001000000;
assign LUT_3[49029] = 32'b00000000000000010001001100011101;
assign LUT_3[49030] = 32'b00000000000000001100101000100100;
assign LUT_3[49031] = 32'b00000000000000010011010100000001;
assign LUT_3[49032] = 32'b00000000000000010010101100010000;
assign LUT_3[49033] = 32'b00000000000000011001010111101101;
assign LUT_3[49034] = 32'b00000000000000010100110011110100;
assign LUT_3[49035] = 32'b00000000000000011011011111010001;
assign LUT_3[49036] = 32'b00000000000000001111111010000110;
assign LUT_3[49037] = 32'b00000000000000010110100101100011;
assign LUT_3[49038] = 32'b00000000000000010010000001101010;
assign LUT_3[49039] = 32'b00000000000000011000101101000111;
assign LUT_3[49040] = 32'b00000000000000010000100110001101;
assign LUT_3[49041] = 32'b00000000000000010111010001101010;
assign LUT_3[49042] = 32'b00000000000000010010101101110001;
assign LUT_3[49043] = 32'b00000000000000011001011001001110;
assign LUT_3[49044] = 32'b00000000000000001101110100000011;
assign LUT_3[49045] = 32'b00000000000000010100011111100000;
assign LUT_3[49046] = 32'b00000000000000001111111011100111;
assign LUT_3[49047] = 32'b00000000000000010110100111000100;
assign LUT_3[49048] = 32'b00000000000000010101111111010011;
assign LUT_3[49049] = 32'b00000000000000011100101010110000;
assign LUT_3[49050] = 32'b00000000000000011000000110110111;
assign LUT_3[49051] = 32'b00000000000000011110110010010100;
assign LUT_3[49052] = 32'b00000000000000010011001101001001;
assign LUT_3[49053] = 32'b00000000000000011001111000100110;
assign LUT_3[49054] = 32'b00000000000000010101010100101101;
assign LUT_3[49055] = 32'b00000000000000011100000000001010;
assign LUT_3[49056] = 32'b00000000000000001110100001101010;
assign LUT_3[49057] = 32'b00000000000000010101001101000111;
assign LUT_3[49058] = 32'b00000000000000010000101001001110;
assign LUT_3[49059] = 32'b00000000000000010111010100101011;
assign LUT_3[49060] = 32'b00000000000000001011101111100000;
assign LUT_3[49061] = 32'b00000000000000010010011010111101;
assign LUT_3[49062] = 32'b00000000000000001101110111000100;
assign LUT_3[49063] = 32'b00000000000000010100100010100001;
assign LUT_3[49064] = 32'b00000000000000010011111010110000;
assign LUT_3[49065] = 32'b00000000000000011010100110001101;
assign LUT_3[49066] = 32'b00000000000000010110000010010100;
assign LUT_3[49067] = 32'b00000000000000011100101101110001;
assign LUT_3[49068] = 32'b00000000000000010001001000100110;
assign LUT_3[49069] = 32'b00000000000000010111110100000011;
assign LUT_3[49070] = 32'b00000000000000010011010000001010;
assign LUT_3[49071] = 32'b00000000000000011001111011100111;
assign LUT_3[49072] = 32'b00000000000000010001110100101101;
assign LUT_3[49073] = 32'b00000000000000011000100000001010;
assign LUT_3[49074] = 32'b00000000000000010011111100010001;
assign LUT_3[49075] = 32'b00000000000000011010100111101110;
assign LUT_3[49076] = 32'b00000000000000001111000010100011;
assign LUT_3[49077] = 32'b00000000000000010101101110000000;
assign LUT_3[49078] = 32'b00000000000000010001001010000111;
assign LUT_3[49079] = 32'b00000000000000010111110101100100;
assign LUT_3[49080] = 32'b00000000000000010111001101110011;
assign LUT_3[49081] = 32'b00000000000000011101111001010000;
assign LUT_3[49082] = 32'b00000000000000011001010101010111;
assign LUT_3[49083] = 32'b00000000000000100000000000110100;
assign LUT_3[49084] = 32'b00000000000000010100011011101001;
assign LUT_3[49085] = 32'b00000000000000011011000111000110;
assign LUT_3[49086] = 32'b00000000000000010110100011001101;
assign LUT_3[49087] = 32'b00000000000000011101001110101010;
assign LUT_3[49088] = 32'b00000000000000001101001011110101;
assign LUT_3[49089] = 32'b00000000000000010011110111010010;
assign LUT_3[49090] = 32'b00000000000000001111010011011001;
assign LUT_3[49091] = 32'b00000000000000010101111110110110;
assign LUT_3[49092] = 32'b00000000000000001010011001101011;
assign LUT_3[49093] = 32'b00000000000000010001000101001000;
assign LUT_3[49094] = 32'b00000000000000001100100001001111;
assign LUT_3[49095] = 32'b00000000000000010011001100101100;
assign LUT_3[49096] = 32'b00000000000000010010100100111011;
assign LUT_3[49097] = 32'b00000000000000011001010000011000;
assign LUT_3[49098] = 32'b00000000000000010100101100011111;
assign LUT_3[49099] = 32'b00000000000000011011010111111100;
assign LUT_3[49100] = 32'b00000000000000001111110010110001;
assign LUT_3[49101] = 32'b00000000000000010110011110001110;
assign LUT_3[49102] = 32'b00000000000000010001111010010101;
assign LUT_3[49103] = 32'b00000000000000011000100101110010;
assign LUT_3[49104] = 32'b00000000000000010000011110111000;
assign LUT_3[49105] = 32'b00000000000000010111001010010101;
assign LUT_3[49106] = 32'b00000000000000010010100110011100;
assign LUT_3[49107] = 32'b00000000000000011001010001111001;
assign LUT_3[49108] = 32'b00000000000000001101101100101110;
assign LUT_3[49109] = 32'b00000000000000010100011000001011;
assign LUT_3[49110] = 32'b00000000000000001111110100010010;
assign LUT_3[49111] = 32'b00000000000000010110011111101111;
assign LUT_3[49112] = 32'b00000000000000010101110111111110;
assign LUT_3[49113] = 32'b00000000000000011100100011011011;
assign LUT_3[49114] = 32'b00000000000000010111111111100010;
assign LUT_3[49115] = 32'b00000000000000011110101010111111;
assign LUT_3[49116] = 32'b00000000000000010011000101110100;
assign LUT_3[49117] = 32'b00000000000000011001110001010001;
assign LUT_3[49118] = 32'b00000000000000010101001101011000;
assign LUT_3[49119] = 32'b00000000000000011011111000110101;
assign LUT_3[49120] = 32'b00000000000000001110011010010101;
assign LUT_3[49121] = 32'b00000000000000010101000101110010;
assign LUT_3[49122] = 32'b00000000000000010000100001111001;
assign LUT_3[49123] = 32'b00000000000000010111001101010110;
assign LUT_3[49124] = 32'b00000000000000001011101000001011;
assign LUT_3[49125] = 32'b00000000000000010010010011101000;
assign LUT_3[49126] = 32'b00000000000000001101101111101111;
assign LUT_3[49127] = 32'b00000000000000010100011011001100;
assign LUT_3[49128] = 32'b00000000000000010011110011011011;
assign LUT_3[49129] = 32'b00000000000000011010011110111000;
assign LUT_3[49130] = 32'b00000000000000010101111010111111;
assign LUT_3[49131] = 32'b00000000000000011100100110011100;
assign LUT_3[49132] = 32'b00000000000000010001000001010001;
assign LUT_3[49133] = 32'b00000000000000010111101100101110;
assign LUT_3[49134] = 32'b00000000000000010011001000110101;
assign LUT_3[49135] = 32'b00000000000000011001110100010010;
assign LUT_3[49136] = 32'b00000000000000010001101101011000;
assign LUT_3[49137] = 32'b00000000000000011000011000110101;
assign LUT_3[49138] = 32'b00000000000000010011110100111100;
assign LUT_3[49139] = 32'b00000000000000011010100000011001;
assign LUT_3[49140] = 32'b00000000000000001110111011001110;
assign LUT_3[49141] = 32'b00000000000000010101100110101011;
assign LUT_3[49142] = 32'b00000000000000010001000010110010;
assign LUT_3[49143] = 32'b00000000000000010111101110001111;
assign LUT_3[49144] = 32'b00000000000000010111000110011110;
assign LUT_3[49145] = 32'b00000000000000011101110001111011;
assign LUT_3[49146] = 32'b00000000000000011001001110000010;
assign LUT_3[49147] = 32'b00000000000000011111111001011111;
assign LUT_3[49148] = 32'b00000000000000010100010100010100;
assign LUT_3[49149] = 32'b00000000000000011010111111110001;
assign LUT_3[49150] = 32'b00000000000000010110011011111000;
assign LUT_3[49151] = 32'b00000000000000011101000111010101;
assign LUT_3[49152] = 32'b11111111111111111101010000000101;
assign LUT_3[49153] = 32'b00000000000000000011111011100010;
assign LUT_3[49154] = 32'b11111111111111111111010111101001;
assign LUT_3[49155] = 32'b00000000000000000110000011000110;
assign LUT_3[49156] = 32'b11111111111111111010011101111011;
assign LUT_3[49157] = 32'b00000000000000000001001001011000;
assign LUT_3[49158] = 32'b11111111111111111100100101011111;
assign LUT_3[49159] = 32'b00000000000000000011010000111100;
assign LUT_3[49160] = 32'b00000000000000000010101001001011;
assign LUT_3[49161] = 32'b00000000000000001001010100101000;
assign LUT_3[49162] = 32'b00000000000000000100110000101111;
assign LUT_3[49163] = 32'b00000000000000001011011100001100;
assign LUT_3[49164] = 32'b11111111111111111111110111000001;
assign LUT_3[49165] = 32'b00000000000000000110100010011110;
assign LUT_3[49166] = 32'b00000000000000000001111110100101;
assign LUT_3[49167] = 32'b00000000000000001000101010000010;
assign LUT_3[49168] = 32'b00000000000000000000100011001000;
assign LUT_3[49169] = 32'b00000000000000000111001110100101;
assign LUT_3[49170] = 32'b00000000000000000010101010101100;
assign LUT_3[49171] = 32'b00000000000000001001010110001001;
assign LUT_3[49172] = 32'b11111111111111111101110000111110;
assign LUT_3[49173] = 32'b00000000000000000100011100011011;
assign LUT_3[49174] = 32'b11111111111111111111111000100010;
assign LUT_3[49175] = 32'b00000000000000000110100011111111;
assign LUT_3[49176] = 32'b00000000000000000101111100001110;
assign LUT_3[49177] = 32'b00000000000000001100100111101011;
assign LUT_3[49178] = 32'b00000000000000001000000011110010;
assign LUT_3[49179] = 32'b00000000000000001110101111001111;
assign LUT_3[49180] = 32'b00000000000000000011001010000100;
assign LUT_3[49181] = 32'b00000000000000001001110101100001;
assign LUT_3[49182] = 32'b00000000000000000101010001101000;
assign LUT_3[49183] = 32'b00000000000000001011111101000101;
assign LUT_3[49184] = 32'b11111111111111111110011110100101;
assign LUT_3[49185] = 32'b00000000000000000101001010000010;
assign LUT_3[49186] = 32'b00000000000000000000100110001001;
assign LUT_3[49187] = 32'b00000000000000000111010001100110;
assign LUT_3[49188] = 32'b11111111111111111011101100011011;
assign LUT_3[49189] = 32'b00000000000000000010010111111000;
assign LUT_3[49190] = 32'b11111111111111111101110011111111;
assign LUT_3[49191] = 32'b00000000000000000100011111011100;
assign LUT_3[49192] = 32'b00000000000000000011110111101011;
assign LUT_3[49193] = 32'b00000000000000001010100011001000;
assign LUT_3[49194] = 32'b00000000000000000101111111001111;
assign LUT_3[49195] = 32'b00000000000000001100101010101100;
assign LUT_3[49196] = 32'b00000000000000000001000101100001;
assign LUT_3[49197] = 32'b00000000000000000111110000111110;
assign LUT_3[49198] = 32'b00000000000000000011001101000101;
assign LUT_3[49199] = 32'b00000000000000001001111000100010;
assign LUT_3[49200] = 32'b00000000000000000001110001101000;
assign LUT_3[49201] = 32'b00000000000000001000011101000101;
assign LUT_3[49202] = 32'b00000000000000000011111001001100;
assign LUT_3[49203] = 32'b00000000000000001010100100101001;
assign LUT_3[49204] = 32'b11111111111111111110111111011110;
assign LUT_3[49205] = 32'b00000000000000000101101010111011;
assign LUT_3[49206] = 32'b00000000000000000001000111000010;
assign LUT_3[49207] = 32'b00000000000000000111110010011111;
assign LUT_3[49208] = 32'b00000000000000000111001010101110;
assign LUT_3[49209] = 32'b00000000000000001101110110001011;
assign LUT_3[49210] = 32'b00000000000000001001010010010010;
assign LUT_3[49211] = 32'b00000000000000001111111101101111;
assign LUT_3[49212] = 32'b00000000000000000100011000100100;
assign LUT_3[49213] = 32'b00000000000000001011000100000001;
assign LUT_3[49214] = 32'b00000000000000000110100000001000;
assign LUT_3[49215] = 32'b00000000000000001101001011100101;
assign LUT_3[49216] = 32'b11111111111111111101001000110000;
assign LUT_3[49217] = 32'b00000000000000000011110100001101;
assign LUT_3[49218] = 32'b11111111111111111111010000010100;
assign LUT_3[49219] = 32'b00000000000000000101111011110001;
assign LUT_3[49220] = 32'b11111111111111111010010110100110;
assign LUT_3[49221] = 32'b00000000000000000001000010000011;
assign LUT_3[49222] = 32'b11111111111111111100011110001010;
assign LUT_3[49223] = 32'b00000000000000000011001001100111;
assign LUT_3[49224] = 32'b00000000000000000010100001110110;
assign LUT_3[49225] = 32'b00000000000000001001001101010011;
assign LUT_3[49226] = 32'b00000000000000000100101001011010;
assign LUT_3[49227] = 32'b00000000000000001011010100110111;
assign LUT_3[49228] = 32'b11111111111111111111101111101100;
assign LUT_3[49229] = 32'b00000000000000000110011011001001;
assign LUT_3[49230] = 32'b00000000000000000001110111010000;
assign LUT_3[49231] = 32'b00000000000000001000100010101101;
assign LUT_3[49232] = 32'b00000000000000000000011011110011;
assign LUT_3[49233] = 32'b00000000000000000111000111010000;
assign LUT_3[49234] = 32'b00000000000000000010100011010111;
assign LUT_3[49235] = 32'b00000000000000001001001110110100;
assign LUT_3[49236] = 32'b11111111111111111101101001101001;
assign LUT_3[49237] = 32'b00000000000000000100010101000110;
assign LUT_3[49238] = 32'b11111111111111111111110001001101;
assign LUT_3[49239] = 32'b00000000000000000110011100101010;
assign LUT_3[49240] = 32'b00000000000000000101110100111001;
assign LUT_3[49241] = 32'b00000000000000001100100000010110;
assign LUT_3[49242] = 32'b00000000000000000111111100011101;
assign LUT_3[49243] = 32'b00000000000000001110100111111010;
assign LUT_3[49244] = 32'b00000000000000000011000010101111;
assign LUT_3[49245] = 32'b00000000000000001001101110001100;
assign LUT_3[49246] = 32'b00000000000000000101001010010011;
assign LUT_3[49247] = 32'b00000000000000001011110101110000;
assign LUT_3[49248] = 32'b11111111111111111110010111010000;
assign LUT_3[49249] = 32'b00000000000000000101000010101101;
assign LUT_3[49250] = 32'b00000000000000000000011110110100;
assign LUT_3[49251] = 32'b00000000000000000111001010010001;
assign LUT_3[49252] = 32'b11111111111111111011100101000110;
assign LUT_3[49253] = 32'b00000000000000000010010000100011;
assign LUT_3[49254] = 32'b11111111111111111101101100101010;
assign LUT_3[49255] = 32'b00000000000000000100011000000111;
assign LUT_3[49256] = 32'b00000000000000000011110000010110;
assign LUT_3[49257] = 32'b00000000000000001010011011110011;
assign LUT_3[49258] = 32'b00000000000000000101110111111010;
assign LUT_3[49259] = 32'b00000000000000001100100011010111;
assign LUT_3[49260] = 32'b00000000000000000000111110001100;
assign LUT_3[49261] = 32'b00000000000000000111101001101001;
assign LUT_3[49262] = 32'b00000000000000000011000101110000;
assign LUT_3[49263] = 32'b00000000000000001001110001001101;
assign LUT_3[49264] = 32'b00000000000000000001101010010011;
assign LUT_3[49265] = 32'b00000000000000001000010101110000;
assign LUT_3[49266] = 32'b00000000000000000011110001110111;
assign LUT_3[49267] = 32'b00000000000000001010011101010100;
assign LUT_3[49268] = 32'b11111111111111111110111000001001;
assign LUT_3[49269] = 32'b00000000000000000101100011100110;
assign LUT_3[49270] = 32'b00000000000000000000111111101101;
assign LUT_3[49271] = 32'b00000000000000000111101011001010;
assign LUT_3[49272] = 32'b00000000000000000111000011011001;
assign LUT_3[49273] = 32'b00000000000000001101101110110110;
assign LUT_3[49274] = 32'b00000000000000001001001010111101;
assign LUT_3[49275] = 32'b00000000000000001111110110011010;
assign LUT_3[49276] = 32'b00000000000000000100010001001111;
assign LUT_3[49277] = 32'b00000000000000001010111100101100;
assign LUT_3[49278] = 32'b00000000000000000110011000110011;
assign LUT_3[49279] = 32'b00000000000000001101000100010000;
assign LUT_3[49280] = 32'b11111111111111111111011011000011;
assign LUT_3[49281] = 32'b00000000000000000110000110100000;
assign LUT_3[49282] = 32'b00000000000000000001100010100111;
assign LUT_3[49283] = 32'b00000000000000001000001110000100;
assign LUT_3[49284] = 32'b11111111111111111100101000111001;
assign LUT_3[49285] = 32'b00000000000000000011010100010110;
assign LUT_3[49286] = 32'b11111111111111111110110000011101;
assign LUT_3[49287] = 32'b00000000000000000101011011111010;
assign LUT_3[49288] = 32'b00000000000000000100110100001001;
assign LUT_3[49289] = 32'b00000000000000001011011111100110;
assign LUT_3[49290] = 32'b00000000000000000110111011101101;
assign LUT_3[49291] = 32'b00000000000000001101100111001010;
assign LUT_3[49292] = 32'b00000000000000000010000001111111;
assign LUT_3[49293] = 32'b00000000000000001000101101011100;
assign LUT_3[49294] = 32'b00000000000000000100001001100011;
assign LUT_3[49295] = 32'b00000000000000001010110101000000;
assign LUT_3[49296] = 32'b00000000000000000010101110000110;
assign LUT_3[49297] = 32'b00000000000000001001011001100011;
assign LUT_3[49298] = 32'b00000000000000000100110101101010;
assign LUT_3[49299] = 32'b00000000000000001011100001000111;
assign LUT_3[49300] = 32'b11111111111111111111111011111100;
assign LUT_3[49301] = 32'b00000000000000000110100111011001;
assign LUT_3[49302] = 32'b00000000000000000010000011100000;
assign LUT_3[49303] = 32'b00000000000000001000101110111101;
assign LUT_3[49304] = 32'b00000000000000001000000111001100;
assign LUT_3[49305] = 32'b00000000000000001110110010101001;
assign LUT_3[49306] = 32'b00000000000000001010001110110000;
assign LUT_3[49307] = 32'b00000000000000010000111010001101;
assign LUT_3[49308] = 32'b00000000000000000101010101000010;
assign LUT_3[49309] = 32'b00000000000000001100000000011111;
assign LUT_3[49310] = 32'b00000000000000000111011100100110;
assign LUT_3[49311] = 32'b00000000000000001110001000000011;
assign LUT_3[49312] = 32'b00000000000000000000101001100011;
assign LUT_3[49313] = 32'b00000000000000000111010101000000;
assign LUT_3[49314] = 32'b00000000000000000010110001000111;
assign LUT_3[49315] = 32'b00000000000000001001011100100100;
assign LUT_3[49316] = 32'b11111111111111111101110111011001;
assign LUT_3[49317] = 32'b00000000000000000100100010110110;
assign LUT_3[49318] = 32'b11111111111111111111111110111101;
assign LUT_3[49319] = 32'b00000000000000000110101010011010;
assign LUT_3[49320] = 32'b00000000000000000110000010101001;
assign LUT_3[49321] = 32'b00000000000000001100101110000110;
assign LUT_3[49322] = 32'b00000000000000001000001010001101;
assign LUT_3[49323] = 32'b00000000000000001110110101101010;
assign LUT_3[49324] = 32'b00000000000000000011010000011111;
assign LUT_3[49325] = 32'b00000000000000001001111011111100;
assign LUT_3[49326] = 32'b00000000000000000101011000000011;
assign LUT_3[49327] = 32'b00000000000000001100000011100000;
assign LUT_3[49328] = 32'b00000000000000000011111100100110;
assign LUT_3[49329] = 32'b00000000000000001010101000000011;
assign LUT_3[49330] = 32'b00000000000000000110000100001010;
assign LUT_3[49331] = 32'b00000000000000001100101111100111;
assign LUT_3[49332] = 32'b00000000000000000001001010011100;
assign LUT_3[49333] = 32'b00000000000000000111110101111001;
assign LUT_3[49334] = 32'b00000000000000000011010010000000;
assign LUT_3[49335] = 32'b00000000000000001001111101011101;
assign LUT_3[49336] = 32'b00000000000000001001010101101100;
assign LUT_3[49337] = 32'b00000000000000010000000001001001;
assign LUT_3[49338] = 32'b00000000000000001011011101010000;
assign LUT_3[49339] = 32'b00000000000000010010001000101101;
assign LUT_3[49340] = 32'b00000000000000000110100011100010;
assign LUT_3[49341] = 32'b00000000000000001101001110111111;
assign LUT_3[49342] = 32'b00000000000000001000101011000110;
assign LUT_3[49343] = 32'b00000000000000001111010110100011;
assign LUT_3[49344] = 32'b11111111111111111111010011101110;
assign LUT_3[49345] = 32'b00000000000000000101111111001011;
assign LUT_3[49346] = 32'b00000000000000000001011011010010;
assign LUT_3[49347] = 32'b00000000000000001000000110101111;
assign LUT_3[49348] = 32'b11111111111111111100100001100100;
assign LUT_3[49349] = 32'b00000000000000000011001101000001;
assign LUT_3[49350] = 32'b11111111111111111110101001001000;
assign LUT_3[49351] = 32'b00000000000000000101010100100101;
assign LUT_3[49352] = 32'b00000000000000000100101100110100;
assign LUT_3[49353] = 32'b00000000000000001011011000010001;
assign LUT_3[49354] = 32'b00000000000000000110110100011000;
assign LUT_3[49355] = 32'b00000000000000001101011111110101;
assign LUT_3[49356] = 32'b00000000000000000001111010101010;
assign LUT_3[49357] = 32'b00000000000000001000100110000111;
assign LUT_3[49358] = 32'b00000000000000000100000010001110;
assign LUT_3[49359] = 32'b00000000000000001010101101101011;
assign LUT_3[49360] = 32'b00000000000000000010100110110001;
assign LUT_3[49361] = 32'b00000000000000001001010010001110;
assign LUT_3[49362] = 32'b00000000000000000100101110010101;
assign LUT_3[49363] = 32'b00000000000000001011011001110010;
assign LUT_3[49364] = 32'b11111111111111111111110100100111;
assign LUT_3[49365] = 32'b00000000000000000110100000000100;
assign LUT_3[49366] = 32'b00000000000000000001111100001011;
assign LUT_3[49367] = 32'b00000000000000001000100111101000;
assign LUT_3[49368] = 32'b00000000000000000111111111110111;
assign LUT_3[49369] = 32'b00000000000000001110101011010100;
assign LUT_3[49370] = 32'b00000000000000001010000111011011;
assign LUT_3[49371] = 32'b00000000000000010000110010111000;
assign LUT_3[49372] = 32'b00000000000000000101001101101101;
assign LUT_3[49373] = 32'b00000000000000001011111001001010;
assign LUT_3[49374] = 32'b00000000000000000111010101010001;
assign LUT_3[49375] = 32'b00000000000000001110000000101110;
assign LUT_3[49376] = 32'b00000000000000000000100010001110;
assign LUT_3[49377] = 32'b00000000000000000111001101101011;
assign LUT_3[49378] = 32'b00000000000000000010101001110010;
assign LUT_3[49379] = 32'b00000000000000001001010101001111;
assign LUT_3[49380] = 32'b11111111111111111101110000000100;
assign LUT_3[49381] = 32'b00000000000000000100011011100001;
assign LUT_3[49382] = 32'b11111111111111111111110111101000;
assign LUT_3[49383] = 32'b00000000000000000110100011000101;
assign LUT_3[49384] = 32'b00000000000000000101111011010100;
assign LUT_3[49385] = 32'b00000000000000001100100110110001;
assign LUT_3[49386] = 32'b00000000000000001000000010111000;
assign LUT_3[49387] = 32'b00000000000000001110101110010101;
assign LUT_3[49388] = 32'b00000000000000000011001001001010;
assign LUT_3[49389] = 32'b00000000000000001001110100100111;
assign LUT_3[49390] = 32'b00000000000000000101010000101110;
assign LUT_3[49391] = 32'b00000000000000001011111100001011;
assign LUT_3[49392] = 32'b00000000000000000011110101010001;
assign LUT_3[49393] = 32'b00000000000000001010100000101110;
assign LUT_3[49394] = 32'b00000000000000000101111100110101;
assign LUT_3[49395] = 32'b00000000000000001100101000010010;
assign LUT_3[49396] = 32'b00000000000000000001000011000111;
assign LUT_3[49397] = 32'b00000000000000000111101110100100;
assign LUT_3[49398] = 32'b00000000000000000011001010101011;
assign LUT_3[49399] = 32'b00000000000000001001110110001000;
assign LUT_3[49400] = 32'b00000000000000001001001110010111;
assign LUT_3[49401] = 32'b00000000000000001111111001110100;
assign LUT_3[49402] = 32'b00000000000000001011010101111011;
assign LUT_3[49403] = 32'b00000000000000010010000001011000;
assign LUT_3[49404] = 32'b00000000000000000110011100001101;
assign LUT_3[49405] = 32'b00000000000000001101000111101010;
assign LUT_3[49406] = 32'b00000000000000001000100011110001;
assign LUT_3[49407] = 32'b00000000000000001111001111001110;
assign LUT_3[49408] = 32'b11111111111111111001011111100110;
assign LUT_3[49409] = 32'b00000000000000000000001011000011;
assign LUT_3[49410] = 32'b11111111111111111011100111001010;
assign LUT_3[49411] = 32'b00000000000000000010010010100111;
assign LUT_3[49412] = 32'b11111111111111110110101101011100;
assign LUT_3[49413] = 32'b11111111111111111101011000111001;
assign LUT_3[49414] = 32'b11111111111111111000110101000000;
assign LUT_3[49415] = 32'b11111111111111111111100000011101;
assign LUT_3[49416] = 32'b11111111111111111110111000101100;
assign LUT_3[49417] = 32'b00000000000000000101100100001001;
assign LUT_3[49418] = 32'b00000000000000000001000000010000;
assign LUT_3[49419] = 32'b00000000000000000111101011101101;
assign LUT_3[49420] = 32'b11111111111111111100000110100010;
assign LUT_3[49421] = 32'b00000000000000000010110001111111;
assign LUT_3[49422] = 32'b11111111111111111110001110000110;
assign LUT_3[49423] = 32'b00000000000000000100111001100011;
assign LUT_3[49424] = 32'b11111111111111111100110010101001;
assign LUT_3[49425] = 32'b00000000000000000011011110000110;
assign LUT_3[49426] = 32'b11111111111111111110111010001101;
assign LUT_3[49427] = 32'b00000000000000000101100101101010;
assign LUT_3[49428] = 32'b11111111111111111010000000011111;
assign LUT_3[49429] = 32'b00000000000000000000101011111100;
assign LUT_3[49430] = 32'b11111111111111111100001000000011;
assign LUT_3[49431] = 32'b00000000000000000010110011100000;
assign LUT_3[49432] = 32'b00000000000000000010001011101111;
assign LUT_3[49433] = 32'b00000000000000001000110111001100;
assign LUT_3[49434] = 32'b00000000000000000100010011010011;
assign LUT_3[49435] = 32'b00000000000000001010111110110000;
assign LUT_3[49436] = 32'b11111111111111111111011001100101;
assign LUT_3[49437] = 32'b00000000000000000110000101000010;
assign LUT_3[49438] = 32'b00000000000000000001100001001001;
assign LUT_3[49439] = 32'b00000000000000001000001100100110;
assign LUT_3[49440] = 32'b11111111111111111010101110000110;
assign LUT_3[49441] = 32'b00000000000000000001011001100011;
assign LUT_3[49442] = 32'b11111111111111111100110101101010;
assign LUT_3[49443] = 32'b00000000000000000011100001000111;
assign LUT_3[49444] = 32'b11111111111111110111111011111100;
assign LUT_3[49445] = 32'b11111111111111111110100111011001;
assign LUT_3[49446] = 32'b11111111111111111010000011100000;
assign LUT_3[49447] = 32'b00000000000000000000101110111101;
assign LUT_3[49448] = 32'b00000000000000000000000111001100;
assign LUT_3[49449] = 32'b00000000000000000110110010101001;
assign LUT_3[49450] = 32'b00000000000000000010001110110000;
assign LUT_3[49451] = 32'b00000000000000001000111010001101;
assign LUT_3[49452] = 32'b11111111111111111101010101000010;
assign LUT_3[49453] = 32'b00000000000000000100000000011111;
assign LUT_3[49454] = 32'b11111111111111111111011100100110;
assign LUT_3[49455] = 32'b00000000000000000110001000000011;
assign LUT_3[49456] = 32'b11111111111111111110000001001001;
assign LUT_3[49457] = 32'b00000000000000000100101100100110;
assign LUT_3[49458] = 32'b00000000000000000000001000101101;
assign LUT_3[49459] = 32'b00000000000000000110110100001010;
assign LUT_3[49460] = 32'b11111111111111111011001110111111;
assign LUT_3[49461] = 32'b00000000000000000001111010011100;
assign LUT_3[49462] = 32'b11111111111111111101010110100011;
assign LUT_3[49463] = 32'b00000000000000000100000010000000;
assign LUT_3[49464] = 32'b00000000000000000011011010001111;
assign LUT_3[49465] = 32'b00000000000000001010000101101100;
assign LUT_3[49466] = 32'b00000000000000000101100001110011;
assign LUT_3[49467] = 32'b00000000000000001100001101010000;
assign LUT_3[49468] = 32'b00000000000000000000101000000101;
assign LUT_3[49469] = 32'b00000000000000000111010011100010;
assign LUT_3[49470] = 32'b00000000000000000010101111101001;
assign LUT_3[49471] = 32'b00000000000000001001011011000110;
assign LUT_3[49472] = 32'b11111111111111111001011000010001;
assign LUT_3[49473] = 32'b00000000000000000000000011101110;
assign LUT_3[49474] = 32'b11111111111111111011011111110101;
assign LUT_3[49475] = 32'b00000000000000000010001011010010;
assign LUT_3[49476] = 32'b11111111111111110110100110000111;
assign LUT_3[49477] = 32'b11111111111111111101010001100100;
assign LUT_3[49478] = 32'b11111111111111111000101101101011;
assign LUT_3[49479] = 32'b11111111111111111111011001001000;
assign LUT_3[49480] = 32'b11111111111111111110110001010111;
assign LUT_3[49481] = 32'b00000000000000000101011100110100;
assign LUT_3[49482] = 32'b00000000000000000000111000111011;
assign LUT_3[49483] = 32'b00000000000000000111100100011000;
assign LUT_3[49484] = 32'b11111111111111111011111111001101;
assign LUT_3[49485] = 32'b00000000000000000010101010101010;
assign LUT_3[49486] = 32'b11111111111111111110000110110001;
assign LUT_3[49487] = 32'b00000000000000000100110010001110;
assign LUT_3[49488] = 32'b11111111111111111100101011010100;
assign LUT_3[49489] = 32'b00000000000000000011010110110001;
assign LUT_3[49490] = 32'b11111111111111111110110010111000;
assign LUT_3[49491] = 32'b00000000000000000101011110010101;
assign LUT_3[49492] = 32'b11111111111111111001111001001010;
assign LUT_3[49493] = 32'b00000000000000000000100100100111;
assign LUT_3[49494] = 32'b11111111111111111100000000101110;
assign LUT_3[49495] = 32'b00000000000000000010101100001011;
assign LUT_3[49496] = 32'b00000000000000000010000100011010;
assign LUT_3[49497] = 32'b00000000000000001000101111110111;
assign LUT_3[49498] = 32'b00000000000000000100001011111110;
assign LUT_3[49499] = 32'b00000000000000001010110111011011;
assign LUT_3[49500] = 32'b11111111111111111111010010010000;
assign LUT_3[49501] = 32'b00000000000000000101111101101101;
assign LUT_3[49502] = 32'b00000000000000000001011001110100;
assign LUT_3[49503] = 32'b00000000000000001000000101010001;
assign LUT_3[49504] = 32'b11111111111111111010100110110001;
assign LUT_3[49505] = 32'b00000000000000000001010010001110;
assign LUT_3[49506] = 32'b11111111111111111100101110010101;
assign LUT_3[49507] = 32'b00000000000000000011011001110010;
assign LUT_3[49508] = 32'b11111111111111110111110100100111;
assign LUT_3[49509] = 32'b11111111111111111110100000000100;
assign LUT_3[49510] = 32'b11111111111111111001111100001011;
assign LUT_3[49511] = 32'b00000000000000000000100111101000;
assign LUT_3[49512] = 32'b11111111111111111111111111110111;
assign LUT_3[49513] = 32'b00000000000000000110101011010100;
assign LUT_3[49514] = 32'b00000000000000000010000111011011;
assign LUT_3[49515] = 32'b00000000000000001000110010111000;
assign LUT_3[49516] = 32'b11111111111111111101001101101101;
assign LUT_3[49517] = 32'b00000000000000000011111001001010;
assign LUT_3[49518] = 32'b11111111111111111111010101010001;
assign LUT_3[49519] = 32'b00000000000000000110000000101110;
assign LUT_3[49520] = 32'b11111111111111111101111001110100;
assign LUT_3[49521] = 32'b00000000000000000100100101010001;
assign LUT_3[49522] = 32'b00000000000000000000000001011000;
assign LUT_3[49523] = 32'b00000000000000000110101100110101;
assign LUT_3[49524] = 32'b11111111111111111011000111101010;
assign LUT_3[49525] = 32'b00000000000000000001110011000111;
assign LUT_3[49526] = 32'b11111111111111111101001111001110;
assign LUT_3[49527] = 32'b00000000000000000011111010101011;
assign LUT_3[49528] = 32'b00000000000000000011010010111010;
assign LUT_3[49529] = 32'b00000000000000001001111110010111;
assign LUT_3[49530] = 32'b00000000000000000101011010011110;
assign LUT_3[49531] = 32'b00000000000000001100000101111011;
assign LUT_3[49532] = 32'b00000000000000000000100000110000;
assign LUT_3[49533] = 32'b00000000000000000111001100001101;
assign LUT_3[49534] = 32'b00000000000000000010101000010100;
assign LUT_3[49535] = 32'b00000000000000001001010011110001;
assign LUT_3[49536] = 32'b11111111111111111011101010100100;
assign LUT_3[49537] = 32'b00000000000000000010010110000001;
assign LUT_3[49538] = 32'b11111111111111111101110010001000;
assign LUT_3[49539] = 32'b00000000000000000100011101100101;
assign LUT_3[49540] = 32'b11111111111111111000111000011010;
assign LUT_3[49541] = 32'b11111111111111111111100011110111;
assign LUT_3[49542] = 32'b11111111111111111010111111111110;
assign LUT_3[49543] = 32'b00000000000000000001101011011011;
assign LUT_3[49544] = 32'b00000000000000000001000011101010;
assign LUT_3[49545] = 32'b00000000000000000111101111000111;
assign LUT_3[49546] = 32'b00000000000000000011001011001110;
assign LUT_3[49547] = 32'b00000000000000001001110110101011;
assign LUT_3[49548] = 32'b11111111111111111110010001100000;
assign LUT_3[49549] = 32'b00000000000000000100111100111101;
assign LUT_3[49550] = 32'b00000000000000000000011001000100;
assign LUT_3[49551] = 32'b00000000000000000111000100100001;
assign LUT_3[49552] = 32'b11111111111111111110111101100111;
assign LUT_3[49553] = 32'b00000000000000000101101001000100;
assign LUT_3[49554] = 32'b00000000000000000001000101001011;
assign LUT_3[49555] = 32'b00000000000000000111110000101000;
assign LUT_3[49556] = 32'b11111111111111111100001011011101;
assign LUT_3[49557] = 32'b00000000000000000010110110111010;
assign LUT_3[49558] = 32'b11111111111111111110010011000001;
assign LUT_3[49559] = 32'b00000000000000000100111110011110;
assign LUT_3[49560] = 32'b00000000000000000100010110101101;
assign LUT_3[49561] = 32'b00000000000000001011000010001010;
assign LUT_3[49562] = 32'b00000000000000000110011110010001;
assign LUT_3[49563] = 32'b00000000000000001101001001101110;
assign LUT_3[49564] = 32'b00000000000000000001100100100011;
assign LUT_3[49565] = 32'b00000000000000001000010000000000;
assign LUT_3[49566] = 32'b00000000000000000011101100000111;
assign LUT_3[49567] = 32'b00000000000000001010010111100100;
assign LUT_3[49568] = 32'b11111111111111111100111001000100;
assign LUT_3[49569] = 32'b00000000000000000011100100100001;
assign LUT_3[49570] = 32'b11111111111111111111000000101000;
assign LUT_3[49571] = 32'b00000000000000000101101100000101;
assign LUT_3[49572] = 32'b11111111111111111010000110111010;
assign LUT_3[49573] = 32'b00000000000000000000110010010111;
assign LUT_3[49574] = 32'b11111111111111111100001110011110;
assign LUT_3[49575] = 32'b00000000000000000010111001111011;
assign LUT_3[49576] = 32'b00000000000000000010010010001010;
assign LUT_3[49577] = 32'b00000000000000001000111101100111;
assign LUT_3[49578] = 32'b00000000000000000100011001101110;
assign LUT_3[49579] = 32'b00000000000000001011000101001011;
assign LUT_3[49580] = 32'b11111111111111111111100000000000;
assign LUT_3[49581] = 32'b00000000000000000110001011011101;
assign LUT_3[49582] = 32'b00000000000000000001100111100100;
assign LUT_3[49583] = 32'b00000000000000001000010011000001;
assign LUT_3[49584] = 32'b00000000000000000000001100000111;
assign LUT_3[49585] = 32'b00000000000000000110110111100100;
assign LUT_3[49586] = 32'b00000000000000000010010011101011;
assign LUT_3[49587] = 32'b00000000000000001000111111001000;
assign LUT_3[49588] = 32'b11111111111111111101011001111101;
assign LUT_3[49589] = 32'b00000000000000000100000101011010;
assign LUT_3[49590] = 32'b11111111111111111111100001100001;
assign LUT_3[49591] = 32'b00000000000000000110001100111110;
assign LUT_3[49592] = 32'b00000000000000000101100101001101;
assign LUT_3[49593] = 32'b00000000000000001100010000101010;
assign LUT_3[49594] = 32'b00000000000000000111101100110001;
assign LUT_3[49595] = 32'b00000000000000001110011000001110;
assign LUT_3[49596] = 32'b00000000000000000010110011000011;
assign LUT_3[49597] = 32'b00000000000000001001011110100000;
assign LUT_3[49598] = 32'b00000000000000000100111010100111;
assign LUT_3[49599] = 32'b00000000000000001011100110000100;
assign LUT_3[49600] = 32'b11111111111111111011100011001111;
assign LUT_3[49601] = 32'b00000000000000000010001110101100;
assign LUT_3[49602] = 32'b11111111111111111101101010110011;
assign LUT_3[49603] = 32'b00000000000000000100010110010000;
assign LUT_3[49604] = 32'b11111111111111111000110001000101;
assign LUT_3[49605] = 32'b11111111111111111111011100100010;
assign LUT_3[49606] = 32'b11111111111111111010111000101001;
assign LUT_3[49607] = 32'b00000000000000000001100100000110;
assign LUT_3[49608] = 32'b00000000000000000000111100010101;
assign LUT_3[49609] = 32'b00000000000000000111100111110010;
assign LUT_3[49610] = 32'b00000000000000000011000011111001;
assign LUT_3[49611] = 32'b00000000000000001001101111010110;
assign LUT_3[49612] = 32'b11111111111111111110001010001011;
assign LUT_3[49613] = 32'b00000000000000000100110101101000;
assign LUT_3[49614] = 32'b00000000000000000000010001101111;
assign LUT_3[49615] = 32'b00000000000000000110111101001100;
assign LUT_3[49616] = 32'b11111111111111111110110110010010;
assign LUT_3[49617] = 32'b00000000000000000101100001101111;
assign LUT_3[49618] = 32'b00000000000000000000111101110110;
assign LUT_3[49619] = 32'b00000000000000000111101001010011;
assign LUT_3[49620] = 32'b11111111111111111100000100001000;
assign LUT_3[49621] = 32'b00000000000000000010101111100101;
assign LUT_3[49622] = 32'b11111111111111111110001011101100;
assign LUT_3[49623] = 32'b00000000000000000100110111001001;
assign LUT_3[49624] = 32'b00000000000000000100001111011000;
assign LUT_3[49625] = 32'b00000000000000001010111010110101;
assign LUT_3[49626] = 32'b00000000000000000110010110111100;
assign LUT_3[49627] = 32'b00000000000000001101000010011001;
assign LUT_3[49628] = 32'b00000000000000000001011101001110;
assign LUT_3[49629] = 32'b00000000000000001000001000101011;
assign LUT_3[49630] = 32'b00000000000000000011100100110010;
assign LUT_3[49631] = 32'b00000000000000001010010000001111;
assign LUT_3[49632] = 32'b11111111111111111100110001101111;
assign LUT_3[49633] = 32'b00000000000000000011011101001100;
assign LUT_3[49634] = 32'b11111111111111111110111001010011;
assign LUT_3[49635] = 32'b00000000000000000101100100110000;
assign LUT_3[49636] = 32'b11111111111111111001111111100101;
assign LUT_3[49637] = 32'b00000000000000000000101011000010;
assign LUT_3[49638] = 32'b11111111111111111100000111001001;
assign LUT_3[49639] = 32'b00000000000000000010110010100110;
assign LUT_3[49640] = 32'b00000000000000000010001010110101;
assign LUT_3[49641] = 32'b00000000000000001000110110010010;
assign LUT_3[49642] = 32'b00000000000000000100010010011001;
assign LUT_3[49643] = 32'b00000000000000001010111101110110;
assign LUT_3[49644] = 32'b11111111111111111111011000101011;
assign LUT_3[49645] = 32'b00000000000000000110000100001000;
assign LUT_3[49646] = 32'b00000000000000000001100000001111;
assign LUT_3[49647] = 32'b00000000000000001000001011101100;
assign LUT_3[49648] = 32'b00000000000000000000000100110010;
assign LUT_3[49649] = 32'b00000000000000000110110000001111;
assign LUT_3[49650] = 32'b00000000000000000010001100010110;
assign LUT_3[49651] = 32'b00000000000000001000110111110011;
assign LUT_3[49652] = 32'b11111111111111111101010010101000;
assign LUT_3[49653] = 32'b00000000000000000011111110000101;
assign LUT_3[49654] = 32'b11111111111111111111011010001100;
assign LUT_3[49655] = 32'b00000000000000000110000101101001;
assign LUT_3[49656] = 32'b00000000000000000101011101111000;
assign LUT_3[49657] = 32'b00000000000000001100001001010101;
assign LUT_3[49658] = 32'b00000000000000000111100101011100;
assign LUT_3[49659] = 32'b00000000000000001110010000111001;
assign LUT_3[49660] = 32'b00000000000000000010101011101110;
assign LUT_3[49661] = 32'b00000000000000001001010111001011;
assign LUT_3[49662] = 32'b00000000000000000100110011010010;
assign LUT_3[49663] = 32'b00000000000000001011011110101111;
assign LUT_3[49664] = 32'b00000000000000000000100101010001;
assign LUT_3[49665] = 32'b00000000000000000111010000101110;
assign LUT_3[49666] = 32'b00000000000000000010101100110101;
assign LUT_3[49667] = 32'b00000000000000001001011000010010;
assign LUT_3[49668] = 32'b11111111111111111101110011000111;
assign LUT_3[49669] = 32'b00000000000000000100011110100100;
assign LUT_3[49670] = 32'b11111111111111111111111010101011;
assign LUT_3[49671] = 32'b00000000000000000110100110001000;
assign LUT_3[49672] = 32'b00000000000000000101111110010111;
assign LUT_3[49673] = 32'b00000000000000001100101001110100;
assign LUT_3[49674] = 32'b00000000000000001000000101111011;
assign LUT_3[49675] = 32'b00000000000000001110110001011000;
assign LUT_3[49676] = 32'b00000000000000000011001100001101;
assign LUT_3[49677] = 32'b00000000000000001001110111101010;
assign LUT_3[49678] = 32'b00000000000000000101010011110001;
assign LUT_3[49679] = 32'b00000000000000001011111111001110;
assign LUT_3[49680] = 32'b00000000000000000011111000010100;
assign LUT_3[49681] = 32'b00000000000000001010100011110001;
assign LUT_3[49682] = 32'b00000000000000000101111111111000;
assign LUT_3[49683] = 32'b00000000000000001100101011010101;
assign LUT_3[49684] = 32'b00000000000000000001000110001010;
assign LUT_3[49685] = 32'b00000000000000000111110001100111;
assign LUT_3[49686] = 32'b00000000000000000011001101101110;
assign LUT_3[49687] = 32'b00000000000000001001111001001011;
assign LUT_3[49688] = 32'b00000000000000001001010001011010;
assign LUT_3[49689] = 32'b00000000000000001111111100110111;
assign LUT_3[49690] = 32'b00000000000000001011011000111110;
assign LUT_3[49691] = 32'b00000000000000010010000100011011;
assign LUT_3[49692] = 32'b00000000000000000110011111010000;
assign LUT_3[49693] = 32'b00000000000000001101001010101101;
assign LUT_3[49694] = 32'b00000000000000001000100110110100;
assign LUT_3[49695] = 32'b00000000000000001111010010010001;
assign LUT_3[49696] = 32'b00000000000000000001110011110001;
assign LUT_3[49697] = 32'b00000000000000001000011111001110;
assign LUT_3[49698] = 32'b00000000000000000011111011010101;
assign LUT_3[49699] = 32'b00000000000000001010100110110010;
assign LUT_3[49700] = 32'b11111111111111111111000001100111;
assign LUT_3[49701] = 32'b00000000000000000101101101000100;
assign LUT_3[49702] = 32'b00000000000000000001001001001011;
assign LUT_3[49703] = 32'b00000000000000000111110100101000;
assign LUT_3[49704] = 32'b00000000000000000111001100110111;
assign LUT_3[49705] = 32'b00000000000000001101111000010100;
assign LUT_3[49706] = 32'b00000000000000001001010100011011;
assign LUT_3[49707] = 32'b00000000000000001111111111111000;
assign LUT_3[49708] = 32'b00000000000000000100011010101101;
assign LUT_3[49709] = 32'b00000000000000001011000110001010;
assign LUT_3[49710] = 32'b00000000000000000110100010010001;
assign LUT_3[49711] = 32'b00000000000000001101001101101110;
assign LUT_3[49712] = 32'b00000000000000000101000110110100;
assign LUT_3[49713] = 32'b00000000000000001011110010010001;
assign LUT_3[49714] = 32'b00000000000000000111001110011000;
assign LUT_3[49715] = 32'b00000000000000001101111001110101;
assign LUT_3[49716] = 32'b00000000000000000010010100101010;
assign LUT_3[49717] = 32'b00000000000000001001000000000111;
assign LUT_3[49718] = 32'b00000000000000000100011100001110;
assign LUT_3[49719] = 32'b00000000000000001011000111101011;
assign LUT_3[49720] = 32'b00000000000000001010011111111010;
assign LUT_3[49721] = 32'b00000000000000010001001011010111;
assign LUT_3[49722] = 32'b00000000000000001100100111011110;
assign LUT_3[49723] = 32'b00000000000000010011010010111011;
assign LUT_3[49724] = 32'b00000000000000000111101101110000;
assign LUT_3[49725] = 32'b00000000000000001110011001001101;
assign LUT_3[49726] = 32'b00000000000000001001110101010100;
assign LUT_3[49727] = 32'b00000000000000010000100000110001;
assign LUT_3[49728] = 32'b00000000000000000000011101111100;
assign LUT_3[49729] = 32'b00000000000000000111001001011001;
assign LUT_3[49730] = 32'b00000000000000000010100101100000;
assign LUT_3[49731] = 32'b00000000000000001001010000111101;
assign LUT_3[49732] = 32'b11111111111111111101101011110010;
assign LUT_3[49733] = 32'b00000000000000000100010111001111;
assign LUT_3[49734] = 32'b11111111111111111111110011010110;
assign LUT_3[49735] = 32'b00000000000000000110011110110011;
assign LUT_3[49736] = 32'b00000000000000000101110111000010;
assign LUT_3[49737] = 32'b00000000000000001100100010011111;
assign LUT_3[49738] = 32'b00000000000000000111111110100110;
assign LUT_3[49739] = 32'b00000000000000001110101010000011;
assign LUT_3[49740] = 32'b00000000000000000011000100111000;
assign LUT_3[49741] = 32'b00000000000000001001110000010101;
assign LUT_3[49742] = 32'b00000000000000000101001100011100;
assign LUT_3[49743] = 32'b00000000000000001011110111111001;
assign LUT_3[49744] = 32'b00000000000000000011110000111111;
assign LUT_3[49745] = 32'b00000000000000001010011100011100;
assign LUT_3[49746] = 32'b00000000000000000101111000100011;
assign LUT_3[49747] = 32'b00000000000000001100100100000000;
assign LUT_3[49748] = 32'b00000000000000000000111110110101;
assign LUT_3[49749] = 32'b00000000000000000111101010010010;
assign LUT_3[49750] = 32'b00000000000000000011000110011001;
assign LUT_3[49751] = 32'b00000000000000001001110001110110;
assign LUT_3[49752] = 32'b00000000000000001001001010000101;
assign LUT_3[49753] = 32'b00000000000000001111110101100010;
assign LUT_3[49754] = 32'b00000000000000001011010001101001;
assign LUT_3[49755] = 32'b00000000000000010001111101000110;
assign LUT_3[49756] = 32'b00000000000000000110010111111011;
assign LUT_3[49757] = 32'b00000000000000001101000011011000;
assign LUT_3[49758] = 32'b00000000000000001000011111011111;
assign LUT_3[49759] = 32'b00000000000000001111001010111100;
assign LUT_3[49760] = 32'b00000000000000000001101100011100;
assign LUT_3[49761] = 32'b00000000000000001000010111111001;
assign LUT_3[49762] = 32'b00000000000000000011110100000000;
assign LUT_3[49763] = 32'b00000000000000001010011111011101;
assign LUT_3[49764] = 32'b11111111111111111110111010010010;
assign LUT_3[49765] = 32'b00000000000000000101100101101111;
assign LUT_3[49766] = 32'b00000000000000000001000001110110;
assign LUT_3[49767] = 32'b00000000000000000111101101010011;
assign LUT_3[49768] = 32'b00000000000000000111000101100010;
assign LUT_3[49769] = 32'b00000000000000001101110000111111;
assign LUT_3[49770] = 32'b00000000000000001001001101000110;
assign LUT_3[49771] = 32'b00000000000000001111111000100011;
assign LUT_3[49772] = 32'b00000000000000000100010011011000;
assign LUT_3[49773] = 32'b00000000000000001010111110110101;
assign LUT_3[49774] = 32'b00000000000000000110011010111100;
assign LUT_3[49775] = 32'b00000000000000001101000110011001;
assign LUT_3[49776] = 32'b00000000000000000100111111011111;
assign LUT_3[49777] = 32'b00000000000000001011101010111100;
assign LUT_3[49778] = 32'b00000000000000000111000111000011;
assign LUT_3[49779] = 32'b00000000000000001101110010100000;
assign LUT_3[49780] = 32'b00000000000000000010001101010101;
assign LUT_3[49781] = 32'b00000000000000001000111000110010;
assign LUT_3[49782] = 32'b00000000000000000100010100111001;
assign LUT_3[49783] = 32'b00000000000000001011000000010110;
assign LUT_3[49784] = 32'b00000000000000001010011000100101;
assign LUT_3[49785] = 32'b00000000000000010001000100000010;
assign LUT_3[49786] = 32'b00000000000000001100100000001001;
assign LUT_3[49787] = 32'b00000000000000010011001011100110;
assign LUT_3[49788] = 32'b00000000000000000111100110011011;
assign LUT_3[49789] = 32'b00000000000000001110010001111000;
assign LUT_3[49790] = 32'b00000000000000001001101101111111;
assign LUT_3[49791] = 32'b00000000000000010000011001011100;
assign LUT_3[49792] = 32'b00000000000000000010110000001111;
assign LUT_3[49793] = 32'b00000000000000001001011011101100;
assign LUT_3[49794] = 32'b00000000000000000100110111110011;
assign LUT_3[49795] = 32'b00000000000000001011100011010000;
assign LUT_3[49796] = 32'b11111111111111111111111110000101;
assign LUT_3[49797] = 32'b00000000000000000110101001100010;
assign LUT_3[49798] = 32'b00000000000000000010000101101001;
assign LUT_3[49799] = 32'b00000000000000001000110001000110;
assign LUT_3[49800] = 32'b00000000000000001000001001010101;
assign LUT_3[49801] = 32'b00000000000000001110110100110010;
assign LUT_3[49802] = 32'b00000000000000001010010000111001;
assign LUT_3[49803] = 32'b00000000000000010000111100010110;
assign LUT_3[49804] = 32'b00000000000000000101010111001011;
assign LUT_3[49805] = 32'b00000000000000001100000010101000;
assign LUT_3[49806] = 32'b00000000000000000111011110101111;
assign LUT_3[49807] = 32'b00000000000000001110001010001100;
assign LUT_3[49808] = 32'b00000000000000000110000011010010;
assign LUT_3[49809] = 32'b00000000000000001100101110101111;
assign LUT_3[49810] = 32'b00000000000000001000001010110110;
assign LUT_3[49811] = 32'b00000000000000001110110110010011;
assign LUT_3[49812] = 32'b00000000000000000011010001001000;
assign LUT_3[49813] = 32'b00000000000000001001111100100101;
assign LUT_3[49814] = 32'b00000000000000000101011000101100;
assign LUT_3[49815] = 32'b00000000000000001100000100001001;
assign LUT_3[49816] = 32'b00000000000000001011011100011000;
assign LUT_3[49817] = 32'b00000000000000010010000111110101;
assign LUT_3[49818] = 32'b00000000000000001101100011111100;
assign LUT_3[49819] = 32'b00000000000000010100001111011001;
assign LUT_3[49820] = 32'b00000000000000001000101010001110;
assign LUT_3[49821] = 32'b00000000000000001111010101101011;
assign LUT_3[49822] = 32'b00000000000000001010110001110010;
assign LUT_3[49823] = 32'b00000000000000010001011101001111;
assign LUT_3[49824] = 32'b00000000000000000011111110101111;
assign LUT_3[49825] = 32'b00000000000000001010101010001100;
assign LUT_3[49826] = 32'b00000000000000000110000110010011;
assign LUT_3[49827] = 32'b00000000000000001100110001110000;
assign LUT_3[49828] = 32'b00000000000000000001001100100101;
assign LUT_3[49829] = 32'b00000000000000000111111000000010;
assign LUT_3[49830] = 32'b00000000000000000011010100001001;
assign LUT_3[49831] = 32'b00000000000000001001111111100110;
assign LUT_3[49832] = 32'b00000000000000001001010111110101;
assign LUT_3[49833] = 32'b00000000000000010000000011010010;
assign LUT_3[49834] = 32'b00000000000000001011011111011001;
assign LUT_3[49835] = 32'b00000000000000010010001010110110;
assign LUT_3[49836] = 32'b00000000000000000110100101101011;
assign LUT_3[49837] = 32'b00000000000000001101010001001000;
assign LUT_3[49838] = 32'b00000000000000001000101101001111;
assign LUT_3[49839] = 32'b00000000000000001111011000101100;
assign LUT_3[49840] = 32'b00000000000000000111010001110010;
assign LUT_3[49841] = 32'b00000000000000001101111101001111;
assign LUT_3[49842] = 32'b00000000000000001001011001010110;
assign LUT_3[49843] = 32'b00000000000000010000000100110011;
assign LUT_3[49844] = 32'b00000000000000000100011111101000;
assign LUT_3[49845] = 32'b00000000000000001011001011000101;
assign LUT_3[49846] = 32'b00000000000000000110100111001100;
assign LUT_3[49847] = 32'b00000000000000001101010010101001;
assign LUT_3[49848] = 32'b00000000000000001100101010111000;
assign LUT_3[49849] = 32'b00000000000000010011010110010101;
assign LUT_3[49850] = 32'b00000000000000001110110010011100;
assign LUT_3[49851] = 32'b00000000000000010101011101111001;
assign LUT_3[49852] = 32'b00000000000000001001111000101110;
assign LUT_3[49853] = 32'b00000000000000010000100100001011;
assign LUT_3[49854] = 32'b00000000000000001100000000010010;
assign LUT_3[49855] = 32'b00000000000000010010101011101111;
assign LUT_3[49856] = 32'b00000000000000000010101000111010;
assign LUT_3[49857] = 32'b00000000000000001001010100010111;
assign LUT_3[49858] = 32'b00000000000000000100110000011110;
assign LUT_3[49859] = 32'b00000000000000001011011011111011;
assign LUT_3[49860] = 32'b11111111111111111111110110110000;
assign LUT_3[49861] = 32'b00000000000000000110100010001101;
assign LUT_3[49862] = 32'b00000000000000000001111110010100;
assign LUT_3[49863] = 32'b00000000000000001000101001110001;
assign LUT_3[49864] = 32'b00000000000000001000000010000000;
assign LUT_3[49865] = 32'b00000000000000001110101101011101;
assign LUT_3[49866] = 32'b00000000000000001010001001100100;
assign LUT_3[49867] = 32'b00000000000000010000110101000001;
assign LUT_3[49868] = 32'b00000000000000000101001111110110;
assign LUT_3[49869] = 32'b00000000000000001011111011010011;
assign LUT_3[49870] = 32'b00000000000000000111010111011010;
assign LUT_3[49871] = 32'b00000000000000001110000010110111;
assign LUT_3[49872] = 32'b00000000000000000101111011111101;
assign LUT_3[49873] = 32'b00000000000000001100100111011010;
assign LUT_3[49874] = 32'b00000000000000001000000011100001;
assign LUT_3[49875] = 32'b00000000000000001110101110111110;
assign LUT_3[49876] = 32'b00000000000000000011001001110011;
assign LUT_3[49877] = 32'b00000000000000001001110101010000;
assign LUT_3[49878] = 32'b00000000000000000101010001010111;
assign LUT_3[49879] = 32'b00000000000000001011111100110100;
assign LUT_3[49880] = 32'b00000000000000001011010101000011;
assign LUT_3[49881] = 32'b00000000000000010010000000100000;
assign LUT_3[49882] = 32'b00000000000000001101011100100111;
assign LUT_3[49883] = 32'b00000000000000010100001000000100;
assign LUT_3[49884] = 32'b00000000000000001000100010111001;
assign LUT_3[49885] = 32'b00000000000000001111001110010110;
assign LUT_3[49886] = 32'b00000000000000001010101010011101;
assign LUT_3[49887] = 32'b00000000000000010001010101111010;
assign LUT_3[49888] = 32'b00000000000000000011110111011010;
assign LUT_3[49889] = 32'b00000000000000001010100010110111;
assign LUT_3[49890] = 32'b00000000000000000101111110111110;
assign LUT_3[49891] = 32'b00000000000000001100101010011011;
assign LUT_3[49892] = 32'b00000000000000000001000101010000;
assign LUT_3[49893] = 32'b00000000000000000111110000101101;
assign LUT_3[49894] = 32'b00000000000000000011001100110100;
assign LUT_3[49895] = 32'b00000000000000001001111000010001;
assign LUT_3[49896] = 32'b00000000000000001001010000100000;
assign LUT_3[49897] = 32'b00000000000000001111111011111101;
assign LUT_3[49898] = 32'b00000000000000001011011000000100;
assign LUT_3[49899] = 32'b00000000000000010010000011100001;
assign LUT_3[49900] = 32'b00000000000000000110011110010110;
assign LUT_3[49901] = 32'b00000000000000001101001001110011;
assign LUT_3[49902] = 32'b00000000000000001000100101111010;
assign LUT_3[49903] = 32'b00000000000000001111010001010111;
assign LUT_3[49904] = 32'b00000000000000000111001010011101;
assign LUT_3[49905] = 32'b00000000000000001101110101111010;
assign LUT_3[49906] = 32'b00000000000000001001010010000001;
assign LUT_3[49907] = 32'b00000000000000001111111101011110;
assign LUT_3[49908] = 32'b00000000000000000100011000010011;
assign LUT_3[49909] = 32'b00000000000000001011000011110000;
assign LUT_3[49910] = 32'b00000000000000000110011111110111;
assign LUT_3[49911] = 32'b00000000000000001101001011010100;
assign LUT_3[49912] = 32'b00000000000000001100100011100011;
assign LUT_3[49913] = 32'b00000000000000010011001111000000;
assign LUT_3[49914] = 32'b00000000000000001110101011000111;
assign LUT_3[49915] = 32'b00000000000000010101010110100100;
assign LUT_3[49916] = 32'b00000000000000001001110001011001;
assign LUT_3[49917] = 32'b00000000000000010000011100110110;
assign LUT_3[49918] = 32'b00000000000000001011111000111101;
assign LUT_3[49919] = 32'b00000000000000010010100100011010;
assign LUT_3[49920] = 32'b11111111111111111100110100110010;
assign LUT_3[49921] = 32'b00000000000000000011100000001111;
assign LUT_3[49922] = 32'b11111111111111111110111100010110;
assign LUT_3[49923] = 32'b00000000000000000101100111110011;
assign LUT_3[49924] = 32'b11111111111111111010000010101000;
assign LUT_3[49925] = 32'b00000000000000000000101110000101;
assign LUT_3[49926] = 32'b11111111111111111100001010001100;
assign LUT_3[49927] = 32'b00000000000000000010110101101001;
assign LUT_3[49928] = 32'b00000000000000000010001101111000;
assign LUT_3[49929] = 32'b00000000000000001000111001010101;
assign LUT_3[49930] = 32'b00000000000000000100010101011100;
assign LUT_3[49931] = 32'b00000000000000001011000000111001;
assign LUT_3[49932] = 32'b11111111111111111111011011101110;
assign LUT_3[49933] = 32'b00000000000000000110000111001011;
assign LUT_3[49934] = 32'b00000000000000000001100011010010;
assign LUT_3[49935] = 32'b00000000000000001000001110101111;
assign LUT_3[49936] = 32'b00000000000000000000000111110101;
assign LUT_3[49937] = 32'b00000000000000000110110011010010;
assign LUT_3[49938] = 32'b00000000000000000010001111011001;
assign LUT_3[49939] = 32'b00000000000000001000111010110110;
assign LUT_3[49940] = 32'b11111111111111111101010101101011;
assign LUT_3[49941] = 32'b00000000000000000100000001001000;
assign LUT_3[49942] = 32'b11111111111111111111011101001111;
assign LUT_3[49943] = 32'b00000000000000000110001000101100;
assign LUT_3[49944] = 32'b00000000000000000101100000111011;
assign LUT_3[49945] = 32'b00000000000000001100001100011000;
assign LUT_3[49946] = 32'b00000000000000000111101000011111;
assign LUT_3[49947] = 32'b00000000000000001110010011111100;
assign LUT_3[49948] = 32'b00000000000000000010101110110001;
assign LUT_3[49949] = 32'b00000000000000001001011010001110;
assign LUT_3[49950] = 32'b00000000000000000100110110010101;
assign LUT_3[49951] = 32'b00000000000000001011100001110010;
assign LUT_3[49952] = 32'b11111111111111111110000011010010;
assign LUT_3[49953] = 32'b00000000000000000100101110101111;
assign LUT_3[49954] = 32'b00000000000000000000001010110110;
assign LUT_3[49955] = 32'b00000000000000000110110110010011;
assign LUT_3[49956] = 32'b11111111111111111011010001001000;
assign LUT_3[49957] = 32'b00000000000000000001111100100101;
assign LUT_3[49958] = 32'b11111111111111111101011000101100;
assign LUT_3[49959] = 32'b00000000000000000100000100001001;
assign LUT_3[49960] = 32'b00000000000000000011011100011000;
assign LUT_3[49961] = 32'b00000000000000001010000111110101;
assign LUT_3[49962] = 32'b00000000000000000101100011111100;
assign LUT_3[49963] = 32'b00000000000000001100001111011001;
assign LUT_3[49964] = 32'b00000000000000000000101010001110;
assign LUT_3[49965] = 32'b00000000000000000111010101101011;
assign LUT_3[49966] = 32'b00000000000000000010110001110010;
assign LUT_3[49967] = 32'b00000000000000001001011101001111;
assign LUT_3[49968] = 32'b00000000000000000001010110010101;
assign LUT_3[49969] = 32'b00000000000000001000000001110010;
assign LUT_3[49970] = 32'b00000000000000000011011101111001;
assign LUT_3[49971] = 32'b00000000000000001010001001010110;
assign LUT_3[49972] = 32'b11111111111111111110100100001011;
assign LUT_3[49973] = 32'b00000000000000000101001111101000;
assign LUT_3[49974] = 32'b00000000000000000000101011101111;
assign LUT_3[49975] = 32'b00000000000000000111010111001100;
assign LUT_3[49976] = 32'b00000000000000000110101111011011;
assign LUT_3[49977] = 32'b00000000000000001101011010111000;
assign LUT_3[49978] = 32'b00000000000000001000110110111111;
assign LUT_3[49979] = 32'b00000000000000001111100010011100;
assign LUT_3[49980] = 32'b00000000000000000011111101010001;
assign LUT_3[49981] = 32'b00000000000000001010101000101110;
assign LUT_3[49982] = 32'b00000000000000000110000100110101;
assign LUT_3[49983] = 32'b00000000000000001100110000010010;
assign LUT_3[49984] = 32'b11111111111111111100101101011101;
assign LUT_3[49985] = 32'b00000000000000000011011000111010;
assign LUT_3[49986] = 32'b11111111111111111110110101000001;
assign LUT_3[49987] = 32'b00000000000000000101100000011110;
assign LUT_3[49988] = 32'b11111111111111111001111011010011;
assign LUT_3[49989] = 32'b00000000000000000000100110110000;
assign LUT_3[49990] = 32'b11111111111111111100000010110111;
assign LUT_3[49991] = 32'b00000000000000000010101110010100;
assign LUT_3[49992] = 32'b00000000000000000010000110100011;
assign LUT_3[49993] = 32'b00000000000000001000110010000000;
assign LUT_3[49994] = 32'b00000000000000000100001110000111;
assign LUT_3[49995] = 32'b00000000000000001010111001100100;
assign LUT_3[49996] = 32'b11111111111111111111010100011001;
assign LUT_3[49997] = 32'b00000000000000000101111111110110;
assign LUT_3[49998] = 32'b00000000000000000001011011111101;
assign LUT_3[49999] = 32'b00000000000000001000000111011010;
assign LUT_3[50000] = 32'b00000000000000000000000000100000;
assign LUT_3[50001] = 32'b00000000000000000110101011111101;
assign LUT_3[50002] = 32'b00000000000000000010001000000100;
assign LUT_3[50003] = 32'b00000000000000001000110011100001;
assign LUT_3[50004] = 32'b11111111111111111101001110010110;
assign LUT_3[50005] = 32'b00000000000000000011111001110011;
assign LUT_3[50006] = 32'b11111111111111111111010101111010;
assign LUT_3[50007] = 32'b00000000000000000110000001010111;
assign LUT_3[50008] = 32'b00000000000000000101011001100110;
assign LUT_3[50009] = 32'b00000000000000001100000101000011;
assign LUT_3[50010] = 32'b00000000000000000111100001001010;
assign LUT_3[50011] = 32'b00000000000000001110001100100111;
assign LUT_3[50012] = 32'b00000000000000000010100111011100;
assign LUT_3[50013] = 32'b00000000000000001001010010111001;
assign LUT_3[50014] = 32'b00000000000000000100101111000000;
assign LUT_3[50015] = 32'b00000000000000001011011010011101;
assign LUT_3[50016] = 32'b11111111111111111101111011111101;
assign LUT_3[50017] = 32'b00000000000000000100100111011010;
assign LUT_3[50018] = 32'b00000000000000000000000011100001;
assign LUT_3[50019] = 32'b00000000000000000110101110111110;
assign LUT_3[50020] = 32'b11111111111111111011001001110011;
assign LUT_3[50021] = 32'b00000000000000000001110101010000;
assign LUT_3[50022] = 32'b11111111111111111101010001010111;
assign LUT_3[50023] = 32'b00000000000000000011111100110100;
assign LUT_3[50024] = 32'b00000000000000000011010101000011;
assign LUT_3[50025] = 32'b00000000000000001010000000100000;
assign LUT_3[50026] = 32'b00000000000000000101011100100111;
assign LUT_3[50027] = 32'b00000000000000001100001000000100;
assign LUT_3[50028] = 32'b00000000000000000000100010111001;
assign LUT_3[50029] = 32'b00000000000000000111001110010110;
assign LUT_3[50030] = 32'b00000000000000000010101010011101;
assign LUT_3[50031] = 32'b00000000000000001001010101111010;
assign LUT_3[50032] = 32'b00000000000000000001001111000000;
assign LUT_3[50033] = 32'b00000000000000000111111010011101;
assign LUT_3[50034] = 32'b00000000000000000011010110100100;
assign LUT_3[50035] = 32'b00000000000000001010000010000001;
assign LUT_3[50036] = 32'b11111111111111111110011100110110;
assign LUT_3[50037] = 32'b00000000000000000101001000010011;
assign LUT_3[50038] = 32'b00000000000000000000100100011010;
assign LUT_3[50039] = 32'b00000000000000000111001111110111;
assign LUT_3[50040] = 32'b00000000000000000110101000000110;
assign LUT_3[50041] = 32'b00000000000000001101010011100011;
assign LUT_3[50042] = 32'b00000000000000001000101111101010;
assign LUT_3[50043] = 32'b00000000000000001111011011000111;
assign LUT_3[50044] = 32'b00000000000000000011110101111100;
assign LUT_3[50045] = 32'b00000000000000001010100001011001;
assign LUT_3[50046] = 32'b00000000000000000101111101100000;
assign LUT_3[50047] = 32'b00000000000000001100101000111101;
assign LUT_3[50048] = 32'b11111111111111111110111111110000;
assign LUT_3[50049] = 32'b00000000000000000101101011001101;
assign LUT_3[50050] = 32'b00000000000000000001000111010100;
assign LUT_3[50051] = 32'b00000000000000000111110010110001;
assign LUT_3[50052] = 32'b11111111111111111100001101100110;
assign LUT_3[50053] = 32'b00000000000000000010111001000011;
assign LUT_3[50054] = 32'b11111111111111111110010101001010;
assign LUT_3[50055] = 32'b00000000000000000101000000100111;
assign LUT_3[50056] = 32'b00000000000000000100011000110110;
assign LUT_3[50057] = 32'b00000000000000001011000100010011;
assign LUT_3[50058] = 32'b00000000000000000110100000011010;
assign LUT_3[50059] = 32'b00000000000000001101001011110111;
assign LUT_3[50060] = 32'b00000000000000000001100110101100;
assign LUT_3[50061] = 32'b00000000000000001000010010001001;
assign LUT_3[50062] = 32'b00000000000000000011101110010000;
assign LUT_3[50063] = 32'b00000000000000001010011001101101;
assign LUT_3[50064] = 32'b00000000000000000010010010110011;
assign LUT_3[50065] = 32'b00000000000000001000111110010000;
assign LUT_3[50066] = 32'b00000000000000000100011010010111;
assign LUT_3[50067] = 32'b00000000000000001011000101110100;
assign LUT_3[50068] = 32'b11111111111111111111100000101001;
assign LUT_3[50069] = 32'b00000000000000000110001100000110;
assign LUT_3[50070] = 32'b00000000000000000001101000001101;
assign LUT_3[50071] = 32'b00000000000000001000010011101010;
assign LUT_3[50072] = 32'b00000000000000000111101011111001;
assign LUT_3[50073] = 32'b00000000000000001110010111010110;
assign LUT_3[50074] = 32'b00000000000000001001110011011101;
assign LUT_3[50075] = 32'b00000000000000010000011110111010;
assign LUT_3[50076] = 32'b00000000000000000100111001101111;
assign LUT_3[50077] = 32'b00000000000000001011100101001100;
assign LUT_3[50078] = 32'b00000000000000000111000001010011;
assign LUT_3[50079] = 32'b00000000000000001101101100110000;
assign LUT_3[50080] = 32'b00000000000000000000001110010000;
assign LUT_3[50081] = 32'b00000000000000000110111001101101;
assign LUT_3[50082] = 32'b00000000000000000010010101110100;
assign LUT_3[50083] = 32'b00000000000000001001000001010001;
assign LUT_3[50084] = 32'b11111111111111111101011100000110;
assign LUT_3[50085] = 32'b00000000000000000100000111100011;
assign LUT_3[50086] = 32'b11111111111111111111100011101010;
assign LUT_3[50087] = 32'b00000000000000000110001111000111;
assign LUT_3[50088] = 32'b00000000000000000101100111010110;
assign LUT_3[50089] = 32'b00000000000000001100010010110011;
assign LUT_3[50090] = 32'b00000000000000000111101110111010;
assign LUT_3[50091] = 32'b00000000000000001110011010010111;
assign LUT_3[50092] = 32'b00000000000000000010110101001100;
assign LUT_3[50093] = 32'b00000000000000001001100000101001;
assign LUT_3[50094] = 32'b00000000000000000100111100110000;
assign LUT_3[50095] = 32'b00000000000000001011101000001101;
assign LUT_3[50096] = 32'b00000000000000000011100001010011;
assign LUT_3[50097] = 32'b00000000000000001010001100110000;
assign LUT_3[50098] = 32'b00000000000000000101101000110111;
assign LUT_3[50099] = 32'b00000000000000001100010100010100;
assign LUT_3[50100] = 32'b00000000000000000000101111001001;
assign LUT_3[50101] = 32'b00000000000000000111011010100110;
assign LUT_3[50102] = 32'b00000000000000000010110110101101;
assign LUT_3[50103] = 32'b00000000000000001001100010001010;
assign LUT_3[50104] = 32'b00000000000000001000111010011001;
assign LUT_3[50105] = 32'b00000000000000001111100101110110;
assign LUT_3[50106] = 32'b00000000000000001011000001111101;
assign LUT_3[50107] = 32'b00000000000000010001101101011010;
assign LUT_3[50108] = 32'b00000000000000000110001000001111;
assign LUT_3[50109] = 32'b00000000000000001100110011101100;
assign LUT_3[50110] = 32'b00000000000000001000001111110011;
assign LUT_3[50111] = 32'b00000000000000001110111011010000;
assign LUT_3[50112] = 32'b11111111111111111110111000011011;
assign LUT_3[50113] = 32'b00000000000000000101100011111000;
assign LUT_3[50114] = 32'b00000000000000000000111111111111;
assign LUT_3[50115] = 32'b00000000000000000111101011011100;
assign LUT_3[50116] = 32'b11111111111111111100000110010001;
assign LUT_3[50117] = 32'b00000000000000000010110001101110;
assign LUT_3[50118] = 32'b11111111111111111110001101110101;
assign LUT_3[50119] = 32'b00000000000000000100111001010010;
assign LUT_3[50120] = 32'b00000000000000000100010001100001;
assign LUT_3[50121] = 32'b00000000000000001010111100111110;
assign LUT_3[50122] = 32'b00000000000000000110011001000101;
assign LUT_3[50123] = 32'b00000000000000001101000100100010;
assign LUT_3[50124] = 32'b00000000000000000001011111010111;
assign LUT_3[50125] = 32'b00000000000000001000001010110100;
assign LUT_3[50126] = 32'b00000000000000000011100110111011;
assign LUT_3[50127] = 32'b00000000000000001010010010011000;
assign LUT_3[50128] = 32'b00000000000000000010001011011110;
assign LUT_3[50129] = 32'b00000000000000001000110110111011;
assign LUT_3[50130] = 32'b00000000000000000100010011000010;
assign LUT_3[50131] = 32'b00000000000000001010111110011111;
assign LUT_3[50132] = 32'b11111111111111111111011001010100;
assign LUT_3[50133] = 32'b00000000000000000110000100110001;
assign LUT_3[50134] = 32'b00000000000000000001100000111000;
assign LUT_3[50135] = 32'b00000000000000001000001100010101;
assign LUT_3[50136] = 32'b00000000000000000111100100100100;
assign LUT_3[50137] = 32'b00000000000000001110010000000001;
assign LUT_3[50138] = 32'b00000000000000001001101100001000;
assign LUT_3[50139] = 32'b00000000000000010000010111100101;
assign LUT_3[50140] = 32'b00000000000000000100110010011010;
assign LUT_3[50141] = 32'b00000000000000001011011101110111;
assign LUT_3[50142] = 32'b00000000000000000110111001111110;
assign LUT_3[50143] = 32'b00000000000000001101100101011011;
assign LUT_3[50144] = 32'b00000000000000000000000110111011;
assign LUT_3[50145] = 32'b00000000000000000110110010011000;
assign LUT_3[50146] = 32'b00000000000000000010001110011111;
assign LUT_3[50147] = 32'b00000000000000001000111001111100;
assign LUT_3[50148] = 32'b11111111111111111101010100110001;
assign LUT_3[50149] = 32'b00000000000000000100000000001110;
assign LUT_3[50150] = 32'b11111111111111111111011100010101;
assign LUT_3[50151] = 32'b00000000000000000110000111110010;
assign LUT_3[50152] = 32'b00000000000000000101100000000001;
assign LUT_3[50153] = 32'b00000000000000001100001011011110;
assign LUT_3[50154] = 32'b00000000000000000111100111100101;
assign LUT_3[50155] = 32'b00000000000000001110010011000010;
assign LUT_3[50156] = 32'b00000000000000000010101101110111;
assign LUT_3[50157] = 32'b00000000000000001001011001010100;
assign LUT_3[50158] = 32'b00000000000000000100110101011011;
assign LUT_3[50159] = 32'b00000000000000001011100000111000;
assign LUT_3[50160] = 32'b00000000000000000011011001111110;
assign LUT_3[50161] = 32'b00000000000000001010000101011011;
assign LUT_3[50162] = 32'b00000000000000000101100001100010;
assign LUT_3[50163] = 32'b00000000000000001100001100111111;
assign LUT_3[50164] = 32'b00000000000000000000100111110100;
assign LUT_3[50165] = 32'b00000000000000000111010011010001;
assign LUT_3[50166] = 32'b00000000000000000010101111011000;
assign LUT_3[50167] = 32'b00000000000000001001011010110101;
assign LUT_3[50168] = 32'b00000000000000001000110011000100;
assign LUT_3[50169] = 32'b00000000000000001111011110100001;
assign LUT_3[50170] = 32'b00000000000000001010111010101000;
assign LUT_3[50171] = 32'b00000000000000010001100110000101;
assign LUT_3[50172] = 32'b00000000000000000110000000111010;
assign LUT_3[50173] = 32'b00000000000000001100101100010111;
assign LUT_3[50174] = 32'b00000000000000001000001000011110;
assign LUT_3[50175] = 32'b00000000000000001110110011111011;
assign LUT_3[50176] = 32'b00000000000000000011110101000010;
assign LUT_3[50177] = 32'b00000000000000001010100000011111;
assign LUT_3[50178] = 32'b00000000000000000101111100100110;
assign LUT_3[50179] = 32'b00000000000000001100101000000011;
assign LUT_3[50180] = 32'b00000000000000000001000010111000;
assign LUT_3[50181] = 32'b00000000000000000111101110010101;
assign LUT_3[50182] = 32'b00000000000000000011001010011100;
assign LUT_3[50183] = 32'b00000000000000001001110101111001;
assign LUT_3[50184] = 32'b00000000000000001001001110001000;
assign LUT_3[50185] = 32'b00000000000000001111111001100101;
assign LUT_3[50186] = 32'b00000000000000001011010101101100;
assign LUT_3[50187] = 32'b00000000000000010010000001001001;
assign LUT_3[50188] = 32'b00000000000000000110011011111110;
assign LUT_3[50189] = 32'b00000000000000001101000111011011;
assign LUT_3[50190] = 32'b00000000000000001000100011100010;
assign LUT_3[50191] = 32'b00000000000000001111001110111111;
assign LUT_3[50192] = 32'b00000000000000000111001000000101;
assign LUT_3[50193] = 32'b00000000000000001101110011100010;
assign LUT_3[50194] = 32'b00000000000000001001001111101001;
assign LUT_3[50195] = 32'b00000000000000001111111011000110;
assign LUT_3[50196] = 32'b00000000000000000100010101111011;
assign LUT_3[50197] = 32'b00000000000000001011000001011000;
assign LUT_3[50198] = 32'b00000000000000000110011101011111;
assign LUT_3[50199] = 32'b00000000000000001101001000111100;
assign LUT_3[50200] = 32'b00000000000000001100100001001011;
assign LUT_3[50201] = 32'b00000000000000010011001100101000;
assign LUT_3[50202] = 32'b00000000000000001110101000101111;
assign LUT_3[50203] = 32'b00000000000000010101010100001100;
assign LUT_3[50204] = 32'b00000000000000001001101111000001;
assign LUT_3[50205] = 32'b00000000000000010000011010011110;
assign LUT_3[50206] = 32'b00000000000000001011110110100101;
assign LUT_3[50207] = 32'b00000000000000010010100010000010;
assign LUT_3[50208] = 32'b00000000000000000101000011100010;
assign LUT_3[50209] = 32'b00000000000000001011101110111111;
assign LUT_3[50210] = 32'b00000000000000000111001011000110;
assign LUT_3[50211] = 32'b00000000000000001101110110100011;
assign LUT_3[50212] = 32'b00000000000000000010010001011000;
assign LUT_3[50213] = 32'b00000000000000001000111100110101;
assign LUT_3[50214] = 32'b00000000000000000100011000111100;
assign LUT_3[50215] = 32'b00000000000000001011000100011001;
assign LUT_3[50216] = 32'b00000000000000001010011100101000;
assign LUT_3[50217] = 32'b00000000000000010001001000000101;
assign LUT_3[50218] = 32'b00000000000000001100100100001100;
assign LUT_3[50219] = 32'b00000000000000010011001111101001;
assign LUT_3[50220] = 32'b00000000000000000111101010011110;
assign LUT_3[50221] = 32'b00000000000000001110010101111011;
assign LUT_3[50222] = 32'b00000000000000001001110010000010;
assign LUT_3[50223] = 32'b00000000000000010000011101011111;
assign LUT_3[50224] = 32'b00000000000000001000010110100101;
assign LUT_3[50225] = 32'b00000000000000001111000010000010;
assign LUT_3[50226] = 32'b00000000000000001010011110001001;
assign LUT_3[50227] = 32'b00000000000000010001001001100110;
assign LUT_3[50228] = 32'b00000000000000000101100100011011;
assign LUT_3[50229] = 32'b00000000000000001100001111111000;
assign LUT_3[50230] = 32'b00000000000000000111101011111111;
assign LUT_3[50231] = 32'b00000000000000001110010111011100;
assign LUT_3[50232] = 32'b00000000000000001101101111101011;
assign LUT_3[50233] = 32'b00000000000000010100011011001000;
assign LUT_3[50234] = 32'b00000000000000001111110111001111;
assign LUT_3[50235] = 32'b00000000000000010110100010101100;
assign LUT_3[50236] = 32'b00000000000000001010111101100001;
assign LUT_3[50237] = 32'b00000000000000010001101000111110;
assign LUT_3[50238] = 32'b00000000000000001101000101000101;
assign LUT_3[50239] = 32'b00000000000000010011110000100010;
assign LUT_3[50240] = 32'b00000000000000000011101101101101;
assign LUT_3[50241] = 32'b00000000000000001010011001001010;
assign LUT_3[50242] = 32'b00000000000000000101110101010001;
assign LUT_3[50243] = 32'b00000000000000001100100000101110;
assign LUT_3[50244] = 32'b00000000000000000000111011100011;
assign LUT_3[50245] = 32'b00000000000000000111100111000000;
assign LUT_3[50246] = 32'b00000000000000000011000011000111;
assign LUT_3[50247] = 32'b00000000000000001001101110100100;
assign LUT_3[50248] = 32'b00000000000000001001000110110011;
assign LUT_3[50249] = 32'b00000000000000001111110010010000;
assign LUT_3[50250] = 32'b00000000000000001011001110010111;
assign LUT_3[50251] = 32'b00000000000000010001111001110100;
assign LUT_3[50252] = 32'b00000000000000000110010100101001;
assign LUT_3[50253] = 32'b00000000000000001101000000000110;
assign LUT_3[50254] = 32'b00000000000000001000011100001101;
assign LUT_3[50255] = 32'b00000000000000001111000111101010;
assign LUT_3[50256] = 32'b00000000000000000111000000110000;
assign LUT_3[50257] = 32'b00000000000000001101101100001101;
assign LUT_3[50258] = 32'b00000000000000001001001000010100;
assign LUT_3[50259] = 32'b00000000000000001111110011110001;
assign LUT_3[50260] = 32'b00000000000000000100001110100110;
assign LUT_3[50261] = 32'b00000000000000001010111010000011;
assign LUT_3[50262] = 32'b00000000000000000110010110001010;
assign LUT_3[50263] = 32'b00000000000000001101000001100111;
assign LUT_3[50264] = 32'b00000000000000001100011001110110;
assign LUT_3[50265] = 32'b00000000000000010011000101010011;
assign LUT_3[50266] = 32'b00000000000000001110100001011010;
assign LUT_3[50267] = 32'b00000000000000010101001100110111;
assign LUT_3[50268] = 32'b00000000000000001001100111101100;
assign LUT_3[50269] = 32'b00000000000000010000010011001001;
assign LUT_3[50270] = 32'b00000000000000001011101111010000;
assign LUT_3[50271] = 32'b00000000000000010010011010101101;
assign LUT_3[50272] = 32'b00000000000000000100111100001101;
assign LUT_3[50273] = 32'b00000000000000001011100111101010;
assign LUT_3[50274] = 32'b00000000000000000111000011110001;
assign LUT_3[50275] = 32'b00000000000000001101101111001110;
assign LUT_3[50276] = 32'b00000000000000000010001010000011;
assign LUT_3[50277] = 32'b00000000000000001000110101100000;
assign LUT_3[50278] = 32'b00000000000000000100010001100111;
assign LUT_3[50279] = 32'b00000000000000001010111101000100;
assign LUT_3[50280] = 32'b00000000000000001010010101010011;
assign LUT_3[50281] = 32'b00000000000000010001000000110000;
assign LUT_3[50282] = 32'b00000000000000001100011100110111;
assign LUT_3[50283] = 32'b00000000000000010011001000010100;
assign LUT_3[50284] = 32'b00000000000000000111100011001001;
assign LUT_3[50285] = 32'b00000000000000001110001110100110;
assign LUT_3[50286] = 32'b00000000000000001001101010101101;
assign LUT_3[50287] = 32'b00000000000000010000010110001010;
assign LUT_3[50288] = 32'b00000000000000001000001111010000;
assign LUT_3[50289] = 32'b00000000000000001110111010101101;
assign LUT_3[50290] = 32'b00000000000000001010010110110100;
assign LUT_3[50291] = 32'b00000000000000010001000010010001;
assign LUT_3[50292] = 32'b00000000000000000101011101000110;
assign LUT_3[50293] = 32'b00000000000000001100001000100011;
assign LUT_3[50294] = 32'b00000000000000000111100100101010;
assign LUT_3[50295] = 32'b00000000000000001110010000000111;
assign LUT_3[50296] = 32'b00000000000000001101101000010110;
assign LUT_3[50297] = 32'b00000000000000010100010011110011;
assign LUT_3[50298] = 32'b00000000000000001111101111111010;
assign LUT_3[50299] = 32'b00000000000000010110011011010111;
assign LUT_3[50300] = 32'b00000000000000001010110110001100;
assign LUT_3[50301] = 32'b00000000000000010001100001101001;
assign LUT_3[50302] = 32'b00000000000000001100111101110000;
assign LUT_3[50303] = 32'b00000000000000010011101001001101;
assign LUT_3[50304] = 32'b00000000000000000110000000000000;
assign LUT_3[50305] = 32'b00000000000000001100101011011101;
assign LUT_3[50306] = 32'b00000000000000001000000111100100;
assign LUT_3[50307] = 32'b00000000000000001110110011000001;
assign LUT_3[50308] = 32'b00000000000000000011001101110110;
assign LUT_3[50309] = 32'b00000000000000001001111001010011;
assign LUT_3[50310] = 32'b00000000000000000101010101011010;
assign LUT_3[50311] = 32'b00000000000000001100000000110111;
assign LUT_3[50312] = 32'b00000000000000001011011001000110;
assign LUT_3[50313] = 32'b00000000000000010010000100100011;
assign LUT_3[50314] = 32'b00000000000000001101100000101010;
assign LUT_3[50315] = 32'b00000000000000010100001100000111;
assign LUT_3[50316] = 32'b00000000000000001000100110111100;
assign LUT_3[50317] = 32'b00000000000000001111010010011001;
assign LUT_3[50318] = 32'b00000000000000001010101110100000;
assign LUT_3[50319] = 32'b00000000000000010001011001111101;
assign LUT_3[50320] = 32'b00000000000000001001010011000011;
assign LUT_3[50321] = 32'b00000000000000001111111110100000;
assign LUT_3[50322] = 32'b00000000000000001011011010100111;
assign LUT_3[50323] = 32'b00000000000000010010000110000100;
assign LUT_3[50324] = 32'b00000000000000000110100000111001;
assign LUT_3[50325] = 32'b00000000000000001101001100010110;
assign LUT_3[50326] = 32'b00000000000000001000101000011101;
assign LUT_3[50327] = 32'b00000000000000001111010011111010;
assign LUT_3[50328] = 32'b00000000000000001110101100001001;
assign LUT_3[50329] = 32'b00000000000000010101010111100110;
assign LUT_3[50330] = 32'b00000000000000010000110011101101;
assign LUT_3[50331] = 32'b00000000000000010111011111001010;
assign LUT_3[50332] = 32'b00000000000000001011111001111111;
assign LUT_3[50333] = 32'b00000000000000010010100101011100;
assign LUT_3[50334] = 32'b00000000000000001110000001100011;
assign LUT_3[50335] = 32'b00000000000000010100101101000000;
assign LUT_3[50336] = 32'b00000000000000000111001110100000;
assign LUT_3[50337] = 32'b00000000000000001101111001111101;
assign LUT_3[50338] = 32'b00000000000000001001010110000100;
assign LUT_3[50339] = 32'b00000000000000010000000001100001;
assign LUT_3[50340] = 32'b00000000000000000100011100010110;
assign LUT_3[50341] = 32'b00000000000000001011000111110011;
assign LUT_3[50342] = 32'b00000000000000000110100011111010;
assign LUT_3[50343] = 32'b00000000000000001101001111010111;
assign LUT_3[50344] = 32'b00000000000000001100100111100110;
assign LUT_3[50345] = 32'b00000000000000010011010011000011;
assign LUT_3[50346] = 32'b00000000000000001110101111001010;
assign LUT_3[50347] = 32'b00000000000000010101011010100111;
assign LUT_3[50348] = 32'b00000000000000001001110101011100;
assign LUT_3[50349] = 32'b00000000000000010000100000111001;
assign LUT_3[50350] = 32'b00000000000000001011111101000000;
assign LUT_3[50351] = 32'b00000000000000010010101000011101;
assign LUT_3[50352] = 32'b00000000000000001010100001100011;
assign LUT_3[50353] = 32'b00000000000000010001001101000000;
assign LUT_3[50354] = 32'b00000000000000001100101001000111;
assign LUT_3[50355] = 32'b00000000000000010011010100100100;
assign LUT_3[50356] = 32'b00000000000000000111101111011001;
assign LUT_3[50357] = 32'b00000000000000001110011010110110;
assign LUT_3[50358] = 32'b00000000000000001001110110111101;
assign LUT_3[50359] = 32'b00000000000000010000100010011010;
assign LUT_3[50360] = 32'b00000000000000001111111010101001;
assign LUT_3[50361] = 32'b00000000000000010110100110000110;
assign LUT_3[50362] = 32'b00000000000000010010000010001101;
assign LUT_3[50363] = 32'b00000000000000011000101101101010;
assign LUT_3[50364] = 32'b00000000000000001101001000011111;
assign LUT_3[50365] = 32'b00000000000000010011110011111100;
assign LUT_3[50366] = 32'b00000000000000001111010000000011;
assign LUT_3[50367] = 32'b00000000000000010101111011100000;
assign LUT_3[50368] = 32'b00000000000000000101111000101011;
assign LUT_3[50369] = 32'b00000000000000001100100100001000;
assign LUT_3[50370] = 32'b00000000000000001000000000001111;
assign LUT_3[50371] = 32'b00000000000000001110101011101100;
assign LUT_3[50372] = 32'b00000000000000000011000110100001;
assign LUT_3[50373] = 32'b00000000000000001001110001111110;
assign LUT_3[50374] = 32'b00000000000000000101001110000101;
assign LUT_3[50375] = 32'b00000000000000001011111001100010;
assign LUT_3[50376] = 32'b00000000000000001011010001110001;
assign LUT_3[50377] = 32'b00000000000000010001111101001110;
assign LUT_3[50378] = 32'b00000000000000001101011001010101;
assign LUT_3[50379] = 32'b00000000000000010100000100110010;
assign LUT_3[50380] = 32'b00000000000000001000011111100111;
assign LUT_3[50381] = 32'b00000000000000001111001011000100;
assign LUT_3[50382] = 32'b00000000000000001010100111001011;
assign LUT_3[50383] = 32'b00000000000000010001010010101000;
assign LUT_3[50384] = 32'b00000000000000001001001011101110;
assign LUT_3[50385] = 32'b00000000000000001111110111001011;
assign LUT_3[50386] = 32'b00000000000000001011010011010010;
assign LUT_3[50387] = 32'b00000000000000010001111110101111;
assign LUT_3[50388] = 32'b00000000000000000110011001100100;
assign LUT_3[50389] = 32'b00000000000000001101000101000001;
assign LUT_3[50390] = 32'b00000000000000001000100001001000;
assign LUT_3[50391] = 32'b00000000000000001111001100100101;
assign LUT_3[50392] = 32'b00000000000000001110100100110100;
assign LUT_3[50393] = 32'b00000000000000010101010000010001;
assign LUT_3[50394] = 32'b00000000000000010000101100011000;
assign LUT_3[50395] = 32'b00000000000000010111010111110101;
assign LUT_3[50396] = 32'b00000000000000001011110010101010;
assign LUT_3[50397] = 32'b00000000000000010010011110000111;
assign LUT_3[50398] = 32'b00000000000000001101111010001110;
assign LUT_3[50399] = 32'b00000000000000010100100101101011;
assign LUT_3[50400] = 32'b00000000000000000111000111001011;
assign LUT_3[50401] = 32'b00000000000000001101110010101000;
assign LUT_3[50402] = 32'b00000000000000001001001110101111;
assign LUT_3[50403] = 32'b00000000000000001111111010001100;
assign LUT_3[50404] = 32'b00000000000000000100010101000001;
assign LUT_3[50405] = 32'b00000000000000001011000000011110;
assign LUT_3[50406] = 32'b00000000000000000110011100100101;
assign LUT_3[50407] = 32'b00000000000000001101001000000010;
assign LUT_3[50408] = 32'b00000000000000001100100000010001;
assign LUT_3[50409] = 32'b00000000000000010011001011101110;
assign LUT_3[50410] = 32'b00000000000000001110100111110101;
assign LUT_3[50411] = 32'b00000000000000010101010011010010;
assign LUT_3[50412] = 32'b00000000000000001001101110000111;
assign LUT_3[50413] = 32'b00000000000000010000011001100100;
assign LUT_3[50414] = 32'b00000000000000001011110101101011;
assign LUT_3[50415] = 32'b00000000000000010010100001001000;
assign LUT_3[50416] = 32'b00000000000000001010011010001110;
assign LUT_3[50417] = 32'b00000000000000010001000101101011;
assign LUT_3[50418] = 32'b00000000000000001100100001110010;
assign LUT_3[50419] = 32'b00000000000000010011001101001111;
assign LUT_3[50420] = 32'b00000000000000000111101000000100;
assign LUT_3[50421] = 32'b00000000000000001110010011100001;
assign LUT_3[50422] = 32'b00000000000000001001101111101000;
assign LUT_3[50423] = 32'b00000000000000010000011011000101;
assign LUT_3[50424] = 32'b00000000000000001111110011010100;
assign LUT_3[50425] = 32'b00000000000000010110011110110001;
assign LUT_3[50426] = 32'b00000000000000010001111010111000;
assign LUT_3[50427] = 32'b00000000000000011000100110010101;
assign LUT_3[50428] = 32'b00000000000000001101000001001010;
assign LUT_3[50429] = 32'b00000000000000010011101100100111;
assign LUT_3[50430] = 32'b00000000000000001111001000101110;
assign LUT_3[50431] = 32'b00000000000000010101110100001011;
assign LUT_3[50432] = 32'b00000000000000000000000100100011;
assign LUT_3[50433] = 32'b00000000000000000110110000000000;
assign LUT_3[50434] = 32'b00000000000000000010001100000111;
assign LUT_3[50435] = 32'b00000000000000001000110111100100;
assign LUT_3[50436] = 32'b11111111111111111101010010011001;
assign LUT_3[50437] = 32'b00000000000000000011111101110110;
assign LUT_3[50438] = 32'b11111111111111111111011001111101;
assign LUT_3[50439] = 32'b00000000000000000110000101011010;
assign LUT_3[50440] = 32'b00000000000000000101011101101001;
assign LUT_3[50441] = 32'b00000000000000001100001001000110;
assign LUT_3[50442] = 32'b00000000000000000111100101001101;
assign LUT_3[50443] = 32'b00000000000000001110010000101010;
assign LUT_3[50444] = 32'b00000000000000000010101011011111;
assign LUT_3[50445] = 32'b00000000000000001001010110111100;
assign LUT_3[50446] = 32'b00000000000000000100110011000011;
assign LUT_3[50447] = 32'b00000000000000001011011110100000;
assign LUT_3[50448] = 32'b00000000000000000011010111100110;
assign LUT_3[50449] = 32'b00000000000000001010000011000011;
assign LUT_3[50450] = 32'b00000000000000000101011111001010;
assign LUT_3[50451] = 32'b00000000000000001100001010100111;
assign LUT_3[50452] = 32'b00000000000000000000100101011100;
assign LUT_3[50453] = 32'b00000000000000000111010000111001;
assign LUT_3[50454] = 32'b00000000000000000010101101000000;
assign LUT_3[50455] = 32'b00000000000000001001011000011101;
assign LUT_3[50456] = 32'b00000000000000001000110000101100;
assign LUT_3[50457] = 32'b00000000000000001111011100001001;
assign LUT_3[50458] = 32'b00000000000000001010111000010000;
assign LUT_3[50459] = 32'b00000000000000010001100011101101;
assign LUT_3[50460] = 32'b00000000000000000101111110100010;
assign LUT_3[50461] = 32'b00000000000000001100101001111111;
assign LUT_3[50462] = 32'b00000000000000001000000110000110;
assign LUT_3[50463] = 32'b00000000000000001110110001100011;
assign LUT_3[50464] = 32'b00000000000000000001010011000011;
assign LUT_3[50465] = 32'b00000000000000000111111110100000;
assign LUT_3[50466] = 32'b00000000000000000011011010100111;
assign LUT_3[50467] = 32'b00000000000000001010000110000100;
assign LUT_3[50468] = 32'b11111111111111111110100000111001;
assign LUT_3[50469] = 32'b00000000000000000101001100010110;
assign LUT_3[50470] = 32'b00000000000000000000101000011101;
assign LUT_3[50471] = 32'b00000000000000000111010011111010;
assign LUT_3[50472] = 32'b00000000000000000110101100001001;
assign LUT_3[50473] = 32'b00000000000000001101010111100110;
assign LUT_3[50474] = 32'b00000000000000001000110011101101;
assign LUT_3[50475] = 32'b00000000000000001111011111001010;
assign LUT_3[50476] = 32'b00000000000000000011111001111111;
assign LUT_3[50477] = 32'b00000000000000001010100101011100;
assign LUT_3[50478] = 32'b00000000000000000110000001100011;
assign LUT_3[50479] = 32'b00000000000000001100101101000000;
assign LUT_3[50480] = 32'b00000000000000000100100110000110;
assign LUT_3[50481] = 32'b00000000000000001011010001100011;
assign LUT_3[50482] = 32'b00000000000000000110101101101010;
assign LUT_3[50483] = 32'b00000000000000001101011001000111;
assign LUT_3[50484] = 32'b00000000000000000001110011111100;
assign LUT_3[50485] = 32'b00000000000000001000011111011001;
assign LUT_3[50486] = 32'b00000000000000000011111011100000;
assign LUT_3[50487] = 32'b00000000000000001010100110111101;
assign LUT_3[50488] = 32'b00000000000000001001111111001100;
assign LUT_3[50489] = 32'b00000000000000010000101010101001;
assign LUT_3[50490] = 32'b00000000000000001100000110110000;
assign LUT_3[50491] = 32'b00000000000000010010110010001101;
assign LUT_3[50492] = 32'b00000000000000000111001101000010;
assign LUT_3[50493] = 32'b00000000000000001101111000011111;
assign LUT_3[50494] = 32'b00000000000000001001010100100110;
assign LUT_3[50495] = 32'b00000000000000010000000000000011;
assign LUT_3[50496] = 32'b11111111111111111111111101001110;
assign LUT_3[50497] = 32'b00000000000000000110101000101011;
assign LUT_3[50498] = 32'b00000000000000000010000100110010;
assign LUT_3[50499] = 32'b00000000000000001000110000001111;
assign LUT_3[50500] = 32'b11111111111111111101001011000100;
assign LUT_3[50501] = 32'b00000000000000000011110110100001;
assign LUT_3[50502] = 32'b11111111111111111111010010101000;
assign LUT_3[50503] = 32'b00000000000000000101111110000101;
assign LUT_3[50504] = 32'b00000000000000000101010110010100;
assign LUT_3[50505] = 32'b00000000000000001100000001110001;
assign LUT_3[50506] = 32'b00000000000000000111011101111000;
assign LUT_3[50507] = 32'b00000000000000001110001001010101;
assign LUT_3[50508] = 32'b00000000000000000010100100001010;
assign LUT_3[50509] = 32'b00000000000000001001001111100111;
assign LUT_3[50510] = 32'b00000000000000000100101011101110;
assign LUT_3[50511] = 32'b00000000000000001011010111001011;
assign LUT_3[50512] = 32'b00000000000000000011010000010001;
assign LUT_3[50513] = 32'b00000000000000001001111011101110;
assign LUT_3[50514] = 32'b00000000000000000101010111110101;
assign LUT_3[50515] = 32'b00000000000000001100000011010010;
assign LUT_3[50516] = 32'b00000000000000000000011110000111;
assign LUT_3[50517] = 32'b00000000000000000111001001100100;
assign LUT_3[50518] = 32'b00000000000000000010100101101011;
assign LUT_3[50519] = 32'b00000000000000001001010001001000;
assign LUT_3[50520] = 32'b00000000000000001000101001010111;
assign LUT_3[50521] = 32'b00000000000000001111010100110100;
assign LUT_3[50522] = 32'b00000000000000001010110000111011;
assign LUT_3[50523] = 32'b00000000000000010001011100011000;
assign LUT_3[50524] = 32'b00000000000000000101110111001101;
assign LUT_3[50525] = 32'b00000000000000001100100010101010;
assign LUT_3[50526] = 32'b00000000000000000111111110110001;
assign LUT_3[50527] = 32'b00000000000000001110101010001110;
assign LUT_3[50528] = 32'b00000000000000000001001011101110;
assign LUT_3[50529] = 32'b00000000000000000111110111001011;
assign LUT_3[50530] = 32'b00000000000000000011010011010010;
assign LUT_3[50531] = 32'b00000000000000001001111110101111;
assign LUT_3[50532] = 32'b11111111111111111110011001100100;
assign LUT_3[50533] = 32'b00000000000000000101000101000001;
assign LUT_3[50534] = 32'b00000000000000000000100001001000;
assign LUT_3[50535] = 32'b00000000000000000111001100100101;
assign LUT_3[50536] = 32'b00000000000000000110100100110100;
assign LUT_3[50537] = 32'b00000000000000001101010000010001;
assign LUT_3[50538] = 32'b00000000000000001000101100011000;
assign LUT_3[50539] = 32'b00000000000000001111010111110101;
assign LUT_3[50540] = 32'b00000000000000000011110010101010;
assign LUT_3[50541] = 32'b00000000000000001010011110000111;
assign LUT_3[50542] = 32'b00000000000000000101111010001110;
assign LUT_3[50543] = 32'b00000000000000001100100101101011;
assign LUT_3[50544] = 32'b00000000000000000100011110110001;
assign LUT_3[50545] = 32'b00000000000000001011001010001110;
assign LUT_3[50546] = 32'b00000000000000000110100110010101;
assign LUT_3[50547] = 32'b00000000000000001101010001110010;
assign LUT_3[50548] = 32'b00000000000000000001101100100111;
assign LUT_3[50549] = 32'b00000000000000001000011000000100;
assign LUT_3[50550] = 32'b00000000000000000011110100001011;
assign LUT_3[50551] = 32'b00000000000000001010011111101000;
assign LUT_3[50552] = 32'b00000000000000001001110111110111;
assign LUT_3[50553] = 32'b00000000000000010000100011010100;
assign LUT_3[50554] = 32'b00000000000000001011111111011011;
assign LUT_3[50555] = 32'b00000000000000010010101010111000;
assign LUT_3[50556] = 32'b00000000000000000111000101101101;
assign LUT_3[50557] = 32'b00000000000000001101110001001010;
assign LUT_3[50558] = 32'b00000000000000001001001101010001;
assign LUT_3[50559] = 32'b00000000000000001111111000101110;
assign LUT_3[50560] = 32'b00000000000000000010001111100001;
assign LUT_3[50561] = 32'b00000000000000001000111010111110;
assign LUT_3[50562] = 32'b00000000000000000100010111000101;
assign LUT_3[50563] = 32'b00000000000000001011000010100010;
assign LUT_3[50564] = 32'b11111111111111111111011101010111;
assign LUT_3[50565] = 32'b00000000000000000110001000110100;
assign LUT_3[50566] = 32'b00000000000000000001100100111011;
assign LUT_3[50567] = 32'b00000000000000001000010000011000;
assign LUT_3[50568] = 32'b00000000000000000111101000100111;
assign LUT_3[50569] = 32'b00000000000000001110010100000100;
assign LUT_3[50570] = 32'b00000000000000001001110000001011;
assign LUT_3[50571] = 32'b00000000000000010000011011101000;
assign LUT_3[50572] = 32'b00000000000000000100110110011101;
assign LUT_3[50573] = 32'b00000000000000001011100001111010;
assign LUT_3[50574] = 32'b00000000000000000110111110000001;
assign LUT_3[50575] = 32'b00000000000000001101101001011110;
assign LUT_3[50576] = 32'b00000000000000000101100010100100;
assign LUT_3[50577] = 32'b00000000000000001100001110000001;
assign LUT_3[50578] = 32'b00000000000000000111101010001000;
assign LUT_3[50579] = 32'b00000000000000001110010101100101;
assign LUT_3[50580] = 32'b00000000000000000010110000011010;
assign LUT_3[50581] = 32'b00000000000000001001011011110111;
assign LUT_3[50582] = 32'b00000000000000000100110111111110;
assign LUT_3[50583] = 32'b00000000000000001011100011011011;
assign LUT_3[50584] = 32'b00000000000000001010111011101010;
assign LUT_3[50585] = 32'b00000000000000010001100111000111;
assign LUT_3[50586] = 32'b00000000000000001101000011001110;
assign LUT_3[50587] = 32'b00000000000000010011101110101011;
assign LUT_3[50588] = 32'b00000000000000001000001001100000;
assign LUT_3[50589] = 32'b00000000000000001110110100111101;
assign LUT_3[50590] = 32'b00000000000000001010010001000100;
assign LUT_3[50591] = 32'b00000000000000010000111100100001;
assign LUT_3[50592] = 32'b00000000000000000011011110000001;
assign LUT_3[50593] = 32'b00000000000000001010001001011110;
assign LUT_3[50594] = 32'b00000000000000000101100101100101;
assign LUT_3[50595] = 32'b00000000000000001100010001000010;
assign LUT_3[50596] = 32'b00000000000000000000101011110111;
assign LUT_3[50597] = 32'b00000000000000000111010111010100;
assign LUT_3[50598] = 32'b00000000000000000010110011011011;
assign LUT_3[50599] = 32'b00000000000000001001011110111000;
assign LUT_3[50600] = 32'b00000000000000001000110111000111;
assign LUT_3[50601] = 32'b00000000000000001111100010100100;
assign LUT_3[50602] = 32'b00000000000000001010111110101011;
assign LUT_3[50603] = 32'b00000000000000010001101010001000;
assign LUT_3[50604] = 32'b00000000000000000110000100111101;
assign LUT_3[50605] = 32'b00000000000000001100110000011010;
assign LUT_3[50606] = 32'b00000000000000001000001100100001;
assign LUT_3[50607] = 32'b00000000000000001110110111111110;
assign LUT_3[50608] = 32'b00000000000000000110110001000100;
assign LUT_3[50609] = 32'b00000000000000001101011100100001;
assign LUT_3[50610] = 32'b00000000000000001000111000101000;
assign LUT_3[50611] = 32'b00000000000000001111100100000101;
assign LUT_3[50612] = 32'b00000000000000000011111110111010;
assign LUT_3[50613] = 32'b00000000000000001010101010010111;
assign LUT_3[50614] = 32'b00000000000000000110000110011110;
assign LUT_3[50615] = 32'b00000000000000001100110001111011;
assign LUT_3[50616] = 32'b00000000000000001100001010001010;
assign LUT_3[50617] = 32'b00000000000000010010110101100111;
assign LUT_3[50618] = 32'b00000000000000001110010001101110;
assign LUT_3[50619] = 32'b00000000000000010100111101001011;
assign LUT_3[50620] = 32'b00000000000000001001011000000000;
assign LUT_3[50621] = 32'b00000000000000010000000011011101;
assign LUT_3[50622] = 32'b00000000000000001011011111100100;
assign LUT_3[50623] = 32'b00000000000000010010001011000001;
assign LUT_3[50624] = 32'b00000000000000000010001000001100;
assign LUT_3[50625] = 32'b00000000000000001000110011101001;
assign LUT_3[50626] = 32'b00000000000000000100001111110000;
assign LUT_3[50627] = 32'b00000000000000001010111011001101;
assign LUT_3[50628] = 32'b11111111111111111111010110000010;
assign LUT_3[50629] = 32'b00000000000000000110000001011111;
assign LUT_3[50630] = 32'b00000000000000000001011101100110;
assign LUT_3[50631] = 32'b00000000000000001000001001000011;
assign LUT_3[50632] = 32'b00000000000000000111100001010010;
assign LUT_3[50633] = 32'b00000000000000001110001100101111;
assign LUT_3[50634] = 32'b00000000000000001001101000110110;
assign LUT_3[50635] = 32'b00000000000000010000010100010011;
assign LUT_3[50636] = 32'b00000000000000000100101111001000;
assign LUT_3[50637] = 32'b00000000000000001011011010100101;
assign LUT_3[50638] = 32'b00000000000000000110110110101100;
assign LUT_3[50639] = 32'b00000000000000001101100010001001;
assign LUT_3[50640] = 32'b00000000000000000101011011001111;
assign LUT_3[50641] = 32'b00000000000000001100000110101100;
assign LUT_3[50642] = 32'b00000000000000000111100010110011;
assign LUT_3[50643] = 32'b00000000000000001110001110010000;
assign LUT_3[50644] = 32'b00000000000000000010101001000101;
assign LUT_3[50645] = 32'b00000000000000001001010100100010;
assign LUT_3[50646] = 32'b00000000000000000100110000101001;
assign LUT_3[50647] = 32'b00000000000000001011011100000110;
assign LUT_3[50648] = 32'b00000000000000001010110100010101;
assign LUT_3[50649] = 32'b00000000000000010001011111110010;
assign LUT_3[50650] = 32'b00000000000000001100111011111001;
assign LUT_3[50651] = 32'b00000000000000010011100111010110;
assign LUT_3[50652] = 32'b00000000000000001000000010001011;
assign LUT_3[50653] = 32'b00000000000000001110101101101000;
assign LUT_3[50654] = 32'b00000000000000001010001001101111;
assign LUT_3[50655] = 32'b00000000000000010000110101001100;
assign LUT_3[50656] = 32'b00000000000000000011010110101100;
assign LUT_3[50657] = 32'b00000000000000001010000010001001;
assign LUT_3[50658] = 32'b00000000000000000101011110010000;
assign LUT_3[50659] = 32'b00000000000000001100001001101101;
assign LUT_3[50660] = 32'b00000000000000000000100100100010;
assign LUT_3[50661] = 32'b00000000000000000111001111111111;
assign LUT_3[50662] = 32'b00000000000000000010101100000110;
assign LUT_3[50663] = 32'b00000000000000001001010111100011;
assign LUT_3[50664] = 32'b00000000000000001000101111110010;
assign LUT_3[50665] = 32'b00000000000000001111011011001111;
assign LUT_3[50666] = 32'b00000000000000001010110111010110;
assign LUT_3[50667] = 32'b00000000000000010001100010110011;
assign LUT_3[50668] = 32'b00000000000000000101111101101000;
assign LUT_3[50669] = 32'b00000000000000001100101001000101;
assign LUT_3[50670] = 32'b00000000000000001000000101001100;
assign LUT_3[50671] = 32'b00000000000000001110110000101001;
assign LUT_3[50672] = 32'b00000000000000000110101001101111;
assign LUT_3[50673] = 32'b00000000000000001101010101001100;
assign LUT_3[50674] = 32'b00000000000000001000110001010011;
assign LUT_3[50675] = 32'b00000000000000001111011100110000;
assign LUT_3[50676] = 32'b00000000000000000011110111100101;
assign LUT_3[50677] = 32'b00000000000000001010100011000010;
assign LUT_3[50678] = 32'b00000000000000000101111111001001;
assign LUT_3[50679] = 32'b00000000000000001100101010100110;
assign LUT_3[50680] = 32'b00000000000000001100000010110101;
assign LUT_3[50681] = 32'b00000000000000010010101110010010;
assign LUT_3[50682] = 32'b00000000000000001110001010011001;
assign LUT_3[50683] = 32'b00000000000000010100110101110110;
assign LUT_3[50684] = 32'b00000000000000001001010000101011;
assign LUT_3[50685] = 32'b00000000000000001111111100001000;
assign LUT_3[50686] = 32'b00000000000000001011011000001111;
assign LUT_3[50687] = 32'b00000000000000010010000011101100;
assign LUT_3[50688] = 32'b00000000000000000111001010001110;
assign LUT_3[50689] = 32'b00000000000000001101110101101011;
assign LUT_3[50690] = 32'b00000000000000001001010001110010;
assign LUT_3[50691] = 32'b00000000000000001111111101001111;
assign LUT_3[50692] = 32'b00000000000000000100011000000100;
assign LUT_3[50693] = 32'b00000000000000001011000011100001;
assign LUT_3[50694] = 32'b00000000000000000110011111101000;
assign LUT_3[50695] = 32'b00000000000000001101001011000101;
assign LUT_3[50696] = 32'b00000000000000001100100011010100;
assign LUT_3[50697] = 32'b00000000000000010011001110110001;
assign LUT_3[50698] = 32'b00000000000000001110101010111000;
assign LUT_3[50699] = 32'b00000000000000010101010110010101;
assign LUT_3[50700] = 32'b00000000000000001001110001001010;
assign LUT_3[50701] = 32'b00000000000000010000011100100111;
assign LUT_3[50702] = 32'b00000000000000001011111000101110;
assign LUT_3[50703] = 32'b00000000000000010010100100001011;
assign LUT_3[50704] = 32'b00000000000000001010011101010001;
assign LUT_3[50705] = 32'b00000000000000010001001000101110;
assign LUT_3[50706] = 32'b00000000000000001100100100110101;
assign LUT_3[50707] = 32'b00000000000000010011010000010010;
assign LUT_3[50708] = 32'b00000000000000000111101011000111;
assign LUT_3[50709] = 32'b00000000000000001110010110100100;
assign LUT_3[50710] = 32'b00000000000000001001110010101011;
assign LUT_3[50711] = 32'b00000000000000010000011110001000;
assign LUT_3[50712] = 32'b00000000000000001111110110010111;
assign LUT_3[50713] = 32'b00000000000000010110100001110100;
assign LUT_3[50714] = 32'b00000000000000010001111101111011;
assign LUT_3[50715] = 32'b00000000000000011000101001011000;
assign LUT_3[50716] = 32'b00000000000000001101000100001101;
assign LUT_3[50717] = 32'b00000000000000010011101111101010;
assign LUT_3[50718] = 32'b00000000000000001111001011110001;
assign LUT_3[50719] = 32'b00000000000000010101110111001110;
assign LUT_3[50720] = 32'b00000000000000001000011000101110;
assign LUT_3[50721] = 32'b00000000000000001111000100001011;
assign LUT_3[50722] = 32'b00000000000000001010100000010010;
assign LUT_3[50723] = 32'b00000000000000010001001011101111;
assign LUT_3[50724] = 32'b00000000000000000101100110100100;
assign LUT_3[50725] = 32'b00000000000000001100010010000001;
assign LUT_3[50726] = 32'b00000000000000000111101110001000;
assign LUT_3[50727] = 32'b00000000000000001110011001100101;
assign LUT_3[50728] = 32'b00000000000000001101110001110100;
assign LUT_3[50729] = 32'b00000000000000010100011101010001;
assign LUT_3[50730] = 32'b00000000000000001111111001011000;
assign LUT_3[50731] = 32'b00000000000000010110100100110101;
assign LUT_3[50732] = 32'b00000000000000001010111111101010;
assign LUT_3[50733] = 32'b00000000000000010001101011000111;
assign LUT_3[50734] = 32'b00000000000000001101000111001110;
assign LUT_3[50735] = 32'b00000000000000010011110010101011;
assign LUT_3[50736] = 32'b00000000000000001011101011110001;
assign LUT_3[50737] = 32'b00000000000000010010010111001110;
assign LUT_3[50738] = 32'b00000000000000001101110011010101;
assign LUT_3[50739] = 32'b00000000000000010100011110110010;
assign LUT_3[50740] = 32'b00000000000000001000111001100111;
assign LUT_3[50741] = 32'b00000000000000001111100101000100;
assign LUT_3[50742] = 32'b00000000000000001011000001001011;
assign LUT_3[50743] = 32'b00000000000000010001101100101000;
assign LUT_3[50744] = 32'b00000000000000010001000100110111;
assign LUT_3[50745] = 32'b00000000000000010111110000010100;
assign LUT_3[50746] = 32'b00000000000000010011001100011011;
assign LUT_3[50747] = 32'b00000000000000011001110111111000;
assign LUT_3[50748] = 32'b00000000000000001110010010101101;
assign LUT_3[50749] = 32'b00000000000000010100111110001010;
assign LUT_3[50750] = 32'b00000000000000010000011010010001;
assign LUT_3[50751] = 32'b00000000000000010111000101101110;
assign LUT_3[50752] = 32'b00000000000000000111000010111001;
assign LUT_3[50753] = 32'b00000000000000001101101110010110;
assign LUT_3[50754] = 32'b00000000000000001001001010011101;
assign LUT_3[50755] = 32'b00000000000000001111110101111010;
assign LUT_3[50756] = 32'b00000000000000000100010000101111;
assign LUT_3[50757] = 32'b00000000000000001010111100001100;
assign LUT_3[50758] = 32'b00000000000000000110011000010011;
assign LUT_3[50759] = 32'b00000000000000001101000011110000;
assign LUT_3[50760] = 32'b00000000000000001100011011111111;
assign LUT_3[50761] = 32'b00000000000000010011000111011100;
assign LUT_3[50762] = 32'b00000000000000001110100011100011;
assign LUT_3[50763] = 32'b00000000000000010101001111000000;
assign LUT_3[50764] = 32'b00000000000000001001101001110101;
assign LUT_3[50765] = 32'b00000000000000010000010101010010;
assign LUT_3[50766] = 32'b00000000000000001011110001011001;
assign LUT_3[50767] = 32'b00000000000000010010011100110110;
assign LUT_3[50768] = 32'b00000000000000001010010101111100;
assign LUT_3[50769] = 32'b00000000000000010001000001011001;
assign LUT_3[50770] = 32'b00000000000000001100011101100000;
assign LUT_3[50771] = 32'b00000000000000010011001000111101;
assign LUT_3[50772] = 32'b00000000000000000111100011110010;
assign LUT_3[50773] = 32'b00000000000000001110001111001111;
assign LUT_3[50774] = 32'b00000000000000001001101011010110;
assign LUT_3[50775] = 32'b00000000000000010000010110110011;
assign LUT_3[50776] = 32'b00000000000000001111101111000010;
assign LUT_3[50777] = 32'b00000000000000010110011010011111;
assign LUT_3[50778] = 32'b00000000000000010001110110100110;
assign LUT_3[50779] = 32'b00000000000000011000100010000011;
assign LUT_3[50780] = 32'b00000000000000001100111100111000;
assign LUT_3[50781] = 32'b00000000000000010011101000010101;
assign LUT_3[50782] = 32'b00000000000000001111000100011100;
assign LUT_3[50783] = 32'b00000000000000010101101111111001;
assign LUT_3[50784] = 32'b00000000000000001000010001011001;
assign LUT_3[50785] = 32'b00000000000000001110111100110110;
assign LUT_3[50786] = 32'b00000000000000001010011000111101;
assign LUT_3[50787] = 32'b00000000000000010001000100011010;
assign LUT_3[50788] = 32'b00000000000000000101011111001111;
assign LUT_3[50789] = 32'b00000000000000001100001010101100;
assign LUT_3[50790] = 32'b00000000000000000111100110110011;
assign LUT_3[50791] = 32'b00000000000000001110010010010000;
assign LUT_3[50792] = 32'b00000000000000001101101010011111;
assign LUT_3[50793] = 32'b00000000000000010100010101111100;
assign LUT_3[50794] = 32'b00000000000000001111110010000011;
assign LUT_3[50795] = 32'b00000000000000010110011101100000;
assign LUT_3[50796] = 32'b00000000000000001010111000010101;
assign LUT_3[50797] = 32'b00000000000000010001100011110010;
assign LUT_3[50798] = 32'b00000000000000001100111111111001;
assign LUT_3[50799] = 32'b00000000000000010011101011010110;
assign LUT_3[50800] = 32'b00000000000000001011100100011100;
assign LUT_3[50801] = 32'b00000000000000010010001111111001;
assign LUT_3[50802] = 32'b00000000000000001101101100000000;
assign LUT_3[50803] = 32'b00000000000000010100010111011101;
assign LUT_3[50804] = 32'b00000000000000001000110010010010;
assign LUT_3[50805] = 32'b00000000000000001111011101101111;
assign LUT_3[50806] = 32'b00000000000000001010111001110110;
assign LUT_3[50807] = 32'b00000000000000010001100101010011;
assign LUT_3[50808] = 32'b00000000000000010000111101100010;
assign LUT_3[50809] = 32'b00000000000000010111101000111111;
assign LUT_3[50810] = 32'b00000000000000010011000101000110;
assign LUT_3[50811] = 32'b00000000000000011001110000100011;
assign LUT_3[50812] = 32'b00000000000000001110001011011000;
assign LUT_3[50813] = 32'b00000000000000010100110110110101;
assign LUT_3[50814] = 32'b00000000000000010000010010111100;
assign LUT_3[50815] = 32'b00000000000000010110111110011001;
assign LUT_3[50816] = 32'b00000000000000001001010101001100;
assign LUT_3[50817] = 32'b00000000000000010000000000101001;
assign LUT_3[50818] = 32'b00000000000000001011011100110000;
assign LUT_3[50819] = 32'b00000000000000010010001000001101;
assign LUT_3[50820] = 32'b00000000000000000110100011000010;
assign LUT_3[50821] = 32'b00000000000000001101001110011111;
assign LUT_3[50822] = 32'b00000000000000001000101010100110;
assign LUT_3[50823] = 32'b00000000000000001111010110000011;
assign LUT_3[50824] = 32'b00000000000000001110101110010010;
assign LUT_3[50825] = 32'b00000000000000010101011001101111;
assign LUT_3[50826] = 32'b00000000000000010000110101110110;
assign LUT_3[50827] = 32'b00000000000000010111100001010011;
assign LUT_3[50828] = 32'b00000000000000001011111100001000;
assign LUT_3[50829] = 32'b00000000000000010010100111100101;
assign LUT_3[50830] = 32'b00000000000000001110000011101100;
assign LUT_3[50831] = 32'b00000000000000010100101111001001;
assign LUT_3[50832] = 32'b00000000000000001100101000001111;
assign LUT_3[50833] = 32'b00000000000000010011010011101100;
assign LUT_3[50834] = 32'b00000000000000001110101111110011;
assign LUT_3[50835] = 32'b00000000000000010101011011010000;
assign LUT_3[50836] = 32'b00000000000000001001110110000101;
assign LUT_3[50837] = 32'b00000000000000010000100001100010;
assign LUT_3[50838] = 32'b00000000000000001011111101101001;
assign LUT_3[50839] = 32'b00000000000000010010101001000110;
assign LUT_3[50840] = 32'b00000000000000010010000001010101;
assign LUT_3[50841] = 32'b00000000000000011000101100110010;
assign LUT_3[50842] = 32'b00000000000000010100001000111001;
assign LUT_3[50843] = 32'b00000000000000011010110100010110;
assign LUT_3[50844] = 32'b00000000000000001111001111001011;
assign LUT_3[50845] = 32'b00000000000000010101111010101000;
assign LUT_3[50846] = 32'b00000000000000010001010110101111;
assign LUT_3[50847] = 32'b00000000000000011000000010001100;
assign LUT_3[50848] = 32'b00000000000000001010100011101100;
assign LUT_3[50849] = 32'b00000000000000010001001111001001;
assign LUT_3[50850] = 32'b00000000000000001100101011010000;
assign LUT_3[50851] = 32'b00000000000000010011010110101101;
assign LUT_3[50852] = 32'b00000000000000000111110001100010;
assign LUT_3[50853] = 32'b00000000000000001110011100111111;
assign LUT_3[50854] = 32'b00000000000000001001111001000110;
assign LUT_3[50855] = 32'b00000000000000010000100100100011;
assign LUT_3[50856] = 32'b00000000000000001111111100110010;
assign LUT_3[50857] = 32'b00000000000000010110101000001111;
assign LUT_3[50858] = 32'b00000000000000010010000100010110;
assign LUT_3[50859] = 32'b00000000000000011000101111110011;
assign LUT_3[50860] = 32'b00000000000000001101001010101000;
assign LUT_3[50861] = 32'b00000000000000010011110110000101;
assign LUT_3[50862] = 32'b00000000000000001111010010001100;
assign LUT_3[50863] = 32'b00000000000000010101111101101001;
assign LUT_3[50864] = 32'b00000000000000001101110110101111;
assign LUT_3[50865] = 32'b00000000000000010100100010001100;
assign LUT_3[50866] = 32'b00000000000000001111111110010011;
assign LUT_3[50867] = 32'b00000000000000010110101001110000;
assign LUT_3[50868] = 32'b00000000000000001011000100100101;
assign LUT_3[50869] = 32'b00000000000000010001110000000010;
assign LUT_3[50870] = 32'b00000000000000001101001100001001;
assign LUT_3[50871] = 32'b00000000000000010011110111100110;
assign LUT_3[50872] = 32'b00000000000000010011001111110101;
assign LUT_3[50873] = 32'b00000000000000011001111011010010;
assign LUT_3[50874] = 32'b00000000000000010101010111011001;
assign LUT_3[50875] = 32'b00000000000000011100000010110110;
assign LUT_3[50876] = 32'b00000000000000010000011101101011;
assign LUT_3[50877] = 32'b00000000000000010111001001001000;
assign LUT_3[50878] = 32'b00000000000000010010100101001111;
assign LUT_3[50879] = 32'b00000000000000011001010000101100;
assign LUT_3[50880] = 32'b00000000000000001001001101110111;
assign LUT_3[50881] = 32'b00000000000000001111111001010100;
assign LUT_3[50882] = 32'b00000000000000001011010101011011;
assign LUT_3[50883] = 32'b00000000000000010010000000111000;
assign LUT_3[50884] = 32'b00000000000000000110011011101101;
assign LUT_3[50885] = 32'b00000000000000001101000111001010;
assign LUT_3[50886] = 32'b00000000000000001000100011010001;
assign LUT_3[50887] = 32'b00000000000000001111001110101110;
assign LUT_3[50888] = 32'b00000000000000001110100110111101;
assign LUT_3[50889] = 32'b00000000000000010101010010011010;
assign LUT_3[50890] = 32'b00000000000000010000101110100001;
assign LUT_3[50891] = 32'b00000000000000010111011001111110;
assign LUT_3[50892] = 32'b00000000000000001011110100110011;
assign LUT_3[50893] = 32'b00000000000000010010100000010000;
assign LUT_3[50894] = 32'b00000000000000001101111100010111;
assign LUT_3[50895] = 32'b00000000000000010100100111110100;
assign LUT_3[50896] = 32'b00000000000000001100100000111010;
assign LUT_3[50897] = 32'b00000000000000010011001100010111;
assign LUT_3[50898] = 32'b00000000000000001110101000011110;
assign LUT_3[50899] = 32'b00000000000000010101010011111011;
assign LUT_3[50900] = 32'b00000000000000001001101110110000;
assign LUT_3[50901] = 32'b00000000000000010000011010001101;
assign LUT_3[50902] = 32'b00000000000000001011110110010100;
assign LUT_3[50903] = 32'b00000000000000010010100001110001;
assign LUT_3[50904] = 32'b00000000000000010001111010000000;
assign LUT_3[50905] = 32'b00000000000000011000100101011101;
assign LUT_3[50906] = 32'b00000000000000010100000001100100;
assign LUT_3[50907] = 32'b00000000000000011010101101000001;
assign LUT_3[50908] = 32'b00000000000000001111000111110110;
assign LUT_3[50909] = 32'b00000000000000010101110011010011;
assign LUT_3[50910] = 32'b00000000000000010001001111011010;
assign LUT_3[50911] = 32'b00000000000000010111111010110111;
assign LUT_3[50912] = 32'b00000000000000001010011100010111;
assign LUT_3[50913] = 32'b00000000000000010001000111110100;
assign LUT_3[50914] = 32'b00000000000000001100100011111011;
assign LUT_3[50915] = 32'b00000000000000010011001111011000;
assign LUT_3[50916] = 32'b00000000000000000111101010001101;
assign LUT_3[50917] = 32'b00000000000000001110010101101010;
assign LUT_3[50918] = 32'b00000000000000001001110001110001;
assign LUT_3[50919] = 32'b00000000000000010000011101001110;
assign LUT_3[50920] = 32'b00000000000000001111110101011101;
assign LUT_3[50921] = 32'b00000000000000010110100000111010;
assign LUT_3[50922] = 32'b00000000000000010001111101000001;
assign LUT_3[50923] = 32'b00000000000000011000101000011110;
assign LUT_3[50924] = 32'b00000000000000001101000011010011;
assign LUT_3[50925] = 32'b00000000000000010011101110110000;
assign LUT_3[50926] = 32'b00000000000000001111001010110111;
assign LUT_3[50927] = 32'b00000000000000010101110110010100;
assign LUT_3[50928] = 32'b00000000000000001101101111011010;
assign LUT_3[50929] = 32'b00000000000000010100011010110111;
assign LUT_3[50930] = 32'b00000000000000001111110110111110;
assign LUT_3[50931] = 32'b00000000000000010110100010011011;
assign LUT_3[50932] = 32'b00000000000000001010111101010000;
assign LUT_3[50933] = 32'b00000000000000010001101000101101;
assign LUT_3[50934] = 32'b00000000000000001101000100110100;
assign LUT_3[50935] = 32'b00000000000000010011110000010001;
assign LUT_3[50936] = 32'b00000000000000010011001000100000;
assign LUT_3[50937] = 32'b00000000000000011001110011111101;
assign LUT_3[50938] = 32'b00000000000000010101010000000100;
assign LUT_3[50939] = 32'b00000000000000011011111011100001;
assign LUT_3[50940] = 32'b00000000000000010000010110010110;
assign LUT_3[50941] = 32'b00000000000000010111000001110011;
assign LUT_3[50942] = 32'b00000000000000010010011101111010;
assign LUT_3[50943] = 32'b00000000000000011001001001010111;
assign LUT_3[50944] = 32'b00000000000000000011011001101111;
assign LUT_3[50945] = 32'b00000000000000001010000101001100;
assign LUT_3[50946] = 32'b00000000000000000101100001010011;
assign LUT_3[50947] = 32'b00000000000000001100001100110000;
assign LUT_3[50948] = 32'b00000000000000000000100111100101;
assign LUT_3[50949] = 32'b00000000000000000111010011000010;
assign LUT_3[50950] = 32'b00000000000000000010101111001001;
assign LUT_3[50951] = 32'b00000000000000001001011010100110;
assign LUT_3[50952] = 32'b00000000000000001000110010110101;
assign LUT_3[50953] = 32'b00000000000000001111011110010010;
assign LUT_3[50954] = 32'b00000000000000001010111010011001;
assign LUT_3[50955] = 32'b00000000000000010001100101110110;
assign LUT_3[50956] = 32'b00000000000000000110000000101011;
assign LUT_3[50957] = 32'b00000000000000001100101100001000;
assign LUT_3[50958] = 32'b00000000000000001000001000001111;
assign LUT_3[50959] = 32'b00000000000000001110110011101100;
assign LUT_3[50960] = 32'b00000000000000000110101100110010;
assign LUT_3[50961] = 32'b00000000000000001101011000001111;
assign LUT_3[50962] = 32'b00000000000000001000110100010110;
assign LUT_3[50963] = 32'b00000000000000001111011111110011;
assign LUT_3[50964] = 32'b00000000000000000011111010101000;
assign LUT_3[50965] = 32'b00000000000000001010100110000101;
assign LUT_3[50966] = 32'b00000000000000000110000010001100;
assign LUT_3[50967] = 32'b00000000000000001100101101101001;
assign LUT_3[50968] = 32'b00000000000000001100000101111000;
assign LUT_3[50969] = 32'b00000000000000010010110001010101;
assign LUT_3[50970] = 32'b00000000000000001110001101011100;
assign LUT_3[50971] = 32'b00000000000000010100111000111001;
assign LUT_3[50972] = 32'b00000000000000001001010011101110;
assign LUT_3[50973] = 32'b00000000000000001111111111001011;
assign LUT_3[50974] = 32'b00000000000000001011011011010010;
assign LUT_3[50975] = 32'b00000000000000010010000110101111;
assign LUT_3[50976] = 32'b00000000000000000100101000001111;
assign LUT_3[50977] = 32'b00000000000000001011010011101100;
assign LUT_3[50978] = 32'b00000000000000000110101111110011;
assign LUT_3[50979] = 32'b00000000000000001101011011010000;
assign LUT_3[50980] = 32'b00000000000000000001110110000101;
assign LUT_3[50981] = 32'b00000000000000001000100001100010;
assign LUT_3[50982] = 32'b00000000000000000011111101101001;
assign LUT_3[50983] = 32'b00000000000000001010101001000110;
assign LUT_3[50984] = 32'b00000000000000001010000001010101;
assign LUT_3[50985] = 32'b00000000000000010000101100110010;
assign LUT_3[50986] = 32'b00000000000000001100001000111001;
assign LUT_3[50987] = 32'b00000000000000010010110100010110;
assign LUT_3[50988] = 32'b00000000000000000111001111001011;
assign LUT_3[50989] = 32'b00000000000000001101111010101000;
assign LUT_3[50990] = 32'b00000000000000001001010110101111;
assign LUT_3[50991] = 32'b00000000000000010000000010001100;
assign LUT_3[50992] = 32'b00000000000000000111111011010010;
assign LUT_3[50993] = 32'b00000000000000001110100110101111;
assign LUT_3[50994] = 32'b00000000000000001010000010110110;
assign LUT_3[50995] = 32'b00000000000000010000101110010011;
assign LUT_3[50996] = 32'b00000000000000000101001001001000;
assign LUT_3[50997] = 32'b00000000000000001011110100100101;
assign LUT_3[50998] = 32'b00000000000000000111010000101100;
assign LUT_3[50999] = 32'b00000000000000001101111100001001;
assign LUT_3[51000] = 32'b00000000000000001101010100011000;
assign LUT_3[51001] = 32'b00000000000000010011111111110101;
assign LUT_3[51002] = 32'b00000000000000001111011011111100;
assign LUT_3[51003] = 32'b00000000000000010110000111011001;
assign LUT_3[51004] = 32'b00000000000000001010100010001110;
assign LUT_3[51005] = 32'b00000000000000010001001101101011;
assign LUT_3[51006] = 32'b00000000000000001100101001110010;
assign LUT_3[51007] = 32'b00000000000000010011010101001111;
assign LUT_3[51008] = 32'b00000000000000000011010010011010;
assign LUT_3[51009] = 32'b00000000000000001001111101110111;
assign LUT_3[51010] = 32'b00000000000000000101011001111110;
assign LUT_3[51011] = 32'b00000000000000001100000101011011;
assign LUT_3[51012] = 32'b00000000000000000000100000010000;
assign LUT_3[51013] = 32'b00000000000000000111001011101101;
assign LUT_3[51014] = 32'b00000000000000000010100111110100;
assign LUT_3[51015] = 32'b00000000000000001001010011010001;
assign LUT_3[51016] = 32'b00000000000000001000101011100000;
assign LUT_3[51017] = 32'b00000000000000001111010110111101;
assign LUT_3[51018] = 32'b00000000000000001010110011000100;
assign LUT_3[51019] = 32'b00000000000000010001011110100001;
assign LUT_3[51020] = 32'b00000000000000000101111001010110;
assign LUT_3[51021] = 32'b00000000000000001100100100110011;
assign LUT_3[51022] = 32'b00000000000000001000000000111010;
assign LUT_3[51023] = 32'b00000000000000001110101100010111;
assign LUT_3[51024] = 32'b00000000000000000110100101011101;
assign LUT_3[51025] = 32'b00000000000000001101010000111010;
assign LUT_3[51026] = 32'b00000000000000001000101101000001;
assign LUT_3[51027] = 32'b00000000000000001111011000011110;
assign LUT_3[51028] = 32'b00000000000000000011110011010011;
assign LUT_3[51029] = 32'b00000000000000001010011110110000;
assign LUT_3[51030] = 32'b00000000000000000101111010110111;
assign LUT_3[51031] = 32'b00000000000000001100100110010100;
assign LUT_3[51032] = 32'b00000000000000001011111110100011;
assign LUT_3[51033] = 32'b00000000000000010010101010000000;
assign LUT_3[51034] = 32'b00000000000000001110000110000111;
assign LUT_3[51035] = 32'b00000000000000010100110001100100;
assign LUT_3[51036] = 32'b00000000000000001001001100011001;
assign LUT_3[51037] = 32'b00000000000000001111110111110110;
assign LUT_3[51038] = 32'b00000000000000001011010011111101;
assign LUT_3[51039] = 32'b00000000000000010001111111011010;
assign LUT_3[51040] = 32'b00000000000000000100100000111010;
assign LUT_3[51041] = 32'b00000000000000001011001100010111;
assign LUT_3[51042] = 32'b00000000000000000110101000011110;
assign LUT_3[51043] = 32'b00000000000000001101010011111011;
assign LUT_3[51044] = 32'b00000000000000000001101110110000;
assign LUT_3[51045] = 32'b00000000000000001000011010001101;
assign LUT_3[51046] = 32'b00000000000000000011110110010100;
assign LUT_3[51047] = 32'b00000000000000001010100001110001;
assign LUT_3[51048] = 32'b00000000000000001001111010000000;
assign LUT_3[51049] = 32'b00000000000000010000100101011101;
assign LUT_3[51050] = 32'b00000000000000001100000001100100;
assign LUT_3[51051] = 32'b00000000000000010010101101000001;
assign LUT_3[51052] = 32'b00000000000000000111000111110110;
assign LUT_3[51053] = 32'b00000000000000001101110011010011;
assign LUT_3[51054] = 32'b00000000000000001001001111011010;
assign LUT_3[51055] = 32'b00000000000000001111111010110111;
assign LUT_3[51056] = 32'b00000000000000000111110011111101;
assign LUT_3[51057] = 32'b00000000000000001110011111011010;
assign LUT_3[51058] = 32'b00000000000000001001111011100001;
assign LUT_3[51059] = 32'b00000000000000010000100110111110;
assign LUT_3[51060] = 32'b00000000000000000101000001110011;
assign LUT_3[51061] = 32'b00000000000000001011101101010000;
assign LUT_3[51062] = 32'b00000000000000000111001001010111;
assign LUT_3[51063] = 32'b00000000000000001101110100110100;
assign LUT_3[51064] = 32'b00000000000000001101001101000011;
assign LUT_3[51065] = 32'b00000000000000010011111000100000;
assign LUT_3[51066] = 32'b00000000000000001111010100100111;
assign LUT_3[51067] = 32'b00000000000000010110000000000100;
assign LUT_3[51068] = 32'b00000000000000001010011010111001;
assign LUT_3[51069] = 32'b00000000000000010001000110010110;
assign LUT_3[51070] = 32'b00000000000000001100100010011101;
assign LUT_3[51071] = 32'b00000000000000010011001101111010;
assign LUT_3[51072] = 32'b00000000000000000101100100101101;
assign LUT_3[51073] = 32'b00000000000000001100010000001010;
assign LUT_3[51074] = 32'b00000000000000000111101100010001;
assign LUT_3[51075] = 32'b00000000000000001110010111101110;
assign LUT_3[51076] = 32'b00000000000000000010110010100011;
assign LUT_3[51077] = 32'b00000000000000001001011110000000;
assign LUT_3[51078] = 32'b00000000000000000100111010000111;
assign LUT_3[51079] = 32'b00000000000000001011100101100100;
assign LUT_3[51080] = 32'b00000000000000001010111101110011;
assign LUT_3[51081] = 32'b00000000000000010001101001010000;
assign LUT_3[51082] = 32'b00000000000000001101000101010111;
assign LUT_3[51083] = 32'b00000000000000010011110000110100;
assign LUT_3[51084] = 32'b00000000000000001000001011101001;
assign LUT_3[51085] = 32'b00000000000000001110110111000110;
assign LUT_3[51086] = 32'b00000000000000001010010011001101;
assign LUT_3[51087] = 32'b00000000000000010000111110101010;
assign LUT_3[51088] = 32'b00000000000000001000110111110000;
assign LUT_3[51089] = 32'b00000000000000001111100011001101;
assign LUT_3[51090] = 32'b00000000000000001010111111010100;
assign LUT_3[51091] = 32'b00000000000000010001101010110001;
assign LUT_3[51092] = 32'b00000000000000000110000101100110;
assign LUT_3[51093] = 32'b00000000000000001100110001000011;
assign LUT_3[51094] = 32'b00000000000000001000001101001010;
assign LUT_3[51095] = 32'b00000000000000001110111000100111;
assign LUT_3[51096] = 32'b00000000000000001110010000110110;
assign LUT_3[51097] = 32'b00000000000000010100111100010011;
assign LUT_3[51098] = 32'b00000000000000010000011000011010;
assign LUT_3[51099] = 32'b00000000000000010111000011110111;
assign LUT_3[51100] = 32'b00000000000000001011011110101100;
assign LUT_3[51101] = 32'b00000000000000010010001010001001;
assign LUT_3[51102] = 32'b00000000000000001101100110010000;
assign LUT_3[51103] = 32'b00000000000000010100010001101101;
assign LUT_3[51104] = 32'b00000000000000000110110011001101;
assign LUT_3[51105] = 32'b00000000000000001101011110101010;
assign LUT_3[51106] = 32'b00000000000000001000111010110001;
assign LUT_3[51107] = 32'b00000000000000001111100110001110;
assign LUT_3[51108] = 32'b00000000000000000100000001000011;
assign LUT_3[51109] = 32'b00000000000000001010101100100000;
assign LUT_3[51110] = 32'b00000000000000000110001000100111;
assign LUT_3[51111] = 32'b00000000000000001100110100000100;
assign LUT_3[51112] = 32'b00000000000000001100001100010011;
assign LUT_3[51113] = 32'b00000000000000010010110111110000;
assign LUT_3[51114] = 32'b00000000000000001110010011110111;
assign LUT_3[51115] = 32'b00000000000000010100111111010100;
assign LUT_3[51116] = 32'b00000000000000001001011010001001;
assign LUT_3[51117] = 32'b00000000000000010000000101100110;
assign LUT_3[51118] = 32'b00000000000000001011100001101101;
assign LUT_3[51119] = 32'b00000000000000010010001101001010;
assign LUT_3[51120] = 32'b00000000000000001010000110010000;
assign LUT_3[51121] = 32'b00000000000000010000110001101101;
assign LUT_3[51122] = 32'b00000000000000001100001101110100;
assign LUT_3[51123] = 32'b00000000000000010010111001010001;
assign LUT_3[51124] = 32'b00000000000000000111010100000110;
assign LUT_3[51125] = 32'b00000000000000001101111111100011;
assign LUT_3[51126] = 32'b00000000000000001001011011101010;
assign LUT_3[51127] = 32'b00000000000000010000000111000111;
assign LUT_3[51128] = 32'b00000000000000001111011111010110;
assign LUT_3[51129] = 32'b00000000000000010110001010110011;
assign LUT_3[51130] = 32'b00000000000000010001100110111010;
assign LUT_3[51131] = 32'b00000000000000011000010010010111;
assign LUT_3[51132] = 32'b00000000000000001100101101001100;
assign LUT_3[51133] = 32'b00000000000000010011011000101001;
assign LUT_3[51134] = 32'b00000000000000001110110100110000;
assign LUT_3[51135] = 32'b00000000000000010101100000001101;
assign LUT_3[51136] = 32'b00000000000000000101011101011000;
assign LUT_3[51137] = 32'b00000000000000001100001000110101;
assign LUT_3[51138] = 32'b00000000000000000111100100111100;
assign LUT_3[51139] = 32'b00000000000000001110010000011001;
assign LUT_3[51140] = 32'b00000000000000000010101011001110;
assign LUT_3[51141] = 32'b00000000000000001001010110101011;
assign LUT_3[51142] = 32'b00000000000000000100110010110010;
assign LUT_3[51143] = 32'b00000000000000001011011110001111;
assign LUT_3[51144] = 32'b00000000000000001010110110011110;
assign LUT_3[51145] = 32'b00000000000000010001100001111011;
assign LUT_3[51146] = 32'b00000000000000001100111110000010;
assign LUT_3[51147] = 32'b00000000000000010011101001011111;
assign LUT_3[51148] = 32'b00000000000000001000000100010100;
assign LUT_3[51149] = 32'b00000000000000001110101111110001;
assign LUT_3[51150] = 32'b00000000000000001010001011111000;
assign LUT_3[51151] = 32'b00000000000000010000110111010101;
assign LUT_3[51152] = 32'b00000000000000001000110000011011;
assign LUT_3[51153] = 32'b00000000000000001111011011111000;
assign LUT_3[51154] = 32'b00000000000000001010110111111111;
assign LUT_3[51155] = 32'b00000000000000010001100011011100;
assign LUT_3[51156] = 32'b00000000000000000101111110010001;
assign LUT_3[51157] = 32'b00000000000000001100101001101110;
assign LUT_3[51158] = 32'b00000000000000001000000101110101;
assign LUT_3[51159] = 32'b00000000000000001110110001010010;
assign LUT_3[51160] = 32'b00000000000000001110001001100001;
assign LUT_3[51161] = 32'b00000000000000010100110100111110;
assign LUT_3[51162] = 32'b00000000000000010000010001000101;
assign LUT_3[51163] = 32'b00000000000000010110111100100010;
assign LUT_3[51164] = 32'b00000000000000001011010111010111;
assign LUT_3[51165] = 32'b00000000000000010010000010110100;
assign LUT_3[51166] = 32'b00000000000000001101011110111011;
assign LUT_3[51167] = 32'b00000000000000010100001010011000;
assign LUT_3[51168] = 32'b00000000000000000110101011111000;
assign LUT_3[51169] = 32'b00000000000000001101010111010101;
assign LUT_3[51170] = 32'b00000000000000001000110011011100;
assign LUT_3[51171] = 32'b00000000000000001111011110111001;
assign LUT_3[51172] = 32'b00000000000000000011111001101110;
assign LUT_3[51173] = 32'b00000000000000001010100101001011;
assign LUT_3[51174] = 32'b00000000000000000110000001010010;
assign LUT_3[51175] = 32'b00000000000000001100101100101111;
assign LUT_3[51176] = 32'b00000000000000001100000100111110;
assign LUT_3[51177] = 32'b00000000000000010010110000011011;
assign LUT_3[51178] = 32'b00000000000000001110001100100010;
assign LUT_3[51179] = 32'b00000000000000010100110111111111;
assign LUT_3[51180] = 32'b00000000000000001001010010110100;
assign LUT_3[51181] = 32'b00000000000000001111111110010001;
assign LUT_3[51182] = 32'b00000000000000001011011010011000;
assign LUT_3[51183] = 32'b00000000000000010010000101110101;
assign LUT_3[51184] = 32'b00000000000000001001111110111011;
assign LUT_3[51185] = 32'b00000000000000010000101010011000;
assign LUT_3[51186] = 32'b00000000000000001100000110011111;
assign LUT_3[51187] = 32'b00000000000000010010110001111100;
assign LUT_3[51188] = 32'b00000000000000000111001100110001;
assign LUT_3[51189] = 32'b00000000000000001101111000001110;
assign LUT_3[51190] = 32'b00000000000000001001010100010101;
assign LUT_3[51191] = 32'b00000000000000001111111111110010;
assign LUT_3[51192] = 32'b00000000000000001111011000000001;
assign LUT_3[51193] = 32'b00000000000000010110000011011110;
assign LUT_3[51194] = 32'b00000000000000010001011111100101;
assign LUT_3[51195] = 32'b00000000000000011000001011000010;
assign LUT_3[51196] = 32'b00000000000000001100100101110111;
assign LUT_3[51197] = 32'b00000000000000010011010001010100;
assign LUT_3[51198] = 32'b00000000000000001110101101011011;
assign LUT_3[51199] = 32'b00000000000000010101011000111000;
assign LUT_3[51200] = 32'b11111111111111111111000110010011;
assign LUT_3[51201] = 32'b00000000000000000101110001110000;
assign LUT_3[51202] = 32'b00000000000000000001001101110111;
assign LUT_3[51203] = 32'b00000000000000000111111001010100;
assign LUT_3[51204] = 32'b11111111111111111100010100001001;
assign LUT_3[51205] = 32'b00000000000000000010111111100110;
assign LUT_3[51206] = 32'b11111111111111111110011011101101;
assign LUT_3[51207] = 32'b00000000000000000101000111001010;
assign LUT_3[51208] = 32'b00000000000000000100011111011001;
assign LUT_3[51209] = 32'b00000000000000001011001010110110;
assign LUT_3[51210] = 32'b00000000000000000110100110111101;
assign LUT_3[51211] = 32'b00000000000000001101010010011010;
assign LUT_3[51212] = 32'b00000000000000000001101101001111;
assign LUT_3[51213] = 32'b00000000000000001000011000101100;
assign LUT_3[51214] = 32'b00000000000000000011110100110011;
assign LUT_3[51215] = 32'b00000000000000001010100000010000;
assign LUT_3[51216] = 32'b00000000000000000010011001010110;
assign LUT_3[51217] = 32'b00000000000000001001000100110011;
assign LUT_3[51218] = 32'b00000000000000000100100000111010;
assign LUT_3[51219] = 32'b00000000000000001011001100010111;
assign LUT_3[51220] = 32'b11111111111111111111100111001100;
assign LUT_3[51221] = 32'b00000000000000000110010010101001;
assign LUT_3[51222] = 32'b00000000000000000001101110110000;
assign LUT_3[51223] = 32'b00000000000000001000011010001101;
assign LUT_3[51224] = 32'b00000000000000000111110010011100;
assign LUT_3[51225] = 32'b00000000000000001110011101111001;
assign LUT_3[51226] = 32'b00000000000000001001111010000000;
assign LUT_3[51227] = 32'b00000000000000010000100101011101;
assign LUT_3[51228] = 32'b00000000000000000101000000010010;
assign LUT_3[51229] = 32'b00000000000000001011101011101111;
assign LUT_3[51230] = 32'b00000000000000000111000111110110;
assign LUT_3[51231] = 32'b00000000000000001101110011010011;
assign LUT_3[51232] = 32'b00000000000000000000010100110011;
assign LUT_3[51233] = 32'b00000000000000000111000000010000;
assign LUT_3[51234] = 32'b00000000000000000010011100010111;
assign LUT_3[51235] = 32'b00000000000000001001000111110100;
assign LUT_3[51236] = 32'b11111111111111111101100010101001;
assign LUT_3[51237] = 32'b00000000000000000100001110000110;
assign LUT_3[51238] = 32'b11111111111111111111101010001101;
assign LUT_3[51239] = 32'b00000000000000000110010101101010;
assign LUT_3[51240] = 32'b00000000000000000101101101111001;
assign LUT_3[51241] = 32'b00000000000000001100011001010110;
assign LUT_3[51242] = 32'b00000000000000000111110101011101;
assign LUT_3[51243] = 32'b00000000000000001110100000111010;
assign LUT_3[51244] = 32'b00000000000000000010111011101111;
assign LUT_3[51245] = 32'b00000000000000001001100111001100;
assign LUT_3[51246] = 32'b00000000000000000101000011010011;
assign LUT_3[51247] = 32'b00000000000000001011101110110000;
assign LUT_3[51248] = 32'b00000000000000000011100111110110;
assign LUT_3[51249] = 32'b00000000000000001010010011010011;
assign LUT_3[51250] = 32'b00000000000000000101101111011010;
assign LUT_3[51251] = 32'b00000000000000001100011010110111;
assign LUT_3[51252] = 32'b00000000000000000000110101101100;
assign LUT_3[51253] = 32'b00000000000000000111100001001001;
assign LUT_3[51254] = 32'b00000000000000000010111101010000;
assign LUT_3[51255] = 32'b00000000000000001001101000101101;
assign LUT_3[51256] = 32'b00000000000000001001000000111100;
assign LUT_3[51257] = 32'b00000000000000001111101100011001;
assign LUT_3[51258] = 32'b00000000000000001011001000100000;
assign LUT_3[51259] = 32'b00000000000000010001110011111101;
assign LUT_3[51260] = 32'b00000000000000000110001110110010;
assign LUT_3[51261] = 32'b00000000000000001100111010001111;
assign LUT_3[51262] = 32'b00000000000000001000010110010110;
assign LUT_3[51263] = 32'b00000000000000001111000001110011;
assign LUT_3[51264] = 32'b11111111111111111110111110111110;
assign LUT_3[51265] = 32'b00000000000000000101101010011011;
assign LUT_3[51266] = 32'b00000000000000000001000110100010;
assign LUT_3[51267] = 32'b00000000000000000111110001111111;
assign LUT_3[51268] = 32'b11111111111111111100001100110100;
assign LUT_3[51269] = 32'b00000000000000000010111000010001;
assign LUT_3[51270] = 32'b11111111111111111110010100011000;
assign LUT_3[51271] = 32'b00000000000000000100111111110101;
assign LUT_3[51272] = 32'b00000000000000000100011000000100;
assign LUT_3[51273] = 32'b00000000000000001011000011100001;
assign LUT_3[51274] = 32'b00000000000000000110011111101000;
assign LUT_3[51275] = 32'b00000000000000001101001011000101;
assign LUT_3[51276] = 32'b00000000000000000001100101111010;
assign LUT_3[51277] = 32'b00000000000000001000010001010111;
assign LUT_3[51278] = 32'b00000000000000000011101101011110;
assign LUT_3[51279] = 32'b00000000000000001010011000111011;
assign LUT_3[51280] = 32'b00000000000000000010010010000001;
assign LUT_3[51281] = 32'b00000000000000001000111101011110;
assign LUT_3[51282] = 32'b00000000000000000100011001100101;
assign LUT_3[51283] = 32'b00000000000000001011000101000010;
assign LUT_3[51284] = 32'b11111111111111111111011111110111;
assign LUT_3[51285] = 32'b00000000000000000110001011010100;
assign LUT_3[51286] = 32'b00000000000000000001100111011011;
assign LUT_3[51287] = 32'b00000000000000001000010010111000;
assign LUT_3[51288] = 32'b00000000000000000111101011000111;
assign LUT_3[51289] = 32'b00000000000000001110010110100100;
assign LUT_3[51290] = 32'b00000000000000001001110010101011;
assign LUT_3[51291] = 32'b00000000000000010000011110001000;
assign LUT_3[51292] = 32'b00000000000000000100111000111101;
assign LUT_3[51293] = 32'b00000000000000001011100100011010;
assign LUT_3[51294] = 32'b00000000000000000111000000100001;
assign LUT_3[51295] = 32'b00000000000000001101101011111110;
assign LUT_3[51296] = 32'b00000000000000000000001101011110;
assign LUT_3[51297] = 32'b00000000000000000110111000111011;
assign LUT_3[51298] = 32'b00000000000000000010010101000010;
assign LUT_3[51299] = 32'b00000000000000001001000000011111;
assign LUT_3[51300] = 32'b11111111111111111101011011010100;
assign LUT_3[51301] = 32'b00000000000000000100000110110001;
assign LUT_3[51302] = 32'b11111111111111111111100010111000;
assign LUT_3[51303] = 32'b00000000000000000110001110010101;
assign LUT_3[51304] = 32'b00000000000000000101100110100100;
assign LUT_3[51305] = 32'b00000000000000001100010010000001;
assign LUT_3[51306] = 32'b00000000000000000111101110001000;
assign LUT_3[51307] = 32'b00000000000000001110011001100101;
assign LUT_3[51308] = 32'b00000000000000000010110100011010;
assign LUT_3[51309] = 32'b00000000000000001001011111110111;
assign LUT_3[51310] = 32'b00000000000000000100111011111110;
assign LUT_3[51311] = 32'b00000000000000001011100111011011;
assign LUT_3[51312] = 32'b00000000000000000011100000100001;
assign LUT_3[51313] = 32'b00000000000000001010001011111110;
assign LUT_3[51314] = 32'b00000000000000000101101000000101;
assign LUT_3[51315] = 32'b00000000000000001100010011100010;
assign LUT_3[51316] = 32'b00000000000000000000101110010111;
assign LUT_3[51317] = 32'b00000000000000000111011001110100;
assign LUT_3[51318] = 32'b00000000000000000010110101111011;
assign LUT_3[51319] = 32'b00000000000000001001100001011000;
assign LUT_3[51320] = 32'b00000000000000001000111001100111;
assign LUT_3[51321] = 32'b00000000000000001111100101000100;
assign LUT_3[51322] = 32'b00000000000000001011000001001011;
assign LUT_3[51323] = 32'b00000000000000010001101100101000;
assign LUT_3[51324] = 32'b00000000000000000110000111011101;
assign LUT_3[51325] = 32'b00000000000000001100110010111010;
assign LUT_3[51326] = 32'b00000000000000001000001111000001;
assign LUT_3[51327] = 32'b00000000000000001110111010011110;
assign LUT_3[51328] = 32'b00000000000000000001010001010001;
assign LUT_3[51329] = 32'b00000000000000000111111100101110;
assign LUT_3[51330] = 32'b00000000000000000011011000110101;
assign LUT_3[51331] = 32'b00000000000000001010000100010010;
assign LUT_3[51332] = 32'b11111111111111111110011111000111;
assign LUT_3[51333] = 32'b00000000000000000101001010100100;
assign LUT_3[51334] = 32'b00000000000000000000100110101011;
assign LUT_3[51335] = 32'b00000000000000000111010010001000;
assign LUT_3[51336] = 32'b00000000000000000110101010010111;
assign LUT_3[51337] = 32'b00000000000000001101010101110100;
assign LUT_3[51338] = 32'b00000000000000001000110001111011;
assign LUT_3[51339] = 32'b00000000000000001111011101011000;
assign LUT_3[51340] = 32'b00000000000000000011111000001101;
assign LUT_3[51341] = 32'b00000000000000001010100011101010;
assign LUT_3[51342] = 32'b00000000000000000101111111110001;
assign LUT_3[51343] = 32'b00000000000000001100101011001110;
assign LUT_3[51344] = 32'b00000000000000000100100100010100;
assign LUT_3[51345] = 32'b00000000000000001011001111110001;
assign LUT_3[51346] = 32'b00000000000000000110101011111000;
assign LUT_3[51347] = 32'b00000000000000001101010111010101;
assign LUT_3[51348] = 32'b00000000000000000001110010001010;
assign LUT_3[51349] = 32'b00000000000000001000011101100111;
assign LUT_3[51350] = 32'b00000000000000000011111001101110;
assign LUT_3[51351] = 32'b00000000000000001010100101001011;
assign LUT_3[51352] = 32'b00000000000000001001111101011010;
assign LUT_3[51353] = 32'b00000000000000010000101000110111;
assign LUT_3[51354] = 32'b00000000000000001100000100111110;
assign LUT_3[51355] = 32'b00000000000000010010110000011011;
assign LUT_3[51356] = 32'b00000000000000000111001011010000;
assign LUT_3[51357] = 32'b00000000000000001101110110101101;
assign LUT_3[51358] = 32'b00000000000000001001010010110100;
assign LUT_3[51359] = 32'b00000000000000001111111110010001;
assign LUT_3[51360] = 32'b00000000000000000010011111110001;
assign LUT_3[51361] = 32'b00000000000000001001001011001110;
assign LUT_3[51362] = 32'b00000000000000000100100111010101;
assign LUT_3[51363] = 32'b00000000000000001011010010110010;
assign LUT_3[51364] = 32'b11111111111111111111101101100111;
assign LUT_3[51365] = 32'b00000000000000000110011001000100;
assign LUT_3[51366] = 32'b00000000000000000001110101001011;
assign LUT_3[51367] = 32'b00000000000000001000100000101000;
assign LUT_3[51368] = 32'b00000000000000000111111000110111;
assign LUT_3[51369] = 32'b00000000000000001110100100010100;
assign LUT_3[51370] = 32'b00000000000000001010000000011011;
assign LUT_3[51371] = 32'b00000000000000010000101011111000;
assign LUT_3[51372] = 32'b00000000000000000101000110101101;
assign LUT_3[51373] = 32'b00000000000000001011110010001010;
assign LUT_3[51374] = 32'b00000000000000000111001110010001;
assign LUT_3[51375] = 32'b00000000000000001101111001101110;
assign LUT_3[51376] = 32'b00000000000000000101110010110100;
assign LUT_3[51377] = 32'b00000000000000001100011110010001;
assign LUT_3[51378] = 32'b00000000000000000111111010011000;
assign LUT_3[51379] = 32'b00000000000000001110100101110101;
assign LUT_3[51380] = 32'b00000000000000000011000000101010;
assign LUT_3[51381] = 32'b00000000000000001001101100000111;
assign LUT_3[51382] = 32'b00000000000000000101001000001110;
assign LUT_3[51383] = 32'b00000000000000001011110011101011;
assign LUT_3[51384] = 32'b00000000000000001011001011111010;
assign LUT_3[51385] = 32'b00000000000000010001110111010111;
assign LUT_3[51386] = 32'b00000000000000001101010011011110;
assign LUT_3[51387] = 32'b00000000000000010011111110111011;
assign LUT_3[51388] = 32'b00000000000000001000011001110000;
assign LUT_3[51389] = 32'b00000000000000001111000101001101;
assign LUT_3[51390] = 32'b00000000000000001010100001010100;
assign LUT_3[51391] = 32'b00000000000000010001001100110001;
assign LUT_3[51392] = 32'b00000000000000000001001001111100;
assign LUT_3[51393] = 32'b00000000000000000111110101011001;
assign LUT_3[51394] = 32'b00000000000000000011010001100000;
assign LUT_3[51395] = 32'b00000000000000001001111100111101;
assign LUT_3[51396] = 32'b11111111111111111110010111110010;
assign LUT_3[51397] = 32'b00000000000000000101000011001111;
assign LUT_3[51398] = 32'b00000000000000000000011111010110;
assign LUT_3[51399] = 32'b00000000000000000111001010110011;
assign LUT_3[51400] = 32'b00000000000000000110100011000010;
assign LUT_3[51401] = 32'b00000000000000001101001110011111;
assign LUT_3[51402] = 32'b00000000000000001000101010100110;
assign LUT_3[51403] = 32'b00000000000000001111010110000011;
assign LUT_3[51404] = 32'b00000000000000000011110000111000;
assign LUT_3[51405] = 32'b00000000000000001010011100010101;
assign LUT_3[51406] = 32'b00000000000000000101111000011100;
assign LUT_3[51407] = 32'b00000000000000001100100011111001;
assign LUT_3[51408] = 32'b00000000000000000100011100111111;
assign LUT_3[51409] = 32'b00000000000000001011001000011100;
assign LUT_3[51410] = 32'b00000000000000000110100100100011;
assign LUT_3[51411] = 32'b00000000000000001101010000000000;
assign LUT_3[51412] = 32'b00000000000000000001101010110101;
assign LUT_3[51413] = 32'b00000000000000001000010110010010;
assign LUT_3[51414] = 32'b00000000000000000011110010011001;
assign LUT_3[51415] = 32'b00000000000000001010011101110110;
assign LUT_3[51416] = 32'b00000000000000001001110110000101;
assign LUT_3[51417] = 32'b00000000000000010000100001100010;
assign LUT_3[51418] = 32'b00000000000000001011111101101001;
assign LUT_3[51419] = 32'b00000000000000010010101001000110;
assign LUT_3[51420] = 32'b00000000000000000111000011111011;
assign LUT_3[51421] = 32'b00000000000000001101101111011000;
assign LUT_3[51422] = 32'b00000000000000001001001011011111;
assign LUT_3[51423] = 32'b00000000000000001111110110111100;
assign LUT_3[51424] = 32'b00000000000000000010011000011100;
assign LUT_3[51425] = 32'b00000000000000001001000011111001;
assign LUT_3[51426] = 32'b00000000000000000100100000000000;
assign LUT_3[51427] = 32'b00000000000000001011001011011101;
assign LUT_3[51428] = 32'b11111111111111111111100110010010;
assign LUT_3[51429] = 32'b00000000000000000110010001101111;
assign LUT_3[51430] = 32'b00000000000000000001101101110110;
assign LUT_3[51431] = 32'b00000000000000001000011001010011;
assign LUT_3[51432] = 32'b00000000000000000111110001100010;
assign LUT_3[51433] = 32'b00000000000000001110011100111111;
assign LUT_3[51434] = 32'b00000000000000001001111001000110;
assign LUT_3[51435] = 32'b00000000000000010000100100100011;
assign LUT_3[51436] = 32'b00000000000000000100111111011000;
assign LUT_3[51437] = 32'b00000000000000001011101010110101;
assign LUT_3[51438] = 32'b00000000000000000111000110111100;
assign LUT_3[51439] = 32'b00000000000000001101110010011001;
assign LUT_3[51440] = 32'b00000000000000000101101011011111;
assign LUT_3[51441] = 32'b00000000000000001100010110111100;
assign LUT_3[51442] = 32'b00000000000000000111110011000011;
assign LUT_3[51443] = 32'b00000000000000001110011110100000;
assign LUT_3[51444] = 32'b00000000000000000010111001010101;
assign LUT_3[51445] = 32'b00000000000000001001100100110010;
assign LUT_3[51446] = 32'b00000000000000000101000000111001;
assign LUT_3[51447] = 32'b00000000000000001011101100010110;
assign LUT_3[51448] = 32'b00000000000000001011000100100101;
assign LUT_3[51449] = 32'b00000000000000010001110000000010;
assign LUT_3[51450] = 32'b00000000000000001101001100001001;
assign LUT_3[51451] = 32'b00000000000000010011110111100110;
assign LUT_3[51452] = 32'b00000000000000001000010010011011;
assign LUT_3[51453] = 32'b00000000000000001110111101111000;
assign LUT_3[51454] = 32'b00000000000000001010011001111111;
assign LUT_3[51455] = 32'b00000000000000010001000101011100;
assign LUT_3[51456] = 32'b11111111111111111011010101110100;
assign LUT_3[51457] = 32'b00000000000000000010000001010001;
assign LUT_3[51458] = 32'b11111111111111111101011101011000;
assign LUT_3[51459] = 32'b00000000000000000100001000110101;
assign LUT_3[51460] = 32'b11111111111111111000100011101010;
assign LUT_3[51461] = 32'b11111111111111111111001111000111;
assign LUT_3[51462] = 32'b11111111111111111010101011001110;
assign LUT_3[51463] = 32'b00000000000000000001010110101011;
assign LUT_3[51464] = 32'b00000000000000000000101110111010;
assign LUT_3[51465] = 32'b00000000000000000111011010010111;
assign LUT_3[51466] = 32'b00000000000000000010110110011110;
assign LUT_3[51467] = 32'b00000000000000001001100001111011;
assign LUT_3[51468] = 32'b11111111111111111101111100110000;
assign LUT_3[51469] = 32'b00000000000000000100101000001101;
assign LUT_3[51470] = 32'b00000000000000000000000100010100;
assign LUT_3[51471] = 32'b00000000000000000110101111110001;
assign LUT_3[51472] = 32'b11111111111111111110101000110111;
assign LUT_3[51473] = 32'b00000000000000000101010100010100;
assign LUT_3[51474] = 32'b00000000000000000000110000011011;
assign LUT_3[51475] = 32'b00000000000000000111011011111000;
assign LUT_3[51476] = 32'b11111111111111111011110110101101;
assign LUT_3[51477] = 32'b00000000000000000010100010001010;
assign LUT_3[51478] = 32'b11111111111111111101111110010001;
assign LUT_3[51479] = 32'b00000000000000000100101001101110;
assign LUT_3[51480] = 32'b00000000000000000100000001111101;
assign LUT_3[51481] = 32'b00000000000000001010101101011010;
assign LUT_3[51482] = 32'b00000000000000000110001001100001;
assign LUT_3[51483] = 32'b00000000000000001100110100111110;
assign LUT_3[51484] = 32'b00000000000000000001001111110011;
assign LUT_3[51485] = 32'b00000000000000000111111011010000;
assign LUT_3[51486] = 32'b00000000000000000011010111010111;
assign LUT_3[51487] = 32'b00000000000000001010000010110100;
assign LUT_3[51488] = 32'b11111111111111111100100100010100;
assign LUT_3[51489] = 32'b00000000000000000011001111110001;
assign LUT_3[51490] = 32'b11111111111111111110101011111000;
assign LUT_3[51491] = 32'b00000000000000000101010111010101;
assign LUT_3[51492] = 32'b11111111111111111001110010001010;
assign LUT_3[51493] = 32'b00000000000000000000011101100111;
assign LUT_3[51494] = 32'b11111111111111111011111001101110;
assign LUT_3[51495] = 32'b00000000000000000010100101001011;
assign LUT_3[51496] = 32'b00000000000000000001111101011010;
assign LUT_3[51497] = 32'b00000000000000001000101000110111;
assign LUT_3[51498] = 32'b00000000000000000100000100111110;
assign LUT_3[51499] = 32'b00000000000000001010110000011011;
assign LUT_3[51500] = 32'b11111111111111111111001011010000;
assign LUT_3[51501] = 32'b00000000000000000101110110101101;
assign LUT_3[51502] = 32'b00000000000000000001010010110100;
assign LUT_3[51503] = 32'b00000000000000000111111110010001;
assign LUT_3[51504] = 32'b11111111111111111111110111010111;
assign LUT_3[51505] = 32'b00000000000000000110100010110100;
assign LUT_3[51506] = 32'b00000000000000000001111110111011;
assign LUT_3[51507] = 32'b00000000000000001000101010011000;
assign LUT_3[51508] = 32'b11111111111111111101000101001101;
assign LUT_3[51509] = 32'b00000000000000000011110000101010;
assign LUT_3[51510] = 32'b11111111111111111111001100110001;
assign LUT_3[51511] = 32'b00000000000000000101111000001110;
assign LUT_3[51512] = 32'b00000000000000000101010000011101;
assign LUT_3[51513] = 32'b00000000000000001011111011111010;
assign LUT_3[51514] = 32'b00000000000000000111011000000001;
assign LUT_3[51515] = 32'b00000000000000001110000011011110;
assign LUT_3[51516] = 32'b00000000000000000010011110010011;
assign LUT_3[51517] = 32'b00000000000000001001001001110000;
assign LUT_3[51518] = 32'b00000000000000000100100101110111;
assign LUT_3[51519] = 32'b00000000000000001011010001010100;
assign LUT_3[51520] = 32'b11111111111111111011001110011111;
assign LUT_3[51521] = 32'b00000000000000000001111001111100;
assign LUT_3[51522] = 32'b11111111111111111101010110000011;
assign LUT_3[51523] = 32'b00000000000000000100000001100000;
assign LUT_3[51524] = 32'b11111111111111111000011100010101;
assign LUT_3[51525] = 32'b11111111111111111111000111110010;
assign LUT_3[51526] = 32'b11111111111111111010100011111001;
assign LUT_3[51527] = 32'b00000000000000000001001111010110;
assign LUT_3[51528] = 32'b00000000000000000000100111100101;
assign LUT_3[51529] = 32'b00000000000000000111010011000010;
assign LUT_3[51530] = 32'b00000000000000000010101111001001;
assign LUT_3[51531] = 32'b00000000000000001001011010100110;
assign LUT_3[51532] = 32'b11111111111111111101110101011011;
assign LUT_3[51533] = 32'b00000000000000000100100000111000;
assign LUT_3[51534] = 32'b11111111111111111111111100111111;
assign LUT_3[51535] = 32'b00000000000000000110101000011100;
assign LUT_3[51536] = 32'b11111111111111111110100001100010;
assign LUT_3[51537] = 32'b00000000000000000101001100111111;
assign LUT_3[51538] = 32'b00000000000000000000101001000110;
assign LUT_3[51539] = 32'b00000000000000000111010100100011;
assign LUT_3[51540] = 32'b11111111111111111011101111011000;
assign LUT_3[51541] = 32'b00000000000000000010011010110101;
assign LUT_3[51542] = 32'b11111111111111111101110110111100;
assign LUT_3[51543] = 32'b00000000000000000100100010011001;
assign LUT_3[51544] = 32'b00000000000000000011111010101000;
assign LUT_3[51545] = 32'b00000000000000001010100110000101;
assign LUT_3[51546] = 32'b00000000000000000110000010001100;
assign LUT_3[51547] = 32'b00000000000000001100101101101001;
assign LUT_3[51548] = 32'b00000000000000000001001000011110;
assign LUT_3[51549] = 32'b00000000000000000111110011111011;
assign LUT_3[51550] = 32'b00000000000000000011010000000010;
assign LUT_3[51551] = 32'b00000000000000001001111011011111;
assign LUT_3[51552] = 32'b11111111111111111100011100111111;
assign LUT_3[51553] = 32'b00000000000000000011001000011100;
assign LUT_3[51554] = 32'b11111111111111111110100100100011;
assign LUT_3[51555] = 32'b00000000000000000101010000000000;
assign LUT_3[51556] = 32'b11111111111111111001101010110101;
assign LUT_3[51557] = 32'b00000000000000000000010110010010;
assign LUT_3[51558] = 32'b11111111111111111011110010011001;
assign LUT_3[51559] = 32'b00000000000000000010011101110110;
assign LUT_3[51560] = 32'b00000000000000000001110110000101;
assign LUT_3[51561] = 32'b00000000000000001000100001100010;
assign LUT_3[51562] = 32'b00000000000000000011111101101001;
assign LUT_3[51563] = 32'b00000000000000001010101001000110;
assign LUT_3[51564] = 32'b11111111111111111111000011111011;
assign LUT_3[51565] = 32'b00000000000000000101101111011000;
assign LUT_3[51566] = 32'b00000000000000000001001011011111;
assign LUT_3[51567] = 32'b00000000000000000111110110111100;
assign LUT_3[51568] = 32'b11111111111111111111110000000010;
assign LUT_3[51569] = 32'b00000000000000000110011011011111;
assign LUT_3[51570] = 32'b00000000000000000001110111100110;
assign LUT_3[51571] = 32'b00000000000000001000100011000011;
assign LUT_3[51572] = 32'b11111111111111111100111101111000;
assign LUT_3[51573] = 32'b00000000000000000011101001010101;
assign LUT_3[51574] = 32'b11111111111111111111000101011100;
assign LUT_3[51575] = 32'b00000000000000000101110000111001;
assign LUT_3[51576] = 32'b00000000000000000101001001001000;
assign LUT_3[51577] = 32'b00000000000000001011110100100101;
assign LUT_3[51578] = 32'b00000000000000000111010000101100;
assign LUT_3[51579] = 32'b00000000000000001101111100001001;
assign LUT_3[51580] = 32'b00000000000000000010010110111110;
assign LUT_3[51581] = 32'b00000000000000001001000010011011;
assign LUT_3[51582] = 32'b00000000000000000100011110100010;
assign LUT_3[51583] = 32'b00000000000000001011001001111111;
assign LUT_3[51584] = 32'b11111111111111111101100000110010;
assign LUT_3[51585] = 32'b00000000000000000100001100001111;
assign LUT_3[51586] = 32'b11111111111111111111101000010110;
assign LUT_3[51587] = 32'b00000000000000000110010011110011;
assign LUT_3[51588] = 32'b11111111111111111010101110101000;
assign LUT_3[51589] = 32'b00000000000000000001011010000101;
assign LUT_3[51590] = 32'b11111111111111111100110110001100;
assign LUT_3[51591] = 32'b00000000000000000011100001101001;
assign LUT_3[51592] = 32'b00000000000000000010111001111000;
assign LUT_3[51593] = 32'b00000000000000001001100101010101;
assign LUT_3[51594] = 32'b00000000000000000101000001011100;
assign LUT_3[51595] = 32'b00000000000000001011101100111001;
assign LUT_3[51596] = 32'b00000000000000000000000111101110;
assign LUT_3[51597] = 32'b00000000000000000110110011001011;
assign LUT_3[51598] = 32'b00000000000000000010001111010010;
assign LUT_3[51599] = 32'b00000000000000001000111010101111;
assign LUT_3[51600] = 32'b00000000000000000000110011110101;
assign LUT_3[51601] = 32'b00000000000000000111011111010010;
assign LUT_3[51602] = 32'b00000000000000000010111011011001;
assign LUT_3[51603] = 32'b00000000000000001001100110110110;
assign LUT_3[51604] = 32'b11111111111111111110000001101011;
assign LUT_3[51605] = 32'b00000000000000000100101101001000;
assign LUT_3[51606] = 32'b00000000000000000000001001001111;
assign LUT_3[51607] = 32'b00000000000000000110110100101100;
assign LUT_3[51608] = 32'b00000000000000000110001100111011;
assign LUT_3[51609] = 32'b00000000000000001100111000011000;
assign LUT_3[51610] = 32'b00000000000000001000010100011111;
assign LUT_3[51611] = 32'b00000000000000001110111111111100;
assign LUT_3[51612] = 32'b00000000000000000011011010110001;
assign LUT_3[51613] = 32'b00000000000000001010000110001110;
assign LUT_3[51614] = 32'b00000000000000000101100010010101;
assign LUT_3[51615] = 32'b00000000000000001100001101110010;
assign LUT_3[51616] = 32'b11111111111111111110101111010010;
assign LUT_3[51617] = 32'b00000000000000000101011010101111;
assign LUT_3[51618] = 32'b00000000000000000000110110110110;
assign LUT_3[51619] = 32'b00000000000000000111100010010011;
assign LUT_3[51620] = 32'b11111111111111111011111101001000;
assign LUT_3[51621] = 32'b00000000000000000010101000100101;
assign LUT_3[51622] = 32'b11111111111111111110000100101100;
assign LUT_3[51623] = 32'b00000000000000000100110000001001;
assign LUT_3[51624] = 32'b00000000000000000100001000011000;
assign LUT_3[51625] = 32'b00000000000000001010110011110101;
assign LUT_3[51626] = 32'b00000000000000000110001111111100;
assign LUT_3[51627] = 32'b00000000000000001100111011011001;
assign LUT_3[51628] = 32'b00000000000000000001010110001110;
assign LUT_3[51629] = 32'b00000000000000001000000001101011;
assign LUT_3[51630] = 32'b00000000000000000011011101110010;
assign LUT_3[51631] = 32'b00000000000000001010001001001111;
assign LUT_3[51632] = 32'b00000000000000000010000010010101;
assign LUT_3[51633] = 32'b00000000000000001000101101110010;
assign LUT_3[51634] = 32'b00000000000000000100001001111001;
assign LUT_3[51635] = 32'b00000000000000001010110101010110;
assign LUT_3[51636] = 32'b11111111111111111111010000001011;
assign LUT_3[51637] = 32'b00000000000000000101111011101000;
assign LUT_3[51638] = 32'b00000000000000000001010111101111;
assign LUT_3[51639] = 32'b00000000000000001000000011001100;
assign LUT_3[51640] = 32'b00000000000000000111011011011011;
assign LUT_3[51641] = 32'b00000000000000001110000110111000;
assign LUT_3[51642] = 32'b00000000000000001001100010111111;
assign LUT_3[51643] = 32'b00000000000000010000001110011100;
assign LUT_3[51644] = 32'b00000000000000000100101001010001;
assign LUT_3[51645] = 32'b00000000000000001011010100101110;
assign LUT_3[51646] = 32'b00000000000000000110110000110101;
assign LUT_3[51647] = 32'b00000000000000001101011100010010;
assign LUT_3[51648] = 32'b11111111111111111101011001011101;
assign LUT_3[51649] = 32'b00000000000000000100000100111010;
assign LUT_3[51650] = 32'b11111111111111111111100001000001;
assign LUT_3[51651] = 32'b00000000000000000110001100011110;
assign LUT_3[51652] = 32'b11111111111111111010100111010011;
assign LUT_3[51653] = 32'b00000000000000000001010010110000;
assign LUT_3[51654] = 32'b11111111111111111100101110110111;
assign LUT_3[51655] = 32'b00000000000000000011011010010100;
assign LUT_3[51656] = 32'b00000000000000000010110010100011;
assign LUT_3[51657] = 32'b00000000000000001001011110000000;
assign LUT_3[51658] = 32'b00000000000000000100111010000111;
assign LUT_3[51659] = 32'b00000000000000001011100101100100;
assign LUT_3[51660] = 32'b00000000000000000000000000011001;
assign LUT_3[51661] = 32'b00000000000000000110101011110110;
assign LUT_3[51662] = 32'b00000000000000000010000111111101;
assign LUT_3[51663] = 32'b00000000000000001000110011011010;
assign LUT_3[51664] = 32'b00000000000000000000101100100000;
assign LUT_3[51665] = 32'b00000000000000000111010111111101;
assign LUT_3[51666] = 32'b00000000000000000010110100000100;
assign LUT_3[51667] = 32'b00000000000000001001011111100001;
assign LUT_3[51668] = 32'b11111111111111111101111010010110;
assign LUT_3[51669] = 32'b00000000000000000100100101110011;
assign LUT_3[51670] = 32'b00000000000000000000000001111010;
assign LUT_3[51671] = 32'b00000000000000000110101101010111;
assign LUT_3[51672] = 32'b00000000000000000110000101100110;
assign LUT_3[51673] = 32'b00000000000000001100110001000011;
assign LUT_3[51674] = 32'b00000000000000001000001101001010;
assign LUT_3[51675] = 32'b00000000000000001110111000100111;
assign LUT_3[51676] = 32'b00000000000000000011010011011100;
assign LUT_3[51677] = 32'b00000000000000001001111110111001;
assign LUT_3[51678] = 32'b00000000000000000101011011000000;
assign LUT_3[51679] = 32'b00000000000000001100000110011101;
assign LUT_3[51680] = 32'b11111111111111111110100111111101;
assign LUT_3[51681] = 32'b00000000000000000101010011011010;
assign LUT_3[51682] = 32'b00000000000000000000101111100001;
assign LUT_3[51683] = 32'b00000000000000000111011010111110;
assign LUT_3[51684] = 32'b11111111111111111011110101110011;
assign LUT_3[51685] = 32'b00000000000000000010100001010000;
assign LUT_3[51686] = 32'b11111111111111111101111101010111;
assign LUT_3[51687] = 32'b00000000000000000100101000110100;
assign LUT_3[51688] = 32'b00000000000000000100000001000011;
assign LUT_3[51689] = 32'b00000000000000001010101100100000;
assign LUT_3[51690] = 32'b00000000000000000110001000100111;
assign LUT_3[51691] = 32'b00000000000000001100110100000100;
assign LUT_3[51692] = 32'b00000000000000000001001110111001;
assign LUT_3[51693] = 32'b00000000000000000111111010010110;
assign LUT_3[51694] = 32'b00000000000000000011010110011101;
assign LUT_3[51695] = 32'b00000000000000001010000001111010;
assign LUT_3[51696] = 32'b00000000000000000001111011000000;
assign LUT_3[51697] = 32'b00000000000000001000100110011101;
assign LUT_3[51698] = 32'b00000000000000000100000010100100;
assign LUT_3[51699] = 32'b00000000000000001010101110000001;
assign LUT_3[51700] = 32'b11111111111111111111001000110110;
assign LUT_3[51701] = 32'b00000000000000000101110100010011;
assign LUT_3[51702] = 32'b00000000000000000001010000011010;
assign LUT_3[51703] = 32'b00000000000000000111111011110111;
assign LUT_3[51704] = 32'b00000000000000000111010100000110;
assign LUT_3[51705] = 32'b00000000000000001101111111100011;
assign LUT_3[51706] = 32'b00000000000000001001011011101010;
assign LUT_3[51707] = 32'b00000000000000010000000111000111;
assign LUT_3[51708] = 32'b00000000000000000100100001111100;
assign LUT_3[51709] = 32'b00000000000000001011001101011001;
assign LUT_3[51710] = 32'b00000000000000000110101001100000;
assign LUT_3[51711] = 32'b00000000000000001101010100111101;
assign LUT_3[51712] = 32'b00000000000000000010011011011111;
assign LUT_3[51713] = 32'b00000000000000001001000110111100;
assign LUT_3[51714] = 32'b00000000000000000100100011000011;
assign LUT_3[51715] = 32'b00000000000000001011001110100000;
assign LUT_3[51716] = 32'b11111111111111111111101001010101;
assign LUT_3[51717] = 32'b00000000000000000110010100110010;
assign LUT_3[51718] = 32'b00000000000000000001110000111001;
assign LUT_3[51719] = 32'b00000000000000001000011100010110;
assign LUT_3[51720] = 32'b00000000000000000111110100100101;
assign LUT_3[51721] = 32'b00000000000000001110100000000010;
assign LUT_3[51722] = 32'b00000000000000001001111100001001;
assign LUT_3[51723] = 32'b00000000000000010000100111100110;
assign LUT_3[51724] = 32'b00000000000000000101000010011011;
assign LUT_3[51725] = 32'b00000000000000001011101101111000;
assign LUT_3[51726] = 32'b00000000000000000111001001111111;
assign LUT_3[51727] = 32'b00000000000000001101110101011100;
assign LUT_3[51728] = 32'b00000000000000000101101110100010;
assign LUT_3[51729] = 32'b00000000000000001100011001111111;
assign LUT_3[51730] = 32'b00000000000000000111110110000110;
assign LUT_3[51731] = 32'b00000000000000001110100001100011;
assign LUT_3[51732] = 32'b00000000000000000010111100011000;
assign LUT_3[51733] = 32'b00000000000000001001100111110101;
assign LUT_3[51734] = 32'b00000000000000000101000011111100;
assign LUT_3[51735] = 32'b00000000000000001011101111011001;
assign LUT_3[51736] = 32'b00000000000000001011000111101000;
assign LUT_3[51737] = 32'b00000000000000010001110011000101;
assign LUT_3[51738] = 32'b00000000000000001101001111001100;
assign LUT_3[51739] = 32'b00000000000000010011111010101001;
assign LUT_3[51740] = 32'b00000000000000001000010101011110;
assign LUT_3[51741] = 32'b00000000000000001111000000111011;
assign LUT_3[51742] = 32'b00000000000000001010011101000010;
assign LUT_3[51743] = 32'b00000000000000010001001000011111;
assign LUT_3[51744] = 32'b00000000000000000011101001111111;
assign LUT_3[51745] = 32'b00000000000000001010010101011100;
assign LUT_3[51746] = 32'b00000000000000000101110001100011;
assign LUT_3[51747] = 32'b00000000000000001100011101000000;
assign LUT_3[51748] = 32'b00000000000000000000110111110101;
assign LUT_3[51749] = 32'b00000000000000000111100011010010;
assign LUT_3[51750] = 32'b00000000000000000010111111011001;
assign LUT_3[51751] = 32'b00000000000000001001101010110110;
assign LUT_3[51752] = 32'b00000000000000001001000011000101;
assign LUT_3[51753] = 32'b00000000000000001111101110100010;
assign LUT_3[51754] = 32'b00000000000000001011001010101001;
assign LUT_3[51755] = 32'b00000000000000010001110110000110;
assign LUT_3[51756] = 32'b00000000000000000110010000111011;
assign LUT_3[51757] = 32'b00000000000000001100111100011000;
assign LUT_3[51758] = 32'b00000000000000001000011000011111;
assign LUT_3[51759] = 32'b00000000000000001111000011111100;
assign LUT_3[51760] = 32'b00000000000000000110111101000010;
assign LUT_3[51761] = 32'b00000000000000001101101000011111;
assign LUT_3[51762] = 32'b00000000000000001001000100100110;
assign LUT_3[51763] = 32'b00000000000000001111110000000011;
assign LUT_3[51764] = 32'b00000000000000000100001010111000;
assign LUT_3[51765] = 32'b00000000000000001010110110010101;
assign LUT_3[51766] = 32'b00000000000000000110010010011100;
assign LUT_3[51767] = 32'b00000000000000001100111101111001;
assign LUT_3[51768] = 32'b00000000000000001100010110001000;
assign LUT_3[51769] = 32'b00000000000000010011000001100101;
assign LUT_3[51770] = 32'b00000000000000001110011101101100;
assign LUT_3[51771] = 32'b00000000000000010101001001001001;
assign LUT_3[51772] = 32'b00000000000000001001100011111110;
assign LUT_3[51773] = 32'b00000000000000010000001111011011;
assign LUT_3[51774] = 32'b00000000000000001011101011100010;
assign LUT_3[51775] = 32'b00000000000000010010010110111111;
assign LUT_3[51776] = 32'b00000000000000000010010100001010;
assign LUT_3[51777] = 32'b00000000000000001000111111100111;
assign LUT_3[51778] = 32'b00000000000000000100011011101110;
assign LUT_3[51779] = 32'b00000000000000001011000111001011;
assign LUT_3[51780] = 32'b11111111111111111111100010000000;
assign LUT_3[51781] = 32'b00000000000000000110001101011101;
assign LUT_3[51782] = 32'b00000000000000000001101001100100;
assign LUT_3[51783] = 32'b00000000000000001000010101000001;
assign LUT_3[51784] = 32'b00000000000000000111101101010000;
assign LUT_3[51785] = 32'b00000000000000001110011000101101;
assign LUT_3[51786] = 32'b00000000000000001001110100110100;
assign LUT_3[51787] = 32'b00000000000000010000100000010001;
assign LUT_3[51788] = 32'b00000000000000000100111011000110;
assign LUT_3[51789] = 32'b00000000000000001011100110100011;
assign LUT_3[51790] = 32'b00000000000000000111000010101010;
assign LUT_3[51791] = 32'b00000000000000001101101110000111;
assign LUT_3[51792] = 32'b00000000000000000101100111001101;
assign LUT_3[51793] = 32'b00000000000000001100010010101010;
assign LUT_3[51794] = 32'b00000000000000000111101110110001;
assign LUT_3[51795] = 32'b00000000000000001110011010001110;
assign LUT_3[51796] = 32'b00000000000000000010110101000011;
assign LUT_3[51797] = 32'b00000000000000001001100000100000;
assign LUT_3[51798] = 32'b00000000000000000100111100100111;
assign LUT_3[51799] = 32'b00000000000000001011101000000100;
assign LUT_3[51800] = 32'b00000000000000001011000000010011;
assign LUT_3[51801] = 32'b00000000000000010001101011110000;
assign LUT_3[51802] = 32'b00000000000000001101000111110111;
assign LUT_3[51803] = 32'b00000000000000010011110011010100;
assign LUT_3[51804] = 32'b00000000000000001000001110001001;
assign LUT_3[51805] = 32'b00000000000000001110111001100110;
assign LUT_3[51806] = 32'b00000000000000001010010101101101;
assign LUT_3[51807] = 32'b00000000000000010001000001001010;
assign LUT_3[51808] = 32'b00000000000000000011100010101010;
assign LUT_3[51809] = 32'b00000000000000001010001110000111;
assign LUT_3[51810] = 32'b00000000000000000101101010001110;
assign LUT_3[51811] = 32'b00000000000000001100010101101011;
assign LUT_3[51812] = 32'b00000000000000000000110000100000;
assign LUT_3[51813] = 32'b00000000000000000111011011111101;
assign LUT_3[51814] = 32'b00000000000000000010111000000100;
assign LUT_3[51815] = 32'b00000000000000001001100011100001;
assign LUT_3[51816] = 32'b00000000000000001000111011110000;
assign LUT_3[51817] = 32'b00000000000000001111100111001101;
assign LUT_3[51818] = 32'b00000000000000001011000011010100;
assign LUT_3[51819] = 32'b00000000000000010001101110110001;
assign LUT_3[51820] = 32'b00000000000000000110001001100110;
assign LUT_3[51821] = 32'b00000000000000001100110101000011;
assign LUT_3[51822] = 32'b00000000000000001000010001001010;
assign LUT_3[51823] = 32'b00000000000000001110111100100111;
assign LUT_3[51824] = 32'b00000000000000000110110101101101;
assign LUT_3[51825] = 32'b00000000000000001101100001001010;
assign LUT_3[51826] = 32'b00000000000000001000111101010001;
assign LUT_3[51827] = 32'b00000000000000001111101000101110;
assign LUT_3[51828] = 32'b00000000000000000100000011100011;
assign LUT_3[51829] = 32'b00000000000000001010101111000000;
assign LUT_3[51830] = 32'b00000000000000000110001011000111;
assign LUT_3[51831] = 32'b00000000000000001100110110100100;
assign LUT_3[51832] = 32'b00000000000000001100001110110011;
assign LUT_3[51833] = 32'b00000000000000010010111010010000;
assign LUT_3[51834] = 32'b00000000000000001110010110010111;
assign LUT_3[51835] = 32'b00000000000000010101000001110100;
assign LUT_3[51836] = 32'b00000000000000001001011100101001;
assign LUT_3[51837] = 32'b00000000000000010000001000000110;
assign LUT_3[51838] = 32'b00000000000000001011100100001101;
assign LUT_3[51839] = 32'b00000000000000010010001111101010;
assign LUT_3[51840] = 32'b00000000000000000100100110011101;
assign LUT_3[51841] = 32'b00000000000000001011010001111010;
assign LUT_3[51842] = 32'b00000000000000000110101110000001;
assign LUT_3[51843] = 32'b00000000000000001101011001011110;
assign LUT_3[51844] = 32'b00000000000000000001110100010011;
assign LUT_3[51845] = 32'b00000000000000001000011111110000;
assign LUT_3[51846] = 32'b00000000000000000011111011110111;
assign LUT_3[51847] = 32'b00000000000000001010100111010100;
assign LUT_3[51848] = 32'b00000000000000001001111111100011;
assign LUT_3[51849] = 32'b00000000000000010000101011000000;
assign LUT_3[51850] = 32'b00000000000000001100000111000111;
assign LUT_3[51851] = 32'b00000000000000010010110010100100;
assign LUT_3[51852] = 32'b00000000000000000111001101011001;
assign LUT_3[51853] = 32'b00000000000000001101111000110110;
assign LUT_3[51854] = 32'b00000000000000001001010100111101;
assign LUT_3[51855] = 32'b00000000000000010000000000011010;
assign LUT_3[51856] = 32'b00000000000000000111111001100000;
assign LUT_3[51857] = 32'b00000000000000001110100100111101;
assign LUT_3[51858] = 32'b00000000000000001010000001000100;
assign LUT_3[51859] = 32'b00000000000000010000101100100001;
assign LUT_3[51860] = 32'b00000000000000000101000111010110;
assign LUT_3[51861] = 32'b00000000000000001011110010110011;
assign LUT_3[51862] = 32'b00000000000000000111001110111010;
assign LUT_3[51863] = 32'b00000000000000001101111010010111;
assign LUT_3[51864] = 32'b00000000000000001101010010100110;
assign LUT_3[51865] = 32'b00000000000000010011111110000011;
assign LUT_3[51866] = 32'b00000000000000001111011010001010;
assign LUT_3[51867] = 32'b00000000000000010110000101100111;
assign LUT_3[51868] = 32'b00000000000000001010100000011100;
assign LUT_3[51869] = 32'b00000000000000010001001011111001;
assign LUT_3[51870] = 32'b00000000000000001100101000000000;
assign LUT_3[51871] = 32'b00000000000000010011010011011101;
assign LUT_3[51872] = 32'b00000000000000000101110100111101;
assign LUT_3[51873] = 32'b00000000000000001100100000011010;
assign LUT_3[51874] = 32'b00000000000000000111111100100001;
assign LUT_3[51875] = 32'b00000000000000001110100111111110;
assign LUT_3[51876] = 32'b00000000000000000011000010110011;
assign LUT_3[51877] = 32'b00000000000000001001101110010000;
assign LUT_3[51878] = 32'b00000000000000000101001010010111;
assign LUT_3[51879] = 32'b00000000000000001011110101110100;
assign LUT_3[51880] = 32'b00000000000000001011001110000011;
assign LUT_3[51881] = 32'b00000000000000010001111001100000;
assign LUT_3[51882] = 32'b00000000000000001101010101100111;
assign LUT_3[51883] = 32'b00000000000000010100000001000100;
assign LUT_3[51884] = 32'b00000000000000001000011011111001;
assign LUT_3[51885] = 32'b00000000000000001111000111010110;
assign LUT_3[51886] = 32'b00000000000000001010100011011101;
assign LUT_3[51887] = 32'b00000000000000010001001110111010;
assign LUT_3[51888] = 32'b00000000000000001001001000000000;
assign LUT_3[51889] = 32'b00000000000000001111110011011101;
assign LUT_3[51890] = 32'b00000000000000001011001111100100;
assign LUT_3[51891] = 32'b00000000000000010001111011000001;
assign LUT_3[51892] = 32'b00000000000000000110010101110110;
assign LUT_3[51893] = 32'b00000000000000001101000001010011;
assign LUT_3[51894] = 32'b00000000000000001000011101011010;
assign LUT_3[51895] = 32'b00000000000000001111001000110111;
assign LUT_3[51896] = 32'b00000000000000001110100001000110;
assign LUT_3[51897] = 32'b00000000000000010101001100100011;
assign LUT_3[51898] = 32'b00000000000000010000101000101010;
assign LUT_3[51899] = 32'b00000000000000010111010100000111;
assign LUT_3[51900] = 32'b00000000000000001011101110111100;
assign LUT_3[51901] = 32'b00000000000000010010011010011001;
assign LUT_3[51902] = 32'b00000000000000001101110110100000;
assign LUT_3[51903] = 32'b00000000000000010100100001111101;
assign LUT_3[51904] = 32'b00000000000000000100011111001000;
assign LUT_3[51905] = 32'b00000000000000001011001010100101;
assign LUT_3[51906] = 32'b00000000000000000110100110101100;
assign LUT_3[51907] = 32'b00000000000000001101010010001001;
assign LUT_3[51908] = 32'b00000000000000000001101100111110;
assign LUT_3[51909] = 32'b00000000000000001000011000011011;
assign LUT_3[51910] = 32'b00000000000000000011110100100010;
assign LUT_3[51911] = 32'b00000000000000001010011111111111;
assign LUT_3[51912] = 32'b00000000000000001001111000001110;
assign LUT_3[51913] = 32'b00000000000000010000100011101011;
assign LUT_3[51914] = 32'b00000000000000001011111111110010;
assign LUT_3[51915] = 32'b00000000000000010010101011001111;
assign LUT_3[51916] = 32'b00000000000000000111000110000100;
assign LUT_3[51917] = 32'b00000000000000001101110001100001;
assign LUT_3[51918] = 32'b00000000000000001001001101101000;
assign LUT_3[51919] = 32'b00000000000000001111111001000101;
assign LUT_3[51920] = 32'b00000000000000000111110010001011;
assign LUT_3[51921] = 32'b00000000000000001110011101101000;
assign LUT_3[51922] = 32'b00000000000000001001111001101111;
assign LUT_3[51923] = 32'b00000000000000010000100101001100;
assign LUT_3[51924] = 32'b00000000000000000101000000000001;
assign LUT_3[51925] = 32'b00000000000000001011101011011110;
assign LUT_3[51926] = 32'b00000000000000000111000111100101;
assign LUT_3[51927] = 32'b00000000000000001101110011000010;
assign LUT_3[51928] = 32'b00000000000000001101001011010001;
assign LUT_3[51929] = 32'b00000000000000010011110110101110;
assign LUT_3[51930] = 32'b00000000000000001111010010110101;
assign LUT_3[51931] = 32'b00000000000000010101111110010010;
assign LUT_3[51932] = 32'b00000000000000001010011001000111;
assign LUT_3[51933] = 32'b00000000000000010001000100100100;
assign LUT_3[51934] = 32'b00000000000000001100100000101011;
assign LUT_3[51935] = 32'b00000000000000010011001100001000;
assign LUT_3[51936] = 32'b00000000000000000101101101101000;
assign LUT_3[51937] = 32'b00000000000000001100011001000101;
assign LUT_3[51938] = 32'b00000000000000000111110101001100;
assign LUT_3[51939] = 32'b00000000000000001110100000101001;
assign LUT_3[51940] = 32'b00000000000000000010111011011110;
assign LUT_3[51941] = 32'b00000000000000001001100110111011;
assign LUT_3[51942] = 32'b00000000000000000101000011000010;
assign LUT_3[51943] = 32'b00000000000000001011101110011111;
assign LUT_3[51944] = 32'b00000000000000001011000110101110;
assign LUT_3[51945] = 32'b00000000000000010001110010001011;
assign LUT_3[51946] = 32'b00000000000000001101001110010010;
assign LUT_3[51947] = 32'b00000000000000010011111001101111;
assign LUT_3[51948] = 32'b00000000000000001000010100100100;
assign LUT_3[51949] = 32'b00000000000000001111000000000001;
assign LUT_3[51950] = 32'b00000000000000001010011100001000;
assign LUT_3[51951] = 32'b00000000000000010001000111100101;
assign LUT_3[51952] = 32'b00000000000000001001000000101011;
assign LUT_3[51953] = 32'b00000000000000001111101100001000;
assign LUT_3[51954] = 32'b00000000000000001011001000001111;
assign LUT_3[51955] = 32'b00000000000000010001110011101100;
assign LUT_3[51956] = 32'b00000000000000000110001110100001;
assign LUT_3[51957] = 32'b00000000000000001100111001111110;
assign LUT_3[51958] = 32'b00000000000000001000010110000101;
assign LUT_3[51959] = 32'b00000000000000001111000001100010;
assign LUT_3[51960] = 32'b00000000000000001110011001110001;
assign LUT_3[51961] = 32'b00000000000000010101000101001110;
assign LUT_3[51962] = 32'b00000000000000010000100001010101;
assign LUT_3[51963] = 32'b00000000000000010111001100110010;
assign LUT_3[51964] = 32'b00000000000000001011100111100111;
assign LUT_3[51965] = 32'b00000000000000010010010011000100;
assign LUT_3[51966] = 32'b00000000000000001101101111001011;
assign LUT_3[51967] = 32'b00000000000000010100011010101000;
assign LUT_3[51968] = 32'b11111111111111111110101011000000;
assign LUT_3[51969] = 32'b00000000000000000101010110011101;
assign LUT_3[51970] = 32'b00000000000000000000110010100100;
assign LUT_3[51971] = 32'b00000000000000000111011110000001;
assign LUT_3[51972] = 32'b11111111111111111011111000110110;
assign LUT_3[51973] = 32'b00000000000000000010100100010011;
assign LUT_3[51974] = 32'b11111111111111111110000000011010;
assign LUT_3[51975] = 32'b00000000000000000100101011110111;
assign LUT_3[51976] = 32'b00000000000000000100000100000110;
assign LUT_3[51977] = 32'b00000000000000001010101111100011;
assign LUT_3[51978] = 32'b00000000000000000110001011101010;
assign LUT_3[51979] = 32'b00000000000000001100110111000111;
assign LUT_3[51980] = 32'b00000000000000000001010001111100;
assign LUT_3[51981] = 32'b00000000000000000111111101011001;
assign LUT_3[51982] = 32'b00000000000000000011011001100000;
assign LUT_3[51983] = 32'b00000000000000001010000100111101;
assign LUT_3[51984] = 32'b00000000000000000001111110000011;
assign LUT_3[51985] = 32'b00000000000000001000101001100000;
assign LUT_3[51986] = 32'b00000000000000000100000101100111;
assign LUT_3[51987] = 32'b00000000000000001010110001000100;
assign LUT_3[51988] = 32'b11111111111111111111001011111001;
assign LUT_3[51989] = 32'b00000000000000000101110111010110;
assign LUT_3[51990] = 32'b00000000000000000001010011011101;
assign LUT_3[51991] = 32'b00000000000000000111111110111010;
assign LUT_3[51992] = 32'b00000000000000000111010111001001;
assign LUT_3[51993] = 32'b00000000000000001110000010100110;
assign LUT_3[51994] = 32'b00000000000000001001011110101101;
assign LUT_3[51995] = 32'b00000000000000010000001010001010;
assign LUT_3[51996] = 32'b00000000000000000100100100111111;
assign LUT_3[51997] = 32'b00000000000000001011010000011100;
assign LUT_3[51998] = 32'b00000000000000000110101100100011;
assign LUT_3[51999] = 32'b00000000000000001101011000000000;
assign LUT_3[52000] = 32'b11111111111111111111111001100000;
assign LUT_3[52001] = 32'b00000000000000000110100100111101;
assign LUT_3[52002] = 32'b00000000000000000010000001000100;
assign LUT_3[52003] = 32'b00000000000000001000101100100001;
assign LUT_3[52004] = 32'b11111111111111111101000111010110;
assign LUT_3[52005] = 32'b00000000000000000011110010110011;
assign LUT_3[52006] = 32'b11111111111111111111001110111010;
assign LUT_3[52007] = 32'b00000000000000000101111010010111;
assign LUT_3[52008] = 32'b00000000000000000101010010100110;
assign LUT_3[52009] = 32'b00000000000000001011111110000011;
assign LUT_3[52010] = 32'b00000000000000000111011010001010;
assign LUT_3[52011] = 32'b00000000000000001110000101100111;
assign LUT_3[52012] = 32'b00000000000000000010100000011100;
assign LUT_3[52013] = 32'b00000000000000001001001011111001;
assign LUT_3[52014] = 32'b00000000000000000100101000000000;
assign LUT_3[52015] = 32'b00000000000000001011010011011101;
assign LUT_3[52016] = 32'b00000000000000000011001100100011;
assign LUT_3[52017] = 32'b00000000000000001001111000000000;
assign LUT_3[52018] = 32'b00000000000000000101010100000111;
assign LUT_3[52019] = 32'b00000000000000001011111111100100;
assign LUT_3[52020] = 32'b00000000000000000000011010011001;
assign LUT_3[52021] = 32'b00000000000000000111000101110110;
assign LUT_3[52022] = 32'b00000000000000000010100001111101;
assign LUT_3[52023] = 32'b00000000000000001001001101011010;
assign LUT_3[52024] = 32'b00000000000000001000100101101001;
assign LUT_3[52025] = 32'b00000000000000001111010001000110;
assign LUT_3[52026] = 32'b00000000000000001010101101001101;
assign LUT_3[52027] = 32'b00000000000000010001011000101010;
assign LUT_3[52028] = 32'b00000000000000000101110011011111;
assign LUT_3[52029] = 32'b00000000000000001100011110111100;
assign LUT_3[52030] = 32'b00000000000000000111111011000011;
assign LUT_3[52031] = 32'b00000000000000001110100110100000;
assign LUT_3[52032] = 32'b11111111111111111110100011101011;
assign LUT_3[52033] = 32'b00000000000000000101001111001000;
assign LUT_3[52034] = 32'b00000000000000000000101011001111;
assign LUT_3[52035] = 32'b00000000000000000111010110101100;
assign LUT_3[52036] = 32'b11111111111111111011110001100001;
assign LUT_3[52037] = 32'b00000000000000000010011100111110;
assign LUT_3[52038] = 32'b11111111111111111101111001000101;
assign LUT_3[52039] = 32'b00000000000000000100100100100010;
assign LUT_3[52040] = 32'b00000000000000000011111100110001;
assign LUT_3[52041] = 32'b00000000000000001010101000001110;
assign LUT_3[52042] = 32'b00000000000000000110000100010101;
assign LUT_3[52043] = 32'b00000000000000001100101111110010;
assign LUT_3[52044] = 32'b00000000000000000001001010100111;
assign LUT_3[52045] = 32'b00000000000000000111110110000100;
assign LUT_3[52046] = 32'b00000000000000000011010010001011;
assign LUT_3[52047] = 32'b00000000000000001001111101101000;
assign LUT_3[52048] = 32'b00000000000000000001110110101110;
assign LUT_3[52049] = 32'b00000000000000001000100010001011;
assign LUT_3[52050] = 32'b00000000000000000011111110010010;
assign LUT_3[52051] = 32'b00000000000000001010101001101111;
assign LUT_3[52052] = 32'b11111111111111111111000100100100;
assign LUT_3[52053] = 32'b00000000000000000101110000000001;
assign LUT_3[52054] = 32'b00000000000000000001001100001000;
assign LUT_3[52055] = 32'b00000000000000000111110111100101;
assign LUT_3[52056] = 32'b00000000000000000111001111110100;
assign LUT_3[52057] = 32'b00000000000000001101111011010001;
assign LUT_3[52058] = 32'b00000000000000001001010111011000;
assign LUT_3[52059] = 32'b00000000000000010000000010110101;
assign LUT_3[52060] = 32'b00000000000000000100011101101010;
assign LUT_3[52061] = 32'b00000000000000001011001001000111;
assign LUT_3[52062] = 32'b00000000000000000110100101001110;
assign LUT_3[52063] = 32'b00000000000000001101010000101011;
assign LUT_3[52064] = 32'b11111111111111111111110010001011;
assign LUT_3[52065] = 32'b00000000000000000110011101101000;
assign LUT_3[52066] = 32'b00000000000000000001111001101111;
assign LUT_3[52067] = 32'b00000000000000001000100101001100;
assign LUT_3[52068] = 32'b11111111111111111101000000000001;
assign LUT_3[52069] = 32'b00000000000000000011101011011110;
assign LUT_3[52070] = 32'b11111111111111111111000111100101;
assign LUT_3[52071] = 32'b00000000000000000101110011000010;
assign LUT_3[52072] = 32'b00000000000000000101001011010001;
assign LUT_3[52073] = 32'b00000000000000001011110110101110;
assign LUT_3[52074] = 32'b00000000000000000111010010110101;
assign LUT_3[52075] = 32'b00000000000000001101111110010010;
assign LUT_3[52076] = 32'b00000000000000000010011001000111;
assign LUT_3[52077] = 32'b00000000000000001001000100100100;
assign LUT_3[52078] = 32'b00000000000000000100100000101011;
assign LUT_3[52079] = 32'b00000000000000001011001100001000;
assign LUT_3[52080] = 32'b00000000000000000011000101001110;
assign LUT_3[52081] = 32'b00000000000000001001110000101011;
assign LUT_3[52082] = 32'b00000000000000000101001100110010;
assign LUT_3[52083] = 32'b00000000000000001011111000001111;
assign LUT_3[52084] = 32'b00000000000000000000010011000100;
assign LUT_3[52085] = 32'b00000000000000000110111110100001;
assign LUT_3[52086] = 32'b00000000000000000010011010101000;
assign LUT_3[52087] = 32'b00000000000000001001000110000101;
assign LUT_3[52088] = 32'b00000000000000001000011110010100;
assign LUT_3[52089] = 32'b00000000000000001111001001110001;
assign LUT_3[52090] = 32'b00000000000000001010100101111000;
assign LUT_3[52091] = 32'b00000000000000010001010001010101;
assign LUT_3[52092] = 32'b00000000000000000101101100001010;
assign LUT_3[52093] = 32'b00000000000000001100010111100111;
assign LUT_3[52094] = 32'b00000000000000000111110011101110;
assign LUT_3[52095] = 32'b00000000000000001110011111001011;
assign LUT_3[52096] = 32'b00000000000000000000110101111110;
assign LUT_3[52097] = 32'b00000000000000000111100001011011;
assign LUT_3[52098] = 32'b00000000000000000010111101100010;
assign LUT_3[52099] = 32'b00000000000000001001101000111111;
assign LUT_3[52100] = 32'b11111111111111111110000011110100;
assign LUT_3[52101] = 32'b00000000000000000100101111010001;
assign LUT_3[52102] = 32'b00000000000000000000001011011000;
assign LUT_3[52103] = 32'b00000000000000000110110110110101;
assign LUT_3[52104] = 32'b00000000000000000110001111000100;
assign LUT_3[52105] = 32'b00000000000000001100111010100001;
assign LUT_3[52106] = 32'b00000000000000001000010110101000;
assign LUT_3[52107] = 32'b00000000000000001111000010000101;
assign LUT_3[52108] = 32'b00000000000000000011011100111010;
assign LUT_3[52109] = 32'b00000000000000001010001000010111;
assign LUT_3[52110] = 32'b00000000000000000101100100011110;
assign LUT_3[52111] = 32'b00000000000000001100001111111011;
assign LUT_3[52112] = 32'b00000000000000000100001001000001;
assign LUT_3[52113] = 32'b00000000000000001010110100011110;
assign LUT_3[52114] = 32'b00000000000000000110010000100101;
assign LUT_3[52115] = 32'b00000000000000001100111100000010;
assign LUT_3[52116] = 32'b00000000000000000001010110110111;
assign LUT_3[52117] = 32'b00000000000000001000000010010100;
assign LUT_3[52118] = 32'b00000000000000000011011110011011;
assign LUT_3[52119] = 32'b00000000000000001010001001111000;
assign LUT_3[52120] = 32'b00000000000000001001100010000111;
assign LUT_3[52121] = 32'b00000000000000010000001101100100;
assign LUT_3[52122] = 32'b00000000000000001011101001101011;
assign LUT_3[52123] = 32'b00000000000000010010010101001000;
assign LUT_3[52124] = 32'b00000000000000000110101111111101;
assign LUT_3[52125] = 32'b00000000000000001101011011011010;
assign LUT_3[52126] = 32'b00000000000000001000110111100001;
assign LUT_3[52127] = 32'b00000000000000001111100010111110;
assign LUT_3[52128] = 32'b00000000000000000010000100011110;
assign LUT_3[52129] = 32'b00000000000000001000101111111011;
assign LUT_3[52130] = 32'b00000000000000000100001100000010;
assign LUT_3[52131] = 32'b00000000000000001010110111011111;
assign LUT_3[52132] = 32'b11111111111111111111010010010100;
assign LUT_3[52133] = 32'b00000000000000000101111101110001;
assign LUT_3[52134] = 32'b00000000000000000001011001111000;
assign LUT_3[52135] = 32'b00000000000000001000000101010101;
assign LUT_3[52136] = 32'b00000000000000000111011101100100;
assign LUT_3[52137] = 32'b00000000000000001110001001000001;
assign LUT_3[52138] = 32'b00000000000000001001100101001000;
assign LUT_3[52139] = 32'b00000000000000010000010000100101;
assign LUT_3[52140] = 32'b00000000000000000100101011011010;
assign LUT_3[52141] = 32'b00000000000000001011010110110111;
assign LUT_3[52142] = 32'b00000000000000000110110010111110;
assign LUT_3[52143] = 32'b00000000000000001101011110011011;
assign LUT_3[52144] = 32'b00000000000000000101010111100001;
assign LUT_3[52145] = 32'b00000000000000001100000010111110;
assign LUT_3[52146] = 32'b00000000000000000111011111000101;
assign LUT_3[52147] = 32'b00000000000000001110001010100010;
assign LUT_3[52148] = 32'b00000000000000000010100101010111;
assign LUT_3[52149] = 32'b00000000000000001001010000110100;
assign LUT_3[52150] = 32'b00000000000000000100101100111011;
assign LUT_3[52151] = 32'b00000000000000001011011000011000;
assign LUT_3[52152] = 32'b00000000000000001010110000100111;
assign LUT_3[52153] = 32'b00000000000000010001011100000100;
assign LUT_3[52154] = 32'b00000000000000001100111000001011;
assign LUT_3[52155] = 32'b00000000000000010011100011101000;
assign LUT_3[52156] = 32'b00000000000000000111111110011101;
assign LUT_3[52157] = 32'b00000000000000001110101001111010;
assign LUT_3[52158] = 32'b00000000000000001010000110000001;
assign LUT_3[52159] = 32'b00000000000000010000110001011110;
assign LUT_3[52160] = 32'b00000000000000000000101110101001;
assign LUT_3[52161] = 32'b00000000000000000111011010000110;
assign LUT_3[52162] = 32'b00000000000000000010110110001101;
assign LUT_3[52163] = 32'b00000000000000001001100001101010;
assign LUT_3[52164] = 32'b11111111111111111101111100011111;
assign LUT_3[52165] = 32'b00000000000000000100100111111100;
assign LUT_3[52166] = 32'b00000000000000000000000100000011;
assign LUT_3[52167] = 32'b00000000000000000110101111100000;
assign LUT_3[52168] = 32'b00000000000000000110000111101111;
assign LUT_3[52169] = 32'b00000000000000001100110011001100;
assign LUT_3[52170] = 32'b00000000000000001000001111010011;
assign LUT_3[52171] = 32'b00000000000000001110111010110000;
assign LUT_3[52172] = 32'b00000000000000000011010101100101;
assign LUT_3[52173] = 32'b00000000000000001010000001000010;
assign LUT_3[52174] = 32'b00000000000000000101011101001001;
assign LUT_3[52175] = 32'b00000000000000001100001000100110;
assign LUT_3[52176] = 32'b00000000000000000100000001101100;
assign LUT_3[52177] = 32'b00000000000000001010101101001001;
assign LUT_3[52178] = 32'b00000000000000000110001001010000;
assign LUT_3[52179] = 32'b00000000000000001100110100101101;
assign LUT_3[52180] = 32'b00000000000000000001001111100010;
assign LUT_3[52181] = 32'b00000000000000000111111010111111;
assign LUT_3[52182] = 32'b00000000000000000011010111000110;
assign LUT_3[52183] = 32'b00000000000000001010000010100011;
assign LUT_3[52184] = 32'b00000000000000001001011010110010;
assign LUT_3[52185] = 32'b00000000000000010000000110001111;
assign LUT_3[52186] = 32'b00000000000000001011100010010110;
assign LUT_3[52187] = 32'b00000000000000010010001101110011;
assign LUT_3[52188] = 32'b00000000000000000110101000101000;
assign LUT_3[52189] = 32'b00000000000000001101010100000101;
assign LUT_3[52190] = 32'b00000000000000001000110000001100;
assign LUT_3[52191] = 32'b00000000000000001111011011101001;
assign LUT_3[52192] = 32'b00000000000000000001111101001001;
assign LUT_3[52193] = 32'b00000000000000001000101000100110;
assign LUT_3[52194] = 32'b00000000000000000100000100101101;
assign LUT_3[52195] = 32'b00000000000000001010110000001010;
assign LUT_3[52196] = 32'b11111111111111111111001010111111;
assign LUT_3[52197] = 32'b00000000000000000101110110011100;
assign LUT_3[52198] = 32'b00000000000000000001010010100011;
assign LUT_3[52199] = 32'b00000000000000000111111110000000;
assign LUT_3[52200] = 32'b00000000000000000111010110001111;
assign LUT_3[52201] = 32'b00000000000000001110000001101100;
assign LUT_3[52202] = 32'b00000000000000001001011101110011;
assign LUT_3[52203] = 32'b00000000000000010000001001010000;
assign LUT_3[52204] = 32'b00000000000000000100100100000101;
assign LUT_3[52205] = 32'b00000000000000001011001111100010;
assign LUT_3[52206] = 32'b00000000000000000110101011101001;
assign LUT_3[52207] = 32'b00000000000000001101010111000110;
assign LUT_3[52208] = 32'b00000000000000000101010000001100;
assign LUT_3[52209] = 32'b00000000000000001011111011101001;
assign LUT_3[52210] = 32'b00000000000000000111010111110000;
assign LUT_3[52211] = 32'b00000000000000001110000011001101;
assign LUT_3[52212] = 32'b00000000000000000010011110000010;
assign LUT_3[52213] = 32'b00000000000000001001001001011111;
assign LUT_3[52214] = 32'b00000000000000000100100101100110;
assign LUT_3[52215] = 32'b00000000000000001011010001000011;
assign LUT_3[52216] = 32'b00000000000000001010101001010010;
assign LUT_3[52217] = 32'b00000000000000010001010100101111;
assign LUT_3[52218] = 32'b00000000000000001100110000110110;
assign LUT_3[52219] = 32'b00000000000000010011011100010011;
assign LUT_3[52220] = 32'b00000000000000000111110111001000;
assign LUT_3[52221] = 32'b00000000000000001110100010100101;
assign LUT_3[52222] = 32'b00000000000000001001111110101100;
assign LUT_3[52223] = 32'b00000000000000010000101010001001;
assign LUT_3[52224] = 32'b00000000000000000101101011010000;
assign LUT_3[52225] = 32'b00000000000000001100010110101101;
assign LUT_3[52226] = 32'b00000000000000000111110010110100;
assign LUT_3[52227] = 32'b00000000000000001110011110010001;
assign LUT_3[52228] = 32'b00000000000000000010111001000110;
assign LUT_3[52229] = 32'b00000000000000001001100100100011;
assign LUT_3[52230] = 32'b00000000000000000101000000101010;
assign LUT_3[52231] = 32'b00000000000000001011101100000111;
assign LUT_3[52232] = 32'b00000000000000001011000100010110;
assign LUT_3[52233] = 32'b00000000000000010001101111110011;
assign LUT_3[52234] = 32'b00000000000000001101001011111010;
assign LUT_3[52235] = 32'b00000000000000010011110111010111;
assign LUT_3[52236] = 32'b00000000000000001000010010001100;
assign LUT_3[52237] = 32'b00000000000000001110111101101001;
assign LUT_3[52238] = 32'b00000000000000001010011001110000;
assign LUT_3[52239] = 32'b00000000000000010001000101001101;
assign LUT_3[52240] = 32'b00000000000000001000111110010011;
assign LUT_3[52241] = 32'b00000000000000001111101001110000;
assign LUT_3[52242] = 32'b00000000000000001011000101110111;
assign LUT_3[52243] = 32'b00000000000000010001110001010100;
assign LUT_3[52244] = 32'b00000000000000000110001100001001;
assign LUT_3[52245] = 32'b00000000000000001100110111100110;
assign LUT_3[52246] = 32'b00000000000000001000010011101101;
assign LUT_3[52247] = 32'b00000000000000001110111111001010;
assign LUT_3[52248] = 32'b00000000000000001110010111011001;
assign LUT_3[52249] = 32'b00000000000000010101000010110110;
assign LUT_3[52250] = 32'b00000000000000010000011110111101;
assign LUT_3[52251] = 32'b00000000000000010111001010011010;
assign LUT_3[52252] = 32'b00000000000000001011100101001111;
assign LUT_3[52253] = 32'b00000000000000010010010000101100;
assign LUT_3[52254] = 32'b00000000000000001101101100110011;
assign LUT_3[52255] = 32'b00000000000000010100011000010000;
assign LUT_3[52256] = 32'b00000000000000000110111001110000;
assign LUT_3[52257] = 32'b00000000000000001101100101001101;
assign LUT_3[52258] = 32'b00000000000000001001000001010100;
assign LUT_3[52259] = 32'b00000000000000001111101100110001;
assign LUT_3[52260] = 32'b00000000000000000100000111100110;
assign LUT_3[52261] = 32'b00000000000000001010110011000011;
assign LUT_3[52262] = 32'b00000000000000000110001111001010;
assign LUT_3[52263] = 32'b00000000000000001100111010100111;
assign LUT_3[52264] = 32'b00000000000000001100010010110110;
assign LUT_3[52265] = 32'b00000000000000010010111110010011;
assign LUT_3[52266] = 32'b00000000000000001110011010011010;
assign LUT_3[52267] = 32'b00000000000000010101000101110111;
assign LUT_3[52268] = 32'b00000000000000001001100000101100;
assign LUT_3[52269] = 32'b00000000000000010000001100001001;
assign LUT_3[52270] = 32'b00000000000000001011101000010000;
assign LUT_3[52271] = 32'b00000000000000010010010011101101;
assign LUT_3[52272] = 32'b00000000000000001010001100110011;
assign LUT_3[52273] = 32'b00000000000000010000111000010000;
assign LUT_3[52274] = 32'b00000000000000001100010100010111;
assign LUT_3[52275] = 32'b00000000000000010010111111110100;
assign LUT_3[52276] = 32'b00000000000000000111011010101001;
assign LUT_3[52277] = 32'b00000000000000001110000110000110;
assign LUT_3[52278] = 32'b00000000000000001001100010001101;
assign LUT_3[52279] = 32'b00000000000000010000001101101010;
assign LUT_3[52280] = 32'b00000000000000001111100101111001;
assign LUT_3[52281] = 32'b00000000000000010110010001010110;
assign LUT_3[52282] = 32'b00000000000000010001101101011101;
assign LUT_3[52283] = 32'b00000000000000011000011000111010;
assign LUT_3[52284] = 32'b00000000000000001100110011101111;
assign LUT_3[52285] = 32'b00000000000000010011011111001100;
assign LUT_3[52286] = 32'b00000000000000001110111011010011;
assign LUT_3[52287] = 32'b00000000000000010101100110110000;
assign LUT_3[52288] = 32'b00000000000000000101100011111011;
assign LUT_3[52289] = 32'b00000000000000001100001111011000;
assign LUT_3[52290] = 32'b00000000000000000111101011011111;
assign LUT_3[52291] = 32'b00000000000000001110010110111100;
assign LUT_3[52292] = 32'b00000000000000000010110001110001;
assign LUT_3[52293] = 32'b00000000000000001001011101001110;
assign LUT_3[52294] = 32'b00000000000000000100111001010101;
assign LUT_3[52295] = 32'b00000000000000001011100100110010;
assign LUT_3[52296] = 32'b00000000000000001010111101000001;
assign LUT_3[52297] = 32'b00000000000000010001101000011110;
assign LUT_3[52298] = 32'b00000000000000001101000100100101;
assign LUT_3[52299] = 32'b00000000000000010011110000000010;
assign LUT_3[52300] = 32'b00000000000000001000001010110111;
assign LUT_3[52301] = 32'b00000000000000001110110110010100;
assign LUT_3[52302] = 32'b00000000000000001010010010011011;
assign LUT_3[52303] = 32'b00000000000000010000111101111000;
assign LUT_3[52304] = 32'b00000000000000001000110110111110;
assign LUT_3[52305] = 32'b00000000000000001111100010011011;
assign LUT_3[52306] = 32'b00000000000000001010111110100010;
assign LUT_3[52307] = 32'b00000000000000010001101001111111;
assign LUT_3[52308] = 32'b00000000000000000110000100110100;
assign LUT_3[52309] = 32'b00000000000000001100110000010001;
assign LUT_3[52310] = 32'b00000000000000001000001100011000;
assign LUT_3[52311] = 32'b00000000000000001110110111110101;
assign LUT_3[52312] = 32'b00000000000000001110010000000100;
assign LUT_3[52313] = 32'b00000000000000010100111011100001;
assign LUT_3[52314] = 32'b00000000000000010000010111101000;
assign LUT_3[52315] = 32'b00000000000000010111000011000101;
assign LUT_3[52316] = 32'b00000000000000001011011101111010;
assign LUT_3[52317] = 32'b00000000000000010010001001010111;
assign LUT_3[52318] = 32'b00000000000000001101100101011110;
assign LUT_3[52319] = 32'b00000000000000010100010000111011;
assign LUT_3[52320] = 32'b00000000000000000110110010011011;
assign LUT_3[52321] = 32'b00000000000000001101011101111000;
assign LUT_3[52322] = 32'b00000000000000001000111001111111;
assign LUT_3[52323] = 32'b00000000000000001111100101011100;
assign LUT_3[52324] = 32'b00000000000000000100000000010001;
assign LUT_3[52325] = 32'b00000000000000001010101011101110;
assign LUT_3[52326] = 32'b00000000000000000110000111110101;
assign LUT_3[52327] = 32'b00000000000000001100110011010010;
assign LUT_3[52328] = 32'b00000000000000001100001011100001;
assign LUT_3[52329] = 32'b00000000000000010010110110111110;
assign LUT_3[52330] = 32'b00000000000000001110010011000101;
assign LUT_3[52331] = 32'b00000000000000010100111110100010;
assign LUT_3[52332] = 32'b00000000000000001001011001010111;
assign LUT_3[52333] = 32'b00000000000000010000000100110100;
assign LUT_3[52334] = 32'b00000000000000001011100000111011;
assign LUT_3[52335] = 32'b00000000000000010010001100011000;
assign LUT_3[52336] = 32'b00000000000000001010000101011110;
assign LUT_3[52337] = 32'b00000000000000010000110000111011;
assign LUT_3[52338] = 32'b00000000000000001100001101000010;
assign LUT_3[52339] = 32'b00000000000000010010111000011111;
assign LUT_3[52340] = 32'b00000000000000000111010011010100;
assign LUT_3[52341] = 32'b00000000000000001101111110110001;
assign LUT_3[52342] = 32'b00000000000000001001011010111000;
assign LUT_3[52343] = 32'b00000000000000010000000110010101;
assign LUT_3[52344] = 32'b00000000000000001111011110100100;
assign LUT_3[52345] = 32'b00000000000000010110001010000001;
assign LUT_3[52346] = 32'b00000000000000010001100110001000;
assign LUT_3[52347] = 32'b00000000000000011000010001100101;
assign LUT_3[52348] = 32'b00000000000000001100101100011010;
assign LUT_3[52349] = 32'b00000000000000010011010111110111;
assign LUT_3[52350] = 32'b00000000000000001110110011111110;
assign LUT_3[52351] = 32'b00000000000000010101011111011011;
assign LUT_3[52352] = 32'b00000000000000000111110110001110;
assign LUT_3[52353] = 32'b00000000000000001110100001101011;
assign LUT_3[52354] = 32'b00000000000000001001111101110010;
assign LUT_3[52355] = 32'b00000000000000010000101001001111;
assign LUT_3[52356] = 32'b00000000000000000101000100000100;
assign LUT_3[52357] = 32'b00000000000000001011101111100001;
assign LUT_3[52358] = 32'b00000000000000000111001011101000;
assign LUT_3[52359] = 32'b00000000000000001101110111000101;
assign LUT_3[52360] = 32'b00000000000000001101001111010100;
assign LUT_3[52361] = 32'b00000000000000010011111010110001;
assign LUT_3[52362] = 32'b00000000000000001111010110111000;
assign LUT_3[52363] = 32'b00000000000000010110000010010101;
assign LUT_3[52364] = 32'b00000000000000001010011101001010;
assign LUT_3[52365] = 32'b00000000000000010001001000100111;
assign LUT_3[52366] = 32'b00000000000000001100100100101110;
assign LUT_3[52367] = 32'b00000000000000010011010000001011;
assign LUT_3[52368] = 32'b00000000000000001011001001010001;
assign LUT_3[52369] = 32'b00000000000000010001110100101110;
assign LUT_3[52370] = 32'b00000000000000001101010000110101;
assign LUT_3[52371] = 32'b00000000000000010011111100010010;
assign LUT_3[52372] = 32'b00000000000000001000010111000111;
assign LUT_3[52373] = 32'b00000000000000001111000010100100;
assign LUT_3[52374] = 32'b00000000000000001010011110101011;
assign LUT_3[52375] = 32'b00000000000000010001001010001000;
assign LUT_3[52376] = 32'b00000000000000010000100010010111;
assign LUT_3[52377] = 32'b00000000000000010111001101110100;
assign LUT_3[52378] = 32'b00000000000000010010101001111011;
assign LUT_3[52379] = 32'b00000000000000011001010101011000;
assign LUT_3[52380] = 32'b00000000000000001101110000001101;
assign LUT_3[52381] = 32'b00000000000000010100011011101010;
assign LUT_3[52382] = 32'b00000000000000001111110111110001;
assign LUT_3[52383] = 32'b00000000000000010110100011001110;
assign LUT_3[52384] = 32'b00000000000000001001000100101110;
assign LUT_3[52385] = 32'b00000000000000001111110000001011;
assign LUT_3[52386] = 32'b00000000000000001011001100010010;
assign LUT_3[52387] = 32'b00000000000000010001110111101111;
assign LUT_3[52388] = 32'b00000000000000000110010010100100;
assign LUT_3[52389] = 32'b00000000000000001100111110000001;
assign LUT_3[52390] = 32'b00000000000000001000011010001000;
assign LUT_3[52391] = 32'b00000000000000001111000101100101;
assign LUT_3[52392] = 32'b00000000000000001110011101110100;
assign LUT_3[52393] = 32'b00000000000000010101001001010001;
assign LUT_3[52394] = 32'b00000000000000010000100101011000;
assign LUT_3[52395] = 32'b00000000000000010111010000110101;
assign LUT_3[52396] = 32'b00000000000000001011101011101010;
assign LUT_3[52397] = 32'b00000000000000010010010111000111;
assign LUT_3[52398] = 32'b00000000000000001101110011001110;
assign LUT_3[52399] = 32'b00000000000000010100011110101011;
assign LUT_3[52400] = 32'b00000000000000001100010111110001;
assign LUT_3[52401] = 32'b00000000000000010011000011001110;
assign LUT_3[52402] = 32'b00000000000000001110011111010101;
assign LUT_3[52403] = 32'b00000000000000010101001010110010;
assign LUT_3[52404] = 32'b00000000000000001001100101100111;
assign LUT_3[52405] = 32'b00000000000000010000010001000100;
assign LUT_3[52406] = 32'b00000000000000001011101101001011;
assign LUT_3[52407] = 32'b00000000000000010010011000101000;
assign LUT_3[52408] = 32'b00000000000000010001110000110111;
assign LUT_3[52409] = 32'b00000000000000011000011100010100;
assign LUT_3[52410] = 32'b00000000000000010011111000011011;
assign LUT_3[52411] = 32'b00000000000000011010100011111000;
assign LUT_3[52412] = 32'b00000000000000001110111110101101;
assign LUT_3[52413] = 32'b00000000000000010101101010001010;
assign LUT_3[52414] = 32'b00000000000000010001000110010001;
assign LUT_3[52415] = 32'b00000000000000010111110001101110;
assign LUT_3[52416] = 32'b00000000000000000111101110111001;
assign LUT_3[52417] = 32'b00000000000000001110011010010110;
assign LUT_3[52418] = 32'b00000000000000001001110110011101;
assign LUT_3[52419] = 32'b00000000000000010000100001111010;
assign LUT_3[52420] = 32'b00000000000000000100111100101111;
assign LUT_3[52421] = 32'b00000000000000001011101000001100;
assign LUT_3[52422] = 32'b00000000000000000111000100010011;
assign LUT_3[52423] = 32'b00000000000000001101101111110000;
assign LUT_3[52424] = 32'b00000000000000001101000111111111;
assign LUT_3[52425] = 32'b00000000000000010011110011011100;
assign LUT_3[52426] = 32'b00000000000000001111001111100011;
assign LUT_3[52427] = 32'b00000000000000010101111011000000;
assign LUT_3[52428] = 32'b00000000000000001010010101110101;
assign LUT_3[52429] = 32'b00000000000000010001000001010010;
assign LUT_3[52430] = 32'b00000000000000001100011101011001;
assign LUT_3[52431] = 32'b00000000000000010011001000110110;
assign LUT_3[52432] = 32'b00000000000000001011000001111100;
assign LUT_3[52433] = 32'b00000000000000010001101101011001;
assign LUT_3[52434] = 32'b00000000000000001101001001100000;
assign LUT_3[52435] = 32'b00000000000000010011110100111101;
assign LUT_3[52436] = 32'b00000000000000001000001111110010;
assign LUT_3[52437] = 32'b00000000000000001110111011001111;
assign LUT_3[52438] = 32'b00000000000000001010010111010110;
assign LUT_3[52439] = 32'b00000000000000010001000010110011;
assign LUT_3[52440] = 32'b00000000000000010000011011000010;
assign LUT_3[52441] = 32'b00000000000000010111000110011111;
assign LUT_3[52442] = 32'b00000000000000010010100010100110;
assign LUT_3[52443] = 32'b00000000000000011001001110000011;
assign LUT_3[52444] = 32'b00000000000000001101101000111000;
assign LUT_3[52445] = 32'b00000000000000010100010100010101;
assign LUT_3[52446] = 32'b00000000000000001111110000011100;
assign LUT_3[52447] = 32'b00000000000000010110011011111001;
assign LUT_3[52448] = 32'b00000000000000001000111101011001;
assign LUT_3[52449] = 32'b00000000000000001111101000110110;
assign LUT_3[52450] = 32'b00000000000000001011000100111101;
assign LUT_3[52451] = 32'b00000000000000010001110000011010;
assign LUT_3[52452] = 32'b00000000000000000110001011001111;
assign LUT_3[52453] = 32'b00000000000000001100110110101100;
assign LUT_3[52454] = 32'b00000000000000001000010010110011;
assign LUT_3[52455] = 32'b00000000000000001110111110010000;
assign LUT_3[52456] = 32'b00000000000000001110010110011111;
assign LUT_3[52457] = 32'b00000000000000010101000001111100;
assign LUT_3[52458] = 32'b00000000000000010000011110000011;
assign LUT_3[52459] = 32'b00000000000000010111001001100000;
assign LUT_3[52460] = 32'b00000000000000001011100100010101;
assign LUT_3[52461] = 32'b00000000000000010010001111110010;
assign LUT_3[52462] = 32'b00000000000000001101101011111001;
assign LUT_3[52463] = 32'b00000000000000010100010111010110;
assign LUT_3[52464] = 32'b00000000000000001100010000011100;
assign LUT_3[52465] = 32'b00000000000000010010111011111001;
assign LUT_3[52466] = 32'b00000000000000001110011000000000;
assign LUT_3[52467] = 32'b00000000000000010101000011011101;
assign LUT_3[52468] = 32'b00000000000000001001011110010010;
assign LUT_3[52469] = 32'b00000000000000010000001001101111;
assign LUT_3[52470] = 32'b00000000000000001011100101110110;
assign LUT_3[52471] = 32'b00000000000000010010010001010011;
assign LUT_3[52472] = 32'b00000000000000010001101001100010;
assign LUT_3[52473] = 32'b00000000000000011000010100111111;
assign LUT_3[52474] = 32'b00000000000000010011110001000110;
assign LUT_3[52475] = 32'b00000000000000011010011100100011;
assign LUT_3[52476] = 32'b00000000000000001110110111011000;
assign LUT_3[52477] = 32'b00000000000000010101100010110101;
assign LUT_3[52478] = 32'b00000000000000010000111110111100;
assign LUT_3[52479] = 32'b00000000000000010111101010011001;
assign LUT_3[52480] = 32'b00000000000000000001111010110001;
assign LUT_3[52481] = 32'b00000000000000001000100110001110;
assign LUT_3[52482] = 32'b00000000000000000100000010010101;
assign LUT_3[52483] = 32'b00000000000000001010101101110010;
assign LUT_3[52484] = 32'b11111111111111111111001000100111;
assign LUT_3[52485] = 32'b00000000000000000101110100000100;
assign LUT_3[52486] = 32'b00000000000000000001010000001011;
assign LUT_3[52487] = 32'b00000000000000000111111011101000;
assign LUT_3[52488] = 32'b00000000000000000111010011110111;
assign LUT_3[52489] = 32'b00000000000000001101111111010100;
assign LUT_3[52490] = 32'b00000000000000001001011011011011;
assign LUT_3[52491] = 32'b00000000000000010000000110111000;
assign LUT_3[52492] = 32'b00000000000000000100100001101101;
assign LUT_3[52493] = 32'b00000000000000001011001101001010;
assign LUT_3[52494] = 32'b00000000000000000110101001010001;
assign LUT_3[52495] = 32'b00000000000000001101010100101110;
assign LUT_3[52496] = 32'b00000000000000000101001101110100;
assign LUT_3[52497] = 32'b00000000000000001011111001010001;
assign LUT_3[52498] = 32'b00000000000000000111010101011000;
assign LUT_3[52499] = 32'b00000000000000001110000000110101;
assign LUT_3[52500] = 32'b00000000000000000010011011101010;
assign LUT_3[52501] = 32'b00000000000000001001000111000111;
assign LUT_3[52502] = 32'b00000000000000000100100011001110;
assign LUT_3[52503] = 32'b00000000000000001011001110101011;
assign LUT_3[52504] = 32'b00000000000000001010100110111010;
assign LUT_3[52505] = 32'b00000000000000010001010010010111;
assign LUT_3[52506] = 32'b00000000000000001100101110011110;
assign LUT_3[52507] = 32'b00000000000000010011011001111011;
assign LUT_3[52508] = 32'b00000000000000000111110100110000;
assign LUT_3[52509] = 32'b00000000000000001110100000001101;
assign LUT_3[52510] = 32'b00000000000000001001111100010100;
assign LUT_3[52511] = 32'b00000000000000010000100111110001;
assign LUT_3[52512] = 32'b00000000000000000011001001010001;
assign LUT_3[52513] = 32'b00000000000000001001110100101110;
assign LUT_3[52514] = 32'b00000000000000000101010000110101;
assign LUT_3[52515] = 32'b00000000000000001011111100010010;
assign LUT_3[52516] = 32'b00000000000000000000010111000111;
assign LUT_3[52517] = 32'b00000000000000000111000010100100;
assign LUT_3[52518] = 32'b00000000000000000010011110101011;
assign LUT_3[52519] = 32'b00000000000000001001001010001000;
assign LUT_3[52520] = 32'b00000000000000001000100010010111;
assign LUT_3[52521] = 32'b00000000000000001111001101110100;
assign LUT_3[52522] = 32'b00000000000000001010101001111011;
assign LUT_3[52523] = 32'b00000000000000010001010101011000;
assign LUT_3[52524] = 32'b00000000000000000101110000001101;
assign LUT_3[52525] = 32'b00000000000000001100011011101010;
assign LUT_3[52526] = 32'b00000000000000000111110111110001;
assign LUT_3[52527] = 32'b00000000000000001110100011001110;
assign LUT_3[52528] = 32'b00000000000000000110011100010100;
assign LUT_3[52529] = 32'b00000000000000001101000111110001;
assign LUT_3[52530] = 32'b00000000000000001000100011111000;
assign LUT_3[52531] = 32'b00000000000000001111001111010101;
assign LUT_3[52532] = 32'b00000000000000000011101010001010;
assign LUT_3[52533] = 32'b00000000000000001010010101100111;
assign LUT_3[52534] = 32'b00000000000000000101110001101110;
assign LUT_3[52535] = 32'b00000000000000001100011101001011;
assign LUT_3[52536] = 32'b00000000000000001011110101011010;
assign LUT_3[52537] = 32'b00000000000000010010100000110111;
assign LUT_3[52538] = 32'b00000000000000001101111100111110;
assign LUT_3[52539] = 32'b00000000000000010100101000011011;
assign LUT_3[52540] = 32'b00000000000000001001000011010000;
assign LUT_3[52541] = 32'b00000000000000001111101110101101;
assign LUT_3[52542] = 32'b00000000000000001011001010110100;
assign LUT_3[52543] = 32'b00000000000000010001110110010001;
assign LUT_3[52544] = 32'b00000000000000000001110011011100;
assign LUT_3[52545] = 32'b00000000000000001000011110111001;
assign LUT_3[52546] = 32'b00000000000000000011111011000000;
assign LUT_3[52547] = 32'b00000000000000001010100110011101;
assign LUT_3[52548] = 32'b11111111111111111111000001010010;
assign LUT_3[52549] = 32'b00000000000000000101101100101111;
assign LUT_3[52550] = 32'b00000000000000000001001000110110;
assign LUT_3[52551] = 32'b00000000000000000111110100010011;
assign LUT_3[52552] = 32'b00000000000000000111001100100010;
assign LUT_3[52553] = 32'b00000000000000001101110111111111;
assign LUT_3[52554] = 32'b00000000000000001001010100000110;
assign LUT_3[52555] = 32'b00000000000000001111111111100011;
assign LUT_3[52556] = 32'b00000000000000000100011010011000;
assign LUT_3[52557] = 32'b00000000000000001011000101110101;
assign LUT_3[52558] = 32'b00000000000000000110100001111100;
assign LUT_3[52559] = 32'b00000000000000001101001101011001;
assign LUT_3[52560] = 32'b00000000000000000101000110011111;
assign LUT_3[52561] = 32'b00000000000000001011110001111100;
assign LUT_3[52562] = 32'b00000000000000000111001110000011;
assign LUT_3[52563] = 32'b00000000000000001101111001100000;
assign LUT_3[52564] = 32'b00000000000000000010010100010101;
assign LUT_3[52565] = 32'b00000000000000001000111111110010;
assign LUT_3[52566] = 32'b00000000000000000100011011111001;
assign LUT_3[52567] = 32'b00000000000000001011000111010110;
assign LUT_3[52568] = 32'b00000000000000001010011111100101;
assign LUT_3[52569] = 32'b00000000000000010001001011000010;
assign LUT_3[52570] = 32'b00000000000000001100100111001001;
assign LUT_3[52571] = 32'b00000000000000010011010010100110;
assign LUT_3[52572] = 32'b00000000000000000111101101011011;
assign LUT_3[52573] = 32'b00000000000000001110011000111000;
assign LUT_3[52574] = 32'b00000000000000001001110100111111;
assign LUT_3[52575] = 32'b00000000000000010000100000011100;
assign LUT_3[52576] = 32'b00000000000000000011000001111100;
assign LUT_3[52577] = 32'b00000000000000001001101101011001;
assign LUT_3[52578] = 32'b00000000000000000101001001100000;
assign LUT_3[52579] = 32'b00000000000000001011110100111101;
assign LUT_3[52580] = 32'b00000000000000000000001111110010;
assign LUT_3[52581] = 32'b00000000000000000110111011001111;
assign LUT_3[52582] = 32'b00000000000000000010010111010110;
assign LUT_3[52583] = 32'b00000000000000001001000010110011;
assign LUT_3[52584] = 32'b00000000000000001000011011000010;
assign LUT_3[52585] = 32'b00000000000000001111000110011111;
assign LUT_3[52586] = 32'b00000000000000001010100010100110;
assign LUT_3[52587] = 32'b00000000000000010001001110000011;
assign LUT_3[52588] = 32'b00000000000000000101101000111000;
assign LUT_3[52589] = 32'b00000000000000001100010100010101;
assign LUT_3[52590] = 32'b00000000000000000111110000011100;
assign LUT_3[52591] = 32'b00000000000000001110011011111001;
assign LUT_3[52592] = 32'b00000000000000000110010100111111;
assign LUT_3[52593] = 32'b00000000000000001101000000011100;
assign LUT_3[52594] = 32'b00000000000000001000011100100011;
assign LUT_3[52595] = 32'b00000000000000001111001000000000;
assign LUT_3[52596] = 32'b00000000000000000011100010110101;
assign LUT_3[52597] = 32'b00000000000000001010001110010010;
assign LUT_3[52598] = 32'b00000000000000000101101010011001;
assign LUT_3[52599] = 32'b00000000000000001100010101110110;
assign LUT_3[52600] = 32'b00000000000000001011101110000101;
assign LUT_3[52601] = 32'b00000000000000010010011001100010;
assign LUT_3[52602] = 32'b00000000000000001101110101101001;
assign LUT_3[52603] = 32'b00000000000000010100100001000110;
assign LUT_3[52604] = 32'b00000000000000001000111011111011;
assign LUT_3[52605] = 32'b00000000000000001111100111011000;
assign LUT_3[52606] = 32'b00000000000000001011000011011111;
assign LUT_3[52607] = 32'b00000000000000010001101110111100;
assign LUT_3[52608] = 32'b00000000000000000100000101101111;
assign LUT_3[52609] = 32'b00000000000000001010110001001100;
assign LUT_3[52610] = 32'b00000000000000000110001101010011;
assign LUT_3[52611] = 32'b00000000000000001100111000110000;
assign LUT_3[52612] = 32'b00000000000000000001010011100101;
assign LUT_3[52613] = 32'b00000000000000000111111111000010;
assign LUT_3[52614] = 32'b00000000000000000011011011001001;
assign LUT_3[52615] = 32'b00000000000000001010000110100110;
assign LUT_3[52616] = 32'b00000000000000001001011110110101;
assign LUT_3[52617] = 32'b00000000000000010000001010010010;
assign LUT_3[52618] = 32'b00000000000000001011100110011001;
assign LUT_3[52619] = 32'b00000000000000010010010001110110;
assign LUT_3[52620] = 32'b00000000000000000110101100101011;
assign LUT_3[52621] = 32'b00000000000000001101011000001000;
assign LUT_3[52622] = 32'b00000000000000001000110100001111;
assign LUT_3[52623] = 32'b00000000000000001111011111101100;
assign LUT_3[52624] = 32'b00000000000000000111011000110010;
assign LUT_3[52625] = 32'b00000000000000001110000100001111;
assign LUT_3[52626] = 32'b00000000000000001001100000010110;
assign LUT_3[52627] = 32'b00000000000000010000001011110011;
assign LUT_3[52628] = 32'b00000000000000000100100110101000;
assign LUT_3[52629] = 32'b00000000000000001011010010000101;
assign LUT_3[52630] = 32'b00000000000000000110101110001100;
assign LUT_3[52631] = 32'b00000000000000001101011001101001;
assign LUT_3[52632] = 32'b00000000000000001100110001111000;
assign LUT_3[52633] = 32'b00000000000000010011011101010101;
assign LUT_3[52634] = 32'b00000000000000001110111001011100;
assign LUT_3[52635] = 32'b00000000000000010101100100111001;
assign LUT_3[52636] = 32'b00000000000000001001111111101110;
assign LUT_3[52637] = 32'b00000000000000010000101011001011;
assign LUT_3[52638] = 32'b00000000000000001100000111010010;
assign LUT_3[52639] = 32'b00000000000000010010110010101111;
assign LUT_3[52640] = 32'b00000000000000000101010100001111;
assign LUT_3[52641] = 32'b00000000000000001011111111101100;
assign LUT_3[52642] = 32'b00000000000000000111011011110011;
assign LUT_3[52643] = 32'b00000000000000001110000111010000;
assign LUT_3[52644] = 32'b00000000000000000010100010000101;
assign LUT_3[52645] = 32'b00000000000000001001001101100010;
assign LUT_3[52646] = 32'b00000000000000000100101001101001;
assign LUT_3[52647] = 32'b00000000000000001011010101000110;
assign LUT_3[52648] = 32'b00000000000000001010101101010101;
assign LUT_3[52649] = 32'b00000000000000010001011000110010;
assign LUT_3[52650] = 32'b00000000000000001100110100111001;
assign LUT_3[52651] = 32'b00000000000000010011100000010110;
assign LUT_3[52652] = 32'b00000000000000000111111011001011;
assign LUT_3[52653] = 32'b00000000000000001110100110101000;
assign LUT_3[52654] = 32'b00000000000000001010000010101111;
assign LUT_3[52655] = 32'b00000000000000010000101110001100;
assign LUT_3[52656] = 32'b00000000000000001000100111010010;
assign LUT_3[52657] = 32'b00000000000000001111010010101111;
assign LUT_3[52658] = 32'b00000000000000001010101110110110;
assign LUT_3[52659] = 32'b00000000000000010001011010010011;
assign LUT_3[52660] = 32'b00000000000000000101110101001000;
assign LUT_3[52661] = 32'b00000000000000001100100000100101;
assign LUT_3[52662] = 32'b00000000000000000111111100101100;
assign LUT_3[52663] = 32'b00000000000000001110101000001001;
assign LUT_3[52664] = 32'b00000000000000001110000000011000;
assign LUT_3[52665] = 32'b00000000000000010100101011110101;
assign LUT_3[52666] = 32'b00000000000000010000000111111100;
assign LUT_3[52667] = 32'b00000000000000010110110011011001;
assign LUT_3[52668] = 32'b00000000000000001011001110001110;
assign LUT_3[52669] = 32'b00000000000000010001111001101011;
assign LUT_3[52670] = 32'b00000000000000001101010101110010;
assign LUT_3[52671] = 32'b00000000000000010100000001001111;
assign LUT_3[52672] = 32'b00000000000000000011111110011010;
assign LUT_3[52673] = 32'b00000000000000001010101001110111;
assign LUT_3[52674] = 32'b00000000000000000110000101111110;
assign LUT_3[52675] = 32'b00000000000000001100110001011011;
assign LUT_3[52676] = 32'b00000000000000000001001100010000;
assign LUT_3[52677] = 32'b00000000000000000111110111101101;
assign LUT_3[52678] = 32'b00000000000000000011010011110100;
assign LUT_3[52679] = 32'b00000000000000001001111111010001;
assign LUT_3[52680] = 32'b00000000000000001001010111100000;
assign LUT_3[52681] = 32'b00000000000000010000000010111101;
assign LUT_3[52682] = 32'b00000000000000001011011111000100;
assign LUT_3[52683] = 32'b00000000000000010010001010100001;
assign LUT_3[52684] = 32'b00000000000000000110100101010110;
assign LUT_3[52685] = 32'b00000000000000001101010000110011;
assign LUT_3[52686] = 32'b00000000000000001000101100111010;
assign LUT_3[52687] = 32'b00000000000000001111011000010111;
assign LUT_3[52688] = 32'b00000000000000000111010001011101;
assign LUT_3[52689] = 32'b00000000000000001101111100111010;
assign LUT_3[52690] = 32'b00000000000000001001011001000001;
assign LUT_3[52691] = 32'b00000000000000010000000100011110;
assign LUT_3[52692] = 32'b00000000000000000100011111010011;
assign LUT_3[52693] = 32'b00000000000000001011001010110000;
assign LUT_3[52694] = 32'b00000000000000000110100110110111;
assign LUT_3[52695] = 32'b00000000000000001101010010010100;
assign LUT_3[52696] = 32'b00000000000000001100101010100011;
assign LUT_3[52697] = 32'b00000000000000010011010110000000;
assign LUT_3[52698] = 32'b00000000000000001110110010000111;
assign LUT_3[52699] = 32'b00000000000000010101011101100100;
assign LUT_3[52700] = 32'b00000000000000001001111000011001;
assign LUT_3[52701] = 32'b00000000000000010000100011110110;
assign LUT_3[52702] = 32'b00000000000000001011111111111101;
assign LUT_3[52703] = 32'b00000000000000010010101011011010;
assign LUT_3[52704] = 32'b00000000000000000101001100111010;
assign LUT_3[52705] = 32'b00000000000000001011111000010111;
assign LUT_3[52706] = 32'b00000000000000000111010100011110;
assign LUT_3[52707] = 32'b00000000000000001101111111111011;
assign LUT_3[52708] = 32'b00000000000000000010011010110000;
assign LUT_3[52709] = 32'b00000000000000001001000110001101;
assign LUT_3[52710] = 32'b00000000000000000100100010010100;
assign LUT_3[52711] = 32'b00000000000000001011001101110001;
assign LUT_3[52712] = 32'b00000000000000001010100110000000;
assign LUT_3[52713] = 32'b00000000000000010001010001011101;
assign LUT_3[52714] = 32'b00000000000000001100101101100100;
assign LUT_3[52715] = 32'b00000000000000010011011001000001;
assign LUT_3[52716] = 32'b00000000000000000111110011110110;
assign LUT_3[52717] = 32'b00000000000000001110011111010011;
assign LUT_3[52718] = 32'b00000000000000001001111011011010;
assign LUT_3[52719] = 32'b00000000000000010000100110110111;
assign LUT_3[52720] = 32'b00000000000000001000011111111101;
assign LUT_3[52721] = 32'b00000000000000001111001011011010;
assign LUT_3[52722] = 32'b00000000000000001010100111100001;
assign LUT_3[52723] = 32'b00000000000000010001010010111110;
assign LUT_3[52724] = 32'b00000000000000000101101101110011;
assign LUT_3[52725] = 32'b00000000000000001100011001010000;
assign LUT_3[52726] = 32'b00000000000000000111110101010111;
assign LUT_3[52727] = 32'b00000000000000001110100000110100;
assign LUT_3[52728] = 32'b00000000000000001101111001000011;
assign LUT_3[52729] = 32'b00000000000000010100100100100000;
assign LUT_3[52730] = 32'b00000000000000010000000000100111;
assign LUT_3[52731] = 32'b00000000000000010110101100000100;
assign LUT_3[52732] = 32'b00000000000000001011000110111001;
assign LUT_3[52733] = 32'b00000000000000010001110010010110;
assign LUT_3[52734] = 32'b00000000000000001101001110011101;
assign LUT_3[52735] = 32'b00000000000000010011111001111010;
assign LUT_3[52736] = 32'b00000000000000001001000000011100;
assign LUT_3[52737] = 32'b00000000000000001111101011111001;
assign LUT_3[52738] = 32'b00000000000000001011001000000000;
assign LUT_3[52739] = 32'b00000000000000010001110011011101;
assign LUT_3[52740] = 32'b00000000000000000110001110010010;
assign LUT_3[52741] = 32'b00000000000000001100111001101111;
assign LUT_3[52742] = 32'b00000000000000001000010101110110;
assign LUT_3[52743] = 32'b00000000000000001111000001010011;
assign LUT_3[52744] = 32'b00000000000000001110011001100010;
assign LUT_3[52745] = 32'b00000000000000010101000100111111;
assign LUT_3[52746] = 32'b00000000000000010000100001000110;
assign LUT_3[52747] = 32'b00000000000000010111001100100011;
assign LUT_3[52748] = 32'b00000000000000001011100111011000;
assign LUT_3[52749] = 32'b00000000000000010010010010110101;
assign LUT_3[52750] = 32'b00000000000000001101101110111100;
assign LUT_3[52751] = 32'b00000000000000010100011010011001;
assign LUT_3[52752] = 32'b00000000000000001100010011011111;
assign LUT_3[52753] = 32'b00000000000000010010111110111100;
assign LUT_3[52754] = 32'b00000000000000001110011011000011;
assign LUT_3[52755] = 32'b00000000000000010101000110100000;
assign LUT_3[52756] = 32'b00000000000000001001100001010101;
assign LUT_3[52757] = 32'b00000000000000010000001100110010;
assign LUT_3[52758] = 32'b00000000000000001011101000111001;
assign LUT_3[52759] = 32'b00000000000000010010010100010110;
assign LUT_3[52760] = 32'b00000000000000010001101100100101;
assign LUT_3[52761] = 32'b00000000000000011000011000000010;
assign LUT_3[52762] = 32'b00000000000000010011110100001001;
assign LUT_3[52763] = 32'b00000000000000011010011111100110;
assign LUT_3[52764] = 32'b00000000000000001110111010011011;
assign LUT_3[52765] = 32'b00000000000000010101100101111000;
assign LUT_3[52766] = 32'b00000000000000010001000001111111;
assign LUT_3[52767] = 32'b00000000000000010111101101011100;
assign LUT_3[52768] = 32'b00000000000000001010001110111100;
assign LUT_3[52769] = 32'b00000000000000010000111010011001;
assign LUT_3[52770] = 32'b00000000000000001100010110100000;
assign LUT_3[52771] = 32'b00000000000000010011000001111101;
assign LUT_3[52772] = 32'b00000000000000000111011100110010;
assign LUT_3[52773] = 32'b00000000000000001110001000001111;
assign LUT_3[52774] = 32'b00000000000000001001100100010110;
assign LUT_3[52775] = 32'b00000000000000010000001111110011;
assign LUT_3[52776] = 32'b00000000000000001111101000000010;
assign LUT_3[52777] = 32'b00000000000000010110010011011111;
assign LUT_3[52778] = 32'b00000000000000010001101111100110;
assign LUT_3[52779] = 32'b00000000000000011000011011000011;
assign LUT_3[52780] = 32'b00000000000000001100110101111000;
assign LUT_3[52781] = 32'b00000000000000010011100001010101;
assign LUT_3[52782] = 32'b00000000000000001110111101011100;
assign LUT_3[52783] = 32'b00000000000000010101101000111001;
assign LUT_3[52784] = 32'b00000000000000001101100001111111;
assign LUT_3[52785] = 32'b00000000000000010100001101011100;
assign LUT_3[52786] = 32'b00000000000000001111101001100011;
assign LUT_3[52787] = 32'b00000000000000010110010101000000;
assign LUT_3[52788] = 32'b00000000000000001010101111110101;
assign LUT_3[52789] = 32'b00000000000000010001011011010010;
assign LUT_3[52790] = 32'b00000000000000001100110111011001;
assign LUT_3[52791] = 32'b00000000000000010011100010110110;
assign LUT_3[52792] = 32'b00000000000000010010111011000101;
assign LUT_3[52793] = 32'b00000000000000011001100110100010;
assign LUT_3[52794] = 32'b00000000000000010101000010101001;
assign LUT_3[52795] = 32'b00000000000000011011101110000110;
assign LUT_3[52796] = 32'b00000000000000010000001000111011;
assign LUT_3[52797] = 32'b00000000000000010110110100011000;
assign LUT_3[52798] = 32'b00000000000000010010010000011111;
assign LUT_3[52799] = 32'b00000000000000011000111011111100;
assign LUT_3[52800] = 32'b00000000000000001000111001000111;
assign LUT_3[52801] = 32'b00000000000000001111100100100100;
assign LUT_3[52802] = 32'b00000000000000001011000000101011;
assign LUT_3[52803] = 32'b00000000000000010001101100001000;
assign LUT_3[52804] = 32'b00000000000000000110000110111101;
assign LUT_3[52805] = 32'b00000000000000001100110010011010;
assign LUT_3[52806] = 32'b00000000000000001000001110100001;
assign LUT_3[52807] = 32'b00000000000000001110111001111110;
assign LUT_3[52808] = 32'b00000000000000001110010010001101;
assign LUT_3[52809] = 32'b00000000000000010100111101101010;
assign LUT_3[52810] = 32'b00000000000000010000011001110001;
assign LUT_3[52811] = 32'b00000000000000010111000101001110;
assign LUT_3[52812] = 32'b00000000000000001011100000000011;
assign LUT_3[52813] = 32'b00000000000000010010001011100000;
assign LUT_3[52814] = 32'b00000000000000001101100111100111;
assign LUT_3[52815] = 32'b00000000000000010100010011000100;
assign LUT_3[52816] = 32'b00000000000000001100001100001010;
assign LUT_3[52817] = 32'b00000000000000010010110111100111;
assign LUT_3[52818] = 32'b00000000000000001110010011101110;
assign LUT_3[52819] = 32'b00000000000000010100111111001011;
assign LUT_3[52820] = 32'b00000000000000001001011010000000;
assign LUT_3[52821] = 32'b00000000000000010000000101011101;
assign LUT_3[52822] = 32'b00000000000000001011100001100100;
assign LUT_3[52823] = 32'b00000000000000010010001101000001;
assign LUT_3[52824] = 32'b00000000000000010001100101010000;
assign LUT_3[52825] = 32'b00000000000000011000010000101101;
assign LUT_3[52826] = 32'b00000000000000010011101100110100;
assign LUT_3[52827] = 32'b00000000000000011010011000010001;
assign LUT_3[52828] = 32'b00000000000000001110110011000110;
assign LUT_3[52829] = 32'b00000000000000010101011110100011;
assign LUT_3[52830] = 32'b00000000000000010000111010101010;
assign LUT_3[52831] = 32'b00000000000000010111100110000111;
assign LUT_3[52832] = 32'b00000000000000001010000111100111;
assign LUT_3[52833] = 32'b00000000000000010000110011000100;
assign LUT_3[52834] = 32'b00000000000000001100001111001011;
assign LUT_3[52835] = 32'b00000000000000010010111010101000;
assign LUT_3[52836] = 32'b00000000000000000111010101011101;
assign LUT_3[52837] = 32'b00000000000000001110000000111010;
assign LUT_3[52838] = 32'b00000000000000001001011101000001;
assign LUT_3[52839] = 32'b00000000000000010000001000011110;
assign LUT_3[52840] = 32'b00000000000000001111100000101101;
assign LUT_3[52841] = 32'b00000000000000010110001100001010;
assign LUT_3[52842] = 32'b00000000000000010001101000010001;
assign LUT_3[52843] = 32'b00000000000000011000010011101110;
assign LUT_3[52844] = 32'b00000000000000001100101110100011;
assign LUT_3[52845] = 32'b00000000000000010011011010000000;
assign LUT_3[52846] = 32'b00000000000000001110110110000111;
assign LUT_3[52847] = 32'b00000000000000010101100001100100;
assign LUT_3[52848] = 32'b00000000000000001101011010101010;
assign LUT_3[52849] = 32'b00000000000000010100000110000111;
assign LUT_3[52850] = 32'b00000000000000001111100010001110;
assign LUT_3[52851] = 32'b00000000000000010110001101101011;
assign LUT_3[52852] = 32'b00000000000000001010101000100000;
assign LUT_3[52853] = 32'b00000000000000010001010011111101;
assign LUT_3[52854] = 32'b00000000000000001100110000000100;
assign LUT_3[52855] = 32'b00000000000000010011011011100001;
assign LUT_3[52856] = 32'b00000000000000010010110011110000;
assign LUT_3[52857] = 32'b00000000000000011001011111001101;
assign LUT_3[52858] = 32'b00000000000000010100111011010100;
assign LUT_3[52859] = 32'b00000000000000011011100110110001;
assign LUT_3[52860] = 32'b00000000000000010000000001100110;
assign LUT_3[52861] = 32'b00000000000000010110101101000011;
assign LUT_3[52862] = 32'b00000000000000010010001001001010;
assign LUT_3[52863] = 32'b00000000000000011000110100100111;
assign LUT_3[52864] = 32'b00000000000000001011001011011010;
assign LUT_3[52865] = 32'b00000000000000010001110110110111;
assign LUT_3[52866] = 32'b00000000000000001101010010111110;
assign LUT_3[52867] = 32'b00000000000000010011111110011011;
assign LUT_3[52868] = 32'b00000000000000001000011001010000;
assign LUT_3[52869] = 32'b00000000000000001111000100101101;
assign LUT_3[52870] = 32'b00000000000000001010100000110100;
assign LUT_3[52871] = 32'b00000000000000010001001100010001;
assign LUT_3[52872] = 32'b00000000000000010000100100100000;
assign LUT_3[52873] = 32'b00000000000000010111001111111101;
assign LUT_3[52874] = 32'b00000000000000010010101100000100;
assign LUT_3[52875] = 32'b00000000000000011001010111100001;
assign LUT_3[52876] = 32'b00000000000000001101110010010110;
assign LUT_3[52877] = 32'b00000000000000010100011101110011;
assign LUT_3[52878] = 32'b00000000000000001111111001111010;
assign LUT_3[52879] = 32'b00000000000000010110100101010111;
assign LUT_3[52880] = 32'b00000000000000001110011110011101;
assign LUT_3[52881] = 32'b00000000000000010101001001111010;
assign LUT_3[52882] = 32'b00000000000000010000100110000001;
assign LUT_3[52883] = 32'b00000000000000010111010001011110;
assign LUT_3[52884] = 32'b00000000000000001011101100010011;
assign LUT_3[52885] = 32'b00000000000000010010010111110000;
assign LUT_3[52886] = 32'b00000000000000001101110011110111;
assign LUT_3[52887] = 32'b00000000000000010100011111010100;
assign LUT_3[52888] = 32'b00000000000000010011110111100011;
assign LUT_3[52889] = 32'b00000000000000011010100011000000;
assign LUT_3[52890] = 32'b00000000000000010101111111000111;
assign LUT_3[52891] = 32'b00000000000000011100101010100100;
assign LUT_3[52892] = 32'b00000000000000010001000101011001;
assign LUT_3[52893] = 32'b00000000000000010111110000110110;
assign LUT_3[52894] = 32'b00000000000000010011001100111101;
assign LUT_3[52895] = 32'b00000000000000011001111000011010;
assign LUT_3[52896] = 32'b00000000000000001100011001111010;
assign LUT_3[52897] = 32'b00000000000000010011000101010111;
assign LUT_3[52898] = 32'b00000000000000001110100001011110;
assign LUT_3[52899] = 32'b00000000000000010101001100111011;
assign LUT_3[52900] = 32'b00000000000000001001100111110000;
assign LUT_3[52901] = 32'b00000000000000010000010011001101;
assign LUT_3[52902] = 32'b00000000000000001011101111010100;
assign LUT_3[52903] = 32'b00000000000000010010011010110001;
assign LUT_3[52904] = 32'b00000000000000010001110011000000;
assign LUT_3[52905] = 32'b00000000000000011000011110011101;
assign LUT_3[52906] = 32'b00000000000000010011111010100100;
assign LUT_3[52907] = 32'b00000000000000011010100110000001;
assign LUT_3[52908] = 32'b00000000000000001111000000110110;
assign LUT_3[52909] = 32'b00000000000000010101101100010011;
assign LUT_3[52910] = 32'b00000000000000010001001000011010;
assign LUT_3[52911] = 32'b00000000000000010111110011110111;
assign LUT_3[52912] = 32'b00000000000000001111101100111101;
assign LUT_3[52913] = 32'b00000000000000010110011000011010;
assign LUT_3[52914] = 32'b00000000000000010001110100100001;
assign LUT_3[52915] = 32'b00000000000000011000011111111110;
assign LUT_3[52916] = 32'b00000000000000001100111010110011;
assign LUT_3[52917] = 32'b00000000000000010011100110010000;
assign LUT_3[52918] = 32'b00000000000000001111000010010111;
assign LUT_3[52919] = 32'b00000000000000010101101101110100;
assign LUT_3[52920] = 32'b00000000000000010101000110000011;
assign LUT_3[52921] = 32'b00000000000000011011110001100000;
assign LUT_3[52922] = 32'b00000000000000010111001101100111;
assign LUT_3[52923] = 32'b00000000000000011101111001000100;
assign LUT_3[52924] = 32'b00000000000000010010010011111001;
assign LUT_3[52925] = 32'b00000000000000011000111111010110;
assign LUT_3[52926] = 32'b00000000000000010100011011011101;
assign LUT_3[52927] = 32'b00000000000000011011000110111010;
assign LUT_3[52928] = 32'b00000000000000001011000100000101;
assign LUT_3[52929] = 32'b00000000000000010001101111100010;
assign LUT_3[52930] = 32'b00000000000000001101001011101001;
assign LUT_3[52931] = 32'b00000000000000010011110111000110;
assign LUT_3[52932] = 32'b00000000000000001000010001111011;
assign LUT_3[52933] = 32'b00000000000000001110111101011000;
assign LUT_3[52934] = 32'b00000000000000001010011001011111;
assign LUT_3[52935] = 32'b00000000000000010001000100111100;
assign LUT_3[52936] = 32'b00000000000000010000011101001011;
assign LUT_3[52937] = 32'b00000000000000010111001000101000;
assign LUT_3[52938] = 32'b00000000000000010010100100101111;
assign LUT_3[52939] = 32'b00000000000000011001010000001100;
assign LUT_3[52940] = 32'b00000000000000001101101011000001;
assign LUT_3[52941] = 32'b00000000000000010100010110011110;
assign LUT_3[52942] = 32'b00000000000000001111110010100101;
assign LUT_3[52943] = 32'b00000000000000010110011110000010;
assign LUT_3[52944] = 32'b00000000000000001110010111001000;
assign LUT_3[52945] = 32'b00000000000000010101000010100101;
assign LUT_3[52946] = 32'b00000000000000010000011110101100;
assign LUT_3[52947] = 32'b00000000000000010111001010001001;
assign LUT_3[52948] = 32'b00000000000000001011100100111110;
assign LUT_3[52949] = 32'b00000000000000010010010000011011;
assign LUT_3[52950] = 32'b00000000000000001101101100100010;
assign LUT_3[52951] = 32'b00000000000000010100010111111111;
assign LUT_3[52952] = 32'b00000000000000010011110000001110;
assign LUT_3[52953] = 32'b00000000000000011010011011101011;
assign LUT_3[52954] = 32'b00000000000000010101110111110010;
assign LUT_3[52955] = 32'b00000000000000011100100011001111;
assign LUT_3[52956] = 32'b00000000000000010000111110000100;
assign LUT_3[52957] = 32'b00000000000000010111101001100001;
assign LUT_3[52958] = 32'b00000000000000010011000101101000;
assign LUT_3[52959] = 32'b00000000000000011001110001000101;
assign LUT_3[52960] = 32'b00000000000000001100010010100101;
assign LUT_3[52961] = 32'b00000000000000010010111110000010;
assign LUT_3[52962] = 32'b00000000000000001110011010001001;
assign LUT_3[52963] = 32'b00000000000000010101000101100110;
assign LUT_3[52964] = 32'b00000000000000001001100000011011;
assign LUT_3[52965] = 32'b00000000000000010000001011111000;
assign LUT_3[52966] = 32'b00000000000000001011100111111111;
assign LUT_3[52967] = 32'b00000000000000010010010011011100;
assign LUT_3[52968] = 32'b00000000000000010001101011101011;
assign LUT_3[52969] = 32'b00000000000000011000010111001000;
assign LUT_3[52970] = 32'b00000000000000010011110011001111;
assign LUT_3[52971] = 32'b00000000000000011010011110101100;
assign LUT_3[52972] = 32'b00000000000000001110111001100001;
assign LUT_3[52973] = 32'b00000000000000010101100100111110;
assign LUT_3[52974] = 32'b00000000000000010001000001000101;
assign LUT_3[52975] = 32'b00000000000000010111101100100010;
assign LUT_3[52976] = 32'b00000000000000001111100101101000;
assign LUT_3[52977] = 32'b00000000000000010110010001000101;
assign LUT_3[52978] = 32'b00000000000000010001101101001100;
assign LUT_3[52979] = 32'b00000000000000011000011000101001;
assign LUT_3[52980] = 32'b00000000000000001100110011011110;
assign LUT_3[52981] = 32'b00000000000000010011011110111011;
assign LUT_3[52982] = 32'b00000000000000001110111011000010;
assign LUT_3[52983] = 32'b00000000000000010101100110011111;
assign LUT_3[52984] = 32'b00000000000000010100111110101110;
assign LUT_3[52985] = 32'b00000000000000011011101010001011;
assign LUT_3[52986] = 32'b00000000000000010111000110010010;
assign LUT_3[52987] = 32'b00000000000000011101110001101111;
assign LUT_3[52988] = 32'b00000000000000010010001100100100;
assign LUT_3[52989] = 32'b00000000000000011000111000000001;
assign LUT_3[52990] = 32'b00000000000000010100010100001000;
assign LUT_3[52991] = 32'b00000000000000011010111111100101;
assign LUT_3[52992] = 32'b00000000000000000101001111111101;
assign LUT_3[52993] = 32'b00000000000000001011111011011010;
assign LUT_3[52994] = 32'b00000000000000000111010111100001;
assign LUT_3[52995] = 32'b00000000000000001110000010111110;
assign LUT_3[52996] = 32'b00000000000000000010011101110011;
assign LUT_3[52997] = 32'b00000000000000001001001001010000;
assign LUT_3[52998] = 32'b00000000000000000100100101010111;
assign LUT_3[52999] = 32'b00000000000000001011010000110100;
assign LUT_3[53000] = 32'b00000000000000001010101001000011;
assign LUT_3[53001] = 32'b00000000000000010001010100100000;
assign LUT_3[53002] = 32'b00000000000000001100110000100111;
assign LUT_3[53003] = 32'b00000000000000010011011100000100;
assign LUT_3[53004] = 32'b00000000000000000111110110111001;
assign LUT_3[53005] = 32'b00000000000000001110100010010110;
assign LUT_3[53006] = 32'b00000000000000001001111110011101;
assign LUT_3[53007] = 32'b00000000000000010000101001111010;
assign LUT_3[53008] = 32'b00000000000000001000100011000000;
assign LUT_3[53009] = 32'b00000000000000001111001110011101;
assign LUT_3[53010] = 32'b00000000000000001010101010100100;
assign LUT_3[53011] = 32'b00000000000000010001010110000001;
assign LUT_3[53012] = 32'b00000000000000000101110000110110;
assign LUT_3[53013] = 32'b00000000000000001100011100010011;
assign LUT_3[53014] = 32'b00000000000000000111111000011010;
assign LUT_3[53015] = 32'b00000000000000001110100011110111;
assign LUT_3[53016] = 32'b00000000000000001101111100000110;
assign LUT_3[53017] = 32'b00000000000000010100100111100011;
assign LUT_3[53018] = 32'b00000000000000010000000011101010;
assign LUT_3[53019] = 32'b00000000000000010110101111000111;
assign LUT_3[53020] = 32'b00000000000000001011001001111100;
assign LUT_3[53021] = 32'b00000000000000010001110101011001;
assign LUT_3[53022] = 32'b00000000000000001101010001100000;
assign LUT_3[53023] = 32'b00000000000000010011111100111101;
assign LUT_3[53024] = 32'b00000000000000000110011110011101;
assign LUT_3[53025] = 32'b00000000000000001101001001111010;
assign LUT_3[53026] = 32'b00000000000000001000100110000001;
assign LUT_3[53027] = 32'b00000000000000001111010001011110;
assign LUT_3[53028] = 32'b00000000000000000011101100010011;
assign LUT_3[53029] = 32'b00000000000000001010010111110000;
assign LUT_3[53030] = 32'b00000000000000000101110011110111;
assign LUT_3[53031] = 32'b00000000000000001100011111010100;
assign LUT_3[53032] = 32'b00000000000000001011110111100011;
assign LUT_3[53033] = 32'b00000000000000010010100011000000;
assign LUT_3[53034] = 32'b00000000000000001101111111000111;
assign LUT_3[53035] = 32'b00000000000000010100101010100100;
assign LUT_3[53036] = 32'b00000000000000001001000101011001;
assign LUT_3[53037] = 32'b00000000000000001111110000110110;
assign LUT_3[53038] = 32'b00000000000000001011001100111101;
assign LUT_3[53039] = 32'b00000000000000010001111000011010;
assign LUT_3[53040] = 32'b00000000000000001001110001100000;
assign LUT_3[53041] = 32'b00000000000000010000011100111101;
assign LUT_3[53042] = 32'b00000000000000001011111001000100;
assign LUT_3[53043] = 32'b00000000000000010010100100100001;
assign LUT_3[53044] = 32'b00000000000000000110111111010110;
assign LUT_3[53045] = 32'b00000000000000001101101010110011;
assign LUT_3[53046] = 32'b00000000000000001001000110111010;
assign LUT_3[53047] = 32'b00000000000000001111110010010111;
assign LUT_3[53048] = 32'b00000000000000001111001010100110;
assign LUT_3[53049] = 32'b00000000000000010101110110000011;
assign LUT_3[53050] = 32'b00000000000000010001010010001010;
assign LUT_3[53051] = 32'b00000000000000010111111101100111;
assign LUT_3[53052] = 32'b00000000000000001100011000011100;
assign LUT_3[53053] = 32'b00000000000000010011000011111001;
assign LUT_3[53054] = 32'b00000000000000001110100000000000;
assign LUT_3[53055] = 32'b00000000000000010101001011011101;
assign LUT_3[53056] = 32'b00000000000000000101001000101000;
assign LUT_3[53057] = 32'b00000000000000001011110100000101;
assign LUT_3[53058] = 32'b00000000000000000111010000001100;
assign LUT_3[53059] = 32'b00000000000000001101111011101001;
assign LUT_3[53060] = 32'b00000000000000000010010110011110;
assign LUT_3[53061] = 32'b00000000000000001001000001111011;
assign LUT_3[53062] = 32'b00000000000000000100011110000010;
assign LUT_3[53063] = 32'b00000000000000001011001001011111;
assign LUT_3[53064] = 32'b00000000000000001010100001101110;
assign LUT_3[53065] = 32'b00000000000000010001001101001011;
assign LUT_3[53066] = 32'b00000000000000001100101001010010;
assign LUT_3[53067] = 32'b00000000000000010011010100101111;
assign LUT_3[53068] = 32'b00000000000000000111101111100100;
assign LUT_3[53069] = 32'b00000000000000001110011011000001;
assign LUT_3[53070] = 32'b00000000000000001001110111001000;
assign LUT_3[53071] = 32'b00000000000000010000100010100101;
assign LUT_3[53072] = 32'b00000000000000001000011011101011;
assign LUT_3[53073] = 32'b00000000000000001111000111001000;
assign LUT_3[53074] = 32'b00000000000000001010100011001111;
assign LUT_3[53075] = 32'b00000000000000010001001110101100;
assign LUT_3[53076] = 32'b00000000000000000101101001100001;
assign LUT_3[53077] = 32'b00000000000000001100010100111110;
assign LUT_3[53078] = 32'b00000000000000000111110001000101;
assign LUT_3[53079] = 32'b00000000000000001110011100100010;
assign LUT_3[53080] = 32'b00000000000000001101110100110001;
assign LUT_3[53081] = 32'b00000000000000010100100000001110;
assign LUT_3[53082] = 32'b00000000000000001111111100010101;
assign LUT_3[53083] = 32'b00000000000000010110100111110010;
assign LUT_3[53084] = 32'b00000000000000001011000010100111;
assign LUT_3[53085] = 32'b00000000000000010001101110000100;
assign LUT_3[53086] = 32'b00000000000000001101001010001011;
assign LUT_3[53087] = 32'b00000000000000010011110101101000;
assign LUT_3[53088] = 32'b00000000000000000110010111001000;
assign LUT_3[53089] = 32'b00000000000000001101000010100101;
assign LUT_3[53090] = 32'b00000000000000001000011110101100;
assign LUT_3[53091] = 32'b00000000000000001111001010001001;
assign LUT_3[53092] = 32'b00000000000000000011100100111110;
assign LUT_3[53093] = 32'b00000000000000001010010000011011;
assign LUT_3[53094] = 32'b00000000000000000101101100100010;
assign LUT_3[53095] = 32'b00000000000000001100010111111111;
assign LUT_3[53096] = 32'b00000000000000001011110000001110;
assign LUT_3[53097] = 32'b00000000000000010010011011101011;
assign LUT_3[53098] = 32'b00000000000000001101110111110010;
assign LUT_3[53099] = 32'b00000000000000010100100011001111;
assign LUT_3[53100] = 32'b00000000000000001000111110000100;
assign LUT_3[53101] = 32'b00000000000000001111101001100001;
assign LUT_3[53102] = 32'b00000000000000001011000101101000;
assign LUT_3[53103] = 32'b00000000000000010001110001000101;
assign LUT_3[53104] = 32'b00000000000000001001101010001011;
assign LUT_3[53105] = 32'b00000000000000010000010101101000;
assign LUT_3[53106] = 32'b00000000000000001011110001101111;
assign LUT_3[53107] = 32'b00000000000000010010011101001100;
assign LUT_3[53108] = 32'b00000000000000000110111000000001;
assign LUT_3[53109] = 32'b00000000000000001101100011011110;
assign LUT_3[53110] = 32'b00000000000000001000111111100101;
assign LUT_3[53111] = 32'b00000000000000001111101011000010;
assign LUT_3[53112] = 32'b00000000000000001111000011010001;
assign LUT_3[53113] = 32'b00000000000000010101101110101110;
assign LUT_3[53114] = 32'b00000000000000010001001010110101;
assign LUT_3[53115] = 32'b00000000000000010111110110010010;
assign LUT_3[53116] = 32'b00000000000000001100010001000111;
assign LUT_3[53117] = 32'b00000000000000010010111100100100;
assign LUT_3[53118] = 32'b00000000000000001110011000101011;
assign LUT_3[53119] = 32'b00000000000000010101000100001000;
assign LUT_3[53120] = 32'b00000000000000000111011010111011;
assign LUT_3[53121] = 32'b00000000000000001110000110011000;
assign LUT_3[53122] = 32'b00000000000000001001100010011111;
assign LUT_3[53123] = 32'b00000000000000010000001101111100;
assign LUT_3[53124] = 32'b00000000000000000100101000110001;
assign LUT_3[53125] = 32'b00000000000000001011010100001110;
assign LUT_3[53126] = 32'b00000000000000000110110000010101;
assign LUT_3[53127] = 32'b00000000000000001101011011110010;
assign LUT_3[53128] = 32'b00000000000000001100110100000001;
assign LUT_3[53129] = 32'b00000000000000010011011111011110;
assign LUT_3[53130] = 32'b00000000000000001110111011100101;
assign LUT_3[53131] = 32'b00000000000000010101100111000010;
assign LUT_3[53132] = 32'b00000000000000001010000001110111;
assign LUT_3[53133] = 32'b00000000000000010000101101010100;
assign LUT_3[53134] = 32'b00000000000000001100001001011011;
assign LUT_3[53135] = 32'b00000000000000010010110100111000;
assign LUT_3[53136] = 32'b00000000000000001010101101111110;
assign LUT_3[53137] = 32'b00000000000000010001011001011011;
assign LUT_3[53138] = 32'b00000000000000001100110101100010;
assign LUT_3[53139] = 32'b00000000000000010011100000111111;
assign LUT_3[53140] = 32'b00000000000000000111111011110100;
assign LUT_3[53141] = 32'b00000000000000001110100111010001;
assign LUT_3[53142] = 32'b00000000000000001010000011011000;
assign LUT_3[53143] = 32'b00000000000000010000101110110101;
assign LUT_3[53144] = 32'b00000000000000010000000111000100;
assign LUT_3[53145] = 32'b00000000000000010110110010100001;
assign LUT_3[53146] = 32'b00000000000000010010001110101000;
assign LUT_3[53147] = 32'b00000000000000011000111010000101;
assign LUT_3[53148] = 32'b00000000000000001101010100111010;
assign LUT_3[53149] = 32'b00000000000000010100000000010111;
assign LUT_3[53150] = 32'b00000000000000001111011100011110;
assign LUT_3[53151] = 32'b00000000000000010110000111111011;
assign LUT_3[53152] = 32'b00000000000000001000101001011011;
assign LUT_3[53153] = 32'b00000000000000001111010100111000;
assign LUT_3[53154] = 32'b00000000000000001010110000111111;
assign LUT_3[53155] = 32'b00000000000000010001011100011100;
assign LUT_3[53156] = 32'b00000000000000000101110111010001;
assign LUT_3[53157] = 32'b00000000000000001100100010101110;
assign LUT_3[53158] = 32'b00000000000000000111111110110101;
assign LUT_3[53159] = 32'b00000000000000001110101010010010;
assign LUT_3[53160] = 32'b00000000000000001110000010100001;
assign LUT_3[53161] = 32'b00000000000000010100101101111110;
assign LUT_3[53162] = 32'b00000000000000010000001010000101;
assign LUT_3[53163] = 32'b00000000000000010110110101100010;
assign LUT_3[53164] = 32'b00000000000000001011010000010111;
assign LUT_3[53165] = 32'b00000000000000010001111011110100;
assign LUT_3[53166] = 32'b00000000000000001101010111111011;
assign LUT_3[53167] = 32'b00000000000000010100000011011000;
assign LUT_3[53168] = 32'b00000000000000001011111100011110;
assign LUT_3[53169] = 32'b00000000000000010010100111111011;
assign LUT_3[53170] = 32'b00000000000000001110000100000010;
assign LUT_3[53171] = 32'b00000000000000010100101111011111;
assign LUT_3[53172] = 32'b00000000000000001001001010010100;
assign LUT_3[53173] = 32'b00000000000000001111110101110001;
assign LUT_3[53174] = 32'b00000000000000001011010001111000;
assign LUT_3[53175] = 32'b00000000000000010001111101010101;
assign LUT_3[53176] = 32'b00000000000000010001010101100100;
assign LUT_3[53177] = 32'b00000000000000011000000001000001;
assign LUT_3[53178] = 32'b00000000000000010011011101001000;
assign LUT_3[53179] = 32'b00000000000000011010001000100101;
assign LUT_3[53180] = 32'b00000000000000001110100011011010;
assign LUT_3[53181] = 32'b00000000000000010101001110110111;
assign LUT_3[53182] = 32'b00000000000000010000101010111110;
assign LUT_3[53183] = 32'b00000000000000010111010110011011;
assign LUT_3[53184] = 32'b00000000000000000111010011100110;
assign LUT_3[53185] = 32'b00000000000000001101111111000011;
assign LUT_3[53186] = 32'b00000000000000001001011011001010;
assign LUT_3[53187] = 32'b00000000000000010000000110100111;
assign LUT_3[53188] = 32'b00000000000000000100100001011100;
assign LUT_3[53189] = 32'b00000000000000001011001100111001;
assign LUT_3[53190] = 32'b00000000000000000110101001000000;
assign LUT_3[53191] = 32'b00000000000000001101010100011101;
assign LUT_3[53192] = 32'b00000000000000001100101100101100;
assign LUT_3[53193] = 32'b00000000000000010011011000001001;
assign LUT_3[53194] = 32'b00000000000000001110110100010000;
assign LUT_3[53195] = 32'b00000000000000010101011111101101;
assign LUT_3[53196] = 32'b00000000000000001001111010100010;
assign LUT_3[53197] = 32'b00000000000000010000100101111111;
assign LUT_3[53198] = 32'b00000000000000001100000010000110;
assign LUT_3[53199] = 32'b00000000000000010010101101100011;
assign LUT_3[53200] = 32'b00000000000000001010100110101001;
assign LUT_3[53201] = 32'b00000000000000010001010010000110;
assign LUT_3[53202] = 32'b00000000000000001100101110001101;
assign LUT_3[53203] = 32'b00000000000000010011011001101010;
assign LUT_3[53204] = 32'b00000000000000000111110100011111;
assign LUT_3[53205] = 32'b00000000000000001110011111111100;
assign LUT_3[53206] = 32'b00000000000000001001111100000011;
assign LUT_3[53207] = 32'b00000000000000010000100111100000;
assign LUT_3[53208] = 32'b00000000000000001111111111101111;
assign LUT_3[53209] = 32'b00000000000000010110101011001100;
assign LUT_3[53210] = 32'b00000000000000010010000111010011;
assign LUT_3[53211] = 32'b00000000000000011000110010110000;
assign LUT_3[53212] = 32'b00000000000000001101001101100101;
assign LUT_3[53213] = 32'b00000000000000010011111001000010;
assign LUT_3[53214] = 32'b00000000000000001111010101001001;
assign LUT_3[53215] = 32'b00000000000000010110000000100110;
assign LUT_3[53216] = 32'b00000000000000001000100010000110;
assign LUT_3[53217] = 32'b00000000000000001111001101100011;
assign LUT_3[53218] = 32'b00000000000000001010101001101010;
assign LUT_3[53219] = 32'b00000000000000010001010101000111;
assign LUT_3[53220] = 32'b00000000000000000101101111111100;
assign LUT_3[53221] = 32'b00000000000000001100011011011001;
assign LUT_3[53222] = 32'b00000000000000000111110111100000;
assign LUT_3[53223] = 32'b00000000000000001110100010111101;
assign LUT_3[53224] = 32'b00000000000000001101111011001100;
assign LUT_3[53225] = 32'b00000000000000010100100110101001;
assign LUT_3[53226] = 32'b00000000000000010000000010110000;
assign LUT_3[53227] = 32'b00000000000000010110101110001101;
assign LUT_3[53228] = 32'b00000000000000001011001001000010;
assign LUT_3[53229] = 32'b00000000000000010001110100011111;
assign LUT_3[53230] = 32'b00000000000000001101010000100110;
assign LUT_3[53231] = 32'b00000000000000010011111100000011;
assign LUT_3[53232] = 32'b00000000000000001011110101001001;
assign LUT_3[53233] = 32'b00000000000000010010100000100110;
assign LUT_3[53234] = 32'b00000000000000001101111100101101;
assign LUT_3[53235] = 32'b00000000000000010100101000001010;
assign LUT_3[53236] = 32'b00000000000000001001000010111111;
assign LUT_3[53237] = 32'b00000000000000001111101110011100;
assign LUT_3[53238] = 32'b00000000000000001011001010100011;
assign LUT_3[53239] = 32'b00000000000000010001110110000000;
assign LUT_3[53240] = 32'b00000000000000010001001110001111;
assign LUT_3[53241] = 32'b00000000000000010111111001101100;
assign LUT_3[53242] = 32'b00000000000000010011010101110011;
assign LUT_3[53243] = 32'b00000000000000011010000001010000;
assign LUT_3[53244] = 32'b00000000000000001110011100000101;
assign LUT_3[53245] = 32'b00000000000000010101000111100010;
assign LUT_3[53246] = 32'b00000000000000010000100011101001;
assign LUT_3[53247] = 32'b00000000000000010111001111000110;
assign LUT_3[53248] = 32'b00000000000000000001100001100000;
assign LUT_3[53249] = 32'b00000000000000001000001100111101;
assign LUT_3[53250] = 32'b00000000000000000011101001000100;
assign LUT_3[53251] = 32'b00000000000000001010010100100001;
assign LUT_3[53252] = 32'b11111111111111111110101111010110;
assign LUT_3[53253] = 32'b00000000000000000101011010110011;
assign LUT_3[53254] = 32'b00000000000000000000110110111010;
assign LUT_3[53255] = 32'b00000000000000000111100010010111;
assign LUT_3[53256] = 32'b00000000000000000110111010100110;
assign LUT_3[53257] = 32'b00000000000000001101100110000011;
assign LUT_3[53258] = 32'b00000000000000001001000010001010;
assign LUT_3[53259] = 32'b00000000000000001111101101100111;
assign LUT_3[53260] = 32'b00000000000000000100001000011100;
assign LUT_3[53261] = 32'b00000000000000001010110011111001;
assign LUT_3[53262] = 32'b00000000000000000110010000000000;
assign LUT_3[53263] = 32'b00000000000000001100111011011101;
assign LUT_3[53264] = 32'b00000000000000000100110100100011;
assign LUT_3[53265] = 32'b00000000000000001011100000000000;
assign LUT_3[53266] = 32'b00000000000000000110111100000111;
assign LUT_3[53267] = 32'b00000000000000001101100111100100;
assign LUT_3[53268] = 32'b00000000000000000010000010011001;
assign LUT_3[53269] = 32'b00000000000000001000101101110110;
assign LUT_3[53270] = 32'b00000000000000000100001001111101;
assign LUT_3[53271] = 32'b00000000000000001010110101011010;
assign LUT_3[53272] = 32'b00000000000000001010001101101001;
assign LUT_3[53273] = 32'b00000000000000010000111001000110;
assign LUT_3[53274] = 32'b00000000000000001100010101001101;
assign LUT_3[53275] = 32'b00000000000000010011000000101010;
assign LUT_3[53276] = 32'b00000000000000000111011011011111;
assign LUT_3[53277] = 32'b00000000000000001110000110111100;
assign LUT_3[53278] = 32'b00000000000000001001100011000011;
assign LUT_3[53279] = 32'b00000000000000010000001110100000;
assign LUT_3[53280] = 32'b00000000000000000010110000000000;
assign LUT_3[53281] = 32'b00000000000000001001011011011101;
assign LUT_3[53282] = 32'b00000000000000000100110111100100;
assign LUT_3[53283] = 32'b00000000000000001011100011000001;
assign LUT_3[53284] = 32'b11111111111111111111111101110110;
assign LUT_3[53285] = 32'b00000000000000000110101001010011;
assign LUT_3[53286] = 32'b00000000000000000010000101011010;
assign LUT_3[53287] = 32'b00000000000000001000110000110111;
assign LUT_3[53288] = 32'b00000000000000001000001001000110;
assign LUT_3[53289] = 32'b00000000000000001110110100100011;
assign LUT_3[53290] = 32'b00000000000000001010010000101010;
assign LUT_3[53291] = 32'b00000000000000010000111100000111;
assign LUT_3[53292] = 32'b00000000000000000101010110111100;
assign LUT_3[53293] = 32'b00000000000000001100000010011001;
assign LUT_3[53294] = 32'b00000000000000000111011110100000;
assign LUT_3[53295] = 32'b00000000000000001110001001111101;
assign LUT_3[53296] = 32'b00000000000000000110000011000011;
assign LUT_3[53297] = 32'b00000000000000001100101110100000;
assign LUT_3[53298] = 32'b00000000000000001000001010100111;
assign LUT_3[53299] = 32'b00000000000000001110110110000100;
assign LUT_3[53300] = 32'b00000000000000000011010000111001;
assign LUT_3[53301] = 32'b00000000000000001001111100010110;
assign LUT_3[53302] = 32'b00000000000000000101011000011101;
assign LUT_3[53303] = 32'b00000000000000001100000011111010;
assign LUT_3[53304] = 32'b00000000000000001011011100001001;
assign LUT_3[53305] = 32'b00000000000000010010000111100110;
assign LUT_3[53306] = 32'b00000000000000001101100011101101;
assign LUT_3[53307] = 32'b00000000000000010100001111001010;
assign LUT_3[53308] = 32'b00000000000000001000101001111111;
assign LUT_3[53309] = 32'b00000000000000001111010101011100;
assign LUT_3[53310] = 32'b00000000000000001010110001100011;
assign LUT_3[53311] = 32'b00000000000000010001011101000000;
assign LUT_3[53312] = 32'b00000000000000000001011010001011;
assign LUT_3[53313] = 32'b00000000000000001000000101101000;
assign LUT_3[53314] = 32'b00000000000000000011100001101111;
assign LUT_3[53315] = 32'b00000000000000001010001101001100;
assign LUT_3[53316] = 32'b11111111111111111110101000000001;
assign LUT_3[53317] = 32'b00000000000000000101010011011110;
assign LUT_3[53318] = 32'b00000000000000000000101111100101;
assign LUT_3[53319] = 32'b00000000000000000111011011000010;
assign LUT_3[53320] = 32'b00000000000000000110110011010001;
assign LUT_3[53321] = 32'b00000000000000001101011110101110;
assign LUT_3[53322] = 32'b00000000000000001000111010110101;
assign LUT_3[53323] = 32'b00000000000000001111100110010010;
assign LUT_3[53324] = 32'b00000000000000000100000001000111;
assign LUT_3[53325] = 32'b00000000000000001010101100100100;
assign LUT_3[53326] = 32'b00000000000000000110001000101011;
assign LUT_3[53327] = 32'b00000000000000001100110100001000;
assign LUT_3[53328] = 32'b00000000000000000100101101001110;
assign LUT_3[53329] = 32'b00000000000000001011011000101011;
assign LUT_3[53330] = 32'b00000000000000000110110100110010;
assign LUT_3[53331] = 32'b00000000000000001101100000001111;
assign LUT_3[53332] = 32'b00000000000000000001111011000100;
assign LUT_3[53333] = 32'b00000000000000001000100110100001;
assign LUT_3[53334] = 32'b00000000000000000100000010101000;
assign LUT_3[53335] = 32'b00000000000000001010101110000101;
assign LUT_3[53336] = 32'b00000000000000001010000110010100;
assign LUT_3[53337] = 32'b00000000000000010000110001110001;
assign LUT_3[53338] = 32'b00000000000000001100001101111000;
assign LUT_3[53339] = 32'b00000000000000010010111001010101;
assign LUT_3[53340] = 32'b00000000000000000111010100001010;
assign LUT_3[53341] = 32'b00000000000000001101111111100111;
assign LUT_3[53342] = 32'b00000000000000001001011011101110;
assign LUT_3[53343] = 32'b00000000000000010000000111001011;
assign LUT_3[53344] = 32'b00000000000000000010101000101011;
assign LUT_3[53345] = 32'b00000000000000001001010100001000;
assign LUT_3[53346] = 32'b00000000000000000100110000001111;
assign LUT_3[53347] = 32'b00000000000000001011011011101100;
assign LUT_3[53348] = 32'b11111111111111111111110110100001;
assign LUT_3[53349] = 32'b00000000000000000110100001111110;
assign LUT_3[53350] = 32'b00000000000000000001111110000101;
assign LUT_3[53351] = 32'b00000000000000001000101001100010;
assign LUT_3[53352] = 32'b00000000000000001000000001110001;
assign LUT_3[53353] = 32'b00000000000000001110101101001110;
assign LUT_3[53354] = 32'b00000000000000001010001001010101;
assign LUT_3[53355] = 32'b00000000000000010000110100110010;
assign LUT_3[53356] = 32'b00000000000000000101001111100111;
assign LUT_3[53357] = 32'b00000000000000001011111011000100;
assign LUT_3[53358] = 32'b00000000000000000111010111001011;
assign LUT_3[53359] = 32'b00000000000000001110000010101000;
assign LUT_3[53360] = 32'b00000000000000000101111011101110;
assign LUT_3[53361] = 32'b00000000000000001100100111001011;
assign LUT_3[53362] = 32'b00000000000000001000000011010010;
assign LUT_3[53363] = 32'b00000000000000001110101110101111;
assign LUT_3[53364] = 32'b00000000000000000011001001100100;
assign LUT_3[53365] = 32'b00000000000000001001110101000001;
assign LUT_3[53366] = 32'b00000000000000000101010001001000;
assign LUT_3[53367] = 32'b00000000000000001011111100100101;
assign LUT_3[53368] = 32'b00000000000000001011010100110100;
assign LUT_3[53369] = 32'b00000000000000010010000000010001;
assign LUT_3[53370] = 32'b00000000000000001101011100011000;
assign LUT_3[53371] = 32'b00000000000000010100000111110101;
assign LUT_3[53372] = 32'b00000000000000001000100010101010;
assign LUT_3[53373] = 32'b00000000000000001111001110000111;
assign LUT_3[53374] = 32'b00000000000000001010101010001110;
assign LUT_3[53375] = 32'b00000000000000010001010101101011;
assign LUT_3[53376] = 32'b00000000000000000011101100011110;
assign LUT_3[53377] = 32'b00000000000000001010010111111011;
assign LUT_3[53378] = 32'b00000000000000000101110100000010;
assign LUT_3[53379] = 32'b00000000000000001100011111011111;
assign LUT_3[53380] = 32'b00000000000000000000111010010100;
assign LUT_3[53381] = 32'b00000000000000000111100101110001;
assign LUT_3[53382] = 32'b00000000000000000011000001111000;
assign LUT_3[53383] = 32'b00000000000000001001101101010101;
assign LUT_3[53384] = 32'b00000000000000001001000101100100;
assign LUT_3[53385] = 32'b00000000000000001111110001000001;
assign LUT_3[53386] = 32'b00000000000000001011001101001000;
assign LUT_3[53387] = 32'b00000000000000010001111000100101;
assign LUT_3[53388] = 32'b00000000000000000110010011011010;
assign LUT_3[53389] = 32'b00000000000000001100111110110111;
assign LUT_3[53390] = 32'b00000000000000001000011010111110;
assign LUT_3[53391] = 32'b00000000000000001111000110011011;
assign LUT_3[53392] = 32'b00000000000000000110111111100001;
assign LUT_3[53393] = 32'b00000000000000001101101010111110;
assign LUT_3[53394] = 32'b00000000000000001001000111000101;
assign LUT_3[53395] = 32'b00000000000000001111110010100010;
assign LUT_3[53396] = 32'b00000000000000000100001101010111;
assign LUT_3[53397] = 32'b00000000000000001010111000110100;
assign LUT_3[53398] = 32'b00000000000000000110010100111011;
assign LUT_3[53399] = 32'b00000000000000001101000000011000;
assign LUT_3[53400] = 32'b00000000000000001100011000100111;
assign LUT_3[53401] = 32'b00000000000000010011000100000100;
assign LUT_3[53402] = 32'b00000000000000001110100000001011;
assign LUT_3[53403] = 32'b00000000000000010101001011101000;
assign LUT_3[53404] = 32'b00000000000000001001100110011101;
assign LUT_3[53405] = 32'b00000000000000010000010001111010;
assign LUT_3[53406] = 32'b00000000000000001011101110000001;
assign LUT_3[53407] = 32'b00000000000000010010011001011110;
assign LUT_3[53408] = 32'b00000000000000000100111010111110;
assign LUT_3[53409] = 32'b00000000000000001011100110011011;
assign LUT_3[53410] = 32'b00000000000000000111000010100010;
assign LUT_3[53411] = 32'b00000000000000001101101101111111;
assign LUT_3[53412] = 32'b00000000000000000010001000110100;
assign LUT_3[53413] = 32'b00000000000000001000110100010001;
assign LUT_3[53414] = 32'b00000000000000000100010000011000;
assign LUT_3[53415] = 32'b00000000000000001010111011110101;
assign LUT_3[53416] = 32'b00000000000000001010010100000100;
assign LUT_3[53417] = 32'b00000000000000010000111111100001;
assign LUT_3[53418] = 32'b00000000000000001100011011101000;
assign LUT_3[53419] = 32'b00000000000000010011000111000101;
assign LUT_3[53420] = 32'b00000000000000000111100001111010;
assign LUT_3[53421] = 32'b00000000000000001110001101010111;
assign LUT_3[53422] = 32'b00000000000000001001101001011110;
assign LUT_3[53423] = 32'b00000000000000010000010100111011;
assign LUT_3[53424] = 32'b00000000000000001000001110000001;
assign LUT_3[53425] = 32'b00000000000000001110111001011110;
assign LUT_3[53426] = 32'b00000000000000001010010101100101;
assign LUT_3[53427] = 32'b00000000000000010001000001000010;
assign LUT_3[53428] = 32'b00000000000000000101011011110111;
assign LUT_3[53429] = 32'b00000000000000001100000111010100;
assign LUT_3[53430] = 32'b00000000000000000111100011011011;
assign LUT_3[53431] = 32'b00000000000000001110001110111000;
assign LUT_3[53432] = 32'b00000000000000001101100111000111;
assign LUT_3[53433] = 32'b00000000000000010100010010100100;
assign LUT_3[53434] = 32'b00000000000000001111101110101011;
assign LUT_3[53435] = 32'b00000000000000010110011010001000;
assign LUT_3[53436] = 32'b00000000000000001010110100111101;
assign LUT_3[53437] = 32'b00000000000000010001100000011010;
assign LUT_3[53438] = 32'b00000000000000001100111100100001;
assign LUT_3[53439] = 32'b00000000000000010011100111111110;
assign LUT_3[53440] = 32'b00000000000000000011100101001001;
assign LUT_3[53441] = 32'b00000000000000001010010000100110;
assign LUT_3[53442] = 32'b00000000000000000101101100101101;
assign LUT_3[53443] = 32'b00000000000000001100011000001010;
assign LUT_3[53444] = 32'b00000000000000000000110010111111;
assign LUT_3[53445] = 32'b00000000000000000111011110011100;
assign LUT_3[53446] = 32'b00000000000000000010111010100011;
assign LUT_3[53447] = 32'b00000000000000001001100110000000;
assign LUT_3[53448] = 32'b00000000000000001000111110001111;
assign LUT_3[53449] = 32'b00000000000000001111101001101100;
assign LUT_3[53450] = 32'b00000000000000001011000101110011;
assign LUT_3[53451] = 32'b00000000000000010001110001010000;
assign LUT_3[53452] = 32'b00000000000000000110001100000101;
assign LUT_3[53453] = 32'b00000000000000001100110111100010;
assign LUT_3[53454] = 32'b00000000000000001000010011101001;
assign LUT_3[53455] = 32'b00000000000000001110111111000110;
assign LUT_3[53456] = 32'b00000000000000000110111000001100;
assign LUT_3[53457] = 32'b00000000000000001101100011101001;
assign LUT_3[53458] = 32'b00000000000000001000111111110000;
assign LUT_3[53459] = 32'b00000000000000001111101011001101;
assign LUT_3[53460] = 32'b00000000000000000100000110000010;
assign LUT_3[53461] = 32'b00000000000000001010110001011111;
assign LUT_3[53462] = 32'b00000000000000000110001101100110;
assign LUT_3[53463] = 32'b00000000000000001100111001000011;
assign LUT_3[53464] = 32'b00000000000000001100010001010010;
assign LUT_3[53465] = 32'b00000000000000010010111100101111;
assign LUT_3[53466] = 32'b00000000000000001110011000110110;
assign LUT_3[53467] = 32'b00000000000000010101000100010011;
assign LUT_3[53468] = 32'b00000000000000001001011111001000;
assign LUT_3[53469] = 32'b00000000000000010000001010100101;
assign LUT_3[53470] = 32'b00000000000000001011100110101100;
assign LUT_3[53471] = 32'b00000000000000010010010010001001;
assign LUT_3[53472] = 32'b00000000000000000100110011101001;
assign LUT_3[53473] = 32'b00000000000000001011011111000110;
assign LUT_3[53474] = 32'b00000000000000000110111011001101;
assign LUT_3[53475] = 32'b00000000000000001101100110101010;
assign LUT_3[53476] = 32'b00000000000000000010000001011111;
assign LUT_3[53477] = 32'b00000000000000001000101100111100;
assign LUT_3[53478] = 32'b00000000000000000100001001000011;
assign LUT_3[53479] = 32'b00000000000000001010110100100000;
assign LUT_3[53480] = 32'b00000000000000001010001100101111;
assign LUT_3[53481] = 32'b00000000000000010000111000001100;
assign LUT_3[53482] = 32'b00000000000000001100010100010011;
assign LUT_3[53483] = 32'b00000000000000010010111111110000;
assign LUT_3[53484] = 32'b00000000000000000111011010100101;
assign LUT_3[53485] = 32'b00000000000000001110000110000010;
assign LUT_3[53486] = 32'b00000000000000001001100010001001;
assign LUT_3[53487] = 32'b00000000000000010000001101100110;
assign LUT_3[53488] = 32'b00000000000000001000000110101100;
assign LUT_3[53489] = 32'b00000000000000001110110010001001;
assign LUT_3[53490] = 32'b00000000000000001010001110010000;
assign LUT_3[53491] = 32'b00000000000000010000111001101101;
assign LUT_3[53492] = 32'b00000000000000000101010100100010;
assign LUT_3[53493] = 32'b00000000000000001011111111111111;
assign LUT_3[53494] = 32'b00000000000000000111011100000110;
assign LUT_3[53495] = 32'b00000000000000001110000111100011;
assign LUT_3[53496] = 32'b00000000000000001101011111110010;
assign LUT_3[53497] = 32'b00000000000000010100001011001111;
assign LUT_3[53498] = 32'b00000000000000001111100111010110;
assign LUT_3[53499] = 32'b00000000000000010110010010110011;
assign LUT_3[53500] = 32'b00000000000000001010101101101000;
assign LUT_3[53501] = 32'b00000000000000010001011001000101;
assign LUT_3[53502] = 32'b00000000000000001100110101001100;
assign LUT_3[53503] = 32'b00000000000000010011100000101001;
assign LUT_3[53504] = 32'b11111111111111111101110001000001;
assign LUT_3[53505] = 32'b00000000000000000100011100011110;
assign LUT_3[53506] = 32'b11111111111111111111111000100101;
assign LUT_3[53507] = 32'b00000000000000000110100100000010;
assign LUT_3[53508] = 32'b11111111111111111010111110110111;
assign LUT_3[53509] = 32'b00000000000000000001101010010100;
assign LUT_3[53510] = 32'b11111111111111111101000110011011;
assign LUT_3[53511] = 32'b00000000000000000011110001111000;
assign LUT_3[53512] = 32'b00000000000000000011001010000111;
assign LUT_3[53513] = 32'b00000000000000001001110101100100;
assign LUT_3[53514] = 32'b00000000000000000101010001101011;
assign LUT_3[53515] = 32'b00000000000000001011111101001000;
assign LUT_3[53516] = 32'b00000000000000000000010111111101;
assign LUT_3[53517] = 32'b00000000000000000111000011011010;
assign LUT_3[53518] = 32'b00000000000000000010011111100001;
assign LUT_3[53519] = 32'b00000000000000001001001010111110;
assign LUT_3[53520] = 32'b00000000000000000001000100000100;
assign LUT_3[53521] = 32'b00000000000000000111101111100001;
assign LUT_3[53522] = 32'b00000000000000000011001011101000;
assign LUT_3[53523] = 32'b00000000000000001001110111000101;
assign LUT_3[53524] = 32'b11111111111111111110010001111010;
assign LUT_3[53525] = 32'b00000000000000000100111101010111;
assign LUT_3[53526] = 32'b00000000000000000000011001011110;
assign LUT_3[53527] = 32'b00000000000000000111000100111011;
assign LUT_3[53528] = 32'b00000000000000000110011101001010;
assign LUT_3[53529] = 32'b00000000000000001101001000100111;
assign LUT_3[53530] = 32'b00000000000000001000100100101110;
assign LUT_3[53531] = 32'b00000000000000001111010000001011;
assign LUT_3[53532] = 32'b00000000000000000011101011000000;
assign LUT_3[53533] = 32'b00000000000000001010010110011101;
assign LUT_3[53534] = 32'b00000000000000000101110010100100;
assign LUT_3[53535] = 32'b00000000000000001100011110000001;
assign LUT_3[53536] = 32'b11111111111111111110111111100001;
assign LUT_3[53537] = 32'b00000000000000000101101010111110;
assign LUT_3[53538] = 32'b00000000000000000001000111000101;
assign LUT_3[53539] = 32'b00000000000000000111110010100010;
assign LUT_3[53540] = 32'b11111111111111111100001101010111;
assign LUT_3[53541] = 32'b00000000000000000010111000110100;
assign LUT_3[53542] = 32'b11111111111111111110010100111011;
assign LUT_3[53543] = 32'b00000000000000000101000000011000;
assign LUT_3[53544] = 32'b00000000000000000100011000100111;
assign LUT_3[53545] = 32'b00000000000000001011000100000100;
assign LUT_3[53546] = 32'b00000000000000000110100000001011;
assign LUT_3[53547] = 32'b00000000000000001101001011101000;
assign LUT_3[53548] = 32'b00000000000000000001100110011101;
assign LUT_3[53549] = 32'b00000000000000001000010001111010;
assign LUT_3[53550] = 32'b00000000000000000011101110000001;
assign LUT_3[53551] = 32'b00000000000000001010011001011110;
assign LUT_3[53552] = 32'b00000000000000000010010010100100;
assign LUT_3[53553] = 32'b00000000000000001000111110000001;
assign LUT_3[53554] = 32'b00000000000000000100011010001000;
assign LUT_3[53555] = 32'b00000000000000001011000101100101;
assign LUT_3[53556] = 32'b11111111111111111111100000011010;
assign LUT_3[53557] = 32'b00000000000000000110001011110111;
assign LUT_3[53558] = 32'b00000000000000000001100111111110;
assign LUT_3[53559] = 32'b00000000000000001000010011011011;
assign LUT_3[53560] = 32'b00000000000000000111101011101010;
assign LUT_3[53561] = 32'b00000000000000001110010111000111;
assign LUT_3[53562] = 32'b00000000000000001001110011001110;
assign LUT_3[53563] = 32'b00000000000000010000011110101011;
assign LUT_3[53564] = 32'b00000000000000000100111001100000;
assign LUT_3[53565] = 32'b00000000000000001011100100111101;
assign LUT_3[53566] = 32'b00000000000000000111000001000100;
assign LUT_3[53567] = 32'b00000000000000001101101100100001;
assign LUT_3[53568] = 32'b11111111111111111101101001101100;
assign LUT_3[53569] = 32'b00000000000000000100010101001001;
assign LUT_3[53570] = 32'b11111111111111111111110001010000;
assign LUT_3[53571] = 32'b00000000000000000110011100101101;
assign LUT_3[53572] = 32'b11111111111111111010110111100010;
assign LUT_3[53573] = 32'b00000000000000000001100010111111;
assign LUT_3[53574] = 32'b11111111111111111100111111000110;
assign LUT_3[53575] = 32'b00000000000000000011101010100011;
assign LUT_3[53576] = 32'b00000000000000000011000010110010;
assign LUT_3[53577] = 32'b00000000000000001001101110001111;
assign LUT_3[53578] = 32'b00000000000000000101001010010110;
assign LUT_3[53579] = 32'b00000000000000001011110101110011;
assign LUT_3[53580] = 32'b00000000000000000000010000101000;
assign LUT_3[53581] = 32'b00000000000000000110111100000101;
assign LUT_3[53582] = 32'b00000000000000000010011000001100;
assign LUT_3[53583] = 32'b00000000000000001001000011101001;
assign LUT_3[53584] = 32'b00000000000000000000111100101111;
assign LUT_3[53585] = 32'b00000000000000000111101000001100;
assign LUT_3[53586] = 32'b00000000000000000011000100010011;
assign LUT_3[53587] = 32'b00000000000000001001101111110000;
assign LUT_3[53588] = 32'b11111111111111111110001010100101;
assign LUT_3[53589] = 32'b00000000000000000100110110000010;
assign LUT_3[53590] = 32'b00000000000000000000010010001001;
assign LUT_3[53591] = 32'b00000000000000000110111101100110;
assign LUT_3[53592] = 32'b00000000000000000110010101110101;
assign LUT_3[53593] = 32'b00000000000000001101000001010010;
assign LUT_3[53594] = 32'b00000000000000001000011101011001;
assign LUT_3[53595] = 32'b00000000000000001111001000110110;
assign LUT_3[53596] = 32'b00000000000000000011100011101011;
assign LUT_3[53597] = 32'b00000000000000001010001111001000;
assign LUT_3[53598] = 32'b00000000000000000101101011001111;
assign LUT_3[53599] = 32'b00000000000000001100010110101100;
assign LUT_3[53600] = 32'b11111111111111111110111000001100;
assign LUT_3[53601] = 32'b00000000000000000101100011101001;
assign LUT_3[53602] = 32'b00000000000000000000111111110000;
assign LUT_3[53603] = 32'b00000000000000000111101011001101;
assign LUT_3[53604] = 32'b11111111111111111100000110000010;
assign LUT_3[53605] = 32'b00000000000000000010110001011111;
assign LUT_3[53606] = 32'b11111111111111111110001101100110;
assign LUT_3[53607] = 32'b00000000000000000100111001000011;
assign LUT_3[53608] = 32'b00000000000000000100010001010010;
assign LUT_3[53609] = 32'b00000000000000001010111100101111;
assign LUT_3[53610] = 32'b00000000000000000110011000110110;
assign LUT_3[53611] = 32'b00000000000000001101000100010011;
assign LUT_3[53612] = 32'b00000000000000000001011111001000;
assign LUT_3[53613] = 32'b00000000000000001000001010100101;
assign LUT_3[53614] = 32'b00000000000000000011100110101100;
assign LUT_3[53615] = 32'b00000000000000001010010010001001;
assign LUT_3[53616] = 32'b00000000000000000010001011001111;
assign LUT_3[53617] = 32'b00000000000000001000110110101100;
assign LUT_3[53618] = 32'b00000000000000000100010010110011;
assign LUT_3[53619] = 32'b00000000000000001010111110010000;
assign LUT_3[53620] = 32'b11111111111111111111011001000101;
assign LUT_3[53621] = 32'b00000000000000000110000100100010;
assign LUT_3[53622] = 32'b00000000000000000001100000101001;
assign LUT_3[53623] = 32'b00000000000000001000001100000110;
assign LUT_3[53624] = 32'b00000000000000000111100100010101;
assign LUT_3[53625] = 32'b00000000000000001110001111110010;
assign LUT_3[53626] = 32'b00000000000000001001101011111001;
assign LUT_3[53627] = 32'b00000000000000010000010111010110;
assign LUT_3[53628] = 32'b00000000000000000100110010001011;
assign LUT_3[53629] = 32'b00000000000000001011011101101000;
assign LUT_3[53630] = 32'b00000000000000000110111001101111;
assign LUT_3[53631] = 32'b00000000000000001101100101001100;
assign LUT_3[53632] = 32'b11111111111111111111111011111111;
assign LUT_3[53633] = 32'b00000000000000000110100111011100;
assign LUT_3[53634] = 32'b00000000000000000010000011100011;
assign LUT_3[53635] = 32'b00000000000000001000101111000000;
assign LUT_3[53636] = 32'b11111111111111111101001001110101;
assign LUT_3[53637] = 32'b00000000000000000011110101010010;
assign LUT_3[53638] = 32'b11111111111111111111010001011001;
assign LUT_3[53639] = 32'b00000000000000000101111100110110;
assign LUT_3[53640] = 32'b00000000000000000101010101000101;
assign LUT_3[53641] = 32'b00000000000000001100000000100010;
assign LUT_3[53642] = 32'b00000000000000000111011100101001;
assign LUT_3[53643] = 32'b00000000000000001110001000000110;
assign LUT_3[53644] = 32'b00000000000000000010100010111011;
assign LUT_3[53645] = 32'b00000000000000001001001110011000;
assign LUT_3[53646] = 32'b00000000000000000100101010011111;
assign LUT_3[53647] = 32'b00000000000000001011010101111100;
assign LUT_3[53648] = 32'b00000000000000000011001111000010;
assign LUT_3[53649] = 32'b00000000000000001001111010011111;
assign LUT_3[53650] = 32'b00000000000000000101010110100110;
assign LUT_3[53651] = 32'b00000000000000001100000010000011;
assign LUT_3[53652] = 32'b00000000000000000000011100111000;
assign LUT_3[53653] = 32'b00000000000000000111001000010101;
assign LUT_3[53654] = 32'b00000000000000000010100100011100;
assign LUT_3[53655] = 32'b00000000000000001001001111111001;
assign LUT_3[53656] = 32'b00000000000000001000101000001000;
assign LUT_3[53657] = 32'b00000000000000001111010011100101;
assign LUT_3[53658] = 32'b00000000000000001010101111101100;
assign LUT_3[53659] = 32'b00000000000000010001011011001001;
assign LUT_3[53660] = 32'b00000000000000000101110101111110;
assign LUT_3[53661] = 32'b00000000000000001100100001011011;
assign LUT_3[53662] = 32'b00000000000000000111111101100010;
assign LUT_3[53663] = 32'b00000000000000001110101000111111;
assign LUT_3[53664] = 32'b00000000000000000001001010011111;
assign LUT_3[53665] = 32'b00000000000000000111110101111100;
assign LUT_3[53666] = 32'b00000000000000000011010010000011;
assign LUT_3[53667] = 32'b00000000000000001001111101100000;
assign LUT_3[53668] = 32'b11111111111111111110011000010101;
assign LUT_3[53669] = 32'b00000000000000000101000011110010;
assign LUT_3[53670] = 32'b00000000000000000000011111111001;
assign LUT_3[53671] = 32'b00000000000000000111001011010110;
assign LUT_3[53672] = 32'b00000000000000000110100011100101;
assign LUT_3[53673] = 32'b00000000000000001101001111000010;
assign LUT_3[53674] = 32'b00000000000000001000101011001001;
assign LUT_3[53675] = 32'b00000000000000001111010110100110;
assign LUT_3[53676] = 32'b00000000000000000011110001011011;
assign LUT_3[53677] = 32'b00000000000000001010011100111000;
assign LUT_3[53678] = 32'b00000000000000000101111000111111;
assign LUT_3[53679] = 32'b00000000000000001100100100011100;
assign LUT_3[53680] = 32'b00000000000000000100011101100010;
assign LUT_3[53681] = 32'b00000000000000001011001000111111;
assign LUT_3[53682] = 32'b00000000000000000110100101000110;
assign LUT_3[53683] = 32'b00000000000000001101010000100011;
assign LUT_3[53684] = 32'b00000000000000000001101011011000;
assign LUT_3[53685] = 32'b00000000000000001000010110110101;
assign LUT_3[53686] = 32'b00000000000000000011110010111100;
assign LUT_3[53687] = 32'b00000000000000001010011110011001;
assign LUT_3[53688] = 32'b00000000000000001001110110101000;
assign LUT_3[53689] = 32'b00000000000000010000100010000101;
assign LUT_3[53690] = 32'b00000000000000001011111110001100;
assign LUT_3[53691] = 32'b00000000000000010010101001101001;
assign LUT_3[53692] = 32'b00000000000000000111000100011110;
assign LUT_3[53693] = 32'b00000000000000001101101111111011;
assign LUT_3[53694] = 32'b00000000000000001001001100000010;
assign LUT_3[53695] = 32'b00000000000000001111110111011111;
assign LUT_3[53696] = 32'b11111111111111111111110100101010;
assign LUT_3[53697] = 32'b00000000000000000110100000000111;
assign LUT_3[53698] = 32'b00000000000000000001111100001110;
assign LUT_3[53699] = 32'b00000000000000001000100111101011;
assign LUT_3[53700] = 32'b11111111111111111101000010100000;
assign LUT_3[53701] = 32'b00000000000000000011101101111101;
assign LUT_3[53702] = 32'b11111111111111111111001010000100;
assign LUT_3[53703] = 32'b00000000000000000101110101100001;
assign LUT_3[53704] = 32'b00000000000000000101001101110000;
assign LUT_3[53705] = 32'b00000000000000001011111001001101;
assign LUT_3[53706] = 32'b00000000000000000111010101010100;
assign LUT_3[53707] = 32'b00000000000000001110000000110001;
assign LUT_3[53708] = 32'b00000000000000000010011011100110;
assign LUT_3[53709] = 32'b00000000000000001001000111000011;
assign LUT_3[53710] = 32'b00000000000000000100100011001010;
assign LUT_3[53711] = 32'b00000000000000001011001110100111;
assign LUT_3[53712] = 32'b00000000000000000011000111101101;
assign LUT_3[53713] = 32'b00000000000000001001110011001010;
assign LUT_3[53714] = 32'b00000000000000000101001111010001;
assign LUT_3[53715] = 32'b00000000000000001011111010101110;
assign LUT_3[53716] = 32'b00000000000000000000010101100011;
assign LUT_3[53717] = 32'b00000000000000000111000001000000;
assign LUT_3[53718] = 32'b00000000000000000010011101000111;
assign LUT_3[53719] = 32'b00000000000000001001001000100100;
assign LUT_3[53720] = 32'b00000000000000001000100000110011;
assign LUT_3[53721] = 32'b00000000000000001111001100010000;
assign LUT_3[53722] = 32'b00000000000000001010101000010111;
assign LUT_3[53723] = 32'b00000000000000010001010011110100;
assign LUT_3[53724] = 32'b00000000000000000101101110101001;
assign LUT_3[53725] = 32'b00000000000000001100011010000110;
assign LUT_3[53726] = 32'b00000000000000000111110110001101;
assign LUT_3[53727] = 32'b00000000000000001110100001101010;
assign LUT_3[53728] = 32'b00000000000000000001000011001010;
assign LUT_3[53729] = 32'b00000000000000000111101110100111;
assign LUT_3[53730] = 32'b00000000000000000011001010101110;
assign LUT_3[53731] = 32'b00000000000000001001110110001011;
assign LUT_3[53732] = 32'b11111111111111111110010001000000;
assign LUT_3[53733] = 32'b00000000000000000100111100011101;
assign LUT_3[53734] = 32'b00000000000000000000011000100100;
assign LUT_3[53735] = 32'b00000000000000000111000100000001;
assign LUT_3[53736] = 32'b00000000000000000110011100010000;
assign LUT_3[53737] = 32'b00000000000000001101000111101101;
assign LUT_3[53738] = 32'b00000000000000001000100011110100;
assign LUT_3[53739] = 32'b00000000000000001111001111010001;
assign LUT_3[53740] = 32'b00000000000000000011101010000110;
assign LUT_3[53741] = 32'b00000000000000001010010101100011;
assign LUT_3[53742] = 32'b00000000000000000101110001101010;
assign LUT_3[53743] = 32'b00000000000000001100011101000111;
assign LUT_3[53744] = 32'b00000000000000000100010110001101;
assign LUT_3[53745] = 32'b00000000000000001011000001101010;
assign LUT_3[53746] = 32'b00000000000000000110011101110001;
assign LUT_3[53747] = 32'b00000000000000001101001001001110;
assign LUT_3[53748] = 32'b00000000000000000001100100000011;
assign LUT_3[53749] = 32'b00000000000000001000001111100000;
assign LUT_3[53750] = 32'b00000000000000000011101011100111;
assign LUT_3[53751] = 32'b00000000000000001010010111000100;
assign LUT_3[53752] = 32'b00000000000000001001101111010011;
assign LUT_3[53753] = 32'b00000000000000010000011010110000;
assign LUT_3[53754] = 32'b00000000000000001011110110110111;
assign LUT_3[53755] = 32'b00000000000000010010100010010100;
assign LUT_3[53756] = 32'b00000000000000000110111101001001;
assign LUT_3[53757] = 32'b00000000000000001101101000100110;
assign LUT_3[53758] = 32'b00000000000000001001000100101101;
assign LUT_3[53759] = 32'b00000000000000001111110000001010;
assign LUT_3[53760] = 32'b00000000000000000100110110101100;
assign LUT_3[53761] = 32'b00000000000000001011100010001001;
assign LUT_3[53762] = 32'b00000000000000000110111110010000;
assign LUT_3[53763] = 32'b00000000000000001101101001101101;
assign LUT_3[53764] = 32'b00000000000000000010000100100010;
assign LUT_3[53765] = 32'b00000000000000001000101111111111;
assign LUT_3[53766] = 32'b00000000000000000100001100000110;
assign LUT_3[53767] = 32'b00000000000000001010110111100011;
assign LUT_3[53768] = 32'b00000000000000001010001111110010;
assign LUT_3[53769] = 32'b00000000000000010000111011001111;
assign LUT_3[53770] = 32'b00000000000000001100010111010110;
assign LUT_3[53771] = 32'b00000000000000010011000010110011;
assign LUT_3[53772] = 32'b00000000000000000111011101101000;
assign LUT_3[53773] = 32'b00000000000000001110001001000101;
assign LUT_3[53774] = 32'b00000000000000001001100101001100;
assign LUT_3[53775] = 32'b00000000000000010000010000101001;
assign LUT_3[53776] = 32'b00000000000000001000001001101111;
assign LUT_3[53777] = 32'b00000000000000001110110101001100;
assign LUT_3[53778] = 32'b00000000000000001010010001010011;
assign LUT_3[53779] = 32'b00000000000000010000111100110000;
assign LUT_3[53780] = 32'b00000000000000000101010111100101;
assign LUT_3[53781] = 32'b00000000000000001100000011000010;
assign LUT_3[53782] = 32'b00000000000000000111011111001001;
assign LUT_3[53783] = 32'b00000000000000001110001010100110;
assign LUT_3[53784] = 32'b00000000000000001101100010110101;
assign LUT_3[53785] = 32'b00000000000000010100001110010010;
assign LUT_3[53786] = 32'b00000000000000001111101010011001;
assign LUT_3[53787] = 32'b00000000000000010110010101110110;
assign LUT_3[53788] = 32'b00000000000000001010110000101011;
assign LUT_3[53789] = 32'b00000000000000010001011100001000;
assign LUT_3[53790] = 32'b00000000000000001100111000001111;
assign LUT_3[53791] = 32'b00000000000000010011100011101100;
assign LUT_3[53792] = 32'b00000000000000000110000101001100;
assign LUT_3[53793] = 32'b00000000000000001100110000101001;
assign LUT_3[53794] = 32'b00000000000000001000001100110000;
assign LUT_3[53795] = 32'b00000000000000001110111000001101;
assign LUT_3[53796] = 32'b00000000000000000011010011000010;
assign LUT_3[53797] = 32'b00000000000000001001111110011111;
assign LUT_3[53798] = 32'b00000000000000000101011010100110;
assign LUT_3[53799] = 32'b00000000000000001100000110000011;
assign LUT_3[53800] = 32'b00000000000000001011011110010010;
assign LUT_3[53801] = 32'b00000000000000010010001001101111;
assign LUT_3[53802] = 32'b00000000000000001101100101110110;
assign LUT_3[53803] = 32'b00000000000000010100010001010011;
assign LUT_3[53804] = 32'b00000000000000001000101100001000;
assign LUT_3[53805] = 32'b00000000000000001111010111100101;
assign LUT_3[53806] = 32'b00000000000000001010110011101100;
assign LUT_3[53807] = 32'b00000000000000010001011111001001;
assign LUT_3[53808] = 32'b00000000000000001001011000001111;
assign LUT_3[53809] = 32'b00000000000000010000000011101100;
assign LUT_3[53810] = 32'b00000000000000001011011111110011;
assign LUT_3[53811] = 32'b00000000000000010010001011010000;
assign LUT_3[53812] = 32'b00000000000000000110100110000101;
assign LUT_3[53813] = 32'b00000000000000001101010001100010;
assign LUT_3[53814] = 32'b00000000000000001000101101101001;
assign LUT_3[53815] = 32'b00000000000000001111011001000110;
assign LUT_3[53816] = 32'b00000000000000001110110001010101;
assign LUT_3[53817] = 32'b00000000000000010101011100110010;
assign LUT_3[53818] = 32'b00000000000000010000111000111001;
assign LUT_3[53819] = 32'b00000000000000010111100100010110;
assign LUT_3[53820] = 32'b00000000000000001011111111001011;
assign LUT_3[53821] = 32'b00000000000000010010101010101000;
assign LUT_3[53822] = 32'b00000000000000001110000110101111;
assign LUT_3[53823] = 32'b00000000000000010100110010001100;
assign LUT_3[53824] = 32'b00000000000000000100101111010111;
assign LUT_3[53825] = 32'b00000000000000001011011010110100;
assign LUT_3[53826] = 32'b00000000000000000110110110111011;
assign LUT_3[53827] = 32'b00000000000000001101100010011000;
assign LUT_3[53828] = 32'b00000000000000000001111101001101;
assign LUT_3[53829] = 32'b00000000000000001000101000101010;
assign LUT_3[53830] = 32'b00000000000000000100000100110001;
assign LUT_3[53831] = 32'b00000000000000001010110000001110;
assign LUT_3[53832] = 32'b00000000000000001010001000011101;
assign LUT_3[53833] = 32'b00000000000000010000110011111010;
assign LUT_3[53834] = 32'b00000000000000001100010000000001;
assign LUT_3[53835] = 32'b00000000000000010010111011011110;
assign LUT_3[53836] = 32'b00000000000000000111010110010011;
assign LUT_3[53837] = 32'b00000000000000001110000001110000;
assign LUT_3[53838] = 32'b00000000000000001001011101110111;
assign LUT_3[53839] = 32'b00000000000000010000001001010100;
assign LUT_3[53840] = 32'b00000000000000001000000010011010;
assign LUT_3[53841] = 32'b00000000000000001110101101110111;
assign LUT_3[53842] = 32'b00000000000000001010001001111110;
assign LUT_3[53843] = 32'b00000000000000010000110101011011;
assign LUT_3[53844] = 32'b00000000000000000101010000010000;
assign LUT_3[53845] = 32'b00000000000000001011111011101101;
assign LUT_3[53846] = 32'b00000000000000000111010111110100;
assign LUT_3[53847] = 32'b00000000000000001110000011010001;
assign LUT_3[53848] = 32'b00000000000000001101011011100000;
assign LUT_3[53849] = 32'b00000000000000010100000110111101;
assign LUT_3[53850] = 32'b00000000000000001111100011000100;
assign LUT_3[53851] = 32'b00000000000000010110001110100001;
assign LUT_3[53852] = 32'b00000000000000001010101001010110;
assign LUT_3[53853] = 32'b00000000000000010001010100110011;
assign LUT_3[53854] = 32'b00000000000000001100110000111010;
assign LUT_3[53855] = 32'b00000000000000010011011100010111;
assign LUT_3[53856] = 32'b00000000000000000101111101110111;
assign LUT_3[53857] = 32'b00000000000000001100101001010100;
assign LUT_3[53858] = 32'b00000000000000001000000101011011;
assign LUT_3[53859] = 32'b00000000000000001110110000111000;
assign LUT_3[53860] = 32'b00000000000000000011001011101101;
assign LUT_3[53861] = 32'b00000000000000001001110111001010;
assign LUT_3[53862] = 32'b00000000000000000101010011010001;
assign LUT_3[53863] = 32'b00000000000000001011111110101110;
assign LUT_3[53864] = 32'b00000000000000001011010110111101;
assign LUT_3[53865] = 32'b00000000000000010010000010011010;
assign LUT_3[53866] = 32'b00000000000000001101011110100001;
assign LUT_3[53867] = 32'b00000000000000010100001001111110;
assign LUT_3[53868] = 32'b00000000000000001000100100110011;
assign LUT_3[53869] = 32'b00000000000000001111010000010000;
assign LUT_3[53870] = 32'b00000000000000001010101100010111;
assign LUT_3[53871] = 32'b00000000000000010001010111110100;
assign LUT_3[53872] = 32'b00000000000000001001010000111010;
assign LUT_3[53873] = 32'b00000000000000001111111100010111;
assign LUT_3[53874] = 32'b00000000000000001011011000011110;
assign LUT_3[53875] = 32'b00000000000000010010000011111011;
assign LUT_3[53876] = 32'b00000000000000000110011110110000;
assign LUT_3[53877] = 32'b00000000000000001101001010001101;
assign LUT_3[53878] = 32'b00000000000000001000100110010100;
assign LUT_3[53879] = 32'b00000000000000001111010001110001;
assign LUT_3[53880] = 32'b00000000000000001110101010000000;
assign LUT_3[53881] = 32'b00000000000000010101010101011101;
assign LUT_3[53882] = 32'b00000000000000010000110001100100;
assign LUT_3[53883] = 32'b00000000000000010111011101000001;
assign LUT_3[53884] = 32'b00000000000000001011110111110110;
assign LUT_3[53885] = 32'b00000000000000010010100011010011;
assign LUT_3[53886] = 32'b00000000000000001101111111011010;
assign LUT_3[53887] = 32'b00000000000000010100101010110111;
assign LUT_3[53888] = 32'b00000000000000000111000001101010;
assign LUT_3[53889] = 32'b00000000000000001101101101000111;
assign LUT_3[53890] = 32'b00000000000000001001001001001110;
assign LUT_3[53891] = 32'b00000000000000001111110100101011;
assign LUT_3[53892] = 32'b00000000000000000100001111100000;
assign LUT_3[53893] = 32'b00000000000000001010111010111101;
assign LUT_3[53894] = 32'b00000000000000000110010111000100;
assign LUT_3[53895] = 32'b00000000000000001101000010100001;
assign LUT_3[53896] = 32'b00000000000000001100011010110000;
assign LUT_3[53897] = 32'b00000000000000010011000110001101;
assign LUT_3[53898] = 32'b00000000000000001110100010010100;
assign LUT_3[53899] = 32'b00000000000000010101001101110001;
assign LUT_3[53900] = 32'b00000000000000001001101000100110;
assign LUT_3[53901] = 32'b00000000000000010000010100000011;
assign LUT_3[53902] = 32'b00000000000000001011110000001010;
assign LUT_3[53903] = 32'b00000000000000010010011011100111;
assign LUT_3[53904] = 32'b00000000000000001010010100101101;
assign LUT_3[53905] = 32'b00000000000000010001000000001010;
assign LUT_3[53906] = 32'b00000000000000001100011100010001;
assign LUT_3[53907] = 32'b00000000000000010011000111101110;
assign LUT_3[53908] = 32'b00000000000000000111100010100011;
assign LUT_3[53909] = 32'b00000000000000001110001110000000;
assign LUT_3[53910] = 32'b00000000000000001001101010000111;
assign LUT_3[53911] = 32'b00000000000000010000010101100100;
assign LUT_3[53912] = 32'b00000000000000001111101101110011;
assign LUT_3[53913] = 32'b00000000000000010110011001010000;
assign LUT_3[53914] = 32'b00000000000000010001110101010111;
assign LUT_3[53915] = 32'b00000000000000011000100000110100;
assign LUT_3[53916] = 32'b00000000000000001100111011101001;
assign LUT_3[53917] = 32'b00000000000000010011100111000110;
assign LUT_3[53918] = 32'b00000000000000001111000011001101;
assign LUT_3[53919] = 32'b00000000000000010101101110101010;
assign LUT_3[53920] = 32'b00000000000000001000010000001010;
assign LUT_3[53921] = 32'b00000000000000001110111011100111;
assign LUT_3[53922] = 32'b00000000000000001010010111101110;
assign LUT_3[53923] = 32'b00000000000000010001000011001011;
assign LUT_3[53924] = 32'b00000000000000000101011110000000;
assign LUT_3[53925] = 32'b00000000000000001100001001011101;
assign LUT_3[53926] = 32'b00000000000000000111100101100100;
assign LUT_3[53927] = 32'b00000000000000001110010001000001;
assign LUT_3[53928] = 32'b00000000000000001101101001010000;
assign LUT_3[53929] = 32'b00000000000000010100010100101101;
assign LUT_3[53930] = 32'b00000000000000001111110000110100;
assign LUT_3[53931] = 32'b00000000000000010110011100010001;
assign LUT_3[53932] = 32'b00000000000000001010110111000110;
assign LUT_3[53933] = 32'b00000000000000010001100010100011;
assign LUT_3[53934] = 32'b00000000000000001100111110101010;
assign LUT_3[53935] = 32'b00000000000000010011101010000111;
assign LUT_3[53936] = 32'b00000000000000001011100011001101;
assign LUT_3[53937] = 32'b00000000000000010010001110101010;
assign LUT_3[53938] = 32'b00000000000000001101101010110001;
assign LUT_3[53939] = 32'b00000000000000010100010110001110;
assign LUT_3[53940] = 32'b00000000000000001000110001000011;
assign LUT_3[53941] = 32'b00000000000000001111011100100000;
assign LUT_3[53942] = 32'b00000000000000001010111000100111;
assign LUT_3[53943] = 32'b00000000000000010001100100000100;
assign LUT_3[53944] = 32'b00000000000000010000111100010011;
assign LUT_3[53945] = 32'b00000000000000010111100111110000;
assign LUT_3[53946] = 32'b00000000000000010011000011110111;
assign LUT_3[53947] = 32'b00000000000000011001101111010100;
assign LUT_3[53948] = 32'b00000000000000001110001010001001;
assign LUT_3[53949] = 32'b00000000000000010100110101100110;
assign LUT_3[53950] = 32'b00000000000000010000010001101101;
assign LUT_3[53951] = 32'b00000000000000010110111101001010;
assign LUT_3[53952] = 32'b00000000000000000110111010010101;
assign LUT_3[53953] = 32'b00000000000000001101100101110010;
assign LUT_3[53954] = 32'b00000000000000001001000001111001;
assign LUT_3[53955] = 32'b00000000000000001111101101010110;
assign LUT_3[53956] = 32'b00000000000000000100001000001011;
assign LUT_3[53957] = 32'b00000000000000001010110011101000;
assign LUT_3[53958] = 32'b00000000000000000110001111101111;
assign LUT_3[53959] = 32'b00000000000000001100111011001100;
assign LUT_3[53960] = 32'b00000000000000001100010011011011;
assign LUT_3[53961] = 32'b00000000000000010010111110111000;
assign LUT_3[53962] = 32'b00000000000000001110011010111111;
assign LUT_3[53963] = 32'b00000000000000010101000110011100;
assign LUT_3[53964] = 32'b00000000000000001001100001010001;
assign LUT_3[53965] = 32'b00000000000000010000001100101110;
assign LUT_3[53966] = 32'b00000000000000001011101000110101;
assign LUT_3[53967] = 32'b00000000000000010010010100010010;
assign LUT_3[53968] = 32'b00000000000000001010001101011000;
assign LUT_3[53969] = 32'b00000000000000010000111000110101;
assign LUT_3[53970] = 32'b00000000000000001100010100111100;
assign LUT_3[53971] = 32'b00000000000000010011000000011001;
assign LUT_3[53972] = 32'b00000000000000000111011011001110;
assign LUT_3[53973] = 32'b00000000000000001110000110101011;
assign LUT_3[53974] = 32'b00000000000000001001100010110010;
assign LUT_3[53975] = 32'b00000000000000010000001110001111;
assign LUT_3[53976] = 32'b00000000000000001111100110011110;
assign LUT_3[53977] = 32'b00000000000000010110010001111011;
assign LUT_3[53978] = 32'b00000000000000010001101110000010;
assign LUT_3[53979] = 32'b00000000000000011000011001011111;
assign LUT_3[53980] = 32'b00000000000000001100110100010100;
assign LUT_3[53981] = 32'b00000000000000010011011111110001;
assign LUT_3[53982] = 32'b00000000000000001110111011111000;
assign LUT_3[53983] = 32'b00000000000000010101100111010101;
assign LUT_3[53984] = 32'b00000000000000001000001000110101;
assign LUT_3[53985] = 32'b00000000000000001110110100010010;
assign LUT_3[53986] = 32'b00000000000000001010010000011001;
assign LUT_3[53987] = 32'b00000000000000010000111011110110;
assign LUT_3[53988] = 32'b00000000000000000101010110101011;
assign LUT_3[53989] = 32'b00000000000000001100000010001000;
assign LUT_3[53990] = 32'b00000000000000000111011110001111;
assign LUT_3[53991] = 32'b00000000000000001110001001101100;
assign LUT_3[53992] = 32'b00000000000000001101100001111011;
assign LUT_3[53993] = 32'b00000000000000010100001101011000;
assign LUT_3[53994] = 32'b00000000000000001111101001011111;
assign LUT_3[53995] = 32'b00000000000000010110010100111100;
assign LUT_3[53996] = 32'b00000000000000001010101111110001;
assign LUT_3[53997] = 32'b00000000000000010001011011001110;
assign LUT_3[53998] = 32'b00000000000000001100110111010101;
assign LUT_3[53999] = 32'b00000000000000010011100010110010;
assign LUT_3[54000] = 32'b00000000000000001011011011111000;
assign LUT_3[54001] = 32'b00000000000000010010000111010101;
assign LUT_3[54002] = 32'b00000000000000001101100011011100;
assign LUT_3[54003] = 32'b00000000000000010100001110111001;
assign LUT_3[54004] = 32'b00000000000000001000101001101110;
assign LUT_3[54005] = 32'b00000000000000001111010101001011;
assign LUT_3[54006] = 32'b00000000000000001010110001010010;
assign LUT_3[54007] = 32'b00000000000000010001011100101111;
assign LUT_3[54008] = 32'b00000000000000010000110100111110;
assign LUT_3[54009] = 32'b00000000000000010111100000011011;
assign LUT_3[54010] = 32'b00000000000000010010111100100010;
assign LUT_3[54011] = 32'b00000000000000011001100111111111;
assign LUT_3[54012] = 32'b00000000000000001110000010110100;
assign LUT_3[54013] = 32'b00000000000000010100101110010001;
assign LUT_3[54014] = 32'b00000000000000010000001010011000;
assign LUT_3[54015] = 32'b00000000000000010110110101110101;
assign LUT_3[54016] = 32'b00000000000000000001000110001101;
assign LUT_3[54017] = 32'b00000000000000000111110001101010;
assign LUT_3[54018] = 32'b00000000000000000011001101110001;
assign LUT_3[54019] = 32'b00000000000000001001111001001110;
assign LUT_3[54020] = 32'b11111111111111111110010100000011;
assign LUT_3[54021] = 32'b00000000000000000100111111100000;
assign LUT_3[54022] = 32'b00000000000000000000011011100111;
assign LUT_3[54023] = 32'b00000000000000000111000111000100;
assign LUT_3[54024] = 32'b00000000000000000110011111010011;
assign LUT_3[54025] = 32'b00000000000000001101001010110000;
assign LUT_3[54026] = 32'b00000000000000001000100110110111;
assign LUT_3[54027] = 32'b00000000000000001111010010010100;
assign LUT_3[54028] = 32'b00000000000000000011101101001001;
assign LUT_3[54029] = 32'b00000000000000001010011000100110;
assign LUT_3[54030] = 32'b00000000000000000101110100101101;
assign LUT_3[54031] = 32'b00000000000000001100100000001010;
assign LUT_3[54032] = 32'b00000000000000000100011001010000;
assign LUT_3[54033] = 32'b00000000000000001011000100101101;
assign LUT_3[54034] = 32'b00000000000000000110100000110100;
assign LUT_3[54035] = 32'b00000000000000001101001100010001;
assign LUT_3[54036] = 32'b00000000000000000001100111000110;
assign LUT_3[54037] = 32'b00000000000000001000010010100011;
assign LUT_3[54038] = 32'b00000000000000000011101110101010;
assign LUT_3[54039] = 32'b00000000000000001010011010000111;
assign LUT_3[54040] = 32'b00000000000000001001110010010110;
assign LUT_3[54041] = 32'b00000000000000010000011101110011;
assign LUT_3[54042] = 32'b00000000000000001011111001111010;
assign LUT_3[54043] = 32'b00000000000000010010100101010111;
assign LUT_3[54044] = 32'b00000000000000000111000000001100;
assign LUT_3[54045] = 32'b00000000000000001101101011101001;
assign LUT_3[54046] = 32'b00000000000000001001000111110000;
assign LUT_3[54047] = 32'b00000000000000001111110011001101;
assign LUT_3[54048] = 32'b00000000000000000010010100101101;
assign LUT_3[54049] = 32'b00000000000000001001000000001010;
assign LUT_3[54050] = 32'b00000000000000000100011100010001;
assign LUT_3[54051] = 32'b00000000000000001011000111101110;
assign LUT_3[54052] = 32'b11111111111111111111100010100011;
assign LUT_3[54053] = 32'b00000000000000000110001110000000;
assign LUT_3[54054] = 32'b00000000000000000001101010000111;
assign LUT_3[54055] = 32'b00000000000000001000010101100100;
assign LUT_3[54056] = 32'b00000000000000000111101101110011;
assign LUT_3[54057] = 32'b00000000000000001110011001010000;
assign LUT_3[54058] = 32'b00000000000000001001110101010111;
assign LUT_3[54059] = 32'b00000000000000010000100000110100;
assign LUT_3[54060] = 32'b00000000000000000100111011101001;
assign LUT_3[54061] = 32'b00000000000000001011100111000110;
assign LUT_3[54062] = 32'b00000000000000000111000011001101;
assign LUT_3[54063] = 32'b00000000000000001101101110101010;
assign LUT_3[54064] = 32'b00000000000000000101100111110000;
assign LUT_3[54065] = 32'b00000000000000001100010011001101;
assign LUT_3[54066] = 32'b00000000000000000111101111010100;
assign LUT_3[54067] = 32'b00000000000000001110011010110001;
assign LUT_3[54068] = 32'b00000000000000000010110101100110;
assign LUT_3[54069] = 32'b00000000000000001001100001000011;
assign LUT_3[54070] = 32'b00000000000000000100111101001010;
assign LUT_3[54071] = 32'b00000000000000001011101000100111;
assign LUT_3[54072] = 32'b00000000000000001011000000110110;
assign LUT_3[54073] = 32'b00000000000000010001101100010011;
assign LUT_3[54074] = 32'b00000000000000001101001000011010;
assign LUT_3[54075] = 32'b00000000000000010011110011110111;
assign LUT_3[54076] = 32'b00000000000000001000001110101100;
assign LUT_3[54077] = 32'b00000000000000001110111010001001;
assign LUT_3[54078] = 32'b00000000000000001010010110010000;
assign LUT_3[54079] = 32'b00000000000000010001000001101101;
assign LUT_3[54080] = 32'b00000000000000000000111110111000;
assign LUT_3[54081] = 32'b00000000000000000111101010010101;
assign LUT_3[54082] = 32'b00000000000000000011000110011100;
assign LUT_3[54083] = 32'b00000000000000001001110001111001;
assign LUT_3[54084] = 32'b11111111111111111110001100101110;
assign LUT_3[54085] = 32'b00000000000000000100111000001011;
assign LUT_3[54086] = 32'b00000000000000000000010100010010;
assign LUT_3[54087] = 32'b00000000000000000110111111101111;
assign LUT_3[54088] = 32'b00000000000000000110010111111110;
assign LUT_3[54089] = 32'b00000000000000001101000011011011;
assign LUT_3[54090] = 32'b00000000000000001000011111100010;
assign LUT_3[54091] = 32'b00000000000000001111001010111111;
assign LUT_3[54092] = 32'b00000000000000000011100101110100;
assign LUT_3[54093] = 32'b00000000000000001010010001010001;
assign LUT_3[54094] = 32'b00000000000000000101101101011000;
assign LUT_3[54095] = 32'b00000000000000001100011000110101;
assign LUT_3[54096] = 32'b00000000000000000100010001111011;
assign LUT_3[54097] = 32'b00000000000000001010111101011000;
assign LUT_3[54098] = 32'b00000000000000000110011001011111;
assign LUT_3[54099] = 32'b00000000000000001101000100111100;
assign LUT_3[54100] = 32'b00000000000000000001011111110001;
assign LUT_3[54101] = 32'b00000000000000001000001011001110;
assign LUT_3[54102] = 32'b00000000000000000011100111010101;
assign LUT_3[54103] = 32'b00000000000000001010010010110010;
assign LUT_3[54104] = 32'b00000000000000001001101011000001;
assign LUT_3[54105] = 32'b00000000000000010000010110011110;
assign LUT_3[54106] = 32'b00000000000000001011110010100101;
assign LUT_3[54107] = 32'b00000000000000010010011110000010;
assign LUT_3[54108] = 32'b00000000000000000110111000110111;
assign LUT_3[54109] = 32'b00000000000000001101100100010100;
assign LUT_3[54110] = 32'b00000000000000001001000000011011;
assign LUT_3[54111] = 32'b00000000000000001111101011111000;
assign LUT_3[54112] = 32'b00000000000000000010001101011000;
assign LUT_3[54113] = 32'b00000000000000001000111000110101;
assign LUT_3[54114] = 32'b00000000000000000100010100111100;
assign LUT_3[54115] = 32'b00000000000000001011000000011001;
assign LUT_3[54116] = 32'b11111111111111111111011011001110;
assign LUT_3[54117] = 32'b00000000000000000110000110101011;
assign LUT_3[54118] = 32'b00000000000000000001100010110010;
assign LUT_3[54119] = 32'b00000000000000001000001110001111;
assign LUT_3[54120] = 32'b00000000000000000111100110011110;
assign LUT_3[54121] = 32'b00000000000000001110010001111011;
assign LUT_3[54122] = 32'b00000000000000001001101110000010;
assign LUT_3[54123] = 32'b00000000000000010000011001011111;
assign LUT_3[54124] = 32'b00000000000000000100110100010100;
assign LUT_3[54125] = 32'b00000000000000001011011111110001;
assign LUT_3[54126] = 32'b00000000000000000110111011111000;
assign LUT_3[54127] = 32'b00000000000000001101100111010101;
assign LUT_3[54128] = 32'b00000000000000000101100000011011;
assign LUT_3[54129] = 32'b00000000000000001100001011111000;
assign LUT_3[54130] = 32'b00000000000000000111100111111111;
assign LUT_3[54131] = 32'b00000000000000001110010011011100;
assign LUT_3[54132] = 32'b00000000000000000010101110010001;
assign LUT_3[54133] = 32'b00000000000000001001011001101110;
assign LUT_3[54134] = 32'b00000000000000000100110101110101;
assign LUT_3[54135] = 32'b00000000000000001011100001010010;
assign LUT_3[54136] = 32'b00000000000000001010111001100001;
assign LUT_3[54137] = 32'b00000000000000010001100100111110;
assign LUT_3[54138] = 32'b00000000000000001101000001000101;
assign LUT_3[54139] = 32'b00000000000000010011101100100010;
assign LUT_3[54140] = 32'b00000000000000001000000111010111;
assign LUT_3[54141] = 32'b00000000000000001110110010110100;
assign LUT_3[54142] = 32'b00000000000000001010001110111011;
assign LUT_3[54143] = 32'b00000000000000010000111010011000;
assign LUT_3[54144] = 32'b00000000000000000011010001001011;
assign LUT_3[54145] = 32'b00000000000000001001111100101000;
assign LUT_3[54146] = 32'b00000000000000000101011000101111;
assign LUT_3[54147] = 32'b00000000000000001100000100001100;
assign LUT_3[54148] = 32'b00000000000000000000011111000001;
assign LUT_3[54149] = 32'b00000000000000000111001010011110;
assign LUT_3[54150] = 32'b00000000000000000010100110100101;
assign LUT_3[54151] = 32'b00000000000000001001010010000010;
assign LUT_3[54152] = 32'b00000000000000001000101010010001;
assign LUT_3[54153] = 32'b00000000000000001111010101101110;
assign LUT_3[54154] = 32'b00000000000000001010110001110101;
assign LUT_3[54155] = 32'b00000000000000010001011101010010;
assign LUT_3[54156] = 32'b00000000000000000101111000000111;
assign LUT_3[54157] = 32'b00000000000000001100100011100100;
assign LUT_3[54158] = 32'b00000000000000000111111111101011;
assign LUT_3[54159] = 32'b00000000000000001110101011001000;
assign LUT_3[54160] = 32'b00000000000000000110100100001110;
assign LUT_3[54161] = 32'b00000000000000001101001111101011;
assign LUT_3[54162] = 32'b00000000000000001000101011110010;
assign LUT_3[54163] = 32'b00000000000000001111010111001111;
assign LUT_3[54164] = 32'b00000000000000000011110010000100;
assign LUT_3[54165] = 32'b00000000000000001010011101100001;
assign LUT_3[54166] = 32'b00000000000000000101111001101000;
assign LUT_3[54167] = 32'b00000000000000001100100101000101;
assign LUT_3[54168] = 32'b00000000000000001011111101010100;
assign LUT_3[54169] = 32'b00000000000000010010101000110001;
assign LUT_3[54170] = 32'b00000000000000001110000100111000;
assign LUT_3[54171] = 32'b00000000000000010100110000010101;
assign LUT_3[54172] = 32'b00000000000000001001001011001010;
assign LUT_3[54173] = 32'b00000000000000001111110110100111;
assign LUT_3[54174] = 32'b00000000000000001011010010101110;
assign LUT_3[54175] = 32'b00000000000000010001111110001011;
assign LUT_3[54176] = 32'b00000000000000000100011111101011;
assign LUT_3[54177] = 32'b00000000000000001011001011001000;
assign LUT_3[54178] = 32'b00000000000000000110100111001111;
assign LUT_3[54179] = 32'b00000000000000001101010010101100;
assign LUT_3[54180] = 32'b00000000000000000001101101100001;
assign LUT_3[54181] = 32'b00000000000000001000011000111110;
assign LUT_3[54182] = 32'b00000000000000000011110101000101;
assign LUT_3[54183] = 32'b00000000000000001010100000100010;
assign LUT_3[54184] = 32'b00000000000000001001111000110001;
assign LUT_3[54185] = 32'b00000000000000010000100100001110;
assign LUT_3[54186] = 32'b00000000000000001100000000010101;
assign LUT_3[54187] = 32'b00000000000000010010101011110010;
assign LUT_3[54188] = 32'b00000000000000000111000110100111;
assign LUT_3[54189] = 32'b00000000000000001101110010000100;
assign LUT_3[54190] = 32'b00000000000000001001001110001011;
assign LUT_3[54191] = 32'b00000000000000001111111001101000;
assign LUT_3[54192] = 32'b00000000000000000111110010101110;
assign LUT_3[54193] = 32'b00000000000000001110011110001011;
assign LUT_3[54194] = 32'b00000000000000001001111010010010;
assign LUT_3[54195] = 32'b00000000000000010000100101101111;
assign LUT_3[54196] = 32'b00000000000000000101000000100100;
assign LUT_3[54197] = 32'b00000000000000001011101100000001;
assign LUT_3[54198] = 32'b00000000000000000111001000001000;
assign LUT_3[54199] = 32'b00000000000000001101110011100101;
assign LUT_3[54200] = 32'b00000000000000001101001011110100;
assign LUT_3[54201] = 32'b00000000000000010011110111010001;
assign LUT_3[54202] = 32'b00000000000000001111010011011000;
assign LUT_3[54203] = 32'b00000000000000010101111110110101;
assign LUT_3[54204] = 32'b00000000000000001010011001101010;
assign LUT_3[54205] = 32'b00000000000000010001000101000111;
assign LUT_3[54206] = 32'b00000000000000001100100001001110;
assign LUT_3[54207] = 32'b00000000000000010011001100101011;
assign LUT_3[54208] = 32'b00000000000000000011001001110110;
assign LUT_3[54209] = 32'b00000000000000001001110101010011;
assign LUT_3[54210] = 32'b00000000000000000101010001011010;
assign LUT_3[54211] = 32'b00000000000000001011111100110111;
assign LUT_3[54212] = 32'b00000000000000000000010111101100;
assign LUT_3[54213] = 32'b00000000000000000111000011001001;
assign LUT_3[54214] = 32'b00000000000000000010011111010000;
assign LUT_3[54215] = 32'b00000000000000001001001010101101;
assign LUT_3[54216] = 32'b00000000000000001000100010111100;
assign LUT_3[54217] = 32'b00000000000000001111001110011001;
assign LUT_3[54218] = 32'b00000000000000001010101010100000;
assign LUT_3[54219] = 32'b00000000000000010001010101111101;
assign LUT_3[54220] = 32'b00000000000000000101110000110010;
assign LUT_3[54221] = 32'b00000000000000001100011100001111;
assign LUT_3[54222] = 32'b00000000000000000111111000010110;
assign LUT_3[54223] = 32'b00000000000000001110100011110011;
assign LUT_3[54224] = 32'b00000000000000000110011100111001;
assign LUT_3[54225] = 32'b00000000000000001101001000010110;
assign LUT_3[54226] = 32'b00000000000000001000100100011101;
assign LUT_3[54227] = 32'b00000000000000001111001111111010;
assign LUT_3[54228] = 32'b00000000000000000011101010101111;
assign LUT_3[54229] = 32'b00000000000000001010010110001100;
assign LUT_3[54230] = 32'b00000000000000000101110010010011;
assign LUT_3[54231] = 32'b00000000000000001100011101110000;
assign LUT_3[54232] = 32'b00000000000000001011110101111111;
assign LUT_3[54233] = 32'b00000000000000010010100001011100;
assign LUT_3[54234] = 32'b00000000000000001101111101100011;
assign LUT_3[54235] = 32'b00000000000000010100101001000000;
assign LUT_3[54236] = 32'b00000000000000001001000011110101;
assign LUT_3[54237] = 32'b00000000000000001111101111010010;
assign LUT_3[54238] = 32'b00000000000000001011001011011001;
assign LUT_3[54239] = 32'b00000000000000010001110110110110;
assign LUT_3[54240] = 32'b00000000000000000100011000010110;
assign LUT_3[54241] = 32'b00000000000000001011000011110011;
assign LUT_3[54242] = 32'b00000000000000000110011111111010;
assign LUT_3[54243] = 32'b00000000000000001101001011010111;
assign LUT_3[54244] = 32'b00000000000000000001100110001100;
assign LUT_3[54245] = 32'b00000000000000001000010001101001;
assign LUT_3[54246] = 32'b00000000000000000011101101110000;
assign LUT_3[54247] = 32'b00000000000000001010011001001101;
assign LUT_3[54248] = 32'b00000000000000001001110001011100;
assign LUT_3[54249] = 32'b00000000000000010000011100111001;
assign LUT_3[54250] = 32'b00000000000000001011111001000000;
assign LUT_3[54251] = 32'b00000000000000010010100100011101;
assign LUT_3[54252] = 32'b00000000000000000110111111010010;
assign LUT_3[54253] = 32'b00000000000000001101101010101111;
assign LUT_3[54254] = 32'b00000000000000001001000110110110;
assign LUT_3[54255] = 32'b00000000000000001111110010010011;
assign LUT_3[54256] = 32'b00000000000000000111101011011001;
assign LUT_3[54257] = 32'b00000000000000001110010110110110;
assign LUT_3[54258] = 32'b00000000000000001001110010111101;
assign LUT_3[54259] = 32'b00000000000000010000011110011010;
assign LUT_3[54260] = 32'b00000000000000000100111001001111;
assign LUT_3[54261] = 32'b00000000000000001011100100101100;
assign LUT_3[54262] = 32'b00000000000000000111000000110011;
assign LUT_3[54263] = 32'b00000000000000001101101100010000;
assign LUT_3[54264] = 32'b00000000000000001101000100011111;
assign LUT_3[54265] = 32'b00000000000000010011101111111100;
assign LUT_3[54266] = 32'b00000000000000001111001100000011;
assign LUT_3[54267] = 32'b00000000000000010101110111100000;
assign LUT_3[54268] = 32'b00000000000000001010010010010101;
assign LUT_3[54269] = 32'b00000000000000010000111101110010;
assign LUT_3[54270] = 32'b00000000000000001100011001111001;
assign LUT_3[54271] = 32'b00000000000000010011000101010110;
assign LUT_3[54272] = 32'b00000000000000001000000110011101;
assign LUT_3[54273] = 32'b00000000000000001110110001111010;
assign LUT_3[54274] = 32'b00000000000000001010001110000001;
assign LUT_3[54275] = 32'b00000000000000010000111001011110;
assign LUT_3[54276] = 32'b00000000000000000101010100010011;
assign LUT_3[54277] = 32'b00000000000000001011111111110000;
assign LUT_3[54278] = 32'b00000000000000000111011011110111;
assign LUT_3[54279] = 32'b00000000000000001110000111010100;
assign LUT_3[54280] = 32'b00000000000000001101011111100011;
assign LUT_3[54281] = 32'b00000000000000010100001011000000;
assign LUT_3[54282] = 32'b00000000000000001111100111000111;
assign LUT_3[54283] = 32'b00000000000000010110010010100100;
assign LUT_3[54284] = 32'b00000000000000001010101101011001;
assign LUT_3[54285] = 32'b00000000000000010001011000110110;
assign LUT_3[54286] = 32'b00000000000000001100110100111101;
assign LUT_3[54287] = 32'b00000000000000010011100000011010;
assign LUT_3[54288] = 32'b00000000000000001011011001100000;
assign LUT_3[54289] = 32'b00000000000000010010000100111101;
assign LUT_3[54290] = 32'b00000000000000001101100001000100;
assign LUT_3[54291] = 32'b00000000000000010100001100100001;
assign LUT_3[54292] = 32'b00000000000000001000100111010110;
assign LUT_3[54293] = 32'b00000000000000001111010010110011;
assign LUT_3[54294] = 32'b00000000000000001010101110111010;
assign LUT_3[54295] = 32'b00000000000000010001011010010111;
assign LUT_3[54296] = 32'b00000000000000010000110010100110;
assign LUT_3[54297] = 32'b00000000000000010111011110000011;
assign LUT_3[54298] = 32'b00000000000000010010111010001010;
assign LUT_3[54299] = 32'b00000000000000011001100101100111;
assign LUT_3[54300] = 32'b00000000000000001110000000011100;
assign LUT_3[54301] = 32'b00000000000000010100101011111001;
assign LUT_3[54302] = 32'b00000000000000010000001000000000;
assign LUT_3[54303] = 32'b00000000000000010110110011011101;
assign LUT_3[54304] = 32'b00000000000000001001010100111101;
assign LUT_3[54305] = 32'b00000000000000010000000000011010;
assign LUT_3[54306] = 32'b00000000000000001011011100100001;
assign LUT_3[54307] = 32'b00000000000000010010000111111110;
assign LUT_3[54308] = 32'b00000000000000000110100010110011;
assign LUT_3[54309] = 32'b00000000000000001101001110010000;
assign LUT_3[54310] = 32'b00000000000000001000101010010111;
assign LUT_3[54311] = 32'b00000000000000001111010101110100;
assign LUT_3[54312] = 32'b00000000000000001110101110000011;
assign LUT_3[54313] = 32'b00000000000000010101011001100000;
assign LUT_3[54314] = 32'b00000000000000010000110101100111;
assign LUT_3[54315] = 32'b00000000000000010111100001000100;
assign LUT_3[54316] = 32'b00000000000000001011111011111001;
assign LUT_3[54317] = 32'b00000000000000010010100111010110;
assign LUT_3[54318] = 32'b00000000000000001110000011011101;
assign LUT_3[54319] = 32'b00000000000000010100101110111010;
assign LUT_3[54320] = 32'b00000000000000001100101000000000;
assign LUT_3[54321] = 32'b00000000000000010011010011011101;
assign LUT_3[54322] = 32'b00000000000000001110101111100100;
assign LUT_3[54323] = 32'b00000000000000010101011011000001;
assign LUT_3[54324] = 32'b00000000000000001001110101110110;
assign LUT_3[54325] = 32'b00000000000000010000100001010011;
assign LUT_3[54326] = 32'b00000000000000001011111101011010;
assign LUT_3[54327] = 32'b00000000000000010010101000110111;
assign LUT_3[54328] = 32'b00000000000000010010000001000110;
assign LUT_3[54329] = 32'b00000000000000011000101100100011;
assign LUT_3[54330] = 32'b00000000000000010100001000101010;
assign LUT_3[54331] = 32'b00000000000000011010110100000111;
assign LUT_3[54332] = 32'b00000000000000001111001110111100;
assign LUT_3[54333] = 32'b00000000000000010101111010011001;
assign LUT_3[54334] = 32'b00000000000000010001010110100000;
assign LUT_3[54335] = 32'b00000000000000011000000001111101;
assign LUT_3[54336] = 32'b00000000000000000111111111001000;
assign LUT_3[54337] = 32'b00000000000000001110101010100101;
assign LUT_3[54338] = 32'b00000000000000001010000110101100;
assign LUT_3[54339] = 32'b00000000000000010000110010001001;
assign LUT_3[54340] = 32'b00000000000000000101001100111110;
assign LUT_3[54341] = 32'b00000000000000001011111000011011;
assign LUT_3[54342] = 32'b00000000000000000111010100100010;
assign LUT_3[54343] = 32'b00000000000000001101111111111111;
assign LUT_3[54344] = 32'b00000000000000001101011000001110;
assign LUT_3[54345] = 32'b00000000000000010100000011101011;
assign LUT_3[54346] = 32'b00000000000000001111011111110010;
assign LUT_3[54347] = 32'b00000000000000010110001011001111;
assign LUT_3[54348] = 32'b00000000000000001010100110000100;
assign LUT_3[54349] = 32'b00000000000000010001010001100001;
assign LUT_3[54350] = 32'b00000000000000001100101101101000;
assign LUT_3[54351] = 32'b00000000000000010011011001000101;
assign LUT_3[54352] = 32'b00000000000000001011010010001011;
assign LUT_3[54353] = 32'b00000000000000010001111101101000;
assign LUT_3[54354] = 32'b00000000000000001101011001101111;
assign LUT_3[54355] = 32'b00000000000000010100000101001100;
assign LUT_3[54356] = 32'b00000000000000001000100000000001;
assign LUT_3[54357] = 32'b00000000000000001111001011011110;
assign LUT_3[54358] = 32'b00000000000000001010100111100101;
assign LUT_3[54359] = 32'b00000000000000010001010011000010;
assign LUT_3[54360] = 32'b00000000000000010000101011010001;
assign LUT_3[54361] = 32'b00000000000000010111010110101110;
assign LUT_3[54362] = 32'b00000000000000010010110010110101;
assign LUT_3[54363] = 32'b00000000000000011001011110010010;
assign LUT_3[54364] = 32'b00000000000000001101111001000111;
assign LUT_3[54365] = 32'b00000000000000010100100100100100;
assign LUT_3[54366] = 32'b00000000000000010000000000101011;
assign LUT_3[54367] = 32'b00000000000000010110101100001000;
assign LUT_3[54368] = 32'b00000000000000001001001101101000;
assign LUT_3[54369] = 32'b00000000000000001111111001000101;
assign LUT_3[54370] = 32'b00000000000000001011010101001100;
assign LUT_3[54371] = 32'b00000000000000010010000000101001;
assign LUT_3[54372] = 32'b00000000000000000110011011011110;
assign LUT_3[54373] = 32'b00000000000000001101000110111011;
assign LUT_3[54374] = 32'b00000000000000001000100011000010;
assign LUT_3[54375] = 32'b00000000000000001111001110011111;
assign LUT_3[54376] = 32'b00000000000000001110100110101110;
assign LUT_3[54377] = 32'b00000000000000010101010010001011;
assign LUT_3[54378] = 32'b00000000000000010000101110010010;
assign LUT_3[54379] = 32'b00000000000000010111011001101111;
assign LUT_3[54380] = 32'b00000000000000001011110100100100;
assign LUT_3[54381] = 32'b00000000000000010010100000000001;
assign LUT_3[54382] = 32'b00000000000000001101111100001000;
assign LUT_3[54383] = 32'b00000000000000010100100111100101;
assign LUT_3[54384] = 32'b00000000000000001100100000101011;
assign LUT_3[54385] = 32'b00000000000000010011001100001000;
assign LUT_3[54386] = 32'b00000000000000001110101000001111;
assign LUT_3[54387] = 32'b00000000000000010101010011101100;
assign LUT_3[54388] = 32'b00000000000000001001101110100001;
assign LUT_3[54389] = 32'b00000000000000010000011001111110;
assign LUT_3[54390] = 32'b00000000000000001011110110000101;
assign LUT_3[54391] = 32'b00000000000000010010100001100010;
assign LUT_3[54392] = 32'b00000000000000010001111001110001;
assign LUT_3[54393] = 32'b00000000000000011000100101001110;
assign LUT_3[54394] = 32'b00000000000000010100000001010101;
assign LUT_3[54395] = 32'b00000000000000011010101100110010;
assign LUT_3[54396] = 32'b00000000000000001111000111100111;
assign LUT_3[54397] = 32'b00000000000000010101110011000100;
assign LUT_3[54398] = 32'b00000000000000010001001111001011;
assign LUT_3[54399] = 32'b00000000000000010111111010101000;
assign LUT_3[54400] = 32'b00000000000000001010010001011011;
assign LUT_3[54401] = 32'b00000000000000010000111100111000;
assign LUT_3[54402] = 32'b00000000000000001100011000111111;
assign LUT_3[54403] = 32'b00000000000000010011000100011100;
assign LUT_3[54404] = 32'b00000000000000000111011111010001;
assign LUT_3[54405] = 32'b00000000000000001110001010101110;
assign LUT_3[54406] = 32'b00000000000000001001100110110101;
assign LUT_3[54407] = 32'b00000000000000010000010010010010;
assign LUT_3[54408] = 32'b00000000000000001111101010100001;
assign LUT_3[54409] = 32'b00000000000000010110010101111110;
assign LUT_3[54410] = 32'b00000000000000010001110010000101;
assign LUT_3[54411] = 32'b00000000000000011000011101100010;
assign LUT_3[54412] = 32'b00000000000000001100111000010111;
assign LUT_3[54413] = 32'b00000000000000010011100011110100;
assign LUT_3[54414] = 32'b00000000000000001110111111111011;
assign LUT_3[54415] = 32'b00000000000000010101101011011000;
assign LUT_3[54416] = 32'b00000000000000001101100100011110;
assign LUT_3[54417] = 32'b00000000000000010100001111111011;
assign LUT_3[54418] = 32'b00000000000000001111101100000010;
assign LUT_3[54419] = 32'b00000000000000010110010111011111;
assign LUT_3[54420] = 32'b00000000000000001010110010010100;
assign LUT_3[54421] = 32'b00000000000000010001011101110001;
assign LUT_3[54422] = 32'b00000000000000001100111001111000;
assign LUT_3[54423] = 32'b00000000000000010011100101010101;
assign LUT_3[54424] = 32'b00000000000000010010111101100100;
assign LUT_3[54425] = 32'b00000000000000011001101001000001;
assign LUT_3[54426] = 32'b00000000000000010101000101001000;
assign LUT_3[54427] = 32'b00000000000000011011110000100101;
assign LUT_3[54428] = 32'b00000000000000010000001011011010;
assign LUT_3[54429] = 32'b00000000000000010110110110110111;
assign LUT_3[54430] = 32'b00000000000000010010010010111110;
assign LUT_3[54431] = 32'b00000000000000011000111110011011;
assign LUT_3[54432] = 32'b00000000000000001011011111111011;
assign LUT_3[54433] = 32'b00000000000000010010001011011000;
assign LUT_3[54434] = 32'b00000000000000001101100111011111;
assign LUT_3[54435] = 32'b00000000000000010100010010111100;
assign LUT_3[54436] = 32'b00000000000000001000101101110001;
assign LUT_3[54437] = 32'b00000000000000001111011001001110;
assign LUT_3[54438] = 32'b00000000000000001010110101010101;
assign LUT_3[54439] = 32'b00000000000000010001100000110010;
assign LUT_3[54440] = 32'b00000000000000010000111001000001;
assign LUT_3[54441] = 32'b00000000000000010111100100011110;
assign LUT_3[54442] = 32'b00000000000000010011000000100101;
assign LUT_3[54443] = 32'b00000000000000011001101100000010;
assign LUT_3[54444] = 32'b00000000000000001110000110110111;
assign LUT_3[54445] = 32'b00000000000000010100110010010100;
assign LUT_3[54446] = 32'b00000000000000010000001110011011;
assign LUT_3[54447] = 32'b00000000000000010110111001111000;
assign LUT_3[54448] = 32'b00000000000000001110110010111110;
assign LUT_3[54449] = 32'b00000000000000010101011110011011;
assign LUT_3[54450] = 32'b00000000000000010000111010100010;
assign LUT_3[54451] = 32'b00000000000000010111100101111111;
assign LUT_3[54452] = 32'b00000000000000001100000000110100;
assign LUT_3[54453] = 32'b00000000000000010010101100010001;
assign LUT_3[54454] = 32'b00000000000000001110001000011000;
assign LUT_3[54455] = 32'b00000000000000010100110011110101;
assign LUT_3[54456] = 32'b00000000000000010100001100000100;
assign LUT_3[54457] = 32'b00000000000000011010110111100001;
assign LUT_3[54458] = 32'b00000000000000010110010011101000;
assign LUT_3[54459] = 32'b00000000000000011100111111000101;
assign LUT_3[54460] = 32'b00000000000000010001011001111010;
assign LUT_3[54461] = 32'b00000000000000011000000101010111;
assign LUT_3[54462] = 32'b00000000000000010011100001011110;
assign LUT_3[54463] = 32'b00000000000000011010001100111011;
assign LUT_3[54464] = 32'b00000000000000001010001010000110;
assign LUT_3[54465] = 32'b00000000000000010000110101100011;
assign LUT_3[54466] = 32'b00000000000000001100010001101010;
assign LUT_3[54467] = 32'b00000000000000010010111101000111;
assign LUT_3[54468] = 32'b00000000000000000111010111111100;
assign LUT_3[54469] = 32'b00000000000000001110000011011001;
assign LUT_3[54470] = 32'b00000000000000001001011111100000;
assign LUT_3[54471] = 32'b00000000000000010000001010111101;
assign LUT_3[54472] = 32'b00000000000000001111100011001100;
assign LUT_3[54473] = 32'b00000000000000010110001110101001;
assign LUT_3[54474] = 32'b00000000000000010001101010110000;
assign LUT_3[54475] = 32'b00000000000000011000010110001101;
assign LUT_3[54476] = 32'b00000000000000001100110001000010;
assign LUT_3[54477] = 32'b00000000000000010011011100011111;
assign LUT_3[54478] = 32'b00000000000000001110111000100110;
assign LUT_3[54479] = 32'b00000000000000010101100100000011;
assign LUT_3[54480] = 32'b00000000000000001101011101001001;
assign LUT_3[54481] = 32'b00000000000000010100001000100110;
assign LUT_3[54482] = 32'b00000000000000001111100100101101;
assign LUT_3[54483] = 32'b00000000000000010110010000001010;
assign LUT_3[54484] = 32'b00000000000000001010101010111111;
assign LUT_3[54485] = 32'b00000000000000010001010110011100;
assign LUT_3[54486] = 32'b00000000000000001100110010100011;
assign LUT_3[54487] = 32'b00000000000000010011011110000000;
assign LUT_3[54488] = 32'b00000000000000010010110110001111;
assign LUT_3[54489] = 32'b00000000000000011001100001101100;
assign LUT_3[54490] = 32'b00000000000000010100111101110011;
assign LUT_3[54491] = 32'b00000000000000011011101001010000;
assign LUT_3[54492] = 32'b00000000000000010000000100000101;
assign LUT_3[54493] = 32'b00000000000000010110101111100010;
assign LUT_3[54494] = 32'b00000000000000010010001011101001;
assign LUT_3[54495] = 32'b00000000000000011000110111000110;
assign LUT_3[54496] = 32'b00000000000000001011011000100110;
assign LUT_3[54497] = 32'b00000000000000010010000100000011;
assign LUT_3[54498] = 32'b00000000000000001101100000001010;
assign LUT_3[54499] = 32'b00000000000000010100001011100111;
assign LUT_3[54500] = 32'b00000000000000001000100110011100;
assign LUT_3[54501] = 32'b00000000000000001111010001111001;
assign LUT_3[54502] = 32'b00000000000000001010101110000000;
assign LUT_3[54503] = 32'b00000000000000010001011001011101;
assign LUT_3[54504] = 32'b00000000000000010000110001101100;
assign LUT_3[54505] = 32'b00000000000000010111011101001001;
assign LUT_3[54506] = 32'b00000000000000010010111001010000;
assign LUT_3[54507] = 32'b00000000000000011001100100101101;
assign LUT_3[54508] = 32'b00000000000000001101111111100010;
assign LUT_3[54509] = 32'b00000000000000010100101010111111;
assign LUT_3[54510] = 32'b00000000000000010000000111000110;
assign LUT_3[54511] = 32'b00000000000000010110110010100011;
assign LUT_3[54512] = 32'b00000000000000001110101011101001;
assign LUT_3[54513] = 32'b00000000000000010101010111000110;
assign LUT_3[54514] = 32'b00000000000000010000110011001101;
assign LUT_3[54515] = 32'b00000000000000010111011110101010;
assign LUT_3[54516] = 32'b00000000000000001011111001011111;
assign LUT_3[54517] = 32'b00000000000000010010100100111100;
assign LUT_3[54518] = 32'b00000000000000001110000001000011;
assign LUT_3[54519] = 32'b00000000000000010100101100100000;
assign LUT_3[54520] = 32'b00000000000000010100000100101111;
assign LUT_3[54521] = 32'b00000000000000011010110000001100;
assign LUT_3[54522] = 32'b00000000000000010110001100010011;
assign LUT_3[54523] = 32'b00000000000000011100110111110000;
assign LUT_3[54524] = 32'b00000000000000010001010010100101;
assign LUT_3[54525] = 32'b00000000000000010111111110000010;
assign LUT_3[54526] = 32'b00000000000000010011011010001001;
assign LUT_3[54527] = 32'b00000000000000011010000101100110;
assign LUT_3[54528] = 32'b00000000000000000100010101111110;
assign LUT_3[54529] = 32'b00000000000000001011000001011011;
assign LUT_3[54530] = 32'b00000000000000000110011101100010;
assign LUT_3[54531] = 32'b00000000000000001101001000111111;
assign LUT_3[54532] = 32'b00000000000000000001100011110100;
assign LUT_3[54533] = 32'b00000000000000001000001111010001;
assign LUT_3[54534] = 32'b00000000000000000011101011011000;
assign LUT_3[54535] = 32'b00000000000000001010010110110101;
assign LUT_3[54536] = 32'b00000000000000001001101111000100;
assign LUT_3[54537] = 32'b00000000000000010000011010100001;
assign LUT_3[54538] = 32'b00000000000000001011110110101000;
assign LUT_3[54539] = 32'b00000000000000010010100010000101;
assign LUT_3[54540] = 32'b00000000000000000110111100111010;
assign LUT_3[54541] = 32'b00000000000000001101101000010111;
assign LUT_3[54542] = 32'b00000000000000001001000100011110;
assign LUT_3[54543] = 32'b00000000000000001111101111111011;
assign LUT_3[54544] = 32'b00000000000000000111101001000001;
assign LUT_3[54545] = 32'b00000000000000001110010100011110;
assign LUT_3[54546] = 32'b00000000000000001001110000100101;
assign LUT_3[54547] = 32'b00000000000000010000011100000010;
assign LUT_3[54548] = 32'b00000000000000000100110110110111;
assign LUT_3[54549] = 32'b00000000000000001011100010010100;
assign LUT_3[54550] = 32'b00000000000000000110111110011011;
assign LUT_3[54551] = 32'b00000000000000001101101001111000;
assign LUT_3[54552] = 32'b00000000000000001101000010000111;
assign LUT_3[54553] = 32'b00000000000000010011101101100100;
assign LUT_3[54554] = 32'b00000000000000001111001001101011;
assign LUT_3[54555] = 32'b00000000000000010101110101001000;
assign LUT_3[54556] = 32'b00000000000000001010001111111101;
assign LUT_3[54557] = 32'b00000000000000010000111011011010;
assign LUT_3[54558] = 32'b00000000000000001100010111100001;
assign LUT_3[54559] = 32'b00000000000000010011000010111110;
assign LUT_3[54560] = 32'b00000000000000000101100100011110;
assign LUT_3[54561] = 32'b00000000000000001100001111111011;
assign LUT_3[54562] = 32'b00000000000000000111101100000010;
assign LUT_3[54563] = 32'b00000000000000001110010111011111;
assign LUT_3[54564] = 32'b00000000000000000010110010010100;
assign LUT_3[54565] = 32'b00000000000000001001011101110001;
assign LUT_3[54566] = 32'b00000000000000000100111001111000;
assign LUT_3[54567] = 32'b00000000000000001011100101010101;
assign LUT_3[54568] = 32'b00000000000000001010111101100100;
assign LUT_3[54569] = 32'b00000000000000010001101001000001;
assign LUT_3[54570] = 32'b00000000000000001101000101001000;
assign LUT_3[54571] = 32'b00000000000000010011110000100101;
assign LUT_3[54572] = 32'b00000000000000001000001011011010;
assign LUT_3[54573] = 32'b00000000000000001110110110110111;
assign LUT_3[54574] = 32'b00000000000000001010010010111110;
assign LUT_3[54575] = 32'b00000000000000010000111110011011;
assign LUT_3[54576] = 32'b00000000000000001000110111100001;
assign LUT_3[54577] = 32'b00000000000000001111100010111110;
assign LUT_3[54578] = 32'b00000000000000001010111111000101;
assign LUT_3[54579] = 32'b00000000000000010001101010100010;
assign LUT_3[54580] = 32'b00000000000000000110000101010111;
assign LUT_3[54581] = 32'b00000000000000001100110000110100;
assign LUT_3[54582] = 32'b00000000000000001000001100111011;
assign LUT_3[54583] = 32'b00000000000000001110111000011000;
assign LUT_3[54584] = 32'b00000000000000001110010000100111;
assign LUT_3[54585] = 32'b00000000000000010100111100000100;
assign LUT_3[54586] = 32'b00000000000000010000011000001011;
assign LUT_3[54587] = 32'b00000000000000010111000011101000;
assign LUT_3[54588] = 32'b00000000000000001011011110011101;
assign LUT_3[54589] = 32'b00000000000000010010001001111010;
assign LUT_3[54590] = 32'b00000000000000001101100110000001;
assign LUT_3[54591] = 32'b00000000000000010100010001011110;
assign LUT_3[54592] = 32'b00000000000000000100001110101001;
assign LUT_3[54593] = 32'b00000000000000001010111010000110;
assign LUT_3[54594] = 32'b00000000000000000110010110001101;
assign LUT_3[54595] = 32'b00000000000000001101000001101010;
assign LUT_3[54596] = 32'b00000000000000000001011100011111;
assign LUT_3[54597] = 32'b00000000000000001000000111111100;
assign LUT_3[54598] = 32'b00000000000000000011100100000011;
assign LUT_3[54599] = 32'b00000000000000001010001111100000;
assign LUT_3[54600] = 32'b00000000000000001001100111101111;
assign LUT_3[54601] = 32'b00000000000000010000010011001100;
assign LUT_3[54602] = 32'b00000000000000001011101111010011;
assign LUT_3[54603] = 32'b00000000000000010010011010110000;
assign LUT_3[54604] = 32'b00000000000000000110110101100101;
assign LUT_3[54605] = 32'b00000000000000001101100001000010;
assign LUT_3[54606] = 32'b00000000000000001000111101001001;
assign LUT_3[54607] = 32'b00000000000000001111101000100110;
assign LUT_3[54608] = 32'b00000000000000000111100001101100;
assign LUT_3[54609] = 32'b00000000000000001110001101001001;
assign LUT_3[54610] = 32'b00000000000000001001101001010000;
assign LUT_3[54611] = 32'b00000000000000010000010100101101;
assign LUT_3[54612] = 32'b00000000000000000100101111100010;
assign LUT_3[54613] = 32'b00000000000000001011011010111111;
assign LUT_3[54614] = 32'b00000000000000000110110111000110;
assign LUT_3[54615] = 32'b00000000000000001101100010100011;
assign LUT_3[54616] = 32'b00000000000000001100111010110010;
assign LUT_3[54617] = 32'b00000000000000010011100110001111;
assign LUT_3[54618] = 32'b00000000000000001111000010010110;
assign LUT_3[54619] = 32'b00000000000000010101101101110011;
assign LUT_3[54620] = 32'b00000000000000001010001000101000;
assign LUT_3[54621] = 32'b00000000000000010000110100000101;
assign LUT_3[54622] = 32'b00000000000000001100010000001100;
assign LUT_3[54623] = 32'b00000000000000010010111011101001;
assign LUT_3[54624] = 32'b00000000000000000101011101001001;
assign LUT_3[54625] = 32'b00000000000000001100001000100110;
assign LUT_3[54626] = 32'b00000000000000000111100100101101;
assign LUT_3[54627] = 32'b00000000000000001110010000001010;
assign LUT_3[54628] = 32'b00000000000000000010101010111111;
assign LUT_3[54629] = 32'b00000000000000001001010110011100;
assign LUT_3[54630] = 32'b00000000000000000100110010100011;
assign LUT_3[54631] = 32'b00000000000000001011011110000000;
assign LUT_3[54632] = 32'b00000000000000001010110110001111;
assign LUT_3[54633] = 32'b00000000000000010001100001101100;
assign LUT_3[54634] = 32'b00000000000000001100111101110011;
assign LUT_3[54635] = 32'b00000000000000010011101001010000;
assign LUT_3[54636] = 32'b00000000000000001000000100000101;
assign LUT_3[54637] = 32'b00000000000000001110101111100010;
assign LUT_3[54638] = 32'b00000000000000001010001011101001;
assign LUT_3[54639] = 32'b00000000000000010000110111000110;
assign LUT_3[54640] = 32'b00000000000000001000110000001100;
assign LUT_3[54641] = 32'b00000000000000001111011011101001;
assign LUT_3[54642] = 32'b00000000000000001010110111110000;
assign LUT_3[54643] = 32'b00000000000000010001100011001101;
assign LUT_3[54644] = 32'b00000000000000000101111110000010;
assign LUT_3[54645] = 32'b00000000000000001100101001011111;
assign LUT_3[54646] = 32'b00000000000000001000000101100110;
assign LUT_3[54647] = 32'b00000000000000001110110001000011;
assign LUT_3[54648] = 32'b00000000000000001110001001010010;
assign LUT_3[54649] = 32'b00000000000000010100110100101111;
assign LUT_3[54650] = 32'b00000000000000010000010000110110;
assign LUT_3[54651] = 32'b00000000000000010110111100010011;
assign LUT_3[54652] = 32'b00000000000000001011010111001000;
assign LUT_3[54653] = 32'b00000000000000010010000010100101;
assign LUT_3[54654] = 32'b00000000000000001101011110101100;
assign LUT_3[54655] = 32'b00000000000000010100001010001001;
assign LUT_3[54656] = 32'b00000000000000000110100000111100;
assign LUT_3[54657] = 32'b00000000000000001101001100011001;
assign LUT_3[54658] = 32'b00000000000000001000101000100000;
assign LUT_3[54659] = 32'b00000000000000001111010011111101;
assign LUT_3[54660] = 32'b00000000000000000011101110110010;
assign LUT_3[54661] = 32'b00000000000000001010011010001111;
assign LUT_3[54662] = 32'b00000000000000000101110110010110;
assign LUT_3[54663] = 32'b00000000000000001100100001110011;
assign LUT_3[54664] = 32'b00000000000000001011111010000010;
assign LUT_3[54665] = 32'b00000000000000010010100101011111;
assign LUT_3[54666] = 32'b00000000000000001110000001100110;
assign LUT_3[54667] = 32'b00000000000000010100101101000011;
assign LUT_3[54668] = 32'b00000000000000001001000111111000;
assign LUT_3[54669] = 32'b00000000000000001111110011010101;
assign LUT_3[54670] = 32'b00000000000000001011001111011100;
assign LUT_3[54671] = 32'b00000000000000010001111010111001;
assign LUT_3[54672] = 32'b00000000000000001001110011111111;
assign LUT_3[54673] = 32'b00000000000000010000011111011100;
assign LUT_3[54674] = 32'b00000000000000001011111011100011;
assign LUT_3[54675] = 32'b00000000000000010010100111000000;
assign LUT_3[54676] = 32'b00000000000000000111000001110101;
assign LUT_3[54677] = 32'b00000000000000001101101101010010;
assign LUT_3[54678] = 32'b00000000000000001001001001011001;
assign LUT_3[54679] = 32'b00000000000000001111110100110110;
assign LUT_3[54680] = 32'b00000000000000001111001101000101;
assign LUT_3[54681] = 32'b00000000000000010101111000100010;
assign LUT_3[54682] = 32'b00000000000000010001010100101001;
assign LUT_3[54683] = 32'b00000000000000011000000000000110;
assign LUT_3[54684] = 32'b00000000000000001100011010111011;
assign LUT_3[54685] = 32'b00000000000000010011000110011000;
assign LUT_3[54686] = 32'b00000000000000001110100010011111;
assign LUT_3[54687] = 32'b00000000000000010101001101111100;
assign LUT_3[54688] = 32'b00000000000000000111101111011100;
assign LUT_3[54689] = 32'b00000000000000001110011010111001;
assign LUT_3[54690] = 32'b00000000000000001001110111000000;
assign LUT_3[54691] = 32'b00000000000000010000100010011101;
assign LUT_3[54692] = 32'b00000000000000000100111101010010;
assign LUT_3[54693] = 32'b00000000000000001011101000101111;
assign LUT_3[54694] = 32'b00000000000000000111000100110110;
assign LUT_3[54695] = 32'b00000000000000001101110000010011;
assign LUT_3[54696] = 32'b00000000000000001101001000100010;
assign LUT_3[54697] = 32'b00000000000000010011110011111111;
assign LUT_3[54698] = 32'b00000000000000001111010000000110;
assign LUT_3[54699] = 32'b00000000000000010101111011100011;
assign LUT_3[54700] = 32'b00000000000000001010010110011000;
assign LUT_3[54701] = 32'b00000000000000010001000001110101;
assign LUT_3[54702] = 32'b00000000000000001100011101111100;
assign LUT_3[54703] = 32'b00000000000000010011001001011001;
assign LUT_3[54704] = 32'b00000000000000001011000010011111;
assign LUT_3[54705] = 32'b00000000000000010001101101111100;
assign LUT_3[54706] = 32'b00000000000000001101001010000011;
assign LUT_3[54707] = 32'b00000000000000010011110101100000;
assign LUT_3[54708] = 32'b00000000000000001000010000010101;
assign LUT_3[54709] = 32'b00000000000000001110111011110010;
assign LUT_3[54710] = 32'b00000000000000001010010111111001;
assign LUT_3[54711] = 32'b00000000000000010001000011010110;
assign LUT_3[54712] = 32'b00000000000000010000011011100101;
assign LUT_3[54713] = 32'b00000000000000010111000111000010;
assign LUT_3[54714] = 32'b00000000000000010010100011001001;
assign LUT_3[54715] = 32'b00000000000000011001001110100110;
assign LUT_3[54716] = 32'b00000000000000001101101001011011;
assign LUT_3[54717] = 32'b00000000000000010100010100111000;
assign LUT_3[54718] = 32'b00000000000000001111110000111111;
assign LUT_3[54719] = 32'b00000000000000010110011100011100;
assign LUT_3[54720] = 32'b00000000000000000110011001100111;
assign LUT_3[54721] = 32'b00000000000000001101000101000100;
assign LUT_3[54722] = 32'b00000000000000001000100001001011;
assign LUT_3[54723] = 32'b00000000000000001111001100101000;
assign LUT_3[54724] = 32'b00000000000000000011100111011101;
assign LUT_3[54725] = 32'b00000000000000001010010010111010;
assign LUT_3[54726] = 32'b00000000000000000101101111000001;
assign LUT_3[54727] = 32'b00000000000000001100011010011110;
assign LUT_3[54728] = 32'b00000000000000001011110010101101;
assign LUT_3[54729] = 32'b00000000000000010010011110001010;
assign LUT_3[54730] = 32'b00000000000000001101111010010001;
assign LUT_3[54731] = 32'b00000000000000010100100101101110;
assign LUT_3[54732] = 32'b00000000000000001001000000100011;
assign LUT_3[54733] = 32'b00000000000000001111101100000000;
assign LUT_3[54734] = 32'b00000000000000001011001000000111;
assign LUT_3[54735] = 32'b00000000000000010001110011100100;
assign LUT_3[54736] = 32'b00000000000000001001101100101010;
assign LUT_3[54737] = 32'b00000000000000010000011000000111;
assign LUT_3[54738] = 32'b00000000000000001011110100001110;
assign LUT_3[54739] = 32'b00000000000000010010011111101011;
assign LUT_3[54740] = 32'b00000000000000000110111010100000;
assign LUT_3[54741] = 32'b00000000000000001101100101111101;
assign LUT_3[54742] = 32'b00000000000000001001000010000100;
assign LUT_3[54743] = 32'b00000000000000001111101101100001;
assign LUT_3[54744] = 32'b00000000000000001111000101110000;
assign LUT_3[54745] = 32'b00000000000000010101110001001101;
assign LUT_3[54746] = 32'b00000000000000010001001101010100;
assign LUT_3[54747] = 32'b00000000000000010111111000110001;
assign LUT_3[54748] = 32'b00000000000000001100010011100110;
assign LUT_3[54749] = 32'b00000000000000010010111111000011;
assign LUT_3[54750] = 32'b00000000000000001110011011001010;
assign LUT_3[54751] = 32'b00000000000000010101000110100111;
assign LUT_3[54752] = 32'b00000000000000000111101000000111;
assign LUT_3[54753] = 32'b00000000000000001110010011100100;
assign LUT_3[54754] = 32'b00000000000000001001101111101011;
assign LUT_3[54755] = 32'b00000000000000010000011011001000;
assign LUT_3[54756] = 32'b00000000000000000100110101111101;
assign LUT_3[54757] = 32'b00000000000000001011100001011010;
assign LUT_3[54758] = 32'b00000000000000000110111101100001;
assign LUT_3[54759] = 32'b00000000000000001101101000111110;
assign LUT_3[54760] = 32'b00000000000000001101000001001101;
assign LUT_3[54761] = 32'b00000000000000010011101100101010;
assign LUT_3[54762] = 32'b00000000000000001111001000110001;
assign LUT_3[54763] = 32'b00000000000000010101110100001110;
assign LUT_3[54764] = 32'b00000000000000001010001111000011;
assign LUT_3[54765] = 32'b00000000000000010000111010100000;
assign LUT_3[54766] = 32'b00000000000000001100010110100111;
assign LUT_3[54767] = 32'b00000000000000010011000010000100;
assign LUT_3[54768] = 32'b00000000000000001010111011001010;
assign LUT_3[54769] = 32'b00000000000000010001100110100111;
assign LUT_3[54770] = 32'b00000000000000001101000010101110;
assign LUT_3[54771] = 32'b00000000000000010011101110001011;
assign LUT_3[54772] = 32'b00000000000000001000001001000000;
assign LUT_3[54773] = 32'b00000000000000001110110100011101;
assign LUT_3[54774] = 32'b00000000000000001010010000100100;
assign LUT_3[54775] = 32'b00000000000000010000111100000001;
assign LUT_3[54776] = 32'b00000000000000010000010100010000;
assign LUT_3[54777] = 32'b00000000000000010110111111101101;
assign LUT_3[54778] = 32'b00000000000000010010011011110100;
assign LUT_3[54779] = 32'b00000000000000011001000111010001;
assign LUT_3[54780] = 32'b00000000000000001101100010000110;
assign LUT_3[54781] = 32'b00000000000000010100001101100011;
assign LUT_3[54782] = 32'b00000000000000001111101001101010;
assign LUT_3[54783] = 32'b00000000000000010110010101000111;
assign LUT_3[54784] = 32'b00000000000000001011011011101001;
assign LUT_3[54785] = 32'b00000000000000010010000111000110;
assign LUT_3[54786] = 32'b00000000000000001101100011001101;
assign LUT_3[54787] = 32'b00000000000000010100001110101010;
assign LUT_3[54788] = 32'b00000000000000001000101001011111;
assign LUT_3[54789] = 32'b00000000000000001111010100111100;
assign LUT_3[54790] = 32'b00000000000000001010110001000011;
assign LUT_3[54791] = 32'b00000000000000010001011100100000;
assign LUT_3[54792] = 32'b00000000000000010000110100101111;
assign LUT_3[54793] = 32'b00000000000000010111100000001100;
assign LUT_3[54794] = 32'b00000000000000010010111100010011;
assign LUT_3[54795] = 32'b00000000000000011001100111110000;
assign LUT_3[54796] = 32'b00000000000000001110000010100101;
assign LUT_3[54797] = 32'b00000000000000010100101110000010;
assign LUT_3[54798] = 32'b00000000000000010000001010001001;
assign LUT_3[54799] = 32'b00000000000000010110110101100110;
assign LUT_3[54800] = 32'b00000000000000001110101110101100;
assign LUT_3[54801] = 32'b00000000000000010101011010001001;
assign LUT_3[54802] = 32'b00000000000000010000110110010000;
assign LUT_3[54803] = 32'b00000000000000010111100001101101;
assign LUT_3[54804] = 32'b00000000000000001011111100100010;
assign LUT_3[54805] = 32'b00000000000000010010100111111111;
assign LUT_3[54806] = 32'b00000000000000001110000100000110;
assign LUT_3[54807] = 32'b00000000000000010100101111100011;
assign LUT_3[54808] = 32'b00000000000000010100000111110010;
assign LUT_3[54809] = 32'b00000000000000011010110011001111;
assign LUT_3[54810] = 32'b00000000000000010110001111010110;
assign LUT_3[54811] = 32'b00000000000000011100111010110011;
assign LUT_3[54812] = 32'b00000000000000010001010101101000;
assign LUT_3[54813] = 32'b00000000000000011000000001000101;
assign LUT_3[54814] = 32'b00000000000000010011011101001100;
assign LUT_3[54815] = 32'b00000000000000011010001000101001;
assign LUT_3[54816] = 32'b00000000000000001100101010001001;
assign LUT_3[54817] = 32'b00000000000000010011010101100110;
assign LUT_3[54818] = 32'b00000000000000001110110001101101;
assign LUT_3[54819] = 32'b00000000000000010101011101001010;
assign LUT_3[54820] = 32'b00000000000000001001110111111111;
assign LUT_3[54821] = 32'b00000000000000010000100011011100;
assign LUT_3[54822] = 32'b00000000000000001011111111100011;
assign LUT_3[54823] = 32'b00000000000000010010101011000000;
assign LUT_3[54824] = 32'b00000000000000010010000011001111;
assign LUT_3[54825] = 32'b00000000000000011000101110101100;
assign LUT_3[54826] = 32'b00000000000000010100001010110011;
assign LUT_3[54827] = 32'b00000000000000011010110110010000;
assign LUT_3[54828] = 32'b00000000000000001111010001000101;
assign LUT_3[54829] = 32'b00000000000000010101111100100010;
assign LUT_3[54830] = 32'b00000000000000010001011000101001;
assign LUT_3[54831] = 32'b00000000000000011000000100000110;
assign LUT_3[54832] = 32'b00000000000000001111111101001100;
assign LUT_3[54833] = 32'b00000000000000010110101000101001;
assign LUT_3[54834] = 32'b00000000000000010010000100110000;
assign LUT_3[54835] = 32'b00000000000000011000110000001101;
assign LUT_3[54836] = 32'b00000000000000001101001011000010;
assign LUT_3[54837] = 32'b00000000000000010011110110011111;
assign LUT_3[54838] = 32'b00000000000000001111010010100110;
assign LUT_3[54839] = 32'b00000000000000010101111110000011;
assign LUT_3[54840] = 32'b00000000000000010101010110010010;
assign LUT_3[54841] = 32'b00000000000000011100000001101111;
assign LUT_3[54842] = 32'b00000000000000010111011101110110;
assign LUT_3[54843] = 32'b00000000000000011110001001010011;
assign LUT_3[54844] = 32'b00000000000000010010100100001000;
assign LUT_3[54845] = 32'b00000000000000011001001111100101;
assign LUT_3[54846] = 32'b00000000000000010100101011101100;
assign LUT_3[54847] = 32'b00000000000000011011010111001001;
assign LUT_3[54848] = 32'b00000000000000001011010100010100;
assign LUT_3[54849] = 32'b00000000000000010001111111110001;
assign LUT_3[54850] = 32'b00000000000000001101011011111000;
assign LUT_3[54851] = 32'b00000000000000010100000111010101;
assign LUT_3[54852] = 32'b00000000000000001000100010001010;
assign LUT_3[54853] = 32'b00000000000000001111001101100111;
assign LUT_3[54854] = 32'b00000000000000001010101001101110;
assign LUT_3[54855] = 32'b00000000000000010001010101001011;
assign LUT_3[54856] = 32'b00000000000000010000101101011010;
assign LUT_3[54857] = 32'b00000000000000010111011000110111;
assign LUT_3[54858] = 32'b00000000000000010010110100111110;
assign LUT_3[54859] = 32'b00000000000000011001100000011011;
assign LUT_3[54860] = 32'b00000000000000001101111011010000;
assign LUT_3[54861] = 32'b00000000000000010100100110101101;
assign LUT_3[54862] = 32'b00000000000000010000000010110100;
assign LUT_3[54863] = 32'b00000000000000010110101110010001;
assign LUT_3[54864] = 32'b00000000000000001110100111010111;
assign LUT_3[54865] = 32'b00000000000000010101010010110100;
assign LUT_3[54866] = 32'b00000000000000010000101110111011;
assign LUT_3[54867] = 32'b00000000000000010111011010011000;
assign LUT_3[54868] = 32'b00000000000000001011110101001101;
assign LUT_3[54869] = 32'b00000000000000010010100000101010;
assign LUT_3[54870] = 32'b00000000000000001101111100110001;
assign LUT_3[54871] = 32'b00000000000000010100101000001110;
assign LUT_3[54872] = 32'b00000000000000010100000000011101;
assign LUT_3[54873] = 32'b00000000000000011010101011111010;
assign LUT_3[54874] = 32'b00000000000000010110001000000001;
assign LUT_3[54875] = 32'b00000000000000011100110011011110;
assign LUT_3[54876] = 32'b00000000000000010001001110010011;
assign LUT_3[54877] = 32'b00000000000000010111111001110000;
assign LUT_3[54878] = 32'b00000000000000010011010101110111;
assign LUT_3[54879] = 32'b00000000000000011010000001010100;
assign LUT_3[54880] = 32'b00000000000000001100100010110100;
assign LUT_3[54881] = 32'b00000000000000010011001110010001;
assign LUT_3[54882] = 32'b00000000000000001110101010011000;
assign LUT_3[54883] = 32'b00000000000000010101010101110101;
assign LUT_3[54884] = 32'b00000000000000001001110000101010;
assign LUT_3[54885] = 32'b00000000000000010000011100000111;
assign LUT_3[54886] = 32'b00000000000000001011111000001110;
assign LUT_3[54887] = 32'b00000000000000010010100011101011;
assign LUT_3[54888] = 32'b00000000000000010001111011111010;
assign LUT_3[54889] = 32'b00000000000000011000100111010111;
assign LUT_3[54890] = 32'b00000000000000010100000011011110;
assign LUT_3[54891] = 32'b00000000000000011010101110111011;
assign LUT_3[54892] = 32'b00000000000000001111001001110000;
assign LUT_3[54893] = 32'b00000000000000010101110101001101;
assign LUT_3[54894] = 32'b00000000000000010001010001010100;
assign LUT_3[54895] = 32'b00000000000000010111111100110001;
assign LUT_3[54896] = 32'b00000000000000001111110101110111;
assign LUT_3[54897] = 32'b00000000000000010110100001010100;
assign LUT_3[54898] = 32'b00000000000000010001111101011011;
assign LUT_3[54899] = 32'b00000000000000011000101000111000;
assign LUT_3[54900] = 32'b00000000000000001101000011101101;
assign LUT_3[54901] = 32'b00000000000000010011101111001010;
assign LUT_3[54902] = 32'b00000000000000001111001011010001;
assign LUT_3[54903] = 32'b00000000000000010101110110101110;
assign LUT_3[54904] = 32'b00000000000000010101001110111101;
assign LUT_3[54905] = 32'b00000000000000011011111010011010;
assign LUT_3[54906] = 32'b00000000000000010111010110100001;
assign LUT_3[54907] = 32'b00000000000000011110000001111110;
assign LUT_3[54908] = 32'b00000000000000010010011100110011;
assign LUT_3[54909] = 32'b00000000000000011001001000010000;
assign LUT_3[54910] = 32'b00000000000000010100100100010111;
assign LUT_3[54911] = 32'b00000000000000011011001111110100;
assign LUT_3[54912] = 32'b00000000000000001101100110100111;
assign LUT_3[54913] = 32'b00000000000000010100010010000100;
assign LUT_3[54914] = 32'b00000000000000001111101110001011;
assign LUT_3[54915] = 32'b00000000000000010110011001101000;
assign LUT_3[54916] = 32'b00000000000000001010110100011101;
assign LUT_3[54917] = 32'b00000000000000010001011111111010;
assign LUT_3[54918] = 32'b00000000000000001100111100000001;
assign LUT_3[54919] = 32'b00000000000000010011100111011110;
assign LUT_3[54920] = 32'b00000000000000010010111111101101;
assign LUT_3[54921] = 32'b00000000000000011001101011001010;
assign LUT_3[54922] = 32'b00000000000000010101000111010001;
assign LUT_3[54923] = 32'b00000000000000011011110010101110;
assign LUT_3[54924] = 32'b00000000000000010000001101100011;
assign LUT_3[54925] = 32'b00000000000000010110111001000000;
assign LUT_3[54926] = 32'b00000000000000010010010101000111;
assign LUT_3[54927] = 32'b00000000000000011001000000100100;
assign LUT_3[54928] = 32'b00000000000000010000111001101010;
assign LUT_3[54929] = 32'b00000000000000010111100101000111;
assign LUT_3[54930] = 32'b00000000000000010011000001001110;
assign LUT_3[54931] = 32'b00000000000000011001101100101011;
assign LUT_3[54932] = 32'b00000000000000001110000111100000;
assign LUT_3[54933] = 32'b00000000000000010100110010111101;
assign LUT_3[54934] = 32'b00000000000000010000001111000100;
assign LUT_3[54935] = 32'b00000000000000010110111010100001;
assign LUT_3[54936] = 32'b00000000000000010110010010110000;
assign LUT_3[54937] = 32'b00000000000000011100111110001101;
assign LUT_3[54938] = 32'b00000000000000011000011010010100;
assign LUT_3[54939] = 32'b00000000000000011111000101110001;
assign LUT_3[54940] = 32'b00000000000000010011100000100110;
assign LUT_3[54941] = 32'b00000000000000011010001100000011;
assign LUT_3[54942] = 32'b00000000000000010101101000001010;
assign LUT_3[54943] = 32'b00000000000000011100010011100111;
assign LUT_3[54944] = 32'b00000000000000001110110101000111;
assign LUT_3[54945] = 32'b00000000000000010101100000100100;
assign LUT_3[54946] = 32'b00000000000000010000111100101011;
assign LUT_3[54947] = 32'b00000000000000010111101000001000;
assign LUT_3[54948] = 32'b00000000000000001100000010111101;
assign LUT_3[54949] = 32'b00000000000000010010101110011010;
assign LUT_3[54950] = 32'b00000000000000001110001010100001;
assign LUT_3[54951] = 32'b00000000000000010100110101111110;
assign LUT_3[54952] = 32'b00000000000000010100001110001101;
assign LUT_3[54953] = 32'b00000000000000011010111001101010;
assign LUT_3[54954] = 32'b00000000000000010110010101110001;
assign LUT_3[54955] = 32'b00000000000000011101000001001110;
assign LUT_3[54956] = 32'b00000000000000010001011100000011;
assign LUT_3[54957] = 32'b00000000000000011000000111100000;
assign LUT_3[54958] = 32'b00000000000000010011100011100111;
assign LUT_3[54959] = 32'b00000000000000011010001111000100;
assign LUT_3[54960] = 32'b00000000000000010010001000001010;
assign LUT_3[54961] = 32'b00000000000000011000110011100111;
assign LUT_3[54962] = 32'b00000000000000010100001111101110;
assign LUT_3[54963] = 32'b00000000000000011010111011001011;
assign LUT_3[54964] = 32'b00000000000000001111010110000000;
assign LUT_3[54965] = 32'b00000000000000010110000001011101;
assign LUT_3[54966] = 32'b00000000000000010001011101100100;
assign LUT_3[54967] = 32'b00000000000000011000001001000001;
assign LUT_3[54968] = 32'b00000000000000010111100001010000;
assign LUT_3[54969] = 32'b00000000000000011110001100101101;
assign LUT_3[54970] = 32'b00000000000000011001101000110100;
assign LUT_3[54971] = 32'b00000000000000100000010100010001;
assign LUT_3[54972] = 32'b00000000000000010100101111000110;
assign LUT_3[54973] = 32'b00000000000000011011011010100011;
assign LUT_3[54974] = 32'b00000000000000010110110110101010;
assign LUT_3[54975] = 32'b00000000000000011101100010000111;
assign LUT_3[54976] = 32'b00000000000000001101011111010010;
assign LUT_3[54977] = 32'b00000000000000010100001010101111;
assign LUT_3[54978] = 32'b00000000000000001111100110110110;
assign LUT_3[54979] = 32'b00000000000000010110010010010011;
assign LUT_3[54980] = 32'b00000000000000001010101101001000;
assign LUT_3[54981] = 32'b00000000000000010001011000100101;
assign LUT_3[54982] = 32'b00000000000000001100110100101100;
assign LUT_3[54983] = 32'b00000000000000010011100000001001;
assign LUT_3[54984] = 32'b00000000000000010010111000011000;
assign LUT_3[54985] = 32'b00000000000000011001100011110101;
assign LUT_3[54986] = 32'b00000000000000010100111111111100;
assign LUT_3[54987] = 32'b00000000000000011011101011011001;
assign LUT_3[54988] = 32'b00000000000000010000000110001110;
assign LUT_3[54989] = 32'b00000000000000010110110001101011;
assign LUT_3[54990] = 32'b00000000000000010010001101110010;
assign LUT_3[54991] = 32'b00000000000000011000111001001111;
assign LUT_3[54992] = 32'b00000000000000010000110010010101;
assign LUT_3[54993] = 32'b00000000000000010111011101110010;
assign LUT_3[54994] = 32'b00000000000000010010111001111001;
assign LUT_3[54995] = 32'b00000000000000011001100101010110;
assign LUT_3[54996] = 32'b00000000000000001110000000001011;
assign LUT_3[54997] = 32'b00000000000000010100101011101000;
assign LUT_3[54998] = 32'b00000000000000010000000111101111;
assign LUT_3[54999] = 32'b00000000000000010110110011001100;
assign LUT_3[55000] = 32'b00000000000000010110001011011011;
assign LUT_3[55001] = 32'b00000000000000011100110110111000;
assign LUT_3[55002] = 32'b00000000000000011000010010111111;
assign LUT_3[55003] = 32'b00000000000000011110111110011100;
assign LUT_3[55004] = 32'b00000000000000010011011001010001;
assign LUT_3[55005] = 32'b00000000000000011010000100101110;
assign LUT_3[55006] = 32'b00000000000000010101100000110101;
assign LUT_3[55007] = 32'b00000000000000011100001100010010;
assign LUT_3[55008] = 32'b00000000000000001110101101110010;
assign LUT_3[55009] = 32'b00000000000000010101011001001111;
assign LUT_3[55010] = 32'b00000000000000010000110101010110;
assign LUT_3[55011] = 32'b00000000000000010111100000110011;
assign LUT_3[55012] = 32'b00000000000000001011111011101000;
assign LUT_3[55013] = 32'b00000000000000010010100111000101;
assign LUT_3[55014] = 32'b00000000000000001110000011001100;
assign LUT_3[55015] = 32'b00000000000000010100101110101001;
assign LUT_3[55016] = 32'b00000000000000010100000110111000;
assign LUT_3[55017] = 32'b00000000000000011010110010010101;
assign LUT_3[55018] = 32'b00000000000000010110001110011100;
assign LUT_3[55019] = 32'b00000000000000011100111001111001;
assign LUT_3[55020] = 32'b00000000000000010001010100101110;
assign LUT_3[55021] = 32'b00000000000000011000000000001011;
assign LUT_3[55022] = 32'b00000000000000010011011100010010;
assign LUT_3[55023] = 32'b00000000000000011010000111101111;
assign LUT_3[55024] = 32'b00000000000000010010000000110101;
assign LUT_3[55025] = 32'b00000000000000011000101100010010;
assign LUT_3[55026] = 32'b00000000000000010100001000011001;
assign LUT_3[55027] = 32'b00000000000000011010110011110110;
assign LUT_3[55028] = 32'b00000000000000001111001110101011;
assign LUT_3[55029] = 32'b00000000000000010101111010001000;
assign LUT_3[55030] = 32'b00000000000000010001010110001111;
assign LUT_3[55031] = 32'b00000000000000011000000001101100;
assign LUT_3[55032] = 32'b00000000000000010111011001111011;
assign LUT_3[55033] = 32'b00000000000000011110000101011000;
assign LUT_3[55034] = 32'b00000000000000011001100001011111;
assign LUT_3[55035] = 32'b00000000000000100000001100111100;
assign LUT_3[55036] = 32'b00000000000000010100100111110001;
assign LUT_3[55037] = 32'b00000000000000011011010011001110;
assign LUT_3[55038] = 32'b00000000000000010110101111010101;
assign LUT_3[55039] = 32'b00000000000000011101011010110010;
assign LUT_3[55040] = 32'b00000000000000000111101011001010;
assign LUT_3[55041] = 32'b00000000000000001110010110100111;
assign LUT_3[55042] = 32'b00000000000000001001110010101110;
assign LUT_3[55043] = 32'b00000000000000010000011110001011;
assign LUT_3[55044] = 32'b00000000000000000100111001000000;
assign LUT_3[55045] = 32'b00000000000000001011100100011101;
assign LUT_3[55046] = 32'b00000000000000000111000000100100;
assign LUT_3[55047] = 32'b00000000000000001101101100000001;
assign LUT_3[55048] = 32'b00000000000000001101000100010000;
assign LUT_3[55049] = 32'b00000000000000010011101111101101;
assign LUT_3[55050] = 32'b00000000000000001111001011110100;
assign LUT_3[55051] = 32'b00000000000000010101110111010001;
assign LUT_3[55052] = 32'b00000000000000001010010010000110;
assign LUT_3[55053] = 32'b00000000000000010000111101100011;
assign LUT_3[55054] = 32'b00000000000000001100011001101010;
assign LUT_3[55055] = 32'b00000000000000010011000101000111;
assign LUT_3[55056] = 32'b00000000000000001010111110001101;
assign LUT_3[55057] = 32'b00000000000000010001101001101010;
assign LUT_3[55058] = 32'b00000000000000001101000101110001;
assign LUT_3[55059] = 32'b00000000000000010011110001001110;
assign LUT_3[55060] = 32'b00000000000000001000001100000011;
assign LUT_3[55061] = 32'b00000000000000001110110111100000;
assign LUT_3[55062] = 32'b00000000000000001010010011100111;
assign LUT_3[55063] = 32'b00000000000000010000111111000100;
assign LUT_3[55064] = 32'b00000000000000010000010111010011;
assign LUT_3[55065] = 32'b00000000000000010111000010110000;
assign LUT_3[55066] = 32'b00000000000000010010011110110111;
assign LUT_3[55067] = 32'b00000000000000011001001010010100;
assign LUT_3[55068] = 32'b00000000000000001101100101001001;
assign LUT_3[55069] = 32'b00000000000000010100010000100110;
assign LUT_3[55070] = 32'b00000000000000001111101100101101;
assign LUT_3[55071] = 32'b00000000000000010110011000001010;
assign LUT_3[55072] = 32'b00000000000000001000111001101010;
assign LUT_3[55073] = 32'b00000000000000001111100101000111;
assign LUT_3[55074] = 32'b00000000000000001011000001001110;
assign LUT_3[55075] = 32'b00000000000000010001101100101011;
assign LUT_3[55076] = 32'b00000000000000000110000111100000;
assign LUT_3[55077] = 32'b00000000000000001100110010111101;
assign LUT_3[55078] = 32'b00000000000000001000001111000100;
assign LUT_3[55079] = 32'b00000000000000001110111010100001;
assign LUT_3[55080] = 32'b00000000000000001110010010110000;
assign LUT_3[55081] = 32'b00000000000000010100111110001101;
assign LUT_3[55082] = 32'b00000000000000010000011010010100;
assign LUT_3[55083] = 32'b00000000000000010111000101110001;
assign LUT_3[55084] = 32'b00000000000000001011100000100110;
assign LUT_3[55085] = 32'b00000000000000010010001100000011;
assign LUT_3[55086] = 32'b00000000000000001101101000001010;
assign LUT_3[55087] = 32'b00000000000000010100010011100111;
assign LUT_3[55088] = 32'b00000000000000001100001100101101;
assign LUT_3[55089] = 32'b00000000000000010010111000001010;
assign LUT_3[55090] = 32'b00000000000000001110010100010001;
assign LUT_3[55091] = 32'b00000000000000010100111111101110;
assign LUT_3[55092] = 32'b00000000000000001001011010100011;
assign LUT_3[55093] = 32'b00000000000000010000000110000000;
assign LUT_3[55094] = 32'b00000000000000001011100010000111;
assign LUT_3[55095] = 32'b00000000000000010010001101100100;
assign LUT_3[55096] = 32'b00000000000000010001100101110011;
assign LUT_3[55097] = 32'b00000000000000011000010001010000;
assign LUT_3[55098] = 32'b00000000000000010011101101010111;
assign LUT_3[55099] = 32'b00000000000000011010011000110100;
assign LUT_3[55100] = 32'b00000000000000001110110011101001;
assign LUT_3[55101] = 32'b00000000000000010101011111000110;
assign LUT_3[55102] = 32'b00000000000000010000111011001101;
assign LUT_3[55103] = 32'b00000000000000010111100110101010;
assign LUT_3[55104] = 32'b00000000000000000111100011110101;
assign LUT_3[55105] = 32'b00000000000000001110001111010010;
assign LUT_3[55106] = 32'b00000000000000001001101011011001;
assign LUT_3[55107] = 32'b00000000000000010000010110110110;
assign LUT_3[55108] = 32'b00000000000000000100110001101011;
assign LUT_3[55109] = 32'b00000000000000001011011101001000;
assign LUT_3[55110] = 32'b00000000000000000110111001001111;
assign LUT_3[55111] = 32'b00000000000000001101100100101100;
assign LUT_3[55112] = 32'b00000000000000001100111100111011;
assign LUT_3[55113] = 32'b00000000000000010011101000011000;
assign LUT_3[55114] = 32'b00000000000000001111000100011111;
assign LUT_3[55115] = 32'b00000000000000010101101111111100;
assign LUT_3[55116] = 32'b00000000000000001010001010110001;
assign LUT_3[55117] = 32'b00000000000000010000110110001110;
assign LUT_3[55118] = 32'b00000000000000001100010010010101;
assign LUT_3[55119] = 32'b00000000000000010010111101110010;
assign LUT_3[55120] = 32'b00000000000000001010110110111000;
assign LUT_3[55121] = 32'b00000000000000010001100010010101;
assign LUT_3[55122] = 32'b00000000000000001100111110011100;
assign LUT_3[55123] = 32'b00000000000000010011101001111001;
assign LUT_3[55124] = 32'b00000000000000001000000100101110;
assign LUT_3[55125] = 32'b00000000000000001110110000001011;
assign LUT_3[55126] = 32'b00000000000000001010001100010010;
assign LUT_3[55127] = 32'b00000000000000010000110111101111;
assign LUT_3[55128] = 32'b00000000000000010000001111111110;
assign LUT_3[55129] = 32'b00000000000000010110111011011011;
assign LUT_3[55130] = 32'b00000000000000010010010111100010;
assign LUT_3[55131] = 32'b00000000000000011001000010111111;
assign LUT_3[55132] = 32'b00000000000000001101011101110100;
assign LUT_3[55133] = 32'b00000000000000010100001001010001;
assign LUT_3[55134] = 32'b00000000000000001111100101011000;
assign LUT_3[55135] = 32'b00000000000000010110010000110101;
assign LUT_3[55136] = 32'b00000000000000001000110010010101;
assign LUT_3[55137] = 32'b00000000000000001111011101110010;
assign LUT_3[55138] = 32'b00000000000000001010111001111001;
assign LUT_3[55139] = 32'b00000000000000010001100101010110;
assign LUT_3[55140] = 32'b00000000000000000110000000001011;
assign LUT_3[55141] = 32'b00000000000000001100101011101000;
assign LUT_3[55142] = 32'b00000000000000001000000111101111;
assign LUT_3[55143] = 32'b00000000000000001110110011001100;
assign LUT_3[55144] = 32'b00000000000000001110001011011011;
assign LUT_3[55145] = 32'b00000000000000010100110110111000;
assign LUT_3[55146] = 32'b00000000000000010000010010111111;
assign LUT_3[55147] = 32'b00000000000000010110111110011100;
assign LUT_3[55148] = 32'b00000000000000001011011001010001;
assign LUT_3[55149] = 32'b00000000000000010010000100101110;
assign LUT_3[55150] = 32'b00000000000000001101100000110101;
assign LUT_3[55151] = 32'b00000000000000010100001100010010;
assign LUT_3[55152] = 32'b00000000000000001100000101011000;
assign LUT_3[55153] = 32'b00000000000000010010110000110101;
assign LUT_3[55154] = 32'b00000000000000001110001100111100;
assign LUT_3[55155] = 32'b00000000000000010100111000011001;
assign LUT_3[55156] = 32'b00000000000000001001010011001110;
assign LUT_3[55157] = 32'b00000000000000001111111110101011;
assign LUT_3[55158] = 32'b00000000000000001011011010110010;
assign LUT_3[55159] = 32'b00000000000000010010000110001111;
assign LUT_3[55160] = 32'b00000000000000010001011110011110;
assign LUT_3[55161] = 32'b00000000000000011000001001111011;
assign LUT_3[55162] = 32'b00000000000000010011100110000010;
assign LUT_3[55163] = 32'b00000000000000011010010001011111;
assign LUT_3[55164] = 32'b00000000000000001110101100010100;
assign LUT_3[55165] = 32'b00000000000000010101010111110001;
assign LUT_3[55166] = 32'b00000000000000010000110011111000;
assign LUT_3[55167] = 32'b00000000000000010111011111010101;
assign LUT_3[55168] = 32'b00000000000000001001110110001000;
assign LUT_3[55169] = 32'b00000000000000010000100001100101;
assign LUT_3[55170] = 32'b00000000000000001011111101101100;
assign LUT_3[55171] = 32'b00000000000000010010101001001001;
assign LUT_3[55172] = 32'b00000000000000000111000011111110;
assign LUT_3[55173] = 32'b00000000000000001101101111011011;
assign LUT_3[55174] = 32'b00000000000000001001001011100010;
assign LUT_3[55175] = 32'b00000000000000001111110110111111;
assign LUT_3[55176] = 32'b00000000000000001111001111001110;
assign LUT_3[55177] = 32'b00000000000000010101111010101011;
assign LUT_3[55178] = 32'b00000000000000010001010110110010;
assign LUT_3[55179] = 32'b00000000000000011000000010001111;
assign LUT_3[55180] = 32'b00000000000000001100011101000100;
assign LUT_3[55181] = 32'b00000000000000010011001000100001;
assign LUT_3[55182] = 32'b00000000000000001110100100101000;
assign LUT_3[55183] = 32'b00000000000000010101010000000101;
assign LUT_3[55184] = 32'b00000000000000001101001001001011;
assign LUT_3[55185] = 32'b00000000000000010011110100101000;
assign LUT_3[55186] = 32'b00000000000000001111010000101111;
assign LUT_3[55187] = 32'b00000000000000010101111100001100;
assign LUT_3[55188] = 32'b00000000000000001010010111000001;
assign LUT_3[55189] = 32'b00000000000000010001000010011110;
assign LUT_3[55190] = 32'b00000000000000001100011110100101;
assign LUT_3[55191] = 32'b00000000000000010011001010000010;
assign LUT_3[55192] = 32'b00000000000000010010100010010001;
assign LUT_3[55193] = 32'b00000000000000011001001101101110;
assign LUT_3[55194] = 32'b00000000000000010100101001110101;
assign LUT_3[55195] = 32'b00000000000000011011010101010010;
assign LUT_3[55196] = 32'b00000000000000001111110000000111;
assign LUT_3[55197] = 32'b00000000000000010110011011100100;
assign LUT_3[55198] = 32'b00000000000000010001110111101011;
assign LUT_3[55199] = 32'b00000000000000011000100011001000;
assign LUT_3[55200] = 32'b00000000000000001011000100101000;
assign LUT_3[55201] = 32'b00000000000000010001110000000101;
assign LUT_3[55202] = 32'b00000000000000001101001100001100;
assign LUT_3[55203] = 32'b00000000000000010011110111101001;
assign LUT_3[55204] = 32'b00000000000000001000010010011110;
assign LUT_3[55205] = 32'b00000000000000001110111101111011;
assign LUT_3[55206] = 32'b00000000000000001010011010000010;
assign LUT_3[55207] = 32'b00000000000000010001000101011111;
assign LUT_3[55208] = 32'b00000000000000010000011101101110;
assign LUT_3[55209] = 32'b00000000000000010111001001001011;
assign LUT_3[55210] = 32'b00000000000000010010100101010010;
assign LUT_3[55211] = 32'b00000000000000011001010000101111;
assign LUT_3[55212] = 32'b00000000000000001101101011100100;
assign LUT_3[55213] = 32'b00000000000000010100010111000001;
assign LUT_3[55214] = 32'b00000000000000001111110011001000;
assign LUT_3[55215] = 32'b00000000000000010110011110100101;
assign LUT_3[55216] = 32'b00000000000000001110010111101011;
assign LUT_3[55217] = 32'b00000000000000010101000011001000;
assign LUT_3[55218] = 32'b00000000000000010000011111001111;
assign LUT_3[55219] = 32'b00000000000000010111001010101100;
assign LUT_3[55220] = 32'b00000000000000001011100101100001;
assign LUT_3[55221] = 32'b00000000000000010010010000111110;
assign LUT_3[55222] = 32'b00000000000000001101101101000101;
assign LUT_3[55223] = 32'b00000000000000010100011000100010;
assign LUT_3[55224] = 32'b00000000000000010011110000110001;
assign LUT_3[55225] = 32'b00000000000000011010011100001110;
assign LUT_3[55226] = 32'b00000000000000010101111000010101;
assign LUT_3[55227] = 32'b00000000000000011100100011110010;
assign LUT_3[55228] = 32'b00000000000000010000111110100111;
assign LUT_3[55229] = 32'b00000000000000010111101010000100;
assign LUT_3[55230] = 32'b00000000000000010011000110001011;
assign LUT_3[55231] = 32'b00000000000000011001110001101000;
assign LUT_3[55232] = 32'b00000000000000001001101110110011;
assign LUT_3[55233] = 32'b00000000000000010000011010010000;
assign LUT_3[55234] = 32'b00000000000000001011110110010111;
assign LUT_3[55235] = 32'b00000000000000010010100001110100;
assign LUT_3[55236] = 32'b00000000000000000110111100101001;
assign LUT_3[55237] = 32'b00000000000000001101101000000110;
assign LUT_3[55238] = 32'b00000000000000001001000100001101;
assign LUT_3[55239] = 32'b00000000000000001111101111101010;
assign LUT_3[55240] = 32'b00000000000000001111000111111001;
assign LUT_3[55241] = 32'b00000000000000010101110011010110;
assign LUT_3[55242] = 32'b00000000000000010001001111011101;
assign LUT_3[55243] = 32'b00000000000000010111111010111010;
assign LUT_3[55244] = 32'b00000000000000001100010101101111;
assign LUT_3[55245] = 32'b00000000000000010011000001001100;
assign LUT_3[55246] = 32'b00000000000000001110011101010011;
assign LUT_3[55247] = 32'b00000000000000010101001000110000;
assign LUT_3[55248] = 32'b00000000000000001101000001110110;
assign LUT_3[55249] = 32'b00000000000000010011101101010011;
assign LUT_3[55250] = 32'b00000000000000001111001001011010;
assign LUT_3[55251] = 32'b00000000000000010101110100110111;
assign LUT_3[55252] = 32'b00000000000000001010001111101100;
assign LUT_3[55253] = 32'b00000000000000010000111011001001;
assign LUT_3[55254] = 32'b00000000000000001100010111010000;
assign LUT_3[55255] = 32'b00000000000000010011000010101101;
assign LUT_3[55256] = 32'b00000000000000010010011010111100;
assign LUT_3[55257] = 32'b00000000000000011001000110011001;
assign LUT_3[55258] = 32'b00000000000000010100100010100000;
assign LUT_3[55259] = 32'b00000000000000011011001101111101;
assign LUT_3[55260] = 32'b00000000000000001111101000110010;
assign LUT_3[55261] = 32'b00000000000000010110010100001111;
assign LUT_3[55262] = 32'b00000000000000010001110000010110;
assign LUT_3[55263] = 32'b00000000000000011000011011110011;
assign LUT_3[55264] = 32'b00000000000000001010111101010011;
assign LUT_3[55265] = 32'b00000000000000010001101000110000;
assign LUT_3[55266] = 32'b00000000000000001101000100110111;
assign LUT_3[55267] = 32'b00000000000000010011110000010100;
assign LUT_3[55268] = 32'b00000000000000001000001011001001;
assign LUT_3[55269] = 32'b00000000000000001110110110100110;
assign LUT_3[55270] = 32'b00000000000000001010010010101101;
assign LUT_3[55271] = 32'b00000000000000010000111110001010;
assign LUT_3[55272] = 32'b00000000000000010000010110011001;
assign LUT_3[55273] = 32'b00000000000000010111000001110110;
assign LUT_3[55274] = 32'b00000000000000010010011101111101;
assign LUT_3[55275] = 32'b00000000000000011001001001011010;
assign LUT_3[55276] = 32'b00000000000000001101100100001111;
assign LUT_3[55277] = 32'b00000000000000010100001111101100;
assign LUT_3[55278] = 32'b00000000000000001111101011110011;
assign LUT_3[55279] = 32'b00000000000000010110010111010000;
assign LUT_3[55280] = 32'b00000000000000001110010000010110;
assign LUT_3[55281] = 32'b00000000000000010100111011110011;
assign LUT_3[55282] = 32'b00000000000000010000010111111010;
assign LUT_3[55283] = 32'b00000000000000010111000011010111;
assign LUT_3[55284] = 32'b00000000000000001011011110001100;
assign LUT_3[55285] = 32'b00000000000000010010001001101001;
assign LUT_3[55286] = 32'b00000000000000001101100101110000;
assign LUT_3[55287] = 32'b00000000000000010100010001001101;
assign LUT_3[55288] = 32'b00000000000000010011101001011100;
assign LUT_3[55289] = 32'b00000000000000011010010100111001;
assign LUT_3[55290] = 32'b00000000000000010101110001000000;
assign LUT_3[55291] = 32'b00000000000000011100011100011101;
assign LUT_3[55292] = 32'b00000000000000010000110111010010;
assign LUT_3[55293] = 32'b00000000000000010111100010101111;
assign LUT_3[55294] = 32'b00000000000000010010111110110110;
assign LUT_3[55295] = 32'b00000000000000011001101010010011;
assign LUT_3[55296] = 32'b00000000000000000011010111101110;
assign LUT_3[55297] = 32'b00000000000000001010000011001011;
assign LUT_3[55298] = 32'b00000000000000000101011111010010;
assign LUT_3[55299] = 32'b00000000000000001100001010101111;
assign LUT_3[55300] = 32'b00000000000000000000100101100100;
assign LUT_3[55301] = 32'b00000000000000000111010001000001;
assign LUT_3[55302] = 32'b00000000000000000010101101001000;
assign LUT_3[55303] = 32'b00000000000000001001011000100101;
assign LUT_3[55304] = 32'b00000000000000001000110000110100;
assign LUT_3[55305] = 32'b00000000000000001111011100010001;
assign LUT_3[55306] = 32'b00000000000000001010111000011000;
assign LUT_3[55307] = 32'b00000000000000010001100011110101;
assign LUT_3[55308] = 32'b00000000000000000101111110101010;
assign LUT_3[55309] = 32'b00000000000000001100101010000111;
assign LUT_3[55310] = 32'b00000000000000001000000110001110;
assign LUT_3[55311] = 32'b00000000000000001110110001101011;
assign LUT_3[55312] = 32'b00000000000000000110101010110001;
assign LUT_3[55313] = 32'b00000000000000001101010110001110;
assign LUT_3[55314] = 32'b00000000000000001000110010010101;
assign LUT_3[55315] = 32'b00000000000000001111011101110010;
assign LUT_3[55316] = 32'b00000000000000000011111000100111;
assign LUT_3[55317] = 32'b00000000000000001010100100000100;
assign LUT_3[55318] = 32'b00000000000000000110000000001011;
assign LUT_3[55319] = 32'b00000000000000001100101011101000;
assign LUT_3[55320] = 32'b00000000000000001100000011110111;
assign LUT_3[55321] = 32'b00000000000000010010101111010100;
assign LUT_3[55322] = 32'b00000000000000001110001011011011;
assign LUT_3[55323] = 32'b00000000000000010100110110111000;
assign LUT_3[55324] = 32'b00000000000000001001010001101101;
assign LUT_3[55325] = 32'b00000000000000001111111101001010;
assign LUT_3[55326] = 32'b00000000000000001011011001010001;
assign LUT_3[55327] = 32'b00000000000000010010000100101110;
assign LUT_3[55328] = 32'b00000000000000000100100110001110;
assign LUT_3[55329] = 32'b00000000000000001011010001101011;
assign LUT_3[55330] = 32'b00000000000000000110101101110010;
assign LUT_3[55331] = 32'b00000000000000001101011001001111;
assign LUT_3[55332] = 32'b00000000000000000001110100000100;
assign LUT_3[55333] = 32'b00000000000000001000011111100001;
assign LUT_3[55334] = 32'b00000000000000000011111011101000;
assign LUT_3[55335] = 32'b00000000000000001010100111000101;
assign LUT_3[55336] = 32'b00000000000000001001111111010100;
assign LUT_3[55337] = 32'b00000000000000010000101010110001;
assign LUT_3[55338] = 32'b00000000000000001100000110111000;
assign LUT_3[55339] = 32'b00000000000000010010110010010101;
assign LUT_3[55340] = 32'b00000000000000000111001101001010;
assign LUT_3[55341] = 32'b00000000000000001101111000100111;
assign LUT_3[55342] = 32'b00000000000000001001010100101110;
assign LUT_3[55343] = 32'b00000000000000010000000000001011;
assign LUT_3[55344] = 32'b00000000000000000111111001010001;
assign LUT_3[55345] = 32'b00000000000000001110100100101110;
assign LUT_3[55346] = 32'b00000000000000001010000000110101;
assign LUT_3[55347] = 32'b00000000000000010000101100010010;
assign LUT_3[55348] = 32'b00000000000000000101000111000111;
assign LUT_3[55349] = 32'b00000000000000001011110010100100;
assign LUT_3[55350] = 32'b00000000000000000111001110101011;
assign LUT_3[55351] = 32'b00000000000000001101111010001000;
assign LUT_3[55352] = 32'b00000000000000001101010010010111;
assign LUT_3[55353] = 32'b00000000000000010011111101110100;
assign LUT_3[55354] = 32'b00000000000000001111011001111011;
assign LUT_3[55355] = 32'b00000000000000010110000101011000;
assign LUT_3[55356] = 32'b00000000000000001010100000001101;
assign LUT_3[55357] = 32'b00000000000000010001001011101010;
assign LUT_3[55358] = 32'b00000000000000001100100111110001;
assign LUT_3[55359] = 32'b00000000000000010011010011001110;
assign LUT_3[55360] = 32'b00000000000000000011010000011001;
assign LUT_3[55361] = 32'b00000000000000001001111011110110;
assign LUT_3[55362] = 32'b00000000000000000101010111111101;
assign LUT_3[55363] = 32'b00000000000000001100000011011010;
assign LUT_3[55364] = 32'b00000000000000000000011110001111;
assign LUT_3[55365] = 32'b00000000000000000111001001101100;
assign LUT_3[55366] = 32'b00000000000000000010100101110011;
assign LUT_3[55367] = 32'b00000000000000001001010001010000;
assign LUT_3[55368] = 32'b00000000000000001000101001011111;
assign LUT_3[55369] = 32'b00000000000000001111010100111100;
assign LUT_3[55370] = 32'b00000000000000001010110001000011;
assign LUT_3[55371] = 32'b00000000000000010001011100100000;
assign LUT_3[55372] = 32'b00000000000000000101110111010101;
assign LUT_3[55373] = 32'b00000000000000001100100010110010;
assign LUT_3[55374] = 32'b00000000000000000111111110111001;
assign LUT_3[55375] = 32'b00000000000000001110101010010110;
assign LUT_3[55376] = 32'b00000000000000000110100011011100;
assign LUT_3[55377] = 32'b00000000000000001101001110111001;
assign LUT_3[55378] = 32'b00000000000000001000101011000000;
assign LUT_3[55379] = 32'b00000000000000001111010110011101;
assign LUT_3[55380] = 32'b00000000000000000011110001010010;
assign LUT_3[55381] = 32'b00000000000000001010011100101111;
assign LUT_3[55382] = 32'b00000000000000000101111000110110;
assign LUT_3[55383] = 32'b00000000000000001100100100010011;
assign LUT_3[55384] = 32'b00000000000000001011111100100010;
assign LUT_3[55385] = 32'b00000000000000010010100111111111;
assign LUT_3[55386] = 32'b00000000000000001110000100000110;
assign LUT_3[55387] = 32'b00000000000000010100101111100011;
assign LUT_3[55388] = 32'b00000000000000001001001010011000;
assign LUT_3[55389] = 32'b00000000000000001111110101110101;
assign LUT_3[55390] = 32'b00000000000000001011010001111100;
assign LUT_3[55391] = 32'b00000000000000010001111101011001;
assign LUT_3[55392] = 32'b00000000000000000100011110111001;
assign LUT_3[55393] = 32'b00000000000000001011001010010110;
assign LUT_3[55394] = 32'b00000000000000000110100110011101;
assign LUT_3[55395] = 32'b00000000000000001101010001111010;
assign LUT_3[55396] = 32'b00000000000000000001101100101111;
assign LUT_3[55397] = 32'b00000000000000001000011000001100;
assign LUT_3[55398] = 32'b00000000000000000011110100010011;
assign LUT_3[55399] = 32'b00000000000000001010011111110000;
assign LUT_3[55400] = 32'b00000000000000001001110111111111;
assign LUT_3[55401] = 32'b00000000000000010000100011011100;
assign LUT_3[55402] = 32'b00000000000000001011111111100011;
assign LUT_3[55403] = 32'b00000000000000010010101011000000;
assign LUT_3[55404] = 32'b00000000000000000111000101110101;
assign LUT_3[55405] = 32'b00000000000000001101110001010010;
assign LUT_3[55406] = 32'b00000000000000001001001101011001;
assign LUT_3[55407] = 32'b00000000000000001111111000110110;
assign LUT_3[55408] = 32'b00000000000000000111110001111100;
assign LUT_3[55409] = 32'b00000000000000001110011101011001;
assign LUT_3[55410] = 32'b00000000000000001001111001100000;
assign LUT_3[55411] = 32'b00000000000000010000100100111101;
assign LUT_3[55412] = 32'b00000000000000000100111111110010;
assign LUT_3[55413] = 32'b00000000000000001011101011001111;
assign LUT_3[55414] = 32'b00000000000000000111000111010110;
assign LUT_3[55415] = 32'b00000000000000001101110010110011;
assign LUT_3[55416] = 32'b00000000000000001101001011000010;
assign LUT_3[55417] = 32'b00000000000000010011110110011111;
assign LUT_3[55418] = 32'b00000000000000001111010010100110;
assign LUT_3[55419] = 32'b00000000000000010101111110000011;
assign LUT_3[55420] = 32'b00000000000000001010011000111000;
assign LUT_3[55421] = 32'b00000000000000010001000100010101;
assign LUT_3[55422] = 32'b00000000000000001100100000011100;
assign LUT_3[55423] = 32'b00000000000000010011001011111001;
assign LUT_3[55424] = 32'b00000000000000000101100010101100;
assign LUT_3[55425] = 32'b00000000000000001100001110001001;
assign LUT_3[55426] = 32'b00000000000000000111101010010000;
assign LUT_3[55427] = 32'b00000000000000001110010101101101;
assign LUT_3[55428] = 32'b00000000000000000010110000100010;
assign LUT_3[55429] = 32'b00000000000000001001011011111111;
assign LUT_3[55430] = 32'b00000000000000000100111000000110;
assign LUT_3[55431] = 32'b00000000000000001011100011100011;
assign LUT_3[55432] = 32'b00000000000000001010111011110010;
assign LUT_3[55433] = 32'b00000000000000010001100111001111;
assign LUT_3[55434] = 32'b00000000000000001101000011010110;
assign LUT_3[55435] = 32'b00000000000000010011101110110011;
assign LUT_3[55436] = 32'b00000000000000001000001001101000;
assign LUT_3[55437] = 32'b00000000000000001110110101000101;
assign LUT_3[55438] = 32'b00000000000000001010010001001100;
assign LUT_3[55439] = 32'b00000000000000010000111100101001;
assign LUT_3[55440] = 32'b00000000000000001000110101101111;
assign LUT_3[55441] = 32'b00000000000000001111100001001100;
assign LUT_3[55442] = 32'b00000000000000001010111101010011;
assign LUT_3[55443] = 32'b00000000000000010001101000110000;
assign LUT_3[55444] = 32'b00000000000000000110000011100101;
assign LUT_3[55445] = 32'b00000000000000001100101111000010;
assign LUT_3[55446] = 32'b00000000000000001000001011001001;
assign LUT_3[55447] = 32'b00000000000000001110110110100110;
assign LUT_3[55448] = 32'b00000000000000001110001110110101;
assign LUT_3[55449] = 32'b00000000000000010100111010010010;
assign LUT_3[55450] = 32'b00000000000000010000010110011001;
assign LUT_3[55451] = 32'b00000000000000010111000001110110;
assign LUT_3[55452] = 32'b00000000000000001011011100101011;
assign LUT_3[55453] = 32'b00000000000000010010001000001000;
assign LUT_3[55454] = 32'b00000000000000001101100100001111;
assign LUT_3[55455] = 32'b00000000000000010100001111101100;
assign LUT_3[55456] = 32'b00000000000000000110110001001100;
assign LUT_3[55457] = 32'b00000000000000001101011100101001;
assign LUT_3[55458] = 32'b00000000000000001000111000110000;
assign LUT_3[55459] = 32'b00000000000000001111100100001101;
assign LUT_3[55460] = 32'b00000000000000000011111111000010;
assign LUT_3[55461] = 32'b00000000000000001010101010011111;
assign LUT_3[55462] = 32'b00000000000000000110000110100110;
assign LUT_3[55463] = 32'b00000000000000001100110010000011;
assign LUT_3[55464] = 32'b00000000000000001100001010010010;
assign LUT_3[55465] = 32'b00000000000000010010110101101111;
assign LUT_3[55466] = 32'b00000000000000001110010001110110;
assign LUT_3[55467] = 32'b00000000000000010100111101010011;
assign LUT_3[55468] = 32'b00000000000000001001011000001000;
assign LUT_3[55469] = 32'b00000000000000010000000011100101;
assign LUT_3[55470] = 32'b00000000000000001011011111101100;
assign LUT_3[55471] = 32'b00000000000000010010001011001001;
assign LUT_3[55472] = 32'b00000000000000001010000100001111;
assign LUT_3[55473] = 32'b00000000000000010000101111101100;
assign LUT_3[55474] = 32'b00000000000000001100001011110011;
assign LUT_3[55475] = 32'b00000000000000010010110111010000;
assign LUT_3[55476] = 32'b00000000000000000111010010000101;
assign LUT_3[55477] = 32'b00000000000000001101111101100010;
assign LUT_3[55478] = 32'b00000000000000001001011001101001;
assign LUT_3[55479] = 32'b00000000000000010000000101000110;
assign LUT_3[55480] = 32'b00000000000000001111011101010101;
assign LUT_3[55481] = 32'b00000000000000010110001000110010;
assign LUT_3[55482] = 32'b00000000000000010001100100111001;
assign LUT_3[55483] = 32'b00000000000000011000010000010110;
assign LUT_3[55484] = 32'b00000000000000001100101011001011;
assign LUT_3[55485] = 32'b00000000000000010011010110101000;
assign LUT_3[55486] = 32'b00000000000000001110110010101111;
assign LUT_3[55487] = 32'b00000000000000010101011110001100;
assign LUT_3[55488] = 32'b00000000000000000101011011010111;
assign LUT_3[55489] = 32'b00000000000000001100000110110100;
assign LUT_3[55490] = 32'b00000000000000000111100010111011;
assign LUT_3[55491] = 32'b00000000000000001110001110011000;
assign LUT_3[55492] = 32'b00000000000000000010101001001101;
assign LUT_3[55493] = 32'b00000000000000001001010100101010;
assign LUT_3[55494] = 32'b00000000000000000100110000110001;
assign LUT_3[55495] = 32'b00000000000000001011011100001110;
assign LUT_3[55496] = 32'b00000000000000001010110100011101;
assign LUT_3[55497] = 32'b00000000000000010001011111111010;
assign LUT_3[55498] = 32'b00000000000000001100111100000001;
assign LUT_3[55499] = 32'b00000000000000010011100111011110;
assign LUT_3[55500] = 32'b00000000000000001000000010010011;
assign LUT_3[55501] = 32'b00000000000000001110101101110000;
assign LUT_3[55502] = 32'b00000000000000001010001001110111;
assign LUT_3[55503] = 32'b00000000000000010000110101010100;
assign LUT_3[55504] = 32'b00000000000000001000101110011010;
assign LUT_3[55505] = 32'b00000000000000001111011001110111;
assign LUT_3[55506] = 32'b00000000000000001010110101111110;
assign LUT_3[55507] = 32'b00000000000000010001100001011011;
assign LUT_3[55508] = 32'b00000000000000000101111100010000;
assign LUT_3[55509] = 32'b00000000000000001100100111101101;
assign LUT_3[55510] = 32'b00000000000000001000000011110100;
assign LUT_3[55511] = 32'b00000000000000001110101111010001;
assign LUT_3[55512] = 32'b00000000000000001110000111100000;
assign LUT_3[55513] = 32'b00000000000000010100110010111101;
assign LUT_3[55514] = 32'b00000000000000010000001111000100;
assign LUT_3[55515] = 32'b00000000000000010110111010100001;
assign LUT_3[55516] = 32'b00000000000000001011010101010110;
assign LUT_3[55517] = 32'b00000000000000010010000000110011;
assign LUT_3[55518] = 32'b00000000000000001101011100111010;
assign LUT_3[55519] = 32'b00000000000000010100001000010111;
assign LUT_3[55520] = 32'b00000000000000000110101001110111;
assign LUT_3[55521] = 32'b00000000000000001101010101010100;
assign LUT_3[55522] = 32'b00000000000000001000110001011011;
assign LUT_3[55523] = 32'b00000000000000001111011100111000;
assign LUT_3[55524] = 32'b00000000000000000011110111101101;
assign LUT_3[55525] = 32'b00000000000000001010100011001010;
assign LUT_3[55526] = 32'b00000000000000000101111111010001;
assign LUT_3[55527] = 32'b00000000000000001100101010101110;
assign LUT_3[55528] = 32'b00000000000000001100000010111101;
assign LUT_3[55529] = 32'b00000000000000010010101110011010;
assign LUT_3[55530] = 32'b00000000000000001110001010100001;
assign LUT_3[55531] = 32'b00000000000000010100110101111110;
assign LUT_3[55532] = 32'b00000000000000001001010000110011;
assign LUT_3[55533] = 32'b00000000000000001111111100010000;
assign LUT_3[55534] = 32'b00000000000000001011011000010111;
assign LUT_3[55535] = 32'b00000000000000010010000011110100;
assign LUT_3[55536] = 32'b00000000000000001001111100111010;
assign LUT_3[55537] = 32'b00000000000000010000101000010111;
assign LUT_3[55538] = 32'b00000000000000001100000100011110;
assign LUT_3[55539] = 32'b00000000000000010010101111111011;
assign LUT_3[55540] = 32'b00000000000000000111001010110000;
assign LUT_3[55541] = 32'b00000000000000001101110110001101;
assign LUT_3[55542] = 32'b00000000000000001001010010010100;
assign LUT_3[55543] = 32'b00000000000000001111111101110001;
assign LUT_3[55544] = 32'b00000000000000001111010110000000;
assign LUT_3[55545] = 32'b00000000000000010110000001011101;
assign LUT_3[55546] = 32'b00000000000000010001011101100100;
assign LUT_3[55547] = 32'b00000000000000011000001001000001;
assign LUT_3[55548] = 32'b00000000000000001100100011110110;
assign LUT_3[55549] = 32'b00000000000000010011001111010011;
assign LUT_3[55550] = 32'b00000000000000001110101011011010;
assign LUT_3[55551] = 32'b00000000000000010101010110110111;
assign LUT_3[55552] = 32'b11111111111111111111100111001111;
assign LUT_3[55553] = 32'b00000000000000000110010010101100;
assign LUT_3[55554] = 32'b00000000000000000001101110110011;
assign LUT_3[55555] = 32'b00000000000000001000011010010000;
assign LUT_3[55556] = 32'b11111111111111111100110101000101;
assign LUT_3[55557] = 32'b00000000000000000011100000100010;
assign LUT_3[55558] = 32'b11111111111111111110111100101001;
assign LUT_3[55559] = 32'b00000000000000000101101000000110;
assign LUT_3[55560] = 32'b00000000000000000101000000010101;
assign LUT_3[55561] = 32'b00000000000000001011101011110010;
assign LUT_3[55562] = 32'b00000000000000000111000111111001;
assign LUT_3[55563] = 32'b00000000000000001101110011010110;
assign LUT_3[55564] = 32'b00000000000000000010001110001011;
assign LUT_3[55565] = 32'b00000000000000001000111001101000;
assign LUT_3[55566] = 32'b00000000000000000100010101101111;
assign LUT_3[55567] = 32'b00000000000000001011000001001100;
assign LUT_3[55568] = 32'b00000000000000000010111010010010;
assign LUT_3[55569] = 32'b00000000000000001001100101101111;
assign LUT_3[55570] = 32'b00000000000000000101000001110110;
assign LUT_3[55571] = 32'b00000000000000001011101101010011;
assign LUT_3[55572] = 32'b00000000000000000000001000001000;
assign LUT_3[55573] = 32'b00000000000000000110110011100101;
assign LUT_3[55574] = 32'b00000000000000000010001111101100;
assign LUT_3[55575] = 32'b00000000000000001000111011001001;
assign LUT_3[55576] = 32'b00000000000000001000010011011000;
assign LUT_3[55577] = 32'b00000000000000001110111110110101;
assign LUT_3[55578] = 32'b00000000000000001010011010111100;
assign LUT_3[55579] = 32'b00000000000000010001000110011001;
assign LUT_3[55580] = 32'b00000000000000000101100001001110;
assign LUT_3[55581] = 32'b00000000000000001100001100101011;
assign LUT_3[55582] = 32'b00000000000000000111101000110010;
assign LUT_3[55583] = 32'b00000000000000001110010100001111;
assign LUT_3[55584] = 32'b00000000000000000000110101101111;
assign LUT_3[55585] = 32'b00000000000000000111100001001100;
assign LUT_3[55586] = 32'b00000000000000000010111101010011;
assign LUT_3[55587] = 32'b00000000000000001001101000110000;
assign LUT_3[55588] = 32'b11111111111111111110000011100101;
assign LUT_3[55589] = 32'b00000000000000000100101111000010;
assign LUT_3[55590] = 32'b00000000000000000000001011001001;
assign LUT_3[55591] = 32'b00000000000000000110110110100110;
assign LUT_3[55592] = 32'b00000000000000000110001110110101;
assign LUT_3[55593] = 32'b00000000000000001100111010010010;
assign LUT_3[55594] = 32'b00000000000000001000010110011001;
assign LUT_3[55595] = 32'b00000000000000001111000001110110;
assign LUT_3[55596] = 32'b00000000000000000011011100101011;
assign LUT_3[55597] = 32'b00000000000000001010001000001000;
assign LUT_3[55598] = 32'b00000000000000000101100100001111;
assign LUT_3[55599] = 32'b00000000000000001100001111101100;
assign LUT_3[55600] = 32'b00000000000000000100001000110010;
assign LUT_3[55601] = 32'b00000000000000001010110100001111;
assign LUT_3[55602] = 32'b00000000000000000110010000010110;
assign LUT_3[55603] = 32'b00000000000000001100111011110011;
assign LUT_3[55604] = 32'b00000000000000000001010110101000;
assign LUT_3[55605] = 32'b00000000000000001000000010000101;
assign LUT_3[55606] = 32'b00000000000000000011011110001100;
assign LUT_3[55607] = 32'b00000000000000001010001001101001;
assign LUT_3[55608] = 32'b00000000000000001001100001111000;
assign LUT_3[55609] = 32'b00000000000000010000001101010101;
assign LUT_3[55610] = 32'b00000000000000001011101001011100;
assign LUT_3[55611] = 32'b00000000000000010010010100111001;
assign LUT_3[55612] = 32'b00000000000000000110101111101110;
assign LUT_3[55613] = 32'b00000000000000001101011011001011;
assign LUT_3[55614] = 32'b00000000000000001000110111010010;
assign LUT_3[55615] = 32'b00000000000000001111100010101111;
assign LUT_3[55616] = 32'b11111111111111111111011111111010;
assign LUT_3[55617] = 32'b00000000000000000110001011010111;
assign LUT_3[55618] = 32'b00000000000000000001100111011110;
assign LUT_3[55619] = 32'b00000000000000001000010010111011;
assign LUT_3[55620] = 32'b11111111111111111100101101110000;
assign LUT_3[55621] = 32'b00000000000000000011011001001101;
assign LUT_3[55622] = 32'b11111111111111111110110101010100;
assign LUT_3[55623] = 32'b00000000000000000101100000110001;
assign LUT_3[55624] = 32'b00000000000000000100111001000000;
assign LUT_3[55625] = 32'b00000000000000001011100100011101;
assign LUT_3[55626] = 32'b00000000000000000111000000100100;
assign LUT_3[55627] = 32'b00000000000000001101101100000001;
assign LUT_3[55628] = 32'b00000000000000000010000110110110;
assign LUT_3[55629] = 32'b00000000000000001000110010010011;
assign LUT_3[55630] = 32'b00000000000000000100001110011010;
assign LUT_3[55631] = 32'b00000000000000001010111001110111;
assign LUT_3[55632] = 32'b00000000000000000010110010111101;
assign LUT_3[55633] = 32'b00000000000000001001011110011010;
assign LUT_3[55634] = 32'b00000000000000000100111010100001;
assign LUT_3[55635] = 32'b00000000000000001011100101111110;
assign LUT_3[55636] = 32'b00000000000000000000000000110011;
assign LUT_3[55637] = 32'b00000000000000000110101100010000;
assign LUT_3[55638] = 32'b00000000000000000010001000010111;
assign LUT_3[55639] = 32'b00000000000000001000110011110100;
assign LUT_3[55640] = 32'b00000000000000001000001100000011;
assign LUT_3[55641] = 32'b00000000000000001110110111100000;
assign LUT_3[55642] = 32'b00000000000000001010010011100111;
assign LUT_3[55643] = 32'b00000000000000010000111111000100;
assign LUT_3[55644] = 32'b00000000000000000101011001111001;
assign LUT_3[55645] = 32'b00000000000000001100000101010110;
assign LUT_3[55646] = 32'b00000000000000000111100001011101;
assign LUT_3[55647] = 32'b00000000000000001110001100111010;
assign LUT_3[55648] = 32'b00000000000000000000101110011010;
assign LUT_3[55649] = 32'b00000000000000000111011001110111;
assign LUT_3[55650] = 32'b00000000000000000010110101111110;
assign LUT_3[55651] = 32'b00000000000000001001100001011011;
assign LUT_3[55652] = 32'b11111111111111111101111100010000;
assign LUT_3[55653] = 32'b00000000000000000100100111101101;
assign LUT_3[55654] = 32'b00000000000000000000000011110100;
assign LUT_3[55655] = 32'b00000000000000000110101111010001;
assign LUT_3[55656] = 32'b00000000000000000110000111100000;
assign LUT_3[55657] = 32'b00000000000000001100110010111101;
assign LUT_3[55658] = 32'b00000000000000001000001111000100;
assign LUT_3[55659] = 32'b00000000000000001110111010100001;
assign LUT_3[55660] = 32'b00000000000000000011010101010110;
assign LUT_3[55661] = 32'b00000000000000001010000000110011;
assign LUT_3[55662] = 32'b00000000000000000101011100111010;
assign LUT_3[55663] = 32'b00000000000000001100001000010111;
assign LUT_3[55664] = 32'b00000000000000000100000001011101;
assign LUT_3[55665] = 32'b00000000000000001010101100111010;
assign LUT_3[55666] = 32'b00000000000000000110001001000001;
assign LUT_3[55667] = 32'b00000000000000001100110100011110;
assign LUT_3[55668] = 32'b00000000000000000001001111010011;
assign LUT_3[55669] = 32'b00000000000000000111111010110000;
assign LUT_3[55670] = 32'b00000000000000000011010110110111;
assign LUT_3[55671] = 32'b00000000000000001010000010010100;
assign LUT_3[55672] = 32'b00000000000000001001011010100011;
assign LUT_3[55673] = 32'b00000000000000010000000110000000;
assign LUT_3[55674] = 32'b00000000000000001011100010000111;
assign LUT_3[55675] = 32'b00000000000000010010001101100100;
assign LUT_3[55676] = 32'b00000000000000000110101000011001;
assign LUT_3[55677] = 32'b00000000000000001101010011110110;
assign LUT_3[55678] = 32'b00000000000000001000101111111101;
assign LUT_3[55679] = 32'b00000000000000001111011011011010;
assign LUT_3[55680] = 32'b00000000000000000001110010001101;
assign LUT_3[55681] = 32'b00000000000000001000011101101010;
assign LUT_3[55682] = 32'b00000000000000000011111001110001;
assign LUT_3[55683] = 32'b00000000000000001010100101001110;
assign LUT_3[55684] = 32'b11111111111111111111000000000011;
assign LUT_3[55685] = 32'b00000000000000000101101011100000;
assign LUT_3[55686] = 32'b00000000000000000001000111100111;
assign LUT_3[55687] = 32'b00000000000000000111110011000100;
assign LUT_3[55688] = 32'b00000000000000000111001011010011;
assign LUT_3[55689] = 32'b00000000000000001101110110110000;
assign LUT_3[55690] = 32'b00000000000000001001010010110111;
assign LUT_3[55691] = 32'b00000000000000001111111110010100;
assign LUT_3[55692] = 32'b00000000000000000100011001001001;
assign LUT_3[55693] = 32'b00000000000000001011000100100110;
assign LUT_3[55694] = 32'b00000000000000000110100000101101;
assign LUT_3[55695] = 32'b00000000000000001101001100001010;
assign LUT_3[55696] = 32'b00000000000000000101000101010000;
assign LUT_3[55697] = 32'b00000000000000001011110000101101;
assign LUT_3[55698] = 32'b00000000000000000111001100110100;
assign LUT_3[55699] = 32'b00000000000000001101111000010001;
assign LUT_3[55700] = 32'b00000000000000000010010011000110;
assign LUT_3[55701] = 32'b00000000000000001000111110100011;
assign LUT_3[55702] = 32'b00000000000000000100011010101010;
assign LUT_3[55703] = 32'b00000000000000001011000110000111;
assign LUT_3[55704] = 32'b00000000000000001010011110010110;
assign LUT_3[55705] = 32'b00000000000000010001001001110011;
assign LUT_3[55706] = 32'b00000000000000001100100101111010;
assign LUT_3[55707] = 32'b00000000000000010011010001010111;
assign LUT_3[55708] = 32'b00000000000000000111101100001100;
assign LUT_3[55709] = 32'b00000000000000001110010111101001;
assign LUT_3[55710] = 32'b00000000000000001001110011110000;
assign LUT_3[55711] = 32'b00000000000000010000011111001101;
assign LUT_3[55712] = 32'b00000000000000000011000000101101;
assign LUT_3[55713] = 32'b00000000000000001001101100001010;
assign LUT_3[55714] = 32'b00000000000000000101001000010001;
assign LUT_3[55715] = 32'b00000000000000001011110011101110;
assign LUT_3[55716] = 32'b00000000000000000000001110100011;
assign LUT_3[55717] = 32'b00000000000000000110111010000000;
assign LUT_3[55718] = 32'b00000000000000000010010110000111;
assign LUT_3[55719] = 32'b00000000000000001001000001100100;
assign LUT_3[55720] = 32'b00000000000000001000011001110011;
assign LUT_3[55721] = 32'b00000000000000001111000101010000;
assign LUT_3[55722] = 32'b00000000000000001010100001010111;
assign LUT_3[55723] = 32'b00000000000000010001001100110100;
assign LUT_3[55724] = 32'b00000000000000000101100111101001;
assign LUT_3[55725] = 32'b00000000000000001100010011000110;
assign LUT_3[55726] = 32'b00000000000000000111101111001101;
assign LUT_3[55727] = 32'b00000000000000001110011010101010;
assign LUT_3[55728] = 32'b00000000000000000110010011110000;
assign LUT_3[55729] = 32'b00000000000000001100111111001101;
assign LUT_3[55730] = 32'b00000000000000001000011011010100;
assign LUT_3[55731] = 32'b00000000000000001111000110110001;
assign LUT_3[55732] = 32'b00000000000000000011100001100110;
assign LUT_3[55733] = 32'b00000000000000001010001101000011;
assign LUT_3[55734] = 32'b00000000000000000101101001001010;
assign LUT_3[55735] = 32'b00000000000000001100010100100111;
assign LUT_3[55736] = 32'b00000000000000001011101100110110;
assign LUT_3[55737] = 32'b00000000000000010010011000010011;
assign LUT_3[55738] = 32'b00000000000000001101110100011010;
assign LUT_3[55739] = 32'b00000000000000010100011111110111;
assign LUT_3[55740] = 32'b00000000000000001000111010101100;
assign LUT_3[55741] = 32'b00000000000000001111100110001001;
assign LUT_3[55742] = 32'b00000000000000001011000010010000;
assign LUT_3[55743] = 32'b00000000000000010001101101101101;
assign LUT_3[55744] = 32'b00000000000000000001101010111000;
assign LUT_3[55745] = 32'b00000000000000001000010110010101;
assign LUT_3[55746] = 32'b00000000000000000011110010011100;
assign LUT_3[55747] = 32'b00000000000000001010011101111001;
assign LUT_3[55748] = 32'b11111111111111111110111000101110;
assign LUT_3[55749] = 32'b00000000000000000101100100001011;
assign LUT_3[55750] = 32'b00000000000000000001000000010010;
assign LUT_3[55751] = 32'b00000000000000000111101011101111;
assign LUT_3[55752] = 32'b00000000000000000111000011111110;
assign LUT_3[55753] = 32'b00000000000000001101101111011011;
assign LUT_3[55754] = 32'b00000000000000001001001011100010;
assign LUT_3[55755] = 32'b00000000000000001111110110111111;
assign LUT_3[55756] = 32'b00000000000000000100010001110100;
assign LUT_3[55757] = 32'b00000000000000001010111101010001;
assign LUT_3[55758] = 32'b00000000000000000110011001011000;
assign LUT_3[55759] = 32'b00000000000000001101000100110101;
assign LUT_3[55760] = 32'b00000000000000000100111101111011;
assign LUT_3[55761] = 32'b00000000000000001011101001011000;
assign LUT_3[55762] = 32'b00000000000000000111000101011111;
assign LUT_3[55763] = 32'b00000000000000001101110000111100;
assign LUT_3[55764] = 32'b00000000000000000010001011110001;
assign LUT_3[55765] = 32'b00000000000000001000110111001110;
assign LUT_3[55766] = 32'b00000000000000000100010011010101;
assign LUT_3[55767] = 32'b00000000000000001010111110110010;
assign LUT_3[55768] = 32'b00000000000000001010010111000001;
assign LUT_3[55769] = 32'b00000000000000010001000010011110;
assign LUT_3[55770] = 32'b00000000000000001100011110100101;
assign LUT_3[55771] = 32'b00000000000000010011001010000010;
assign LUT_3[55772] = 32'b00000000000000000111100100110111;
assign LUT_3[55773] = 32'b00000000000000001110010000010100;
assign LUT_3[55774] = 32'b00000000000000001001101100011011;
assign LUT_3[55775] = 32'b00000000000000010000010111111000;
assign LUT_3[55776] = 32'b00000000000000000010111001011000;
assign LUT_3[55777] = 32'b00000000000000001001100100110101;
assign LUT_3[55778] = 32'b00000000000000000101000000111100;
assign LUT_3[55779] = 32'b00000000000000001011101100011001;
assign LUT_3[55780] = 32'b00000000000000000000000111001110;
assign LUT_3[55781] = 32'b00000000000000000110110010101011;
assign LUT_3[55782] = 32'b00000000000000000010001110110010;
assign LUT_3[55783] = 32'b00000000000000001000111010001111;
assign LUT_3[55784] = 32'b00000000000000001000010010011110;
assign LUT_3[55785] = 32'b00000000000000001110111101111011;
assign LUT_3[55786] = 32'b00000000000000001010011010000010;
assign LUT_3[55787] = 32'b00000000000000010001000101011111;
assign LUT_3[55788] = 32'b00000000000000000101100000010100;
assign LUT_3[55789] = 32'b00000000000000001100001011110001;
assign LUT_3[55790] = 32'b00000000000000000111100111111000;
assign LUT_3[55791] = 32'b00000000000000001110010011010101;
assign LUT_3[55792] = 32'b00000000000000000110001100011011;
assign LUT_3[55793] = 32'b00000000000000001100110111111000;
assign LUT_3[55794] = 32'b00000000000000001000010011111111;
assign LUT_3[55795] = 32'b00000000000000001110111111011100;
assign LUT_3[55796] = 32'b00000000000000000011011010010001;
assign LUT_3[55797] = 32'b00000000000000001010000101101110;
assign LUT_3[55798] = 32'b00000000000000000101100001110101;
assign LUT_3[55799] = 32'b00000000000000001100001101010010;
assign LUT_3[55800] = 32'b00000000000000001011100101100001;
assign LUT_3[55801] = 32'b00000000000000010010010000111110;
assign LUT_3[55802] = 32'b00000000000000001101101101000101;
assign LUT_3[55803] = 32'b00000000000000010100011000100010;
assign LUT_3[55804] = 32'b00000000000000001000110011010111;
assign LUT_3[55805] = 32'b00000000000000001111011110110100;
assign LUT_3[55806] = 32'b00000000000000001010111010111011;
assign LUT_3[55807] = 32'b00000000000000010001100110011000;
assign LUT_3[55808] = 32'b00000000000000000110101100111010;
assign LUT_3[55809] = 32'b00000000000000001101011000010111;
assign LUT_3[55810] = 32'b00000000000000001000110100011110;
assign LUT_3[55811] = 32'b00000000000000001111011111111011;
assign LUT_3[55812] = 32'b00000000000000000011111010110000;
assign LUT_3[55813] = 32'b00000000000000001010100110001101;
assign LUT_3[55814] = 32'b00000000000000000110000010010100;
assign LUT_3[55815] = 32'b00000000000000001100101101110001;
assign LUT_3[55816] = 32'b00000000000000001100000110000000;
assign LUT_3[55817] = 32'b00000000000000010010110001011101;
assign LUT_3[55818] = 32'b00000000000000001110001101100100;
assign LUT_3[55819] = 32'b00000000000000010100111001000001;
assign LUT_3[55820] = 32'b00000000000000001001010011110110;
assign LUT_3[55821] = 32'b00000000000000001111111111010011;
assign LUT_3[55822] = 32'b00000000000000001011011011011010;
assign LUT_3[55823] = 32'b00000000000000010010000110110111;
assign LUT_3[55824] = 32'b00000000000000001001111111111101;
assign LUT_3[55825] = 32'b00000000000000010000101011011010;
assign LUT_3[55826] = 32'b00000000000000001100000111100001;
assign LUT_3[55827] = 32'b00000000000000010010110010111110;
assign LUT_3[55828] = 32'b00000000000000000111001101110011;
assign LUT_3[55829] = 32'b00000000000000001101111001010000;
assign LUT_3[55830] = 32'b00000000000000001001010101010111;
assign LUT_3[55831] = 32'b00000000000000010000000000110100;
assign LUT_3[55832] = 32'b00000000000000001111011001000011;
assign LUT_3[55833] = 32'b00000000000000010110000100100000;
assign LUT_3[55834] = 32'b00000000000000010001100000100111;
assign LUT_3[55835] = 32'b00000000000000011000001100000100;
assign LUT_3[55836] = 32'b00000000000000001100100110111001;
assign LUT_3[55837] = 32'b00000000000000010011010010010110;
assign LUT_3[55838] = 32'b00000000000000001110101110011101;
assign LUT_3[55839] = 32'b00000000000000010101011001111010;
assign LUT_3[55840] = 32'b00000000000000000111111011011010;
assign LUT_3[55841] = 32'b00000000000000001110100110110111;
assign LUT_3[55842] = 32'b00000000000000001010000010111110;
assign LUT_3[55843] = 32'b00000000000000010000101110011011;
assign LUT_3[55844] = 32'b00000000000000000101001001010000;
assign LUT_3[55845] = 32'b00000000000000001011110100101101;
assign LUT_3[55846] = 32'b00000000000000000111010000110100;
assign LUT_3[55847] = 32'b00000000000000001101111100010001;
assign LUT_3[55848] = 32'b00000000000000001101010100100000;
assign LUT_3[55849] = 32'b00000000000000010011111111111101;
assign LUT_3[55850] = 32'b00000000000000001111011100000100;
assign LUT_3[55851] = 32'b00000000000000010110000111100001;
assign LUT_3[55852] = 32'b00000000000000001010100010010110;
assign LUT_3[55853] = 32'b00000000000000010001001101110011;
assign LUT_3[55854] = 32'b00000000000000001100101001111010;
assign LUT_3[55855] = 32'b00000000000000010011010101010111;
assign LUT_3[55856] = 32'b00000000000000001011001110011101;
assign LUT_3[55857] = 32'b00000000000000010001111001111010;
assign LUT_3[55858] = 32'b00000000000000001101010110000001;
assign LUT_3[55859] = 32'b00000000000000010100000001011110;
assign LUT_3[55860] = 32'b00000000000000001000011100010011;
assign LUT_3[55861] = 32'b00000000000000001111000111110000;
assign LUT_3[55862] = 32'b00000000000000001010100011110111;
assign LUT_3[55863] = 32'b00000000000000010001001111010100;
assign LUT_3[55864] = 32'b00000000000000010000100111100011;
assign LUT_3[55865] = 32'b00000000000000010111010011000000;
assign LUT_3[55866] = 32'b00000000000000010010101111000111;
assign LUT_3[55867] = 32'b00000000000000011001011010100100;
assign LUT_3[55868] = 32'b00000000000000001101110101011001;
assign LUT_3[55869] = 32'b00000000000000010100100000110110;
assign LUT_3[55870] = 32'b00000000000000001111111100111101;
assign LUT_3[55871] = 32'b00000000000000010110101000011010;
assign LUT_3[55872] = 32'b00000000000000000110100101100101;
assign LUT_3[55873] = 32'b00000000000000001101010001000010;
assign LUT_3[55874] = 32'b00000000000000001000101101001001;
assign LUT_3[55875] = 32'b00000000000000001111011000100110;
assign LUT_3[55876] = 32'b00000000000000000011110011011011;
assign LUT_3[55877] = 32'b00000000000000001010011110111000;
assign LUT_3[55878] = 32'b00000000000000000101111010111111;
assign LUT_3[55879] = 32'b00000000000000001100100110011100;
assign LUT_3[55880] = 32'b00000000000000001011111110101011;
assign LUT_3[55881] = 32'b00000000000000010010101010001000;
assign LUT_3[55882] = 32'b00000000000000001110000110001111;
assign LUT_3[55883] = 32'b00000000000000010100110001101100;
assign LUT_3[55884] = 32'b00000000000000001001001100100001;
assign LUT_3[55885] = 32'b00000000000000001111110111111110;
assign LUT_3[55886] = 32'b00000000000000001011010100000101;
assign LUT_3[55887] = 32'b00000000000000010001111111100010;
assign LUT_3[55888] = 32'b00000000000000001001111000101000;
assign LUT_3[55889] = 32'b00000000000000010000100100000101;
assign LUT_3[55890] = 32'b00000000000000001100000000001100;
assign LUT_3[55891] = 32'b00000000000000010010101011101001;
assign LUT_3[55892] = 32'b00000000000000000111000110011110;
assign LUT_3[55893] = 32'b00000000000000001101110001111011;
assign LUT_3[55894] = 32'b00000000000000001001001110000010;
assign LUT_3[55895] = 32'b00000000000000001111111001011111;
assign LUT_3[55896] = 32'b00000000000000001111010001101110;
assign LUT_3[55897] = 32'b00000000000000010101111101001011;
assign LUT_3[55898] = 32'b00000000000000010001011001010010;
assign LUT_3[55899] = 32'b00000000000000011000000100101111;
assign LUT_3[55900] = 32'b00000000000000001100011111100100;
assign LUT_3[55901] = 32'b00000000000000010011001011000001;
assign LUT_3[55902] = 32'b00000000000000001110100111001000;
assign LUT_3[55903] = 32'b00000000000000010101010010100101;
assign LUT_3[55904] = 32'b00000000000000000111110100000101;
assign LUT_3[55905] = 32'b00000000000000001110011111100010;
assign LUT_3[55906] = 32'b00000000000000001001111011101001;
assign LUT_3[55907] = 32'b00000000000000010000100111000110;
assign LUT_3[55908] = 32'b00000000000000000101000001111011;
assign LUT_3[55909] = 32'b00000000000000001011101101011000;
assign LUT_3[55910] = 32'b00000000000000000111001001011111;
assign LUT_3[55911] = 32'b00000000000000001101110100111100;
assign LUT_3[55912] = 32'b00000000000000001101001101001011;
assign LUT_3[55913] = 32'b00000000000000010011111000101000;
assign LUT_3[55914] = 32'b00000000000000001111010100101111;
assign LUT_3[55915] = 32'b00000000000000010110000000001100;
assign LUT_3[55916] = 32'b00000000000000001010011011000001;
assign LUT_3[55917] = 32'b00000000000000010001000110011110;
assign LUT_3[55918] = 32'b00000000000000001100100010100101;
assign LUT_3[55919] = 32'b00000000000000010011001110000010;
assign LUT_3[55920] = 32'b00000000000000001011000111001000;
assign LUT_3[55921] = 32'b00000000000000010001110010100101;
assign LUT_3[55922] = 32'b00000000000000001101001110101100;
assign LUT_3[55923] = 32'b00000000000000010011111010001001;
assign LUT_3[55924] = 32'b00000000000000001000010100111110;
assign LUT_3[55925] = 32'b00000000000000001111000000011011;
assign LUT_3[55926] = 32'b00000000000000001010011100100010;
assign LUT_3[55927] = 32'b00000000000000010001000111111111;
assign LUT_3[55928] = 32'b00000000000000010000100000001110;
assign LUT_3[55929] = 32'b00000000000000010111001011101011;
assign LUT_3[55930] = 32'b00000000000000010010100111110010;
assign LUT_3[55931] = 32'b00000000000000011001010011001111;
assign LUT_3[55932] = 32'b00000000000000001101101110000100;
assign LUT_3[55933] = 32'b00000000000000010100011001100001;
assign LUT_3[55934] = 32'b00000000000000001111110101101000;
assign LUT_3[55935] = 32'b00000000000000010110100001000101;
assign LUT_3[55936] = 32'b00000000000000001000110111111000;
assign LUT_3[55937] = 32'b00000000000000001111100011010101;
assign LUT_3[55938] = 32'b00000000000000001010111111011100;
assign LUT_3[55939] = 32'b00000000000000010001101010111001;
assign LUT_3[55940] = 32'b00000000000000000110000101101110;
assign LUT_3[55941] = 32'b00000000000000001100110001001011;
assign LUT_3[55942] = 32'b00000000000000001000001101010010;
assign LUT_3[55943] = 32'b00000000000000001110111000101111;
assign LUT_3[55944] = 32'b00000000000000001110010000111110;
assign LUT_3[55945] = 32'b00000000000000010100111100011011;
assign LUT_3[55946] = 32'b00000000000000010000011000100010;
assign LUT_3[55947] = 32'b00000000000000010111000011111111;
assign LUT_3[55948] = 32'b00000000000000001011011110110100;
assign LUT_3[55949] = 32'b00000000000000010010001010010001;
assign LUT_3[55950] = 32'b00000000000000001101100110011000;
assign LUT_3[55951] = 32'b00000000000000010100010001110101;
assign LUT_3[55952] = 32'b00000000000000001100001010111011;
assign LUT_3[55953] = 32'b00000000000000010010110110011000;
assign LUT_3[55954] = 32'b00000000000000001110010010011111;
assign LUT_3[55955] = 32'b00000000000000010100111101111100;
assign LUT_3[55956] = 32'b00000000000000001001011000110001;
assign LUT_3[55957] = 32'b00000000000000010000000100001110;
assign LUT_3[55958] = 32'b00000000000000001011100000010101;
assign LUT_3[55959] = 32'b00000000000000010010001011110010;
assign LUT_3[55960] = 32'b00000000000000010001100100000001;
assign LUT_3[55961] = 32'b00000000000000011000001111011110;
assign LUT_3[55962] = 32'b00000000000000010011101011100101;
assign LUT_3[55963] = 32'b00000000000000011010010111000010;
assign LUT_3[55964] = 32'b00000000000000001110110001110111;
assign LUT_3[55965] = 32'b00000000000000010101011101010100;
assign LUT_3[55966] = 32'b00000000000000010000111001011011;
assign LUT_3[55967] = 32'b00000000000000010111100100111000;
assign LUT_3[55968] = 32'b00000000000000001010000110011000;
assign LUT_3[55969] = 32'b00000000000000010000110001110101;
assign LUT_3[55970] = 32'b00000000000000001100001101111100;
assign LUT_3[55971] = 32'b00000000000000010010111001011001;
assign LUT_3[55972] = 32'b00000000000000000111010100001110;
assign LUT_3[55973] = 32'b00000000000000001101111111101011;
assign LUT_3[55974] = 32'b00000000000000001001011011110010;
assign LUT_3[55975] = 32'b00000000000000010000000111001111;
assign LUT_3[55976] = 32'b00000000000000001111011111011110;
assign LUT_3[55977] = 32'b00000000000000010110001010111011;
assign LUT_3[55978] = 32'b00000000000000010001100111000010;
assign LUT_3[55979] = 32'b00000000000000011000010010011111;
assign LUT_3[55980] = 32'b00000000000000001100101101010100;
assign LUT_3[55981] = 32'b00000000000000010011011000110001;
assign LUT_3[55982] = 32'b00000000000000001110110100111000;
assign LUT_3[55983] = 32'b00000000000000010101100000010101;
assign LUT_3[55984] = 32'b00000000000000001101011001011011;
assign LUT_3[55985] = 32'b00000000000000010100000100111000;
assign LUT_3[55986] = 32'b00000000000000001111100000111111;
assign LUT_3[55987] = 32'b00000000000000010110001100011100;
assign LUT_3[55988] = 32'b00000000000000001010100111010001;
assign LUT_3[55989] = 32'b00000000000000010001010010101110;
assign LUT_3[55990] = 32'b00000000000000001100101110110101;
assign LUT_3[55991] = 32'b00000000000000010011011010010010;
assign LUT_3[55992] = 32'b00000000000000010010110010100001;
assign LUT_3[55993] = 32'b00000000000000011001011101111110;
assign LUT_3[55994] = 32'b00000000000000010100111010000101;
assign LUT_3[55995] = 32'b00000000000000011011100101100010;
assign LUT_3[55996] = 32'b00000000000000010000000000010111;
assign LUT_3[55997] = 32'b00000000000000010110101011110100;
assign LUT_3[55998] = 32'b00000000000000010010000111111011;
assign LUT_3[55999] = 32'b00000000000000011000110011011000;
assign LUT_3[56000] = 32'b00000000000000001000110000100011;
assign LUT_3[56001] = 32'b00000000000000001111011100000000;
assign LUT_3[56002] = 32'b00000000000000001010111000000111;
assign LUT_3[56003] = 32'b00000000000000010001100011100100;
assign LUT_3[56004] = 32'b00000000000000000101111110011001;
assign LUT_3[56005] = 32'b00000000000000001100101001110110;
assign LUT_3[56006] = 32'b00000000000000001000000101111101;
assign LUT_3[56007] = 32'b00000000000000001110110001011010;
assign LUT_3[56008] = 32'b00000000000000001110001001101001;
assign LUT_3[56009] = 32'b00000000000000010100110101000110;
assign LUT_3[56010] = 32'b00000000000000010000010001001101;
assign LUT_3[56011] = 32'b00000000000000010110111100101010;
assign LUT_3[56012] = 32'b00000000000000001011010111011111;
assign LUT_3[56013] = 32'b00000000000000010010000010111100;
assign LUT_3[56014] = 32'b00000000000000001101011111000011;
assign LUT_3[56015] = 32'b00000000000000010100001010100000;
assign LUT_3[56016] = 32'b00000000000000001100000011100110;
assign LUT_3[56017] = 32'b00000000000000010010101111000011;
assign LUT_3[56018] = 32'b00000000000000001110001011001010;
assign LUT_3[56019] = 32'b00000000000000010100110110100111;
assign LUT_3[56020] = 32'b00000000000000001001010001011100;
assign LUT_3[56021] = 32'b00000000000000001111111100111001;
assign LUT_3[56022] = 32'b00000000000000001011011001000000;
assign LUT_3[56023] = 32'b00000000000000010010000100011101;
assign LUT_3[56024] = 32'b00000000000000010001011100101100;
assign LUT_3[56025] = 32'b00000000000000011000001000001001;
assign LUT_3[56026] = 32'b00000000000000010011100100010000;
assign LUT_3[56027] = 32'b00000000000000011010001111101101;
assign LUT_3[56028] = 32'b00000000000000001110101010100010;
assign LUT_3[56029] = 32'b00000000000000010101010101111111;
assign LUT_3[56030] = 32'b00000000000000010000110010000110;
assign LUT_3[56031] = 32'b00000000000000010111011101100011;
assign LUT_3[56032] = 32'b00000000000000001001111111000011;
assign LUT_3[56033] = 32'b00000000000000010000101010100000;
assign LUT_3[56034] = 32'b00000000000000001100000110100111;
assign LUT_3[56035] = 32'b00000000000000010010110010000100;
assign LUT_3[56036] = 32'b00000000000000000111001100111001;
assign LUT_3[56037] = 32'b00000000000000001101111000010110;
assign LUT_3[56038] = 32'b00000000000000001001010100011101;
assign LUT_3[56039] = 32'b00000000000000001111111111111010;
assign LUT_3[56040] = 32'b00000000000000001111011000001001;
assign LUT_3[56041] = 32'b00000000000000010110000011100110;
assign LUT_3[56042] = 32'b00000000000000010001011111101101;
assign LUT_3[56043] = 32'b00000000000000011000001011001010;
assign LUT_3[56044] = 32'b00000000000000001100100101111111;
assign LUT_3[56045] = 32'b00000000000000010011010001011100;
assign LUT_3[56046] = 32'b00000000000000001110101101100011;
assign LUT_3[56047] = 32'b00000000000000010101011001000000;
assign LUT_3[56048] = 32'b00000000000000001101010010000110;
assign LUT_3[56049] = 32'b00000000000000010011111101100011;
assign LUT_3[56050] = 32'b00000000000000001111011001101010;
assign LUT_3[56051] = 32'b00000000000000010110000101000111;
assign LUT_3[56052] = 32'b00000000000000001010011111111100;
assign LUT_3[56053] = 32'b00000000000000010001001011011001;
assign LUT_3[56054] = 32'b00000000000000001100100111100000;
assign LUT_3[56055] = 32'b00000000000000010011010010111101;
assign LUT_3[56056] = 32'b00000000000000010010101011001100;
assign LUT_3[56057] = 32'b00000000000000011001010110101001;
assign LUT_3[56058] = 32'b00000000000000010100110010110000;
assign LUT_3[56059] = 32'b00000000000000011011011110001101;
assign LUT_3[56060] = 32'b00000000000000001111111001000010;
assign LUT_3[56061] = 32'b00000000000000010110100100011111;
assign LUT_3[56062] = 32'b00000000000000010010000000100110;
assign LUT_3[56063] = 32'b00000000000000011000101100000011;
assign LUT_3[56064] = 32'b00000000000000000010111100011011;
assign LUT_3[56065] = 32'b00000000000000001001100111111000;
assign LUT_3[56066] = 32'b00000000000000000101000011111111;
assign LUT_3[56067] = 32'b00000000000000001011101111011100;
assign LUT_3[56068] = 32'b00000000000000000000001010010001;
assign LUT_3[56069] = 32'b00000000000000000110110101101110;
assign LUT_3[56070] = 32'b00000000000000000010010001110101;
assign LUT_3[56071] = 32'b00000000000000001000111101010010;
assign LUT_3[56072] = 32'b00000000000000001000010101100001;
assign LUT_3[56073] = 32'b00000000000000001111000000111110;
assign LUT_3[56074] = 32'b00000000000000001010011101000101;
assign LUT_3[56075] = 32'b00000000000000010001001000100010;
assign LUT_3[56076] = 32'b00000000000000000101100011010111;
assign LUT_3[56077] = 32'b00000000000000001100001110110100;
assign LUT_3[56078] = 32'b00000000000000000111101010111011;
assign LUT_3[56079] = 32'b00000000000000001110010110011000;
assign LUT_3[56080] = 32'b00000000000000000110001111011110;
assign LUT_3[56081] = 32'b00000000000000001100111010111011;
assign LUT_3[56082] = 32'b00000000000000001000010111000010;
assign LUT_3[56083] = 32'b00000000000000001111000010011111;
assign LUT_3[56084] = 32'b00000000000000000011011101010100;
assign LUT_3[56085] = 32'b00000000000000001010001000110001;
assign LUT_3[56086] = 32'b00000000000000000101100100111000;
assign LUT_3[56087] = 32'b00000000000000001100010000010101;
assign LUT_3[56088] = 32'b00000000000000001011101000100100;
assign LUT_3[56089] = 32'b00000000000000010010010100000001;
assign LUT_3[56090] = 32'b00000000000000001101110000001000;
assign LUT_3[56091] = 32'b00000000000000010100011011100101;
assign LUT_3[56092] = 32'b00000000000000001000110110011010;
assign LUT_3[56093] = 32'b00000000000000001111100001110111;
assign LUT_3[56094] = 32'b00000000000000001010111101111110;
assign LUT_3[56095] = 32'b00000000000000010001101001011011;
assign LUT_3[56096] = 32'b00000000000000000100001010111011;
assign LUT_3[56097] = 32'b00000000000000001010110110011000;
assign LUT_3[56098] = 32'b00000000000000000110010010011111;
assign LUT_3[56099] = 32'b00000000000000001100111101111100;
assign LUT_3[56100] = 32'b00000000000000000001011000110001;
assign LUT_3[56101] = 32'b00000000000000001000000100001110;
assign LUT_3[56102] = 32'b00000000000000000011100000010101;
assign LUT_3[56103] = 32'b00000000000000001010001011110010;
assign LUT_3[56104] = 32'b00000000000000001001100100000001;
assign LUT_3[56105] = 32'b00000000000000010000001111011110;
assign LUT_3[56106] = 32'b00000000000000001011101011100101;
assign LUT_3[56107] = 32'b00000000000000010010010111000010;
assign LUT_3[56108] = 32'b00000000000000000110110001110111;
assign LUT_3[56109] = 32'b00000000000000001101011101010100;
assign LUT_3[56110] = 32'b00000000000000001000111001011011;
assign LUT_3[56111] = 32'b00000000000000001111100100111000;
assign LUT_3[56112] = 32'b00000000000000000111011101111110;
assign LUT_3[56113] = 32'b00000000000000001110001001011011;
assign LUT_3[56114] = 32'b00000000000000001001100101100010;
assign LUT_3[56115] = 32'b00000000000000010000010000111111;
assign LUT_3[56116] = 32'b00000000000000000100101011110100;
assign LUT_3[56117] = 32'b00000000000000001011010111010001;
assign LUT_3[56118] = 32'b00000000000000000110110011011000;
assign LUT_3[56119] = 32'b00000000000000001101011110110101;
assign LUT_3[56120] = 32'b00000000000000001100110111000100;
assign LUT_3[56121] = 32'b00000000000000010011100010100001;
assign LUT_3[56122] = 32'b00000000000000001110111110101000;
assign LUT_3[56123] = 32'b00000000000000010101101010000101;
assign LUT_3[56124] = 32'b00000000000000001010000100111010;
assign LUT_3[56125] = 32'b00000000000000010000110000010111;
assign LUT_3[56126] = 32'b00000000000000001100001100011110;
assign LUT_3[56127] = 32'b00000000000000010010110111111011;
assign LUT_3[56128] = 32'b00000000000000000010110101000110;
assign LUT_3[56129] = 32'b00000000000000001001100000100011;
assign LUT_3[56130] = 32'b00000000000000000100111100101010;
assign LUT_3[56131] = 32'b00000000000000001011101000000111;
assign LUT_3[56132] = 32'b00000000000000000000000010111100;
assign LUT_3[56133] = 32'b00000000000000000110101110011001;
assign LUT_3[56134] = 32'b00000000000000000010001010100000;
assign LUT_3[56135] = 32'b00000000000000001000110101111101;
assign LUT_3[56136] = 32'b00000000000000001000001110001100;
assign LUT_3[56137] = 32'b00000000000000001110111001101001;
assign LUT_3[56138] = 32'b00000000000000001010010101110000;
assign LUT_3[56139] = 32'b00000000000000010001000001001101;
assign LUT_3[56140] = 32'b00000000000000000101011100000010;
assign LUT_3[56141] = 32'b00000000000000001100000111011111;
assign LUT_3[56142] = 32'b00000000000000000111100011100110;
assign LUT_3[56143] = 32'b00000000000000001110001111000011;
assign LUT_3[56144] = 32'b00000000000000000110001000001001;
assign LUT_3[56145] = 32'b00000000000000001100110011100110;
assign LUT_3[56146] = 32'b00000000000000001000001111101101;
assign LUT_3[56147] = 32'b00000000000000001110111011001010;
assign LUT_3[56148] = 32'b00000000000000000011010101111111;
assign LUT_3[56149] = 32'b00000000000000001010000001011100;
assign LUT_3[56150] = 32'b00000000000000000101011101100011;
assign LUT_3[56151] = 32'b00000000000000001100001001000000;
assign LUT_3[56152] = 32'b00000000000000001011100001001111;
assign LUT_3[56153] = 32'b00000000000000010010001100101100;
assign LUT_3[56154] = 32'b00000000000000001101101000110011;
assign LUT_3[56155] = 32'b00000000000000010100010100010000;
assign LUT_3[56156] = 32'b00000000000000001000101111000101;
assign LUT_3[56157] = 32'b00000000000000001111011010100010;
assign LUT_3[56158] = 32'b00000000000000001010110110101001;
assign LUT_3[56159] = 32'b00000000000000010001100010000110;
assign LUT_3[56160] = 32'b00000000000000000100000011100110;
assign LUT_3[56161] = 32'b00000000000000001010101111000011;
assign LUT_3[56162] = 32'b00000000000000000110001011001010;
assign LUT_3[56163] = 32'b00000000000000001100110110100111;
assign LUT_3[56164] = 32'b00000000000000000001010001011100;
assign LUT_3[56165] = 32'b00000000000000000111111100111001;
assign LUT_3[56166] = 32'b00000000000000000011011001000000;
assign LUT_3[56167] = 32'b00000000000000001010000100011101;
assign LUT_3[56168] = 32'b00000000000000001001011100101100;
assign LUT_3[56169] = 32'b00000000000000010000001000001001;
assign LUT_3[56170] = 32'b00000000000000001011100100010000;
assign LUT_3[56171] = 32'b00000000000000010010001111101101;
assign LUT_3[56172] = 32'b00000000000000000110101010100010;
assign LUT_3[56173] = 32'b00000000000000001101010101111111;
assign LUT_3[56174] = 32'b00000000000000001000110010000110;
assign LUT_3[56175] = 32'b00000000000000001111011101100011;
assign LUT_3[56176] = 32'b00000000000000000111010110101001;
assign LUT_3[56177] = 32'b00000000000000001110000010000110;
assign LUT_3[56178] = 32'b00000000000000001001011110001101;
assign LUT_3[56179] = 32'b00000000000000010000001001101010;
assign LUT_3[56180] = 32'b00000000000000000100100100011111;
assign LUT_3[56181] = 32'b00000000000000001011001111111100;
assign LUT_3[56182] = 32'b00000000000000000110101100000011;
assign LUT_3[56183] = 32'b00000000000000001101010111100000;
assign LUT_3[56184] = 32'b00000000000000001100101111101111;
assign LUT_3[56185] = 32'b00000000000000010011011011001100;
assign LUT_3[56186] = 32'b00000000000000001110110111010011;
assign LUT_3[56187] = 32'b00000000000000010101100010110000;
assign LUT_3[56188] = 32'b00000000000000001001111101100101;
assign LUT_3[56189] = 32'b00000000000000010000101001000010;
assign LUT_3[56190] = 32'b00000000000000001100000101001001;
assign LUT_3[56191] = 32'b00000000000000010010110000100110;
assign LUT_3[56192] = 32'b00000000000000000101000111011001;
assign LUT_3[56193] = 32'b00000000000000001011110010110110;
assign LUT_3[56194] = 32'b00000000000000000111001110111101;
assign LUT_3[56195] = 32'b00000000000000001101111010011010;
assign LUT_3[56196] = 32'b00000000000000000010010101001111;
assign LUT_3[56197] = 32'b00000000000000001001000000101100;
assign LUT_3[56198] = 32'b00000000000000000100011100110011;
assign LUT_3[56199] = 32'b00000000000000001011001000010000;
assign LUT_3[56200] = 32'b00000000000000001010100000011111;
assign LUT_3[56201] = 32'b00000000000000010001001011111100;
assign LUT_3[56202] = 32'b00000000000000001100101000000011;
assign LUT_3[56203] = 32'b00000000000000010011010011100000;
assign LUT_3[56204] = 32'b00000000000000000111101110010101;
assign LUT_3[56205] = 32'b00000000000000001110011001110010;
assign LUT_3[56206] = 32'b00000000000000001001110101111001;
assign LUT_3[56207] = 32'b00000000000000010000100001010110;
assign LUT_3[56208] = 32'b00000000000000001000011010011100;
assign LUT_3[56209] = 32'b00000000000000001111000101111001;
assign LUT_3[56210] = 32'b00000000000000001010100010000000;
assign LUT_3[56211] = 32'b00000000000000010001001101011101;
assign LUT_3[56212] = 32'b00000000000000000101101000010010;
assign LUT_3[56213] = 32'b00000000000000001100010011101111;
assign LUT_3[56214] = 32'b00000000000000000111101111110110;
assign LUT_3[56215] = 32'b00000000000000001110011011010011;
assign LUT_3[56216] = 32'b00000000000000001101110011100010;
assign LUT_3[56217] = 32'b00000000000000010100011110111111;
assign LUT_3[56218] = 32'b00000000000000001111111011000110;
assign LUT_3[56219] = 32'b00000000000000010110100110100011;
assign LUT_3[56220] = 32'b00000000000000001011000001011000;
assign LUT_3[56221] = 32'b00000000000000010001101100110101;
assign LUT_3[56222] = 32'b00000000000000001101001000111100;
assign LUT_3[56223] = 32'b00000000000000010011110100011001;
assign LUT_3[56224] = 32'b00000000000000000110010101111001;
assign LUT_3[56225] = 32'b00000000000000001101000001010110;
assign LUT_3[56226] = 32'b00000000000000001000011101011101;
assign LUT_3[56227] = 32'b00000000000000001111001000111010;
assign LUT_3[56228] = 32'b00000000000000000011100011101111;
assign LUT_3[56229] = 32'b00000000000000001010001111001100;
assign LUT_3[56230] = 32'b00000000000000000101101011010011;
assign LUT_3[56231] = 32'b00000000000000001100010110110000;
assign LUT_3[56232] = 32'b00000000000000001011101110111111;
assign LUT_3[56233] = 32'b00000000000000010010011010011100;
assign LUT_3[56234] = 32'b00000000000000001101110110100011;
assign LUT_3[56235] = 32'b00000000000000010100100010000000;
assign LUT_3[56236] = 32'b00000000000000001000111100110101;
assign LUT_3[56237] = 32'b00000000000000001111101000010010;
assign LUT_3[56238] = 32'b00000000000000001011000100011001;
assign LUT_3[56239] = 32'b00000000000000010001101111110110;
assign LUT_3[56240] = 32'b00000000000000001001101000111100;
assign LUT_3[56241] = 32'b00000000000000010000010100011001;
assign LUT_3[56242] = 32'b00000000000000001011110000100000;
assign LUT_3[56243] = 32'b00000000000000010010011011111101;
assign LUT_3[56244] = 32'b00000000000000000110110110110010;
assign LUT_3[56245] = 32'b00000000000000001101100010001111;
assign LUT_3[56246] = 32'b00000000000000001000111110010110;
assign LUT_3[56247] = 32'b00000000000000001111101001110011;
assign LUT_3[56248] = 32'b00000000000000001111000010000010;
assign LUT_3[56249] = 32'b00000000000000010101101101011111;
assign LUT_3[56250] = 32'b00000000000000010001001001100110;
assign LUT_3[56251] = 32'b00000000000000010111110101000011;
assign LUT_3[56252] = 32'b00000000000000001100001111111000;
assign LUT_3[56253] = 32'b00000000000000010010111011010101;
assign LUT_3[56254] = 32'b00000000000000001110010111011100;
assign LUT_3[56255] = 32'b00000000000000010101000010111001;
assign LUT_3[56256] = 32'b00000000000000000101000000000100;
assign LUT_3[56257] = 32'b00000000000000001011101011100001;
assign LUT_3[56258] = 32'b00000000000000000111000111101000;
assign LUT_3[56259] = 32'b00000000000000001101110011000101;
assign LUT_3[56260] = 32'b00000000000000000010001101111010;
assign LUT_3[56261] = 32'b00000000000000001000111001010111;
assign LUT_3[56262] = 32'b00000000000000000100010101011110;
assign LUT_3[56263] = 32'b00000000000000001011000000111011;
assign LUT_3[56264] = 32'b00000000000000001010011001001010;
assign LUT_3[56265] = 32'b00000000000000010001000100100111;
assign LUT_3[56266] = 32'b00000000000000001100100000101110;
assign LUT_3[56267] = 32'b00000000000000010011001100001011;
assign LUT_3[56268] = 32'b00000000000000000111100111000000;
assign LUT_3[56269] = 32'b00000000000000001110010010011101;
assign LUT_3[56270] = 32'b00000000000000001001101110100100;
assign LUT_3[56271] = 32'b00000000000000010000011010000001;
assign LUT_3[56272] = 32'b00000000000000001000010011000111;
assign LUT_3[56273] = 32'b00000000000000001110111110100100;
assign LUT_3[56274] = 32'b00000000000000001010011010101011;
assign LUT_3[56275] = 32'b00000000000000010001000110001000;
assign LUT_3[56276] = 32'b00000000000000000101100000111101;
assign LUT_3[56277] = 32'b00000000000000001100001100011010;
assign LUT_3[56278] = 32'b00000000000000000111101000100001;
assign LUT_3[56279] = 32'b00000000000000001110010011111110;
assign LUT_3[56280] = 32'b00000000000000001101101100001101;
assign LUT_3[56281] = 32'b00000000000000010100010111101010;
assign LUT_3[56282] = 32'b00000000000000001111110011110001;
assign LUT_3[56283] = 32'b00000000000000010110011111001110;
assign LUT_3[56284] = 32'b00000000000000001010111010000011;
assign LUT_3[56285] = 32'b00000000000000010001100101100000;
assign LUT_3[56286] = 32'b00000000000000001101000001100111;
assign LUT_3[56287] = 32'b00000000000000010011101101000100;
assign LUT_3[56288] = 32'b00000000000000000110001110100100;
assign LUT_3[56289] = 32'b00000000000000001100111010000001;
assign LUT_3[56290] = 32'b00000000000000001000010110001000;
assign LUT_3[56291] = 32'b00000000000000001111000001100101;
assign LUT_3[56292] = 32'b00000000000000000011011100011010;
assign LUT_3[56293] = 32'b00000000000000001010000111110111;
assign LUT_3[56294] = 32'b00000000000000000101100011111110;
assign LUT_3[56295] = 32'b00000000000000001100001111011011;
assign LUT_3[56296] = 32'b00000000000000001011100111101010;
assign LUT_3[56297] = 32'b00000000000000010010010011000111;
assign LUT_3[56298] = 32'b00000000000000001101101111001110;
assign LUT_3[56299] = 32'b00000000000000010100011010101011;
assign LUT_3[56300] = 32'b00000000000000001000110101100000;
assign LUT_3[56301] = 32'b00000000000000001111100000111101;
assign LUT_3[56302] = 32'b00000000000000001010111101000100;
assign LUT_3[56303] = 32'b00000000000000010001101000100001;
assign LUT_3[56304] = 32'b00000000000000001001100001100111;
assign LUT_3[56305] = 32'b00000000000000010000001101000100;
assign LUT_3[56306] = 32'b00000000000000001011101001001011;
assign LUT_3[56307] = 32'b00000000000000010010010100101000;
assign LUT_3[56308] = 32'b00000000000000000110101111011101;
assign LUT_3[56309] = 32'b00000000000000001101011010111010;
assign LUT_3[56310] = 32'b00000000000000001000110111000001;
assign LUT_3[56311] = 32'b00000000000000001111100010011110;
assign LUT_3[56312] = 32'b00000000000000001110111010101101;
assign LUT_3[56313] = 32'b00000000000000010101100110001010;
assign LUT_3[56314] = 32'b00000000000000010001000010010001;
assign LUT_3[56315] = 32'b00000000000000010111101101101110;
assign LUT_3[56316] = 32'b00000000000000001100001000100011;
assign LUT_3[56317] = 32'b00000000000000010010110100000000;
assign LUT_3[56318] = 32'b00000000000000001110010000000111;
assign LUT_3[56319] = 32'b00000000000000010100111011100100;
assign LUT_3[56320] = 32'b00000000000000001001111100101011;
assign LUT_3[56321] = 32'b00000000000000010000101000001000;
assign LUT_3[56322] = 32'b00000000000000001100000100001111;
assign LUT_3[56323] = 32'b00000000000000010010101111101100;
assign LUT_3[56324] = 32'b00000000000000000111001010100001;
assign LUT_3[56325] = 32'b00000000000000001101110101111110;
assign LUT_3[56326] = 32'b00000000000000001001010010000101;
assign LUT_3[56327] = 32'b00000000000000001111111101100010;
assign LUT_3[56328] = 32'b00000000000000001111010101110001;
assign LUT_3[56329] = 32'b00000000000000010110000001001110;
assign LUT_3[56330] = 32'b00000000000000010001011101010101;
assign LUT_3[56331] = 32'b00000000000000011000001000110010;
assign LUT_3[56332] = 32'b00000000000000001100100011100111;
assign LUT_3[56333] = 32'b00000000000000010011001111000100;
assign LUT_3[56334] = 32'b00000000000000001110101011001011;
assign LUT_3[56335] = 32'b00000000000000010101010110101000;
assign LUT_3[56336] = 32'b00000000000000001101001111101110;
assign LUT_3[56337] = 32'b00000000000000010011111011001011;
assign LUT_3[56338] = 32'b00000000000000001111010111010010;
assign LUT_3[56339] = 32'b00000000000000010110000010101111;
assign LUT_3[56340] = 32'b00000000000000001010011101100100;
assign LUT_3[56341] = 32'b00000000000000010001001001000001;
assign LUT_3[56342] = 32'b00000000000000001100100101001000;
assign LUT_3[56343] = 32'b00000000000000010011010000100101;
assign LUT_3[56344] = 32'b00000000000000010010101000110100;
assign LUT_3[56345] = 32'b00000000000000011001010100010001;
assign LUT_3[56346] = 32'b00000000000000010100110000011000;
assign LUT_3[56347] = 32'b00000000000000011011011011110101;
assign LUT_3[56348] = 32'b00000000000000001111110110101010;
assign LUT_3[56349] = 32'b00000000000000010110100010000111;
assign LUT_3[56350] = 32'b00000000000000010001111110001110;
assign LUT_3[56351] = 32'b00000000000000011000101001101011;
assign LUT_3[56352] = 32'b00000000000000001011001011001011;
assign LUT_3[56353] = 32'b00000000000000010001110110101000;
assign LUT_3[56354] = 32'b00000000000000001101010010101111;
assign LUT_3[56355] = 32'b00000000000000010011111110001100;
assign LUT_3[56356] = 32'b00000000000000001000011001000001;
assign LUT_3[56357] = 32'b00000000000000001111000100011110;
assign LUT_3[56358] = 32'b00000000000000001010100000100101;
assign LUT_3[56359] = 32'b00000000000000010001001100000010;
assign LUT_3[56360] = 32'b00000000000000010000100100010001;
assign LUT_3[56361] = 32'b00000000000000010111001111101110;
assign LUT_3[56362] = 32'b00000000000000010010101011110101;
assign LUT_3[56363] = 32'b00000000000000011001010111010010;
assign LUT_3[56364] = 32'b00000000000000001101110010000111;
assign LUT_3[56365] = 32'b00000000000000010100011101100100;
assign LUT_3[56366] = 32'b00000000000000001111111001101011;
assign LUT_3[56367] = 32'b00000000000000010110100101001000;
assign LUT_3[56368] = 32'b00000000000000001110011110001110;
assign LUT_3[56369] = 32'b00000000000000010101001001101011;
assign LUT_3[56370] = 32'b00000000000000010000100101110010;
assign LUT_3[56371] = 32'b00000000000000010111010001001111;
assign LUT_3[56372] = 32'b00000000000000001011101100000100;
assign LUT_3[56373] = 32'b00000000000000010010010111100001;
assign LUT_3[56374] = 32'b00000000000000001101110011101000;
assign LUT_3[56375] = 32'b00000000000000010100011111000101;
assign LUT_3[56376] = 32'b00000000000000010011110111010100;
assign LUT_3[56377] = 32'b00000000000000011010100010110001;
assign LUT_3[56378] = 32'b00000000000000010101111110111000;
assign LUT_3[56379] = 32'b00000000000000011100101010010101;
assign LUT_3[56380] = 32'b00000000000000010001000101001010;
assign LUT_3[56381] = 32'b00000000000000010111110000100111;
assign LUT_3[56382] = 32'b00000000000000010011001100101110;
assign LUT_3[56383] = 32'b00000000000000011001111000001011;
assign LUT_3[56384] = 32'b00000000000000001001110101010110;
assign LUT_3[56385] = 32'b00000000000000010000100000110011;
assign LUT_3[56386] = 32'b00000000000000001011111100111010;
assign LUT_3[56387] = 32'b00000000000000010010101000010111;
assign LUT_3[56388] = 32'b00000000000000000111000011001100;
assign LUT_3[56389] = 32'b00000000000000001101101110101001;
assign LUT_3[56390] = 32'b00000000000000001001001010110000;
assign LUT_3[56391] = 32'b00000000000000001111110110001101;
assign LUT_3[56392] = 32'b00000000000000001111001110011100;
assign LUT_3[56393] = 32'b00000000000000010101111001111001;
assign LUT_3[56394] = 32'b00000000000000010001010110000000;
assign LUT_3[56395] = 32'b00000000000000011000000001011101;
assign LUT_3[56396] = 32'b00000000000000001100011100010010;
assign LUT_3[56397] = 32'b00000000000000010011000111101111;
assign LUT_3[56398] = 32'b00000000000000001110100011110110;
assign LUT_3[56399] = 32'b00000000000000010101001111010011;
assign LUT_3[56400] = 32'b00000000000000001101001000011001;
assign LUT_3[56401] = 32'b00000000000000010011110011110110;
assign LUT_3[56402] = 32'b00000000000000001111001111111101;
assign LUT_3[56403] = 32'b00000000000000010101111011011010;
assign LUT_3[56404] = 32'b00000000000000001010010110001111;
assign LUT_3[56405] = 32'b00000000000000010001000001101100;
assign LUT_3[56406] = 32'b00000000000000001100011101110011;
assign LUT_3[56407] = 32'b00000000000000010011001001010000;
assign LUT_3[56408] = 32'b00000000000000010010100001011111;
assign LUT_3[56409] = 32'b00000000000000011001001100111100;
assign LUT_3[56410] = 32'b00000000000000010100101001000011;
assign LUT_3[56411] = 32'b00000000000000011011010100100000;
assign LUT_3[56412] = 32'b00000000000000001111101111010101;
assign LUT_3[56413] = 32'b00000000000000010110011010110010;
assign LUT_3[56414] = 32'b00000000000000010001110110111001;
assign LUT_3[56415] = 32'b00000000000000011000100010010110;
assign LUT_3[56416] = 32'b00000000000000001011000011110110;
assign LUT_3[56417] = 32'b00000000000000010001101111010011;
assign LUT_3[56418] = 32'b00000000000000001101001011011010;
assign LUT_3[56419] = 32'b00000000000000010011110110110111;
assign LUT_3[56420] = 32'b00000000000000001000010001101100;
assign LUT_3[56421] = 32'b00000000000000001110111101001001;
assign LUT_3[56422] = 32'b00000000000000001010011001010000;
assign LUT_3[56423] = 32'b00000000000000010001000100101101;
assign LUT_3[56424] = 32'b00000000000000010000011100111100;
assign LUT_3[56425] = 32'b00000000000000010111001000011001;
assign LUT_3[56426] = 32'b00000000000000010010100100100000;
assign LUT_3[56427] = 32'b00000000000000011001001111111101;
assign LUT_3[56428] = 32'b00000000000000001101101010110010;
assign LUT_3[56429] = 32'b00000000000000010100010110001111;
assign LUT_3[56430] = 32'b00000000000000001111110010010110;
assign LUT_3[56431] = 32'b00000000000000010110011101110011;
assign LUT_3[56432] = 32'b00000000000000001110010110111001;
assign LUT_3[56433] = 32'b00000000000000010101000010010110;
assign LUT_3[56434] = 32'b00000000000000010000011110011101;
assign LUT_3[56435] = 32'b00000000000000010111001001111010;
assign LUT_3[56436] = 32'b00000000000000001011100100101111;
assign LUT_3[56437] = 32'b00000000000000010010010000001100;
assign LUT_3[56438] = 32'b00000000000000001101101100010011;
assign LUT_3[56439] = 32'b00000000000000010100010111110000;
assign LUT_3[56440] = 32'b00000000000000010011101111111111;
assign LUT_3[56441] = 32'b00000000000000011010011011011100;
assign LUT_3[56442] = 32'b00000000000000010101110111100011;
assign LUT_3[56443] = 32'b00000000000000011100100011000000;
assign LUT_3[56444] = 32'b00000000000000010000111101110101;
assign LUT_3[56445] = 32'b00000000000000010111101001010010;
assign LUT_3[56446] = 32'b00000000000000010011000101011001;
assign LUT_3[56447] = 32'b00000000000000011001110000110110;
assign LUT_3[56448] = 32'b00000000000000001100000111101001;
assign LUT_3[56449] = 32'b00000000000000010010110011000110;
assign LUT_3[56450] = 32'b00000000000000001110001111001101;
assign LUT_3[56451] = 32'b00000000000000010100111010101010;
assign LUT_3[56452] = 32'b00000000000000001001010101011111;
assign LUT_3[56453] = 32'b00000000000000010000000000111100;
assign LUT_3[56454] = 32'b00000000000000001011011101000011;
assign LUT_3[56455] = 32'b00000000000000010010001000100000;
assign LUT_3[56456] = 32'b00000000000000010001100000101111;
assign LUT_3[56457] = 32'b00000000000000011000001100001100;
assign LUT_3[56458] = 32'b00000000000000010011101000010011;
assign LUT_3[56459] = 32'b00000000000000011010010011110000;
assign LUT_3[56460] = 32'b00000000000000001110101110100101;
assign LUT_3[56461] = 32'b00000000000000010101011010000010;
assign LUT_3[56462] = 32'b00000000000000010000110110001001;
assign LUT_3[56463] = 32'b00000000000000010111100001100110;
assign LUT_3[56464] = 32'b00000000000000001111011010101100;
assign LUT_3[56465] = 32'b00000000000000010110000110001001;
assign LUT_3[56466] = 32'b00000000000000010001100010010000;
assign LUT_3[56467] = 32'b00000000000000011000001101101101;
assign LUT_3[56468] = 32'b00000000000000001100101000100010;
assign LUT_3[56469] = 32'b00000000000000010011010011111111;
assign LUT_3[56470] = 32'b00000000000000001110110000000110;
assign LUT_3[56471] = 32'b00000000000000010101011011100011;
assign LUT_3[56472] = 32'b00000000000000010100110011110010;
assign LUT_3[56473] = 32'b00000000000000011011011111001111;
assign LUT_3[56474] = 32'b00000000000000010110111011010110;
assign LUT_3[56475] = 32'b00000000000000011101100110110011;
assign LUT_3[56476] = 32'b00000000000000010010000001101000;
assign LUT_3[56477] = 32'b00000000000000011000101101000101;
assign LUT_3[56478] = 32'b00000000000000010100001001001100;
assign LUT_3[56479] = 32'b00000000000000011010110100101001;
assign LUT_3[56480] = 32'b00000000000000001101010110001001;
assign LUT_3[56481] = 32'b00000000000000010100000001100110;
assign LUT_3[56482] = 32'b00000000000000001111011101101101;
assign LUT_3[56483] = 32'b00000000000000010110001001001010;
assign LUT_3[56484] = 32'b00000000000000001010100011111111;
assign LUT_3[56485] = 32'b00000000000000010001001111011100;
assign LUT_3[56486] = 32'b00000000000000001100101011100011;
assign LUT_3[56487] = 32'b00000000000000010011010111000000;
assign LUT_3[56488] = 32'b00000000000000010010101111001111;
assign LUT_3[56489] = 32'b00000000000000011001011010101100;
assign LUT_3[56490] = 32'b00000000000000010100110110110011;
assign LUT_3[56491] = 32'b00000000000000011011100010010000;
assign LUT_3[56492] = 32'b00000000000000001111111101000101;
assign LUT_3[56493] = 32'b00000000000000010110101000100010;
assign LUT_3[56494] = 32'b00000000000000010010000100101001;
assign LUT_3[56495] = 32'b00000000000000011000110000000110;
assign LUT_3[56496] = 32'b00000000000000010000101001001100;
assign LUT_3[56497] = 32'b00000000000000010111010100101001;
assign LUT_3[56498] = 32'b00000000000000010010110000110000;
assign LUT_3[56499] = 32'b00000000000000011001011100001101;
assign LUT_3[56500] = 32'b00000000000000001101110111000010;
assign LUT_3[56501] = 32'b00000000000000010100100010011111;
assign LUT_3[56502] = 32'b00000000000000001111111110100110;
assign LUT_3[56503] = 32'b00000000000000010110101010000011;
assign LUT_3[56504] = 32'b00000000000000010110000010010010;
assign LUT_3[56505] = 32'b00000000000000011100101101101111;
assign LUT_3[56506] = 32'b00000000000000011000001001110110;
assign LUT_3[56507] = 32'b00000000000000011110110101010011;
assign LUT_3[56508] = 32'b00000000000000010011010000001000;
assign LUT_3[56509] = 32'b00000000000000011001111011100101;
assign LUT_3[56510] = 32'b00000000000000010101010111101100;
assign LUT_3[56511] = 32'b00000000000000011100000011001001;
assign LUT_3[56512] = 32'b00000000000000001100000000010100;
assign LUT_3[56513] = 32'b00000000000000010010101011110001;
assign LUT_3[56514] = 32'b00000000000000001110000111111000;
assign LUT_3[56515] = 32'b00000000000000010100110011010101;
assign LUT_3[56516] = 32'b00000000000000001001001110001010;
assign LUT_3[56517] = 32'b00000000000000001111111001100111;
assign LUT_3[56518] = 32'b00000000000000001011010101101110;
assign LUT_3[56519] = 32'b00000000000000010010000001001011;
assign LUT_3[56520] = 32'b00000000000000010001011001011010;
assign LUT_3[56521] = 32'b00000000000000011000000100110111;
assign LUT_3[56522] = 32'b00000000000000010011100000111110;
assign LUT_3[56523] = 32'b00000000000000011010001100011011;
assign LUT_3[56524] = 32'b00000000000000001110100111010000;
assign LUT_3[56525] = 32'b00000000000000010101010010101101;
assign LUT_3[56526] = 32'b00000000000000010000101110110100;
assign LUT_3[56527] = 32'b00000000000000010111011010010001;
assign LUT_3[56528] = 32'b00000000000000001111010011010111;
assign LUT_3[56529] = 32'b00000000000000010101111110110100;
assign LUT_3[56530] = 32'b00000000000000010001011010111011;
assign LUT_3[56531] = 32'b00000000000000011000000110011000;
assign LUT_3[56532] = 32'b00000000000000001100100001001101;
assign LUT_3[56533] = 32'b00000000000000010011001100101010;
assign LUT_3[56534] = 32'b00000000000000001110101000110001;
assign LUT_3[56535] = 32'b00000000000000010101010100001110;
assign LUT_3[56536] = 32'b00000000000000010100101100011101;
assign LUT_3[56537] = 32'b00000000000000011011010111111010;
assign LUT_3[56538] = 32'b00000000000000010110110100000001;
assign LUT_3[56539] = 32'b00000000000000011101011111011110;
assign LUT_3[56540] = 32'b00000000000000010001111010010011;
assign LUT_3[56541] = 32'b00000000000000011000100101110000;
assign LUT_3[56542] = 32'b00000000000000010100000001110111;
assign LUT_3[56543] = 32'b00000000000000011010101101010100;
assign LUT_3[56544] = 32'b00000000000000001101001110110100;
assign LUT_3[56545] = 32'b00000000000000010011111010010001;
assign LUT_3[56546] = 32'b00000000000000001111010110011000;
assign LUT_3[56547] = 32'b00000000000000010110000001110101;
assign LUT_3[56548] = 32'b00000000000000001010011100101010;
assign LUT_3[56549] = 32'b00000000000000010001001000000111;
assign LUT_3[56550] = 32'b00000000000000001100100100001110;
assign LUT_3[56551] = 32'b00000000000000010011001111101011;
assign LUT_3[56552] = 32'b00000000000000010010100111111010;
assign LUT_3[56553] = 32'b00000000000000011001010011010111;
assign LUT_3[56554] = 32'b00000000000000010100101111011110;
assign LUT_3[56555] = 32'b00000000000000011011011010111011;
assign LUT_3[56556] = 32'b00000000000000001111110101110000;
assign LUT_3[56557] = 32'b00000000000000010110100001001101;
assign LUT_3[56558] = 32'b00000000000000010001111101010100;
assign LUT_3[56559] = 32'b00000000000000011000101000110001;
assign LUT_3[56560] = 32'b00000000000000010000100001110111;
assign LUT_3[56561] = 32'b00000000000000010111001101010100;
assign LUT_3[56562] = 32'b00000000000000010010101001011011;
assign LUT_3[56563] = 32'b00000000000000011001010100111000;
assign LUT_3[56564] = 32'b00000000000000001101101111101101;
assign LUT_3[56565] = 32'b00000000000000010100011011001010;
assign LUT_3[56566] = 32'b00000000000000001111110111010001;
assign LUT_3[56567] = 32'b00000000000000010110100010101110;
assign LUT_3[56568] = 32'b00000000000000010101111010111101;
assign LUT_3[56569] = 32'b00000000000000011100100110011010;
assign LUT_3[56570] = 32'b00000000000000011000000010100001;
assign LUT_3[56571] = 32'b00000000000000011110101101111110;
assign LUT_3[56572] = 32'b00000000000000010011001000110011;
assign LUT_3[56573] = 32'b00000000000000011001110100010000;
assign LUT_3[56574] = 32'b00000000000000010101010000010111;
assign LUT_3[56575] = 32'b00000000000000011011111011110100;
assign LUT_3[56576] = 32'b00000000000000000110001100001100;
assign LUT_3[56577] = 32'b00000000000000001100110111101001;
assign LUT_3[56578] = 32'b00000000000000001000010011110000;
assign LUT_3[56579] = 32'b00000000000000001110111111001101;
assign LUT_3[56580] = 32'b00000000000000000011011010000010;
assign LUT_3[56581] = 32'b00000000000000001010000101011111;
assign LUT_3[56582] = 32'b00000000000000000101100001100110;
assign LUT_3[56583] = 32'b00000000000000001100001101000011;
assign LUT_3[56584] = 32'b00000000000000001011100101010010;
assign LUT_3[56585] = 32'b00000000000000010010010000101111;
assign LUT_3[56586] = 32'b00000000000000001101101100110110;
assign LUT_3[56587] = 32'b00000000000000010100011000010011;
assign LUT_3[56588] = 32'b00000000000000001000110011001000;
assign LUT_3[56589] = 32'b00000000000000001111011110100101;
assign LUT_3[56590] = 32'b00000000000000001010111010101100;
assign LUT_3[56591] = 32'b00000000000000010001100110001001;
assign LUT_3[56592] = 32'b00000000000000001001011111001111;
assign LUT_3[56593] = 32'b00000000000000010000001010101100;
assign LUT_3[56594] = 32'b00000000000000001011100110110011;
assign LUT_3[56595] = 32'b00000000000000010010010010010000;
assign LUT_3[56596] = 32'b00000000000000000110101101000101;
assign LUT_3[56597] = 32'b00000000000000001101011000100010;
assign LUT_3[56598] = 32'b00000000000000001000110100101001;
assign LUT_3[56599] = 32'b00000000000000001111100000000110;
assign LUT_3[56600] = 32'b00000000000000001110111000010101;
assign LUT_3[56601] = 32'b00000000000000010101100011110010;
assign LUT_3[56602] = 32'b00000000000000010000111111111001;
assign LUT_3[56603] = 32'b00000000000000010111101011010110;
assign LUT_3[56604] = 32'b00000000000000001100000110001011;
assign LUT_3[56605] = 32'b00000000000000010010110001101000;
assign LUT_3[56606] = 32'b00000000000000001110001101101111;
assign LUT_3[56607] = 32'b00000000000000010100111001001100;
assign LUT_3[56608] = 32'b00000000000000000111011010101100;
assign LUT_3[56609] = 32'b00000000000000001110000110001001;
assign LUT_3[56610] = 32'b00000000000000001001100010010000;
assign LUT_3[56611] = 32'b00000000000000010000001101101101;
assign LUT_3[56612] = 32'b00000000000000000100101000100010;
assign LUT_3[56613] = 32'b00000000000000001011010011111111;
assign LUT_3[56614] = 32'b00000000000000000110110000000110;
assign LUT_3[56615] = 32'b00000000000000001101011011100011;
assign LUT_3[56616] = 32'b00000000000000001100110011110010;
assign LUT_3[56617] = 32'b00000000000000010011011111001111;
assign LUT_3[56618] = 32'b00000000000000001110111011010110;
assign LUT_3[56619] = 32'b00000000000000010101100110110011;
assign LUT_3[56620] = 32'b00000000000000001010000001101000;
assign LUT_3[56621] = 32'b00000000000000010000101101000101;
assign LUT_3[56622] = 32'b00000000000000001100001001001100;
assign LUT_3[56623] = 32'b00000000000000010010110100101001;
assign LUT_3[56624] = 32'b00000000000000001010101101101111;
assign LUT_3[56625] = 32'b00000000000000010001011001001100;
assign LUT_3[56626] = 32'b00000000000000001100110101010011;
assign LUT_3[56627] = 32'b00000000000000010011100000110000;
assign LUT_3[56628] = 32'b00000000000000000111111011100101;
assign LUT_3[56629] = 32'b00000000000000001110100111000010;
assign LUT_3[56630] = 32'b00000000000000001010000011001001;
assign LUT_3[56631] = 32'b00000000000000010000101110100110;
assign LUT_3[56632] = 32'b00000000000000010000000110110101;
assign LUT_3[56633] = 32'b00000000000000010110110010010010;
assign LUT_3[56634] = 32'b00000000000000010010001110011001;
assign LUT_3[56635] = 32'b00000000000000011000111001110110;
assign LUT_3[56636] = 32'b00000000000000001101010100101011;
assign LUT_3[56637] = 32'b00000000000000010100000000001000;
assign LUT_3[56638] = 32'b00000000000000001111011100001111;
assign LUT_3[56639] = 32'b00000000000000010110000111101100;
assign LUT_3[56640] = 32'b00000000000000000110000100110111;
assign LUT_3[56641] = 32'b00000000000000001100110000010100;
assign LUT_3[56642] = 32'b00000000000000001000001100011011;
assign LUT_3[56643] = 32'b00000000000000001110110111111000;
assign LUT_3[56644] = 32'b00000000000000000011010010101101;
assign LUT_3[56645] = 32'b00000000000000001001111110001010;
assign LUT_3[56646] = 32'b00000000000000000101011010010001;
assign LUT_3[56647] = 32'b00000000000000001100000101101110;
assign LUT_3[56648] = 32'b00000000000000001011011101111101;
assign LUT_3[56649] = 32'b00000000000000010010001001011010;
assign LUT_3[56650] = 32'b00000000000000001101100101100001;
assign LUT_3[56651] = 32'b00000000000000010100010000111110;
assign LUT_3[56652] = 32'b00000000000000001000101011110011;
assign LUT_3[56653] = 32'b00000000000000001111010111010000;
assign LUT_3[56654] = 32'b00000000000000001010110011010111;
assign LUT_3[56655] = 32'b00000000000000010001011110110100;
assign LUT_3[56656] = 32'b00000000000000001001010111111010;
assign LUT_3[56657] = 32'b00000000000000010000000011010111;
assign LUT_3[56658] = 32'b00000000000000001011011111011110;
assign LUT_3[56659] = 32'b00000000000000010010001010111011;
assign LUT_3[56660] = 32'b00000000000000000110100101110000;
assign LUT_3[56661] = 32'b00000000000000001101010001001101;
assign LUT_3[56662] = 32'b00000000000000001000101101010100;
assign LUT_3[56663] = 32'b00000000000000001111011000110001;
assign LUT_3[56664] = 32'b00000000000000001110110001000000;
assign LUT_3[56665] = 32'b00000000000000010101011100011101;
assign LUT_3[56666] = 32'b00000000000000010000111000100100;
assign LUT_3[56667] = 32'b00000000000000010111100100000001;
assign LUT_3[56668] = 32'b00000000000000001011111110110110;
assign LUT_3[56669] = 32'b00000000000000010010101010010011;
assign LUT_3[56670] = 32'b00000000000000001110000110011010;
assign LUT_3[56671] = 32'b00000000000000010100110001110111;
assign LUT_3[56672] = 32'b00000000000000000111010011010111;
assign LUT_3[56673] = 32'b00000000000000001101111110110100;
assign LUT_3[56674] = 32'b00000000000000001001011010111011;
assign LUT_3[56675] = 32'b00000000000000010000000110011000;
assign LUT_3[56676] = 32'b00000000000000000100100001001101;
assign LUT_3[56677] = 32'b00000000000000001011001100101010;
assign LUT_3[56678] = 32'b00000000000000000110101000110001;
assign LUT_3[56679] = 32'b00000000000000001101010100001110;
assign LUT_3[56680] = 32'b00000000000000001100101100011101;
assign LUT_3[56681] = 32'b00000000000000010011010111111010;
assign LUT_3[56682] = 32'b00000000000000001110110100000001;
assign LUT_3[56683] = 32'b00000000000000010101011111011110;
assign LUT_3[56684] = 32'b00000000000000001001111010010011;
assign LUT_3[56685] = 32'b00000000000000010000100101110000;
assign LUT_3[56686] = 32'b00000000000000001100000001110111;
assign LUT_3[56687] = 32'b00000000000000010010101101010100;
assign LUT_3[56688] = 32'b00000000000000001010100110011010;
assign LUT_3[56689] = 32'b00000000000000010001010001110111;
assign LUT_3[56690] = 32'b00000000000000001100101101111110;
assign LUT_3[56691] = 32'b00000000000000010011011001011011;
assign LUT_3[56692] = 32'b00000000000000000111110100010000;
assign LUT_3[56693] = 32'b00000000000000001110011111101101;
assign LUT_3[56694] = 32'b00000000000000001001111011110100;
assign LUT_3[56695] = 32'b00000000000000010000100111010001;
assign LUT_3[56696] = 32'b00000000000000001111111111100000;
assign LUT_3[56697] = 32'b00000000000000010110101010111101;
assign LUT_3[56698] = 32'b00000000000000010010000111000100;
assign LUT_3[56699] = 32'b00000000000000011000110010100001;
assign LUT_3[56700] = 32'b00000000000000001101001101010110;
assign LUT_3[56701] = 32'b00000000000000010011111000110011;
assign LUT_3[56702] = 32'b00000000000000001111010100111010;
assign LUT_3[56703] = 32'b00000000000000010110000000010111;
assign LUT_3[56704] = 32'b00000000000000001000010111001010;
assign LUT_3[56705] = 32'b00000000000000001111000010100111;
assign LUT_3[56706] = 32'b00000000000000001010011110101110;
assign LUT_3[56707] = 32'b00000000000000010001001010001011;
assign LUT_3[56708] = 32'b00000000000000000101100101000000;
assign LUT_3[56709] = 32'b00000000000000001100010000011101;
assign LUT_3[56710] = 32'b00000000000000000111101100100100;
assign LUT_3[56711] = 32'b00000000000000001110011000000001;
assign LUT_3[56712] = 32'b00000000000000001101110000010000;
assign LUT_3[56713] = 32'b00000000000000010100011011101101;
assign LUT_3[56714] = 32'b00000000000000001111110111110100;
assign LUT_3[56715] = 32'b00000000000000010110100011010001;
assign LUT_3[56716] = 32'b00000000000000001010111110000110;
assign LUT_3[56717] = 32'b00000000000000010001101001100011;
assign LUT_3[56718] = 32'b00000000000000001101000101101010;
assign LUT_3[56719] = 32'b00000000000000010011110001000111;
assign LUT_3[56720] = 32'b00000000000000001011101010001101;
assign LUT_3[56721] = 32'b00000000000000010010010101101010;
assign LUT_3[56722] = 32'b00000000000000001101110001110001;
assign LUT_3[56723] = 32'b00000000000000010100011101001110;
assign LUT_3[56724] = 32'b00000000000000001000111000000011;
assign LUT_3[56725] = 32'b00000000000000001111100011100000;
assign LUT_3[56726] = 32'b00000000000000001010111111100111;
assign LUT_3[56727] = 32'b00000000000000010001101011000100;
assign LUT_3[56728] = 32'b00000000000000010001000011010011;
assign LUT_3[56729] = 32'b00000000000000010111101110110000;
assign LUT_3[56730] = 32'b00000000000000010011001010110111;
assign LUT_3[56731] = 32'b00000000000000011001110110010100;
assign LUT_3[56732] = 32'b00000000000000001110010001001001;
assign LUT_3[56733] = 32'b00000000000000010100111100100110;
assign LUT_3[56734] = 32'b00000000000000010000011000101101;
assign LUT_3[56735] = 32'b00000000000000010111000100001010;
assign LUT_3[56736] = 32'b00000000000000001001100101101010;
assign LUT_3[56737] = 32'b00000000000000010000010001000111;
assign LUT_3[56738] = 32'b00000000000000001011101101001110;
assign LUT_3[56739] = 32'b00000000000000010010011000101011;
assign LUT_3[56740] = 32'b00000000000000000110110011100000;
assign LUT_3[56741] = 32'b00000000000000001101011110111101;
assign LUT_3[56742] = 32'b00000000000000001000111011000100;
assign LUT_3[56743] = 32'b00000000000000001111100110100001;
assign LUT_3[56744] = 32'b00000000000000001110111110110000;
assign LUT_3[56745] = 32'b00000000000000010101101010001101;
assign LUT_3[56746] = 32'b00000000000000010001000110010100;
assign LUT_3[56747] = 32'b00000000000000010111110001110001;
assign LUT_3[56748] = 32'b00000000000000001100001100100110;
assign LUT_3[56749] = 32'b00000000000000010010111000000011;
assign LUT_3[56750] = 32'b00000000000000001110010100001010;
assign LUT_3[56751] = 32'b00000000000000010100111111100111;
assign LUT_3[56752] = 32'b00000000000000001100111000101101;
assign LUT_3[56753] = 32'b00000000000000010011100100001010;
assign LUT_3[56754] = 32'b00000000000000001111000000010001;
assign LUT_3[56755] = 32'b00000000000000010101101011101110;
assign LUT_3[56756] = 32'b00000000000000001010000110100011;
assign LUT_3[56757] = 32'b00000000000000010000110010000000;
assign LUT_3[56758] = 32'b00000000000000001100001110000111;
assign LUT_3[56759] = 32'b00000000000000010010111001100100;
assign LUT_3[56760] = 32'b00000000000000010010010001110011;
assign LUT_3[56761] = 32'b00000000000000011000111101010000;
assign LUT_3[56762] = 32'b00000000000000010100011001010111;
assign LUT_3[56763] = 32'b00000000000000011011000100110100;
assign LUT_3[56764] = 32'b00000000000000001111011111101001;
assign LUT_3[56765] = 32'b00000000000000010110001011000110;
assign LUT_3[56766] = 32'b00000000000000010001100111001101;
assign LUT_3[56767] = 32'b00000000000000011000010010101010;
assign LUT_3[56768] = 32'b00000000000000001000001111110101;
assign LUT_3[56769] = 32'b00000000000000001110111011010010;
assign LUT_3[56770] = 32'b00000000000000001010010111011001;
assign LUT_3[56771] = 32'b00000000000000010001000010110110;
assign LUT_3[56772] = 32'b00000000000000000101011101101011;
assign LUT_3[56773] = 32'b00000000000000001100001001001000;
assign LUT_3[56774] = 32'b00000000000000000111100101001111;
assign LUT_3[56775] = 32'b00000000000000001110010000101100;
assign LUT_3[56776] = 32'b00000000000000001101101000111011;
assign LUT_3[56777] = 32'b00000000000000010100010100011000;
assign LUT_3[56778] = 32'b00000000000000001111110000011111;
assign LUT_3[56779] = 32'b00000000000000010110011011111100;
assign LUT_3[56780] = 32'b00000000000000001010110110110001;
assign LUT_3[56781] = 32'b00000000000000010001100010001110;
assign LUT_3[56782] = 32'b00000000000000001100111110010101;
assign LUT_3[56783] = 32'b00000000000000010011101001110010;
assign LUT_3[56784] = 32'b00000000000000001011100010111000;
assign LUT_3[56785] = 32'b00000000000000010010001110010101;
assign LUT_3[56786] = 32'b00000000000000001101101010011100;
assign LUT_3[56787] = 32'b00000000000000010100010101111001;
assign LUT_3[56788] = 32'b00000000000000001000110000101110;
assign LUT_3[56789] = 32'b00000000000000001111011100001011;
assign LUT_3[56790] = 32'b00000000000000001010111000010010;
assign LUT_3[56791] = 32'b00000000000000010001100011101111;
assign LUT_3[56792] = 32'b00000000000000010000111011111110;
assign LUT_3[56793] = 32'b00000000000000010111100111011011;
assign LUT_3[56794] = 32'b00000000000000010011000011100010;
assign LUT_3[56795] = 32'b00000000000000011001101110111111;
assign LUT_3[56796] = 32'b00000000000000001110001001110100;
assign LUT_3[56797] = 32'b00000000000000010100110101010001;
assign LUT_3[56798] = 32'b00000000000000010000010001011000;
assign LUT_3[56799] = 32'b00000000000000010110111100110101;
assign LUT_3[56800] = 32'b00000000000000001001011110010101;
assign LUT_3[56801] = 32'b00000000000000010000001001110010;
assign LUT_3[56802] = 32'b00000000000000001011100101111001;
assign LUT_3[56803] = 32'b00000000000000010010010001010110;
assign LUT_3[56804] = 32'b00000000000000000110101100001011;
assign LUT_3[56805] = 32'b00000000000000001101010111101000;
assign LUT_3[56806] = 32'b00000000000000001000110011101111;
assign LUT_3[56807] = 32'b00000000000000001111011111001100;
assign LUT_3[56808] = 32'b00000000000000001110110111011011;
assign LUT_3[56809] = 32'b00000000000000010101100010111000;
assign LUT_3[56810] = 32'b00000000000000010000111110111111;
assign LUT_3[56811] = 32'b00000000000000010111101010011100;
assign LUT_3[56812] = 32'b00000000000000001100000101010001;
assign LUT_3[56813] = 32'b00000000000000010010110000101110;
assign LUT_3[56814] = 32'b00000000000000001110001100110101;
assign LUT_3[56815] = 32'b00000000000000010100111000010010;
assign LUT_3[56816] = 32'b00000000000000001100110001011000;
assign LUT_3[56817] = 32'b00000000000000010011011100110101;
assign LUT_3[56818] = 32'b00000000000000001110111000111100;
assign LUT_3[56819] = 32'b00000000000000010101100100011001;
assign LUT_3[56820] = 32'b00000000000000001001111111001110;
assign LUT_3[56821] = 32'b00000000000000010000101010101011;
assign LUT_3[56822] = 32'b00000000000000001100000110110010;
assign LUT_3[56823] = 32'b00000000000000010010110010001111;
assign LUT_3[56824] = 32'b00000000000000010010001010011110;
assign LUT_3[56825] = 32'b00000000000000011000110101111011;
assign LUT_3[56826] = 32'b00000000000000010100010010000010;
assign LUT_3[56827] = 32'b00000000000000011010111101011111;
assign LUT_3[56828] = 32'b00000000000000001111011000010100;
assign LUT_3[56829] = 32'b00000000000000010110000011110001;
assign LUT_3[56830] = 32'b00000000000000010001011111111000;
assign LUT_3[56831] = 32'b00000000000000011000001011010101;
assign LUT_3[56832] = 32'b00000000000000001101010001110111;
assign LUT_3[56833] = 32'b00000000000000010011111101010100;
assign LUT_3[56834] = 32'b00000000000000001111011001011011;
assign LUT_3[56835] = 32'b00000000000000010110000100111000;
assign LUT_3[56836] = 32'b00000000000000001010011111101101;
assign LUT_3[56837] = 32'b00000000000000010001001011001010;
assign LUT_3[56838] = 32'b00000000000000001100100111010001;
assign LUT_3[56839] = 32'b00000000000000010011010010101110;
assign LUT_3[56840] = 32'b00000000000000010010101010111101;
assign LUT_3[56841] = 32'b00000000000000011001010110011010;
assign LUT_3[56842] = 32'b00000000000000010100110010100001;
assign LUT_3[56843] = 32'b00000000000000011011011101111110;
assign LUT_3[56844] = 32'b00000000000000001111111000110011;
assign LUT_3[56845] = 32'b00000000000000010110100100010000;
assign LUT_3[56846] = 32'b00000000000000010010000000010111;
assign LUT_3[56847] = 32'b00000000000000011000101011110100;
assign LUT_3[56848] = 32'b00000000000000010000100100111010;
assign LUT_3[56849] = 32'b00000000000000010111010000010111;
assign LUT_3[56850] = 32'b00000000000000010010101100011110;
assign LUT_3[56851] = 32'b00000000000000011001010111111011;
assign LUT_3[56852] = 32'b00000000000000001101110010110000;
assign LUT_3[56853] = 32'b00000000000000010100011110001101;
assign LUT_3[56854] = 32'b00000000000000001111111010010100;
assign LUT_3[56855] = 32'b00000000000000010110100101110001;
assign LUT_3[56856] = 32'b00000000000000010101111110000000;
assign LUT_3[56857] = 32'b00000000000000011100101001011101;
assign LUT_3[56858] = 32'b00000000000000011000000101100100;
assign LUT_3[56859] = 32'b00000000000000011110110001000001;
assign LUT_3[56860] = 32'b00000000000000010011001011110110;
assign LUT_3[56861] = 32'b00000000000000011001110111010011;
assign LUT_3[56862] = 32'b00000000000000010101010011011010;
assign LUT_3[56863] = 32'b00000000000000011011111110110111;
assign LUT_3[56864] = 32'b00000000000000001110100000010111;
assign LUT_3[56865] = 32'b00000000000000010101001011110100;
assign LUT_3[56866] = 32'b00000000000000010000100111111011;
assign LUT_3[56867] = 32'b00000000000000010111010011011000;
assign LUT_3[56868] = 32'b00000000000000001011101110001101;
assign LUT_3[56869] = 32'b00000000000000010010011001101010;
assign LUT_3[56870] = 32'b00000000000000001101110101110001;
assign LUT_3[56871] = 32'b00000000000000010100100001001110;
assign LUT_3[56872] = 32'b00000000000000010011111001011101;
assign LUT_3[56873] = 32'b00000000000000011010100100111010;
assign LUT_3[56874] = 32'b00000000000000010110000001000001;
assign LUT_3[56875] = 32'b00000000000000011100101100011110;
assign LUT_3[56876] = 32'b00000000000000010001000111010011;
assign LUT_3[56877] = 32'b00000000000000010111110010110000;
assign LUT_3[56878] = 32'b00000000000000010011001110110111;
assign LUT_3[56879] = 32'b00000000000000011001111010010100;
assign LUT_3[56880] = 32'b00000000000000010001110011011010;
assign LUT_3[56881] = 32'b00000000000000011000011110110111;
assign LUT_3[56882] = 32'b00000000000000010011111010111110;
assign LUT_3[56883] = 32'b00000000000000011010100110011011;
assign LUT_3[56884] = 32'b00000000000000001111000001010000;
assign LUT_3[56885] = 32'b00000000000000010101101100101101;
assign LUT_3[56886] = 32'b00000000000000010001001000110100;
assign LUT_3[56887] = 32'b00000000000000010111110100010001;
assign LUT_3[56888] = 32'b00000000000000010111001100100000;
assign LUT_3[56889] = 32'b00000000000000011101110111111101;
assign LUT_3[56890] = 32'b00000000000000011001010100000100;
assign LUT_3[56891] = 32'b00000000000000011111111111100001;
assign LUT_3[56892] = 32'b00000000000000010100011010010110;
assign LUT_3[56893] = 32'b00000000000000011011000101110011;
assign LUT_3[56894] = 32'b00000000000000010110100001111010;
assign LUT_3[56895] = 32'b00000000000000011101001101010111;
assign LUT_3[56896] = 32'b00000000000000001101001010100010;
assign LUT_3[56897] = 32'b00000000000000010011110101111111;
assign LUT_3[56898] = 32'b00000000000000001111010010000110;
assign LUT_3[56899] = 32'b00000000000000010101111101100011;
assign LUT_3[56900] = 32'b00000000000000001010011000011000;
assign LUT_3[56901] = 32'b00000000000000010001000011110101;
assign LUT_3[56902] = 32'b00000000000000001100011111111100;
assign LUT_3[56903] = 32'b00000000000000010011001011011001;
assign LUT_3[56904] = 32'b00000000000000010010100011101000;
assign LUT_3[56905] = 32'b00000000000000011001001111000101;
assign LUT_3[56906] = 32'b00000000000000010100101011001100;
assign LUT_3[56907] = 32'b00000000000000011011010110101001;
assign LUT_3[56908] = 32'b00000000000000001111110001011110;
assign LUT_3[56909] = 32'b00000000000000010110011100111011;
assign LUT_3[56910] = 32'b00000000000000010001111001000010;
assign LUT_3[56911] = 32'b00000000000000011000100100011111;
assign LUT_3[56912] = 32'b00000000000000010000011101100101;
assign LUT_3[56913] = 32'b00000000000000010111001001000010;
assign LUT_3[56914] = 32'b00000000000000010010100101001001;
assign LUT_3[56915] = 32'b00000000000000011001010000100110;
assign LUT_3[56916] = 32'b00000000000000001101101011011011;
assign LUT_3[56917] = 32'b00000000000000010100010110111000;
assign LUT_3[56918] = 32'b00000000000000001111110010111111;
assign LUT_3[56919] = 32'b00000000000000010110011110011100;
assign LUT_3[56920] = 32'b00000000000000010101110110101011;
assign LUT_3[56921] = 32'b00000000000000011100100010001000;
assign LUT_3[56922] = 32'b00000000000000010111111110001111;
assign LUT_3[56923] = 32'b00000000000000011110101001101100;
assign LUT_3[56924] = 32'b00000000000000010011000100100001;
assign LUT_3[56925] = 32'b00000000000000011001101111111110;
assign LUT_3[56926] = 32'b00000000000000010101001100000101;
assign LUT_3[56927] = 32'b00000000000000011011110111100010;
assign LUT_3[56928] = 32'b00000000000000001110011001000010;
assign LUT_3[56929] = 32'b00000000000000010101000100011111;
assign LUT_3[56930] = 32'b00000000000000010000100000100110;
assign LUT_3[56931] = 32'b00000000000000010111001100000011;
assign LUT_3[56932] = 32'b00000000000000001011100110111000;
assign LUT_3[56933] = 32'b00000000000000010010010010010101;
assign LUT_3[56934] = 32'b00000000000000001101101110011100;
assign LUT_3[56935] = 32'b00000000000000010100011001111001;
assign LUT_3[56936] = 32'b00000000000000010011110010001000;
assign LUT_3[56937] = 32'b00000000000000011010011101100101;
assign LUT_3[56938] = 32'b00000000000000010101111001101100;
assign LUT_3[56939] = 32'b00000000000000011100100101001001;
assign LUT_3[56940] = 32'b00000000000000010000111111111110;
assign LUT_3[56941] = 32'b00000000000000010111101011011011;
assign LUT_3[56942] = 32'b00000000000000010011000111100010;
assign LUT_3[56943] = 32'b00000000000000011001110010111111;
assign LUT_3[56944] = 32'b00000000000000010001101100000101;
assign LUT_3[56945] = 32'b00000000000000011000010111100010;
assign LUT_3[56946] = 32'b00000000000000010011110011101001;
assign LUT_3[56947] = 32'b00000000000000011010011111000110;
assign LUT_3[56948] = 32'b00000000000000001110111001111011;
assign LUT_3[56949] = 32'b00000000000000010101100101011000;
assign LUT_3[56950] = 32'b00000000000000010001000001011111;
assign LUT_3[56951] = 32'b00000000000000010111101100111100;
assign LUT_3[56952] = 32'b00000000000000010111000101001011;
assign LUT_3[56953] = 32'b00000000000000011101110000101000;
assign LUT_3[56954] = 32'b00000000000000011001001100101111;
assign LUT_3[56955] = 32'b00000000000000011111111000001100;
assign LUT_3[56956] = 32'b00000000000000010100010011000001;
assign LUT_3[56957] = 32'b00000000000000011010111110011110;
assign LUT_3[56958] = 32'b00000000000000010110011010100101;
assign LUT_3[56959] = 32'b00000000000000011101000110000010;
assign LUT_3[56960] = 32'b00000000000000001111011100110101;
assign LUT_3[56961] = 32'b00000000000000010110001000010010;
assign LUT_3[56962] = 32'b00000000000000010001100100011001;
assign LUT_3[56963] = 32'b00000000000000011000001111110110;
assign LUT_3[56964] = 32'b00000000000000001100101010101011;
assign LUT_3[56965] = 32'b00000000000000010011010110001000;
assign LUT_3[56966] = 32'b00000000000000001110110010001111;
assign LUT_3[56967] = 32'b00000000000000010101011101101100;
assign LUT_3[56968] = 32'b00000000000000010100110101111011;
assign LUT_3[56969] = 32'b00000000000000011011100001011000;
assign LUT_3[56970] = 32'b00000000000000010110111101011111;
assign LUT_3[56971] = 32'b00000000000000011101101000111100;
assign LUT_3[56972] = 32'b00000000000000010010000011110001;
assign LUT_3[56973] = 32'b00000000000000011000101111001110;
assign LUT_3[56974] = 32'b00000000000000010100001011010101;
assign LUT_3[56975] = 32'b00000000000000011010110110110010;
assign LUT_3[56976] = 32'b00000000000000010010101111111000;
assign LUT_3[56977] = 32'b00000000000000011001011011010101;
assign LUT_3[56978] = 32'b00000000000000010100110111011100;
assign LUT_3[56979] = 32'b00000000000000011011100010111001;
assign LUT_3[56980] = 32'b00000000000000001111111101101110;
assign LUT_3[56981] = 32'b00000000000000010110101001001011;
assign LUT_3[56982] = 32'b00000000000000010010000101010010;
assign LUT_3[56983] = 32'b00000000000000011000110000101111;
assign LUT_3[56984] = 32'b00000000000000011000001000111110;
assign LUT_3[56985] = 32'b00000000000000011110110100011011;
assign LUT_3[56986] = 32'b00000000000000011010010000100010;
assign LUT_3[56987] = 32'b00000000000000100000111011111111;
assign LUT_3[56988] = 32'b00000000000000010101010110110100;
assign LUT_3[56989] = 32'b00000000000000011100000010010001;
assign LUT_3[56990] = 32'b00000000000000010111011110011000;
assign LUT_3[56991] = 32'b00000000000000011110001001110101;
assign LUT_3[56992] = 32'b00000000000000010000101011010101;
assign LUT_3[56993] = 32'b00000000000000010111010110110010;
assign LUT_3[56994] = 32'b00000000000000010010110010111001;
assign LUT_3[56995] = 32'b00000000000000011001011110010110;
assign LUT_3[56996] = 32'b00000000000000001101111001001011;
assign LUT_3[56997] = 32'b00000000000000010100100100101000;
assign LUT_3[56998] = 32'b00000000000000010000000000101111;
assign LUT_3[56999] = 32'b00000000000000010110101100001100;
assign LUT_3[57000] = 32'b00000000000000010110000100011011;
assign LUT_3[57001] = 32'b00000000000000011100101111111000;
assign LUT_3[57002] = 32'b00000000000000011000001011111111;
assign LUT_3[57003] = 32'b00000000000000011110110111011100;
assign LUT_3[57004] = 32'b00000000000000010011010010010001;
assign LUT_3[57005] = 32'b00000000000000011001111101101110;
assign LUT_3[57006] = 32'b00000000000000010101011001110101;
assign LUT_3[57007] = 32'b00000000000000011100000101010010;
assign LUT_3[57008] = 32'b00000000000000010011111110011000;
assign LUT_3[57009] = 32'b00000000000000011010101001110101;
assign LUT_3[57010] = 32'b00000000000000010110000101111100;
assign LUT_3[57011] = 32'b00000000000000011100110001011001;
assign LUT_3[57012] = 32'b00000000000000010001001100001110;
assign LUT_3[57013] = 32'b00000000000000010111110111101011;
assign LUT_3[57014] = 32'b00000000000000010011010011110010;
assign LUT_3[57015] = 32'b00000000000000011001111111001111;
assign LUT_3[57016] = 32'b00000000000000011001010111011110;
assign LUT_3[57017] = 32'b00000000000000100000000010111011;
assign LUT_3[57018] = 32'b00000000000000011011011111000010;
assign LUT_3[57019] = 32'b00000000000000100010001010011111;
assign LUT_3[57020] = 32'b00000000000000010110100101010100;
assign LUT_3[57021] = 32'b00000000000000011101010000110001;
assign LUT_3[57022] = 32'b00000000000000011000101100111000;
assign LUT_3[57023] = 32'b00000000000000011111011000010101;
assign LUT_3[57024] = 32'b00000000000000001111010101100000;
assign LUT_3[57025] = 32'b00000000000000010110000000111101;
assign LUT_3[57026] = 32'b00000000000000010001011101000100;
assign LUT_3[57027] = 32'b00000000000000011000001000100001;
assign LUT_3[57028] = 32'b00000000000000001100100011010110;
assign LUT_3[57029] = 32'b00000000000000010011001110110011;
assign LUT_3[57030] = 32'b00000000000000001110101010111010;
assign LUT_3[57031] = 32'b00000000000000010101010110010111;
assign LUT_3[57032] = 32'b00000000000000010100101110100110;
assign LUT_3[57033] = 32'b00000000000000011011011010000011;
assign LUT_3[57034] = 32'b00000000000000010110110110001010;
assign LUT_3[57035] = 32'b00000000000000011101100001100111;
assign LUT_3[57036] = 32'b00000000000000010001111100011100;
assign LUT_3[57037] = 32'b00000000000000011000100111111001;
assign LUT_3[57038] = 32'b00000000000000010100000100000000;
assign LUT_3[57039] = 32'b00000000000000011010101111011101;
assign LUT_3[57040] = 32'b00000000000000010010101000100011;
assign LUT_3[57041] = 32'b00000000000000011001010100000000;
assign LUT_3[57042] = 32'b00000000000000010100110000000111;
assign LUT_3[57043] = 32'b00000000000000011011011011100100;
assign LUT_3[57044] = 32'b00000000000000001111110110011001;
assign LUT_3[57045] = 32'b00000000000000010110100001110110;
assign LUT_3[57046] = 32'b00000000000000010001111101111101;
assign LUT_3[57047] = 32'b00000000000000011000101001011010;
assign LUT_3[57048] = 32'b00000000000000011000000001101001;
assign LUT_3[57049] = 32'b00000000000000011110101101000110;
assign LUT_3[57050] = 32'b00000000000000011010001001001101;
assign LUT_3[57051] = 32'b00000000000000100000110100101010;
assign LUT_3[57052] = 32'b00000000000000010101001111011111;
assign LUT_3[57053] = 32'b00000000000000011011111010111100;
assign LUT_3[57054] = 32'b00000000000000010111010111000011;
assign LUT_3[57055] = 32'b00000000000000011110000010100000;
assign LUT_3[57056] = 32'b00000000000000010000100100000000;
assign LUT_3[57057] = 32'b00000000000000010111001111011101;
assign LUT_3[57058] = 32'b00000000000000010010101011100100;
assign LUT_3[57059] = 32'b00000000000000011001010111000001;
assign LUT_3[57060] = 32'b00000000000000001101110001110110;
assign LUT_3[57061] = 32'b00000000000000010100011101010011;
assign LUT_3[57062] = 32'b00000000000000001111111001011010;
assign LUT_3[57063] = 32'b00000000000000010110100100110111;
assign LUT_3[57064] = 32'b00000000000000010101111101000110;
assign LUT_3[57065] = 32'b00000000000000011100101000100011;
assign LUT_3[57066] = 32'b00000000000000011000000100101010;
assign LUT_3[57067] = 32'b00000000000000011110110000000111;
assign LUT_3[57068] = 32'b00000000000000010011001010111100;
assign LUT_3[57069] = 32'b00000000000000011001110110011001;
assign LUT_3[57070] = 32'b00000000000000010101010010100000;
assign LUT_3[57071] = 32'b00000000000000011011111101111101;
assign LUT_3[57072] = 32'b00000000000000010011110111000011;
assign LUT_3[57073] = 32'b00000000000000011010100010100000;
assign LUT_3[57074] = 32'b00000000000000010101111110100111;
assign LUT_3[57075] = 32'b00000000000000011100101010000100;
assign LUT_3[57076] = 32'b00000000000000010001000100111001;
assign LUT_3[57077] = 32'b00000000000000010111110000010110;
assign LUT_3[57078] = 32'b00000000000000010011001100011101;
assign LUT_3[57079] = 32'b00000000000000011001110111111010;
assign LUT_3[57080] = 32'b00000000000000011001010000001001;
assign LUT_3[57081] = 32'b00000000000000011111111011100110;
assign LUT_3[57082] = 32'b00000000000000011011010111101101;
assign LUT_3[57083] = 32'b00000000000000100010000011001010;
assign LUT_3[57084] = 32'b00000000000000010110011101111111;
assign LUT_3[57085] = 32'b00000000000000011101001001011100;
assign LUT_3[57086] = 32'b00000000000000011000100101100011;
assign LUT_3[57087] = 32'b00000000000000011111010001000000;
assign LUT_3[57088] = 32'b00000000000000001001100001011000;
assign LUT_3[57089] = 32'b00000000000000010000001100110101;
assign LUT_3[57090] = 32'b00000000000000001011101000111100;
assign LUT_3[57091] = 32'b00000000000000010010010100011001;
assign LUT_3[57092] = 32'b00000000000000000110101111001110;
assign LUT_3[57093] = 32'b00000000000000001101011010101011;
assign LUT_3[57094] = 32'b00000000000000001000110110110010;
assign LUT_3[57095] = 32'b00000000000000001111100010001111;
assign LUT_3[57096] = 32'b00000000000000001110111010011110;
assign LUT_3[57097] = 32'b00000000000000010101100101111011;
assign LUT_3[57098] = 32'b00000000000000010001000010000010;
assign LUT_3[57099] = 32'b00000000000000010111101101011111;
assign LUT_3[57100] = 32'b00000000000000001100001000010100;
assign LUT_3[57101] = 32'b00000000000000010010110011110001;
assign LUT_3[57102] = 32'b00000000000000001110001111111000;
assign LUT_3[57103] = 32'b00000000000000010100111011010101;
assign LUT_3[57104] = 32'b00000000000000001100110100011011;
assign LUT_3[57105] = 32'b00000000000000010011011111111000;
assign LUT_3[57106] = 32'b00000000000000001110111011111111;
assign LUT_3[57107] = 32'b00000000000000010101100111011100;
assign LUT_3[57108] = 32'b00000000000000001010000010010001;
assign LUT_3[57109] = 32'b00000000000000010000101101101110;
assign LUT_3[57110] = 32'b00000000000000001100001001110101;
assign LUT_3[57111] = 32'b00000000000000010010110101010010;
assign LUT_3[57112] = 32'b00000000000000010010001101100001;
assign LUT_3[57113] = 32'b00000000000000011000111000111110;
assign LUT_3[57114] = 32'b00000000000000010100010101000101;
assign LUT_3[57115] = 32'b00000000000000011011000000100010;
assign LUT_3[57116] = 32'b00000000000000001111011011010111;
assign LUT_3[57117] = 32'b00000000000000010110000110110100;
assign LUT_3[57118] = 32'b00000000000000010001100010111011;
assign LUT_3[57119] = 32'b00000000000000011000001110011000;
assign LUT_3[57120] = 32'b00000000000000001010101111111000;
assign LUT_3[57121] = 32'b00000000000000010001011011010101;
assign LUT_3[57122] = 32'b00000000000000001100110111011100;
assign LUT_3[57123] = 32'b00000000000000010011100010111001;
assign LUT_3[57124] = 32'b00000000000000000111111101101110;
assign LUT_3[57125] = 32'b00000000000000001110101001001011;
assign LUT_3[57126] = 32'b00000000000000001010000101010010;
assign LUT_3[57127] = 32'b00000000000000010000110000101111;
assign LUT_3[57128] = 32'b00000000000000010000001000111110;
assign LUT_3[57129] = 32'b00000000000000010110110100011011;
assign LUT_3[57130] = 32'b00000000000000010010010000100010;
assign LUT_3[57131] = 32'b00000000000000011000111011111111;
assign LUT_3[57132] = 32'b00000000000000001101010110110100;
assign LUT_3[57133] = 32'b00000000000000010100000010010001;
assign LUT_3[57134] = 32'b00000000000000001111011110011000;
assign LUT_3[57135] = 32'b00000000000000010110001001110101;
assign LUT_3[57136] = 32'b00000000000000001110000010111011;
assign LUT_3[57137] = 32'b00000000000000010100101110011000;
assign LUT_3[57138] = 32'b00000000000000010000001010011111;
assign LUT_3[57139] = 32'b00000000000000010110110101111100;
assign LUT_3[57140] = 32'b00000000000000001011010000110001;
assign LUT_3[57141] = 32'b00000000000000010001111100001110;
assign LUT_3[57142] = 32'b00000000000000001101011000010101;
assign LUT_3[57143] = 32'b00000000000000010100000011110010;
assign LUT_3[57144] = 32'b00000000000000010011011100000001;
assign LUT_3[57145] = 32'b00000000000000011010000111011110;
assign LUT_3[57146] = 32'b00000000000000010101100011100101;
assign LUT_3[57147] = 32'b00000000000000011100001111000010;
assign LUT_3[57148] = 32'b00000000000000010000101001110111;
assign LUT_3[57149] = 32'b00000000000000010111010101010100;
assign LUT_3[57150] = 32'b00000000000000010010110001011011;
assign LUT_3[57151] = 32'b00000000000000011001011100111000;
assign LUT_3[57152] = 32'b00000000000000001001011010000011;
assign LUT_3[57153] = 32'b00000000000000010000000101100000;
assign LUT_3[57154] = 32'b00000000000000001011100001100111;
assign LUT_3[57155] = 32'b00000000000000010010001101000100;
assign LUT_3[57156] = 32'b00000000000000000110100111111001;
assign LUT_3[57157] = 32'b00000000000000001101010011010110;
assign LUT_3[57158] = 32'b00000000000000001000101111011101;
assign LUT_3[57159] = 32'b00000000000000001111011010111010;
assign LUT_3[57160] = 32'b00000000000000001110110011001001;
assign LUT_3[57161] = 32'b00000000000000010101011110100110;
assign LUT_3[57162] = 32'b00000000000000010000111010101101;
assign LUT_3[57163] = 32'b00000000000000010111100110001010;
assign LUT_3[57164] = 32'b00000000000000001100000000111111;
assign LUT_3[57165] = 32'b00000000000000010010101100011100;
assign LUT_3[57166] = 32'b00000000000000001110001000100011;
assign LUT_3[57167] = 32'b00000000000000010100110100000000;
assign LUT_3[57168] = 32'b00000000000000001100101101000110;
assign LUT_3[57169] = 32'b00000000000000010011011000100011;
assign LUT_3[57170] = 32'b00000000000000001110110100101010;
assign LUT_3[57171] = 32'b00000000000000010101100000000111;
assign LUT_3[57172] = 32'b00000000000000001001111010111100;
assign LUT_3[57173] = 32'b00000000000000010000100110011001;
assign LUT_3[57174] = 32'b00000000000000001100000010100000;
assign LUT_3[57175] = 32'b00000000000000010010101101111101;
assign LUT_3[57176] = 32'b00000000000000010010000110001100;
assign LUT_3[57177] = 32'b00000000000000011000110001101001;
assign LUT_3[57178] = 32'b00000000000000010100001101110000;
assign LUT_3[57179] = 32'b00000000000000011010111001001101;
assign LUT_3[57180] = 32'b00000000000000001111010100000010;
assign LUT_3[57181] = 32'b00000000000000010101111111011111;
assign LUT_3[57182] = 32'b00000000000000010001011011100110;
assign LUT_3[57183] = 32'b00000000000000011000000111000011;
assign LUT_3[57184] = 32'b00000000000000001010101000100011;
assign LUT_3[57185] = 32'b00000000000000010001010100000000;
assign LUT_3[57186] = 32'b00000000000000001100110000000111;
assign LUT_3[57187] = 32'b00000000000000010011011011100100;
assign LUT_3[57188] = 32'b00000000000000000111110110011001;
assign LUT_3[57189] = 32'b00000000000000001110100001110110;
assign LUT_3[57190] = 32'b00000000000000001001111101111101;
assign LUT_3[57191] = 32'b00000000000000010000101001011010;
assign LUT_3[57192] = 32'b00000000000000010000000001101001;
assign LUT_3[57193] = 32'b00000000000000010110101101000110;
assign LUT_3[57194] = 32'b00000000000000010010001001001101;
assign LUT_3[57195] = 32'b00000000000000011000110100101010;
assign LUT_3[57196] = 32'b00000000000000001101001111011111;
assign LUT_3[57197] = 32'b00000000000000010011111010111100;
assign LUT_3[57198] = 32'b00000000000000001111010111000011;
assign LUT_3[57199] = 32'b00000000000000010110000010100000;
assign LUT_3[57200] = 32'b00000000000000001101111011100110;
assign LUT_3[57201] = 32'b00000000000000010100100111000011;
assign LUT_3[57202] = 32'b00000000000000010000000011001010;
assign LUT_3[57203] = 32'b00000000000000010110101110100111;
assign LUT_3[57204] = 32'b00000000000000001011001001011100;
assign LUT_3[57205] = 32'b00000000000000010001110100111001;
assign LUT_3[57206] = 32'b00000000000000001101010001000000;
assign LUT_3[57207] = 32'b00000000000000010011111100011101;
assign LUT_3[57208] = 32'b00000000000000010011010100101100;
assign LUT_3[57209] = 32'b00000000000000011010000000001001;
assign LUT_3[57210] = 32'b00000000000000010101011100010000;
assign LUT_3[57211] = 32'b00000000000000011100000111101101;
assign LUT_3[57212] = 32'b00000000000000010000100010100010;
assign LUT_3[57213] = 32'b00000000000000010111001101111111;
assign LUT_3[57214] = 32'b00000000000000010010101010000110;
assign LUT_3[57215] = 32'b00000000000000011001010101100011;
assign LUT_3[57216] = 32'b00000000000000001011101100010110;
assign LUT_3[57217] = 32'b00000000000000010010010111110011;
assign LUT_3[57218] = 32'b00000000000000001101110011111010;
assign LUT_3[57219] = 32'b00000000000000010100011111010111;
assign LUT_3[57220] = 32'b00000000000000001000111010001100;
assign LUT_3[57221] = 32'b00000000000000001111100101101001;
assign LUT_3[57222] = 32'b00000000000000001011000001110000;
assign LUT_3[57223] = 32'b00000000000000010001101101001101;
assign LUT_3[57224] = 32'b00000000000000010001000101011100;
assign LUT_3[57225] = 32'b00000000000000010111110000111001;
assign LUT_3[57226] = 32'b00000000000000010011001101000000;
assign LUT_3[57227] = 32'b00000000000000011001111000011101;
assign LUT_3[57228] = 32'b00000000000000001110010011010010;
assign LUT_3[57229] = 32'b00000000000000010100111110101111;
assign LUT_3[57230] = 32'b00000000000000010000011010110110;
assign LUT_3[57231] = 32'b00000000000000010111000110010011;
assign LUT_3[57232] = 32'b00000000000000001110111111011001;
assign LUT_3[57233] = 32'b00000000000000010101101010110110;
assign LUT_3[57234] = 32'b00000000000000010001000110111101;
assign LUT_3[57235] = 32'b00000000000000010111110010011010;
assign LUT_3[57236] = 32'b00000000000000001100001101001111;
assign LUT_3[57237] = 32'b00000000000000010010111000101100;
assign LUT_3[57238] = 32'b00000000000000001110010100110011;
assign LUT_3[57239] = 32'b00000000000000010101000000010000;
assign LUT_3[57240] = 32'b00000000000000010100011000011111;
assign LUT_3[57241] = 32'b00000000000000011011000011111100;
assign LUT_3[57242] = 32'b00000000000000010110100000000011;
assign LUT_3[57243] = 32'b00000000000000011101001011100000;
assign LUT_3[57244] = 32'b00000000000000010001100110010101;
assign LUT_3[57245] = 32'b00000000000000011000010001110010;
assign LUT_3[57246] = 32'b00000000000000010011101101111001;
assign LUT_3[57247] = 32'b00000000000000011010011001010110;
assign LUT_3[57248] = 32'b00000000000000001100111010110110;
assign LUT_3[57249] = 32'b00000000000000010011100110010011;
assign LUT_3[57250] = 32'b00000000000000001111000010011010;
assign LUT_3[57251] = 32'b00000000000000010101101101110111;
assign LUT_3[57252] = 32'b00000000000000001010001000101100;
assign LUT_3[57253] = 32'b00000000000000010000110100001001;
assign LUT_3[57254] = 32'b00000000000000001100010000010000;
assign LUT_3[57255] = 32'b00000000000000010010111011101101;
assign LUT_3[57256] = 32'b00000000000000010010010011111100;
assign LUT_3[57257] = 32'b00000000000000011000111111011001;
assign LUT_3[57258] = 32'b00000000000000010100011011100000;
assign LUT_3[57259] = 32'b00000000000000011011000110111101;
assign LUT_3[57260] = 32'b00000000000000001111100001110010;
assign LUT_3[57261] = 32'b00000000000000010110001101001111;
assign LUT_3[57262] = 32'b00000000000000010001101001010110;
assign LUT_3[57263] = 32'b00000000000000011000010100110011;
assign LUT_3[57264] = 32'b00000000000000010000001101111001;
assign LUT_3[57265] = 32'b00000000000000010110111001010110;
assign LUT_3[57266] = 32'b00000000000000010010010101011101;
assign LUT_3[57267] = 32'b00000000000000011001000000111010;
assign LUT_3[57268] = 32'b00000000000000001101011011101111;
assign LUT_3[57269] = 32'b00000000000000010100000111001100;
assign LUT_3[57270] = 32'b00000000000000001111100011010011;
assign LUT_3[57271] = 32'b00000000000000010110001110110000;
assign LUT_3[57272] = 32'b00000000000000010101100110111111;
assign LUT_3[57273] = 32'b00000000000000011100010010011100;
assign LUT_3[57274] = 32'b00000000000000010111101110100011;
assign LUT_3[57275] = 32'b00000000000000011110011010000000;
assign LUT_3[57276] = 32'b00000000000000010010110100110101;
assign LUT_3[57277] = 32'b00000000000000011001100000010010;
assign LUT_3[57278] = 32'b00000000000000010100111100011001;
assign LUT_3[57279] = 32'b00000000000000011011100111110110;
assign LUT_3[57280] = 32'b00000000000000001011100101000001;
assign LUT_3[57281] = 32'b00000000000000010010010000011110;
assign LUT_3[57282] = 32'b00000000000000001101101100100101;
assign LUT_3[57283] = 32'b00000000000000010100011000000010;
assign LUT_3[57284] = 32'b00000000000000001000110010110111;
assign LUT_3[57285] = 32'b00000000000000001111011110010100;
assign LUT_3[57286] = 32'b00000000000000001010111010011011;
assign LUT_3[57287] = 32'b00000000000000010001100101111000;
assign LUT_3[57288] = 32'b00000000000000010000111110000111;
assign LUT_3[57289] = 32'b00000000000000010111101001100100;
assign LUT_3[57290] = 32'b00000000000000010011000101101011;
assign LUT_3[57291] = 32'b00000000000000011001110001001000;
assign LUT_3[57292] = 32'b00000000000000001110001011111101;
assign LUT_3[57293] = 32'b00000000000000010100110111011010;
assign LUT_3[57294] = 32'b00000000000000010000010011100001;
assign LUT_3[57295] = 32'b00000000000000010110111110111110;
assign LUT_3[57296] = 32'b00000000000000001110111000000100;
assign LUT_3[57297] = 32'b00000000000000010101100011100001;
assign LUT_3[57298] = 32'b00000000000000010000111111101000;
assign LUT_3[57299] = 32'b00000000000000010111101011000101;
assign LUT_3[57300] = 32'b00000000000000001100000101111010;
assign LUT_3[57301] = 32'b00000000000000010010110001010111;
assign LUT_3[57302] = 32'b00000000000000001110001101011110;
assign LUT_3[57303] = 32'b00000000000000010100111000111011;
assign LUT_3[57304] = 32'b00000000000000010100010001001010;
assign LUT_3[57305] = 32'b00000000000000011010111100100111;
assign LUT_3[57306] = 32'b00000000000000010110011000101110;
assign LUT_3[57307] = 32'b00000000000000011101000100001011;
assign LUT_3[57308] = 32'b00000000000000010001011111000000;
assign LUT_3[57309] = 32'b00000000000000011000001010011101;
assign LUT_3[57310] = 32'b00000000000000010011100110100100;
assign LUT_3[57311] = 32'b00000000000000011010010010000001;
assign LUT_3[57312] = 32'b00000000000000001100110011100001;
assign LUT_3[57313] = 32'b00000000000000010011011110111110;
assign LUT_3[57314] = 32'b00000000000000001110111011000101;
assign LUT_3[57315] = 32'b00000000000000010101100110100010;
assign LUT_3[57316] = 32'b00000000000000001010000001010111;
assign LUT_3[57317] = 32'b00000000000000010000101100110100;
assign LUT_3[57318] = 32'b00000000000000001100001000111011;
assign LUT_3[57319] = 32'b00000000000000010010110100011000;
assign LUT_3[57320] = 32'b00000000000000010010001100100111;
assign LUT_3[57321] = 32'b00000000000000011000111000000100;
assign LUT_3[57322] = 32'b00000000000000010100010100001011;
assign LUT_3[57323] = 32'b00000000000000011010111111101000;
assign LUT_3[57324] = 32'b00000000000000001111011010011101;
assign LUT_3[57325] = 32'b00000000000000010110000101111010;
assign LUT_3[57326] = 32'b00000000000000010001100010000001;
assign LUT_3[57327] = 32'b00000000000000011000001101011110;
assign LUT_3[57328] = 32'b00000000000000010000000110100100;
assign LUT_3[57329] = 32'b00000000000000010110110010000001;
assign LUT_3[57330] = 32'b00000000000000010010001110001000;
assign LUT_3[57331] = 32'b00000000000000011000111001100101;
assign LUT_3[57332] = 32'b00000000000000001101010100011010;
assign LUT_3[57333] = 32'b00000000000000010011111111110111;
assign LUT_3[57334] = 32'b00000000000000001111011011111110;
assign LUT_3[57335] = 32'b00000000000000010110000111011011;
assign LUT_3[57336] = 32'b00000000000000010101011111101010;
assign LUT_3[57337] = 32'b00000000000000011100001011000111;
assign LUT_3[57338] = 32'b00000000000000010111100111001110;
assign LUT_3[57339] = 32'b00000000000000011110010010101011;
assign LUT_3[57340] = 32'b00000000000000010010101101100000;
assign LUT_3[57341] = 32'b00000000000000011001011000111101;
assign LUT_3[57342] = 32'b00000000000000010100110101000100;
assign LUT_3[57343] = 32'b00000000000000011011100000100001;
assign LUT_3[57344] = 32'b00000000000000000011100101100000;
assign LUT_3[57345] = 32'b00000000000000001010010000111101;
assign LUT_3[57346] = 32'b00000000000000000101101101000100;
assign LUT_3[57347] = 32'b00000000000000001100011000100001;
assign LUT_3[57348] = 32'b00000000000000000000110011010110;
assign LUT_3[57349] = 32'b00000000000000000111011110110011;
assign LUT_3[57350] = 32'b00000000000000000010111010111010;
assign LUT_3[57351] = 32'b00000000000000001001100110010111;
assign LUT_3[57352] = 32'b00000000000000001000111110100110;
assign LUT_3[57353] = 32'b00000000000000001111101010000011;
assign LUT_3[57354] = 32'b00000000000000001011000110001010;
assign LUT_3[57355] = 32'b00000000000000010001110001100111;
assign LUT_3[57356] = 32'b00000000000000000110001100011100;
assign LUT_3[57357] = 32'b00000000000000001100110111111001;
assign LUT_3[57358] = 32'b00000000000000001000010100000000;
assign LUT_3[57359] = 32'b00000000000000001110111111011101;
assign LUT_3[57360] = 32'b00000000000000000110111000100011;
assign LUT_3[57361] = 32'b00000000000000001101100100000000;
assign LUT_3[57362] = 32'b00000000000000001001000000000111;
assign LUT_3[57363] = 32'b00000000000000001111101011100100;
assign LUT_3[57364] = 32'b00000000000000000100000110011001;
assign LUT_3[57365] = 32'b00000000000000001010110001110110;
assign LUT_3[57366] = 32'b00000000000000000110001101111101;
assign LUT_3[57367] = 32'b00000000000000001100111001011010;
assign LUT_3[57368] = 32'b00000000000000001100010001101001;
assign LUT_3[57369] = 32'b00000000000000010010111101000110;
assign LUT_3[57370] = 32'b00000000000000001110011001001101;
assign LUT_3[57371] = 32'b00000000000000010101000100101010;
assign LUT_3[57372] = 32'b00000000000000001001011111011111;
assign LUT_3[57373] = 32'b00000000000000010000001010111100;
assign LUT_3[57374] = 32'b00000000000000001011100111000011;
assign LUT_3[57375] = 32'b00000000000000010010010010100000;
assign LUT_3[57376] = 32'b00000000000000000100110100000000;
assign LUT_3[57377] = 32'b00000000000000001011011111011101;
assign LUT_3[57378] = 32'b00000000000000000110111011100100;
assign LUT_3[57379] = 32'b00000000000000001101100111000001;
assign LUT_3[57380] = 32'b00000000000000000010000001110110;
assign LUT_3[57381] = 32'b00000000000000001000101101010011;
assign LUT_3[57382] = 32'b00000000000000000100001001011010;
assign LUT_3[57383] = 32'b00000000000000001010110100110111;
assign LUT_3[57384] = 32'b00000000000000001010001101000110;
assign LUT_3[57385] = 32'b00000000000000010000111000100011;
assign LUT_3[57386] = 32'b00000000000000001100010100101010;
assign LUT_3[57387] = 32'b00000000000000010011000000000111;
assign LUT_3[57388] = 32'b00000000000000000111011010111100;
assign LUT_3[57389] = 32'b00000000000000001110000110011001;
assign LUT_3[57390] = 32'b00000000000000001001100010100000;
assign LUT_3[57391] = 32'b00000000000000010000001101111101;
assign LUT_3[57392] = 32'b00000000000000001000000111000011;
assign LUT_3[57393] = 32'b00000000000000001110110010100000;
assign LUT_3[57394] = 32'b00000000000000001010001110100111;
assign LUT_3[57395] = 32'b00000000000000010000111010000100;
assign LUT_3[57396] = 32'b00000000000000000101010100111001;
assign LUT_3[57397] = 32'b00000000000000001100000000010110;
assign LUT_3[57398] = 32'b00000000000000000111011100011101;
assign LUT_3[57399] = 32'b00000000000000001110000111111010;
assign LUT_3[57400] = 32'b00000000000000001101100000001001;
assign LUT_3[57401] = 32'b00000000000000010100001011100110;
assign LUT_3[57402] = 32'b00000000000000001111100111101101;
assign LUT_3[57403] = 32'b00000000000000010110010011001010;
assign LUT_3[57404] = 32'b00000000000000001010101101111111;
assign LUT_3[57405] = 32'b00000000000000010001011001011100;
assign LUT_3[57406] = 32'b00000000000000001100110101100011;
assign LUT_3[57407] = 32'b00000000000000010011100001000000;
assign LUT_3[57408] = 32'b00000000000000000011011110001011;
assign LUT_3[57409] = 32'b00000000000000001010001001101000;
assign LUT_3[57410] = 32'b00000000000000000101100101101111;
assign LUT_3[57411] = 32'b00000000000000001100010001001100;
assign LUT_3[57412] = 32'b00000000000000000000101100000001;
assign LUT_3[57413] = 32'b00000000000000000111010111011110;
assign LUT_3[57414] = 32'b00000000000000000010110011100101;
assign LUT_3[57415] = 32'b00000000000000001001011111000010;
assign LUT_3[57416] = 32'b00000000000000001000110111010001;
assign LUT_3[57417] = 32'b00000000000000001111100010101110;
assign LUT_3[57418] = 32'b00000000000000001010111110110101;
assign LUT_3[57419] = 32'b00000000000000010001101010010010;
assign LUT_3[57420] = 32'b00000000000000000110000101000111;
assign LUT_3[57421] = 32'b00000000000000001100110000100100;
assign LUT_3[57422] = 32'b00000000000000001000001100101011;
assign LUT_3[57423] = 32'b00000000000000001110111000001000;
assign LUT_3[57424] = 32'b00000000000000000110110001001110;
assign LUT_3[57425] = 32'b00000000000000001101011100101011;
assign LUT_3[57426] = 32'b00000000000000001000111000110010;
assign LUT_3[57427] = 32'b00000000000000001111100100001111;
assign LUT_3[57428] = 32'b00000000000000000011111111000100;
assign LUT_3[57429] = 32'b00000000000000001010101010100001;
assign LUT_3[57430] = 32'b00000000000000000110000110101000;
assign LUT_3[57431] = 32'b00000000000000001100110010000101;
assign LUT_3[57432] = 32'b00000000000000001100001010010100;
assign LUT_3[57433] = 32'b00000000000000010010110101110001;
assign LUT_3[57434] = 32'b00000000000000001110010001111000;
assign LUT_3[57435] = 32'b00000000000000010100111101010101;
assign LUT_3[57436] = 32'b00000000000000001001011000001010;
assign LUT_3[57437] = 32'b00000000000000010000000011100111;
assign LUT_3[57438] = 32'b00000000000000001011011111101110;
assign LUT_3[57439] = 32'b00000000000000010010001011001011;
assign LUT_3[57440] = 32'b00000000000000000100101100101011;
assign LUT_3[57441] = 32'b00000000000000001011011000001000;
assign LUT_3[57442] = 32'b00000000000000000110110100001111;
assign LUT_3[57443] = 32'b00000000000000001101011111101100;
assign LUT_3[57444] = 32'b00000000000000000001111010100001;
assign LUT_3[57445] = 32'b00000000000000001000100101111110;
assign LUT_3[57446] = 32'b00000000000000000100000010000101;
assign LUT_3[57447] = 32'b00000000000000001010101101100010;
assign LUT_3[57448] = 32'b00000000000000001010000101110001;
assign LUT_3[57449] = 32'b00000000000000010000110001001110;
assign LUT_3[57450] = 32'b00000000000000001100001101010101;
assign LUT_3[57451] = 32'b00000000000000010010111000110010;
assign LUT_3[57452] = 32'b00000000000000000111010011100111;
assign LUT_3[57453] = 32'b00000000000000001101111111000100;
assign LUT_3[57454] = 32'b00000000000000001001011011001011;
assign LUT_3[57455] = 32'b00000000000000010000000110101000;
assign LUT_3[57456] = 32'b00000000000000000111111111101110;
assign LUT_3[57457] = 32'b00000000000000001110101011001011;
assign LUT_3[57458] = 32'b00000000000000001010000111010010;
assign LUT_3[57459] = 32'b00000000000000010000110010101111;
assign LUT_3[57460] = 32'b00000000000000000101001101100100;
assign LUT_3[57461] = 32'b00000000000000001011111001000001;
assign LUT_3[57462] = 32'b00000000000000000111010101001000;
assign LUT_3[57463] = 32'b00000000000000001110000000100101;
assign LUT_3[57464] = 32'b00000000000000001101011000110100;
assign LUT_3[57465] = 32'b00000000000000010100000100010001;
assign LUT_3[57466] = 32'b00000000000000001111100000011000;
assign LUT_3[57467] = 32'b00000000000000010110001011110101;
assign LUT_3[57468] = 32'b00000000000000001010100110101010;
assign LUT_3[57469] = 32'b00000000000000010001010010000111;
assign LUT_3[57470] = 32'b00000000000000001100101110001110;
assign LUT_3[57471] = 32'b00000000000000010011011001101011;
assign LUT_3[57472] = 32'b00000000000000000101110000011110;
assign LUT_3[57473] = 32'b00000000000000001100011011111011;
assign LUT_3[57474] = 32'b00000000000000000111111000000010;
assign LUT_3[57475] = 32'b00000000000000001110100011011111;
assign LUT_3[57476] = 32'b00000000000000000010111110010100;
assign LUT_3[57477] = 32'b00000000000000001001101001110001;
assign LUT_3[57478] = 32'b00000000000000000101000101111000;
assign LUT_3[57479] = 32'b00000000000000001011110001010101;
assign LUT_3[57480] = 32'b00000000000000001011001001100100;
assign LUT_3[57481] = 32'b00000000000000010001110101000001;
assign LUT_3[57482] = 32'b00000000000000001101010001001000;
assign LUT_3[57483] = 32'b00000000000000010011111100100101;
assign LUT_3[57484] = 32'b00000000000000001000010111011010;
assign LUT_3[57485] = 32'b00000000000000001111000010110111;
assign LUT_3[57486] = 32'b00000000000000001010011110111110;
assign LUT_3[57487] = 32'b00000000000000010001001010011011;
assign LUT_3[57488] = 32'b00000000000000001001000011100001;
assign LUT_3[57489] = 32'b00000000000000001111101110111110;
assign LUT_3[57490] = 32'b00000000000000001011001011000101;
assign LUT_3[57491] = 32'b00000000000000010001110110100010;
assign LUT_3[57492] = 32'b00000000000000000110010001010111;
assign LUT_3[57493] = 32'b00000000000000001100111100110100;
assign LUT_3[57494] = 32'b00000000000000001000011000111011;
assign LUT_3[57495] = 32'b00000000000000001111000100011000;
assign LUT_3[57496] = 32'b00000000000000001110011100100111;
assign LUT_3[57497] = 32'b00000000000000010101001000000100;
assign LUT_3[57498] = 32'b00000000000000010000100100001011;
assign LUT_3[57499] = 32'b00000000000000010111001111101000;
assign LUT_3[57500] = 32'b00000000000000001011101010011101;
assign LUT_3[57501] = 32'b00000000000000010010010101111010;
assign LUT_3[57502] = 32'b00000000000000001101110010000001;
assign LUT_3[57503] = 32'b00000000000000010100011101011110;
assign LUT_3[57504] = 32'b00000000000000000110111110111110;
assign LUT_3[57505] = 32'b00000000000000001101101010011011;
assign LUT_3[57506] = 32'b00000000000000001001000110100010;
assign LUT_3[57507] = 32'b00000000000000001111110001111111;
assign LUT_3[57508] = 32'b00000000000000000100001100110100;
assign LUT_3[57509] = 32'b00000000000000001010111000010001;
assign LUT_3[57510] = 32'b00000000000000000110010100011000;
assign LUT_3[57511] = 32'b00000000000000001100111111110101;
assign LUT_3[57512] = 32'b00000000000000001100011000000100;
assign LUT_3[57513] = 32'b00000000000000010011000011100001;
assign LUT_3[57514] = 32'b00000000000000001110011111101000;
assign LUT_3[57515] = 32'b00000000000000010101001011000101;
assign LUT_3[57516] = 32'b00000000000000001001100101111010;
assign LUT_3[57517] = 32'b00000000000000010000010001010111;
assign LUT_3[57518] = 32'b00000000000000001011101101011110;
assign LUT_3[57519] = 32'b00000000000000010010011000111011;
assign LUT_3[57520] = 32'b00000000000000001010010010000001;
assign LUT_3[57521] = 32'b00000000000000010000111101011110;
assign LUT_3[57522] = 32'b00000000000000001100011001100101;
assign LUT_3[57523] = 32'b00000000000000010011000101000010;
assign LUT_3[57524] = 32'b00000000000000000111011111110111;
assign LUT_3[57525] = 32'b00000000000000001110001011010100;
assign LUT_3[57526] = 32'b00000000000000001001100111011011;
assign LUT_3[57527] = 32'b00000000000000010000010010111000;
assign LUT_3[57528] = 32'b00000000000000001111101011000111;
assign LUT_3[57529] = 32'b00000000000000010110010110100100;
assign LUT_3[57530] = 32'b00000000000000010001110010101011;
assign LUT_3[57531] = 32'b00000000000000011000011110001000;
assign LUT_3[57532] = 32'b00000000000000001100111000111101;
assign LUT_3[57533] = 32'b00000000000000010011100100011010;
assign LUT_3[57534] = 32'b00000000000000001111000000100001;
assign LUT_3[57535] = 32'b00000000000000010101101011111110;
assign LUT_3[57536] = 32'b00000000000000000101101001001001;
assign LUT_3[57537] = 32'b00000000000000001100010100100110;
assign LUT_3[57538] = 32'b00000000000000000111110000101101;
assign LUT_3[57539] = 32'b00000000000000001110011100001010;
assign LUT_3[57540] = 32'b00000000000000000010110110111111;
assign LUT_3[57541] = 32'b00000000000000001001100010011100;
assign LUT_3[57542] = 32'b00000000000000000100111110100011;
assign LUT_3[57543] = 32'b00000000000000001011101010000000;
assign LUT_3[57544] = 32'b00000000000000001011000010001111;
assign LUT_3[57545] = 32'b00000000000000010001101101101100;
assign LUT_3[57546] = 32'b00000000000000001101001001110011;
assign LUT_3[57547] = 32'b00000000000000010011110101010000;
assign LUT_3[57548] = 32'b00000000000000001000010000000101;
assign LUT_3[57549] = 32'b00000000000000001110111011100010;
assign LUT_3[57550] = 32'b00000000000000001010010111101001;
assign LUT_3[57551] = 32'b00000000000000010001000011000110;
assign LUT_3[57552] = 32'b00000000000000001000111100001100;
assign LUT_3[57553] = 32'b00000000000000001111100111101001;
assign LUT_3[57554] = 32'b00000000000000001011000011110000;
assign LUT_3[57555] = 32'b00000000000000010001101111001101;
assign LUT_3[57556] = 32'b00000000000000000110001010000010;
assign LUT_3[57557] = 32'b00000000000000001100110101011111;
assign LUT_3[57558] = 32'b00000000000000001000010001100110;
assign LUT_3[57559] = 32'b00000000000000001110111101000011;
assign LUT_3[57560] = 32'b00000000000000001110010101010010;
assign LUT_3[57561] = 32'b00000000000000010101000000101111;
assign LUT_3[57562] = 32'b00000000000000010000011100110110;
assign LUT_3[57563] = 32'b00000000000000010111001000010011;
assign LUT_3[57564] = 32'b00000000000000001011100011001000;
assign LUT_3[57565] = 32'b00000000000000010010001110100101;
assign LUT_3[57566] = 32'b00000000000000001101101010101100;
assign LUT_3[57567] = 32'b00000000000000010100010110001001;
assign LUT_3[57568] = 32'b00000000000000000110110111101001;
assign LUT_3[57569] = 32'b00000000000000001101100011000110;
assign LUT_3[57570] = 32'b00000000000000001000111111001101;
assign LUT_3[57571] = 32'b00000000000000001111101010101010;
assign LUT_3[57572] = 32'b00000000000000000100000101011111;
assign LUT_3[57573] = 32'b00000000000000001010110000111100;
assign LUT_3[57574] = 32'b00000000000000000110001101000011;
assign LUT_3[57575] = 32'b00000000000000001100111000100000;
assign LUT_3[57576] = 32'b00000000000000001100010000101111;
assign LUT_3[57577] = 32'b00000000000000010010111100001100;
assign LUT_3[57578] = 32'b00000000000000001110011000010011;
assign LUT_3[57579] = 32'b00000000000000010101000011110000;
assign LUT_3[57580] = 32'b00000000000000001001011110100101;
assign LUT_3[57581] = 32'b00000000000000010000001010000010;
assign LUT_3[57582] = 32'b00000000000000001011100110001001;
assign LUT_3[57583] = 32'b00000000000000010010010001100110;
assign LUT_3[57584] = 32'b00000000000000001010001010101100;
assign LUT_3[57585] = 32'b00000000000000010000110110001001;
assign LUT_3[57586] = 32'b00000000000000001100010010010000;
assign LUT_3[57587] = 32'b00000000000000010010111101101101;
assign LUT_3[57588] = 32'b00000000000000000111011000100010;
assign LUT_3[57589] = 32'b00000000000000001110000011111111;
assign LUT_3[57590] = 32'b00000000000000001001100000000110;
assign LUT_3[57591] = 32'b00000000000000010000001011100011;
assign LUT_3[57592] = 32'b00000000000000001111100011110010;
assign LUT_3[57593] = 32'b00000000000000010110001111001111;
assign LUT_3[57594] = 32'b00000000000000010001101011010110;
assign LUT_3[57595] = 32'b00000000000000011000010110110011;
assign LUT_3[57596] = 32'b00000000000000001100110001101000;
assign LUT_3[57597] = 32'b00000000000000010011011101000101;
assign LUT_3[57598] = 32'b00000000000000001110111001001100;
assign LUT_3[57599] = 32'b00000000000000010101100100101001;
assign LUT_3[57600] = 32'b11111111111111111111110101000001;
assign LUT_3[57601] = 32'b00000000000000000110100000011110;
assign LUT_3[57602] = 32'b00000000000000000001111100100101;
assign LUT_3[57603] = 32'b00000000000000001000101000000010;
assign LUT_3[57604] = 32'b11111111111111111101000010110111;
assign LUT_3[57605] = 32'b00000000000000000011101110010100;
assign LUT_3[57606] = 32'b11111111111111111111001010011011;
assign LUT_3[57607] = 32'b00000000000000000101110101111000;
assign LUT_3[57608] = 32'b00000000000000000101001110000111;
assign LUT_3[57609] = 32'b00000000000000001011111001100100;
assign LUT_3[57610] = 32'b00000000000000000111010101101011;
assign LUT_3[57611] = 32'b00000000000000001110000001001000;
assign LUT_3[57612] = 32'b00000000000000000010011011111101;
assign LUT_3[57613] = 32'b00000000000000001001000111011010;
assign LUT_3[57614] = 32'b00000000000000000100100011100001;
assign LUT_3[57615] = 32'b00000000000000001011001110111110;
assign LUT_3[57616] = 32'b00000000000000000011001000000100;
assign LUT_3[57617] = 32'b00000000000000001001110011100001;
assign LUT_3[57618] = 32'b00000000000000000101001111101000;
assign LUT_3[57619] = 32'b00000000000000001011111011000101;
assign LUT_3[57620] = 32'b00000000000000000000010101111010;
assign LUT_3[57621] = 32'b00000000000000000111000001010111;
assign LUT_3[57622] = 32'b00000000000000000010011101011110;
assign LUT_3[57623] = 32'b00000000000000001001001000111011;
assign LUT_3[57624] = 32'b00000000000000001000100001001010;
assign LUT_3[57625] = 32'b00000000000000001111001100100111;
assign LUT_3[57626] = 32'b00000000000000001010101000101110;
assign LUT_3[57627] = 32'b00000000000000010001010100001011;
assign LUT_3[57628] = 32'b00000000000000000101101111000000;
assign LUT_3[57629] = 32'b00000000000000001100011010011101;
assign LUT_3[57630] = 32'b00000000000000000111110110100100;
assign LUT_3[57631] = 32'b00000000000000001110100010000001;
assign LUT_3[57632] = 32'b00000000000000000001000011100001;
assign LUT_3[57633] = 32'b00000000000000000111101110111110;
assign LUT_3[57634] = 32'b00000000000000000011001011000101;
assign LUT_3[57635] = 32'b00000000000000001001110110100010;
assign LUT_3[57636] = 32'b11111111111111111110010001010111;
assign LUT_3[57637] = 32'b00000000000000000100111100110100;
assign LUT_3[57638] = 32'b00000000000000000000011000111011;
assign LUT_3[57639] = 32'b00000000000000000111000100011000;
assign LUT_3[57640] = 32'b00000000000000000110011100100111;
assign LUT_3[57641] = 32'b00000000000000001101001000000100;
assign LUT_3[57642] = 32'b00000000000000001000100100001011;
assign LUT_3[57643] = 32'b00000000000000001111001111101000;
assign LUT_3[57644] = 32'b00000000000000000011101010011101;
assign LUT_3[57645] = 32'b00000000000000001010010101111010;
assign LUT_3[57646] = 32'b00000000000000000101110010000001;
assign LUT_3[57647] = 32'b00000000000000001100011101011110;
assign LUT_3[57648] = 32'b00000000000000000100010110100100;
assign LUT_3[57649] = 32'b00000000000000001011000010000001;
assign LUT_3[57650] = 32'b00000000000000000110011110001000;
assign LUT_3[57651] = 32'b00000000000000001101001001100101;
assign LUT_3[57652] = 32'b00000000000000000001100100011010;
assign LUT_3[57653] = 32'b00000000000000001000001111110111;
assign LUT_3[57654] = 32'b00000000000000000011101011111110;
assign LUT_3[57655] = 32'b00000000000000001010010111011011;
assign LUT_3[57656] = 32'b00000000000000001001101111101010;
assign LUT_3[57657] = 32'b00000000000000010000011011000111;
assign LUT_3[57658] = 32'b00000000000000001011110111001110;
assign LUT_3[57659] = 32'b00000000000000010010100010101011;
assign LUT_3[57660] = 32'b00000000000000000110111101100000;
assign LUT_3[57661] = 32'b00000000000000001101101000111101;
assign LUT_3[57662] = 32'b00000000000000001001000101000100;
assign LUT_3[57663] = 32'b00000000000000001111110000100001;
assign LUT_3[57664] = 32'b11111111111111111111101101101100;
assign LUT_3[57665] = 32'b00000000000000000110011001001001;
assign LUT_3[57666] = 32'b00000000000000000001110101010000;
assign LUT_3[57667] = 32'b00000000000000001000100000101101;
assign LUT_3[57668] = 32'b11111111111111111100111011100010;
assign LUT_3[57669] = 32'b00000000000000000011100110111111;
assign LUT_3[57670] = 32'b11111111111111111111000011000110;
assign LUT_3[57671] = 32'b00000000000000000101101110100011;
assign LUT_3[57672] = 32'b00000000000000000101000110110010;
assign LUT_3[57673] = 32'b00000000000000001011110010001111;
assign LUT_3[57674] = 32'b00000000000000000111001110010110;
assign LUT_3[57675] = 32'b00000000000000001101111001110011;
assign LUT_3[57676] = 32'b00000000000000000010010100101000;
assign LUT_3[57677] = 32'b00000000000000001001000000000101;
assign LUT_3[57678] = 32'b00000000000000000100011100001100;
assign LUT_3[57679] = 32'b00000000000000001011000111101001;
assign LUT_3[57680] = 32'b00000000000000000011000000101111;
assign LUT_3[57681] = 32'b00000000000000001001101100001100;
assign LUT_3[57682] = 32'b00000000000000000101001000010011;
assign LUT_3[57683] = 32'b00000000000000001011110011110000;
assign LUT_3[57684] = 32'b00000000000000000000001110100101;
assign LUT_3[57685] = 32'b00000000000000000110111010000010;
assign LUT_3[57686] = 32'b00000000000000000010010110001001;
assign LUT_3[57687] = 32'b00000000000000001001000001100110;
assign LUT_3[57688] = 32'b00000000000000001000011001110101;
assign LUT_3[57689] = 32'b00000000000000001111000101010010;
assign LUT_3[57690] = 32'b00000000000000001010100001011001;
assign LUT_3[57691] = 32'b00000000000000010001001100110110;
assign LUT_3[57692] = 32'b00000000000000000101100111101011;
assign LUT_3[57693] = 32'b00000000000000001100010011001000;
assign LUT_3[57694] = 32'b00000000000000000111101111001111;
assign LUT_3[57695] = 32'b00000000000000001110011010101100;
assign LUT_3[57696] = 32'b00000000000000000000111100001100;
assign LUT_3[57697] = 32'b00000000000000000111100111101001;
assign LUT_3[57698] = 32'b00000000000000000011000011110000;
assign LUT_3[57699] = 32'b00000000000000001001101111001101;
assign LUT_3[57700] = 32'b11111111111111111110001010000010;
assign LUT_3[57701] = 32'b00000000000000000100110101011111;
assign LUT_3[57702] = 32'b00000000000000000000010001100110;
assign LUT_3[57703] = 32'b00000000000000000110111101000011;
assign LUT_3[57704] = 32'b00000000000000000110010101010010;
assign LUT_3[57705] = 32'b00000000000000001101000000101111;
assign LUT_3[57706] = 32'b00000000000000001000011100110110;
assign LUT_3[57707] = 32'b00000000000000001111001000010011;
assign LUT_3[57708] = 32'b00000000000000000011100011001000;
assign LUT_3[57709] = 32'b00000000000000001010001110100101;
assign LUT_3[57710] = 32'b00000000000000000101101010101100;
assign LUT_3[57711] = 32'b00000000000000001100010110001001;
assign LUT_3[57712] = 32'b00000000000000000100001111001111;
assign LUT_3[57713] = 32'b00000000000000001010111010101100;
assign LUT_3[57714] = 32'b00000000000000000110010110110011;
assign LUT_3[57715] = 32'b00000000000000001101000010010000;
assign LUT_3[57716] = 32'b00000000000000000001011101000101;
assign LUT_3[57717] = 32'b00000000000000001000001000100010;
assign LUT_3[57718] = 32'b00000000000000000011100100101001;
assign LUT_3[57719] = 32'b00000000000000001010010000000110;
assign LUT_3[57720] = 32'b00000000000000001001101000010101;
assign LUT_3[57721] = 32'b00000000000000010000010011110010;
assign LUT_3[57722] = 32'b00000000000000001011101111111001;
assign LUT_3[57723] = 32'b00000000000000010010011011010110;
assign LUT_3[57724] = 32'b00000000000000000110110110001011;
assign LUT_3[57725] = 32'b00000000000000001101100001101000;
assign LUT_3[57726] = 32'b00000000000000001000111101101111;
assign LUT_3[57727] = 32'b00000000000000001111101001001100;
assign LUT_3[57728] = 32'b00000000000000000001111111111111;
assign LUT_3[57729] = 32'b00000000000000001000101011011100;
assign LUT_3[57730] = 32'b00000000000000000100000111100011;
assign LUT_3[57731] = 32'b00000000000000001010110011000000;
assign LUT_3[57732] = 32'b11111111111111111111001101110101;
assign LUT_3[57733] = 32'b00000000000000000101111001010010;
assign LUT_3[57734] = 32'b00000000000000000001010101011001;
assign LUT_3[57735] = 32'b00000000000000001000000000110110;
assign LUT_3[57736] = 32'b00000000000000000111011001000101;
assign LUT_3[57737] = 32'b00000000000000001110000100100010;
assign LUT_3[57738] = 32'b00000000000000001001100000101001;
assign LUT_3[57739] = 32'b00000000000000010000001100000110;
assign LUT_3[57740] = 32'b00000000000000000100100110111011;
assign LUT_3[57741] = 32'b00000000000000001011010010011000;
assign LUT_3[57742] = 32'b00000000000000000110101110011111;
assign LUT_3[57743] = 32'b00000000000000001101011001111100;
assign LUT_3[57744] = 32'b00000000000000000101010011000010;
assign LUT_3[57745] = 32'b00000000000000001011111110011111;
assign LUT_3[57746] = 32'b00000000000000000111011010100110;
assign LUT_3[57747] = 32'b00000000000000001110000110000011;
assign LUT_3[57748] = 32'b00000000000000000010100000111000;
assign LUT_3[57749] = 32'b00000000000000001001001100010101;
assign LUT_3[57750] = 32'b00000000000000000100101000011100;
assign LUT_3[57751] = 32'b00000000000000001011010011111001;
assign LUT_3[57752] = 32'b00000000000000001010101100001000;
assign LUT_3[57753] = 32'b00000000000000010001010111100101;
assign LUT_3[57754] = 32'b00000000000000001100110011101100;
assign LUT_3[57755] = 32'b00000000000000010011011111001001;
assign LUT_3[57756] = 32'b00000000000000000111111001111110;
assign LUT_3[57757] = 32'b00000000000000001110100101011011;
assign LUT_3[57758] = 32'b00000000000000001010000001100010;
assign LUT_3[57759] = 32'b00000000000000010000101100111111;
assign LUT_3[57760] = 32'b00000000000000000011001110011111;
assign LUT_3[57761] = 32'b00000000000000001001111001111100;
assign LUT_3[57762] = 32'b00000000000000000101010110000011;
assign LUT_3[57763] = 32'b00000000000000001100000001100000;
assign LUT_3[57764] = 32'b00000000000000000000011100010101;
assign LUT_3[57765] = 32'b00000000000000000111000111110010;
assign LUT_3[57766] = 32'b00000000000000000010100011111001;
assign LUT_3[57767] = 32'b00000000000000001001001111010110;
assign LUT_3[57768] = 32'b00000000000000001000100111100101;
assign LUT_3[57769] = 32'b00000000000000001111010011000010;
assign LUT_3[57770] = 32'b00000000000000001010101111001001;
assign LUT_3[57771] = 32'b00000000000000010001011010100110;
assign LUT_3[57772] = 32'b00000000000000000101110101011011;
assign LUT_3[57773] = 32'b00000000000000001100100000111000;
assign LUT_3[57774] = 32'b00000000000000000111111100111111;
assign LUT_3[57775] = 32'b00000000000000001110101000011100;
assign LUT_3[57776] = 32'b00000000000000000110100001100010;
assign LUT_3[57777] = 32'b00000000000000001101001100111111;
assign LUT_3[57778] = 32'b00000000000000001000101001000110;
assign LUT_3[57779] = 32'b00000000000000001111010100100011;
assign LUT_3[57780] = 32'b00000000000000000011101111011000;
assign LUT_3[57781] = 32'b00000000000000001010011010110101;
assign LUT_3[57782] = 32'b00000000000000000101110110111100;
assign LUT_3[57783] = 32'b00000000000000001100100010011001;
assign LUT_3[57784] = 32'b00000000000000001011111010101000;
assign LUT_3[57785] = 32'b00000000000000010010100110000101;
assign LUT_3[57786] = 32'b00000000000000001110000010001100;
assign LUT_3[57787] = 32'b00000000000000010100101101101001;
assign LUT_3[57788] = 32'b00000000000000001001001000011110;
assign LUT_3[57789] = 32'b00000000000000001111110011111011;
assign LUT_3[57790] = 32'b00000000000000001011010000000010;
assign LUT_3[57791] = 32'b00000000000000010001111011011111;
assign LUT_3[57792] = 32'b00000000000000000001111000101010;
assign LUT_3[57793] = 32'b00000000000000001000100100000111;
assign LUT_3[57794] = 32'b00000000000000000100000000001110;
assign LUT_3[57795] = 32'b00000000000000001010101011101011;
assign LUT_3[57796] = 32'b11111111111111111111000110100000;
assign LUT_3[57797] = 32'b00000000000000000101110001111101;
assign LUT_3[57798] = 32'b00000000000000000001001110000100;
assign LUT_3[57799] = 32'b00000000000000000111111001100001;
assign LUT_3[57800] = 32'b00000000000000000111010001110000;
assign LUT_3[57801] = 32'b00000000000000001101111101001101;
assign LUT_3[57802] = 32'b00000000000000001001011001010100;
assign LUT_3[57803] = 32'b00000000000000010000000100110001;
assign LUT_3[57804] = 32'b00000000000000000100011111100110;
assign LUT_3[57805] = 32'b00000000000000001011001011000011;
assign LUT_3[57806] = 32'b00000000000000000110100111001010;
assign LUT_3[57807] = 32'b00000000000000001101010010100111;
assign LUT_3[57808] = 32'b00000000000000000101001011101101;
assign LUT_3[57809] = 32'b00000000000000001011110111001010;
assign LUT_3[57810] = 32'b00000000000000000111010011010001;
assign LUT_3[57811] = 32'b00000000000000001101111110101110;
assign LUT_3[57812] = 32'b00000000000000000010011001100011;
assign LUT_3[57813] = 32'b00000000000000001001000101000000;
assign LUT_3[57814] = 32'b00000000000000000100100001000111;
assign LUT_3[57815] = 32'b00000000000000001011001100100100;
assign LUT_3[57816] = 32'b00000000000000001010100100110011;
assign LUT_3[57817] = 32'b00000000000000010001010000010000;
assign LUT_3[57818] = 32'b00000000000000001100101100010111;
assign LUT_3[57819] = 32'b00000000000000010011010111110100;
assign LUT_3[57820] = 32'b00000000000000000111110010101001;
assign LUT_3[57821] = 32'b00000000000000001110011110000110;
assign LUT_3[57822] = 32'b00000000000000001001111010001101;
assign LUT_3[57823] = 32'b00000000000000010000100101101010;
assign LUT_3[57824] = 32'b00000000000000000011000111001010;
assign LUT_3[57825] = 32'b00000000000000001001110010100111;
assign LUT_3[57826] = 32'b00000000000000000101001110101110;
assign LUT_3[57827] = 32'b00000000000000001011111010001011;
assign LUT_3[57828] = 32'b00000000000000000000010101000000;
assign LUT_3[57829] = 32'b00000000000000000111000000011101;
assign LUT_3[57830] = 32'b00000000000000000010011100100100;
assign LUT_3[57831] = 32'b00000000000000001001001000000001;
assign LUT_3[57832] = 32'b00000000000000001000100000010000;
assign LUT_3[57833] = 32'b00000000000000001111001011101101;
assign LUT_3[57834] = 32'b00000000000000001010100111110100;
assign LUT_3[57835] = 32'b00000000000000010001010011010001;
assign LUT_3[57836] = 32'b00000000000000000101101110000110;
assign LUT_3[57837] = 32'b00000000000000001100011001100011;
assign LUT_3[57838] = 32'b00000000000000000111110101101010;
assign LUT_3[57839] = 32'b00000000000000001110100001000111;
assign LUT_3[57840] = 32'b00000000000000000110011010001101;
assign LUT_3[57841] = 32'b00000000000000001101000101101010;
assign LUT_3[57842] = 32'b00000000000000001000100001110001;
assign LUT_3[57843] = 32'b00000000000000001111001101001110;
assign LUT_3[57844] = 32'b00000000000000000011101000000011;
assign LUT_3[57845] = 32'b00000000000000001010010011100000;
assign LUT_3[57846] = 32'b00000000000000000101101111100111;
assign LUT_3[57847] = 32'b00000000000000001100011011000100;
assign LUT_3[57848] = 32'b00000000000000001011110011010011;
assign LUT_3[57849] = 32'b00000000000000010010011110110000;
assign LUT_3[57850] = 32'b00000000000000001101111010110111;
assign LUT_3[57851] = 32'b00000000000000010100100110010100;
assign LUT_3[57852] = 32'b00000000000000001001000001001001;
assign LUT_3[57853] = 32'b00000000000000001111101100100110;
assign LUT_3[57854] = 32'b00000000000000001011001000101101;
assign LUT_3[57855] = 32'b00000000000000010001110100001010;
assign LUT_3[57856] = 32'b00000000000000000110111010101100;
assign LUT_3[57857] = 32'b00000000000000001101100110001001;
assign LUT_3[57858] = 32'b00000000000000001001000010010000;
assign LUT_3[57859] = 32'b00000000000000001111101101101101;
assign LUT_3[57860] = 32'b00000000000000000100001000100010;
assign LUT_3[57861] = 32'b00000000000000001010110011111111;
assign LUT_3[57862] = 32'b00000000000000000110010000000110;
assign LUT_3[57863] = 32'b00000000000000001100111011100011;
assign LUT_3[57864] = 32'b00000000000000001100010011110010;
assign LUT_3[57865] = 32'b00000000000000010010111111001111;
assign LUT_3[57866] = 32'b00000000000000001110011011010110;
assign LUT_3[57867] = 32'b00000000000000010101000110110011;
assign LUT_3[57868] = 32'b00000000000000001001100001101000;
assign LUT_3[57869] = 32'b00000000000000010000001101000101;
assign LUT_3[57870] = 32'b00000000000000001011101001001100;
assign LUT_3[57871] = 32'b00000000000000010010010100101001;
assign LUT_3[57872] = 32'b00000000000000001010001101101111;
assign LUT_3[57873] = 32'b00000000000000010000111001001100;
assign LUT_3[57874] = 32'b00000000000000001100010101010011;
assign LUT_3[57875] = 32'b00000000000000010011000000110000;
assign LUT_3[57876] = 32'b00000000000000000111011011100101;
assign LUT_3[57877] = 32'b00000000000000001110000111000010;
assign LUT_3[57878] = 32'b00000000000000001001100011001001;
assign LUT_3[57879] = 32'b00000000000000010000001110100110;
assign LUT_3[57880] = 32'b00000000000000001111100110110101;
assign LUT_3[57881] = 32'b00000000000000010110010010010010;
assign LUT_3[57882] = 32'b00000000000000010001101110011001;
assign LUT_3[57883] = 32'b00000000000000011000011001110110;
assign LUT_3[57884] = 32'b00000000000000001100110100101011;
assign LUT_3[57885] = 32'b00000000000000010011100000001000;
assign LUT_3[57886] = 32'b00000000000000001110111100001111;
assign LUT_3[57887] = 32'b00000000000000010101100111101100;
assign LUT_3[57888] = 32'b00000000000000001000001001001100;
assign LUT_3[57889] = 32'b00000000000000001110110100101001;
assign LUT_3[57890] = 32'b00000000000000001010010000110000;
assign LUT_3[57891] = 32'b00000000000000010000111100001101;
assign LUT_3[57892] = 32'b00000000000000000101010111000010;
assign LUT_3[57893] = 32'b00000000000000001100000010011111;
assign LUT_3[57894] = 32'b00000000000000000111011110100110;
assign LUT_3[57895] = 32'b00000000000000001110001010000011;
assign LUT_3[57896] = 32'b00000000000000001101100010010010;
assign LUT_3[57897] = 32'b00000000000000010100001101101111;
assign LUT_3[57898] = 32'b00000000000000001111101001110110;
assign LUT_3[57899] = 32'b00000000000000010110010101010011;
assign LUT_3[57900] = 32'b00000000000000001010110000001000;
assign LUT_3[57901] = 32'b00000000000000010001011011100101;
assign LUT_3[57902] = 32'b00000000000000001100110111101100;
assign LUT_3[57903] = 32'b00000000000000010011100011001001;
assign LUT_3[57904] = 32'b00000000000000001011011100001111;
assign LUT_3[57905] = 32'b00000000000000010010000111101100;
assign LUT_3[57906] = 32'b00000000000000001101100011110011;
assign LUT_3[57907] = 32'b00000000000000010100001111010000;
assign LUT_3[57908] = 32'b00000000000000001000101010000101;
assign LUT_3[57909] = 32'b00000000000000001111010101100010;
assign LUT_3[57910] = 32'b00000000000000001010110001101001;
assign LUT_3[57911] = 32'b00000000000000010001011101000110;
assign LUT_3[57912] = 32'b00000000000000010000110101010101;
assign LUT_3[57913] = 32'b00000000000000010111100000110010;
assign LUT_3[57914] = 32'b00000000000000010010111100111001;
assign LUT_3[57915] = 32'b00000000000000011001101000010110;
assign LUT_3[57916] = 32'b00000000000000001110000011001011;
assign LUT_3[57917] = 32'b00000000000000010100101110101000;
assign LUT_3[57918] = 32'b00000000000000010000001010101111;
assign LUT_3[57919] = 32'b00000000000000010110110110001100;
assign LUT_3[57920] = 32'b00000000000000000110110011010111;
assign LUT_3[57921] = 32'b00000000000000001101011110110100;
assign LUT_3[57922] = 32'b00000000000000001000111010111011;
assign LUT_3[57923] = 32'b00000000000000001111100110011000;
assign LUT_3[57924] = 32'b00000000000000000100000001001101;
assign LUT_3[57925] = 32'b00000000000000001010101100101010;
assign LUT_3[57926] = 32'b00000000000000000110001000110001;
assign LUT_3[57927] = 32'b00000000000000001100110100001110;
assign LUT_3[57928] = 32'b00000000000000001100001100011101;
assign LUT_3[57929] = 32'b00000000000000010010110111111010;
assign LUT_3[57930] = 32'b00000000000000001110010100000001;
assign LUT_3[57931] = 32'b00000000000000010100111111011110;
assign LUT_3[57932] = 32'b00000000000000001001011010010011;
assign LUT_3[57933] = 32'b00000000000000010000000101110000;
assign LUT_3[57934] = 32'b00000000000000001011100001110111;
assign LUT_3[57935] = 32'b00000000000000010010001101010100;
assign LUT_3[57936] = 32'b00000000000000001010000110011010;
assign LUT_3[57937] = 32'b00000000000000010000110001110111;
assign LUT_3[57938] = 32'b00000000000000001100001101111110;
assign LUT_3[57939] = 32'b00000000000000010010111001011011;
assign LUT_3[57940] = 32'b00000000000000000111010100010000;
assign LUT_3[57941] = 32'b00000000000000001101111111101101;
assign LUT_3[57942] = 32'b00000000000000001001011011110100;
assign LUT_3[57943] = 32'b00000000000000010000000111010001;
assign LUT_3[57944] = 32'b00000000000000001111011111100000;
assign LUT_3[57945] = 32'b00000000000000010110001010111101;
assign LUT_3[57946] = 32'b00000000000000010001100111000100;
assign LUT_3[57947] = 32'b00000000000000011000010010100001;
assign LUT_3[57948] = 32'b00000000000000001100101101010110;
assign LUT_3[57949] = 32'b00000000000000010011011000110011;
assign LUT_3[57950] = 32'b00000000000000001110110100111010;
assign LUT_3[57951] = 32'b00000000000000010101100000010111;
assign LUT_3[57952] = 32'b00000000000000001000000001110111;
assign LUT_3[57953] = 32'b00000000000000001110101101010100;
assign LUT_3[57954] = 32'b00000000000000001010001001011011;
assign LUT_3[57955] = 32'b00000000000000010000110100111000;
assign LUT_3[57956] = 32'b00000000000000000101001111101101;
assign LUT_3[57957] = 32'b00000000000000001011111011001010;
assign LUT_3[57958] = 32'b00000000000000000111010111010001;
assign LUT_3[57959] = 32'b00000000000000001110000010101110;
assign LUT_3[57960] = 32'b00000000000000001101011010111101;
assign LUT_3[57961] = 32'b00000000000000010100000110011010;
assign LUT_3[57962] = 32'b00000000000000001111100010100001;
assign LUT_3[57963] = 32'b00000000000000010110001101111110;
assign LUT_3[57964] = 32'b00000000000000001010101000110011;
assign LUT_3[57965] = 32'b00000000000000010001010100010000;
assign LUT_3[57966] = 32'b00000000000000001100110000010111;
assign LUT_3[57967] = 32'b00000000000000010011011011110100;
assign LUT_3[57968] = 32'b00000000000000001011010100111010;
assign LUT_3[57969] = 32'b00000000000000010010000000010111;
assign LUT_3[57970] = 32'b00000000000000001101011100011110;
assign LUT_3[57971] = 32'b00000000000000010100000111111011;
assign LUT_3[57972] = 32'b00000000000000001000100010110000;
assign LUT_3[57973] = 32'b00000000000000001111001110001101;
assign LUT_3[57974] = 32'b00000000000000001010101010010100;
assign LUT_3[57975] = 32'b00000000000000010001010101110001;
assign LUT_3[57976] = 32'b00000000000000010000101110000000;
assign LUT_3[57977] = 32'b00000000000000010111011001011101;
assign LUT_3[57978] = 32'b00000000000000010010110101100100;
assign LUT_3[57979] = 32'b00000000000000011001100001000001;
assign LUT_3[57980] = 32'b00000000000000001101111011110110;
assign LUT_3[57981] = 32'b00000000000000010100100111010011;
assign LUT_3[57982] = 32'b00000000000000010000000011011010;
assign LUT_3[57983] = 32'b00000000000000010110101110110111;
assign LUT_3[57984] = 32'b00000000000000001001000101101010;
assign LUT_3[57985] = 32'b00000000000000001111110001000111;
assign LUT_3[57986] = 32'b00000000000000001011001101001110;
assign LUT_3[57987] = 32'b00000000000000010001111000101011;
assign LUT_3[57988] = 32'b00000000000000000110010011100000;
assign LUT_3[57989] = 32'b00000000000000001100111110111101;
assign LUT_3[57990] = 32'b00000000000000001000011011000100;
assign LUT_3[57991] = 32'b00000000000000001111000110100001;
assign LUT_3[57992] = 32'b00000000000000001110011110110000;
assign LUT_3[57993] = 32'b00000000000000010101001010001101;
assign LUT_3[57994] = 32'b00000000000000010000100110010100;
assign LUT_3[57995] = 32'b00000000000000010111010001110001;
assign LUT_3[57996] = 32'b00000000000000001011101100100110;
assign LUT_3[57997] = 32'b00000000000000010010011000000011;
assign LUT_3[57998] = 32'b00000000000000001101110100001010;
assign LUT_3[57999] = 32'b00000000000000010100011111100111;
assign LUT_3[58000] = 32'b00000000000000001100011000101101;
assign LUT_3[58001] = 32'b00000000000000010011000100001010;
assign LUT_3[58002] = 32'b00000000000000001110100000010001;
assign LUT_3[58003] = 32'b00000000000000010101001011101110;
assign LUT_3[58004] = 32'b00000000000000001001100110100011;
assign LUT_3[58005] = 32'b00000000000000010000010010000000;
assign LUT_3[58006] = 32'b00000000000000001011101110000111;
assign LUT_3[58007] = 32'b00000000000000010010011001100100;
assign LUT_3[58008] = 32'b00000000000000010001110001110011;
assign LUT_3[58009] = 32'b00000000000000011000011101010000;
assign LUT_3[58010] = 32'b00000000000000010011111001010111;
assign LUT_3[58011] = 32'b00000000000000011010100100110100;
assign LUT_3[58012] = 32'b00000000000000001110111111101001;
assign LUT_3[58013] = 32'b00000000000000010101101011000110;
assign LUT_3[58014] = 32'b00000000000000010001000111001101;
assign LUT_3[58015] = 32'b00000000000000010111110010101010;
assign LUT_3[58016] = 32'b00000000000000001010010100001010;
assign LUT_3[58017] = 32'b00000000000000010000111111100111;
assign LUT_3[58018] = 32'b00000000000000001100011011101110;
assign LUT_3[58019] = 32'b00000000000000010011000111001011;
assign LUT_3[58020] = 32'b00000000000000000111100010000000;
assign LUT_3[58021] = 32'b00000000000000001110001101011101;
assign LUT_3[58022] = 32'b00000000000000001001101001100100;
assign LUT_3[58023] = 32'b00000000000000010000010101000001;
assign LUT_3[58024] = 32'b00000000000000001111101101010000;
assign LUT_3[58025] = 32'b00000000000000010110011000101101;
assign LUT_3[58026] = 32'b00000000000000010001110100110100;
assign LUT_3[58027] = 32'b00000000000000011000100000010001;
assign LUT_3[58028] = 32'b00000000000000001100111011000110;
assign LUT_3[58029] = 32'b00000000000000010011100110100011;
assign LUT_3[58030] = 32'b00000000000000001111000010101010;
assign LUT_3[58031] = 32'b00000000000000010101101110000111;
assign LUT_3[58032] = 32'b00000000000000001101100111001101;
assign LUT_3[58033] = 32'b00000000000000010100010010101010;
assign LUT_3[58034] = 32'b00000000000000001111101110110001;
assign LUT_3[58035] = 32'b00000000000000010110011010001110;
assign LUT_3[58036] = 32'b00000000000000001010110101000011;
assign LUT_3[58037] = 32'b00000000000000010001100000100000;
assign LUT_3[58038] = 32'b00000000000000001100111100100111;
assign LUT_3[58039] = 32'b00000000000000010011101000000100;
assign LUT_3[58040] = 32'b00000000000000010011000000010011;
assign LUT_3[58041] = 32'b00000000000000011001101011110000;
assign LUT_3[58042] = 32'b00000000000000010101000111110111;
assign LUT_3[58043] = 32'b00000000000000011011110011010100;
assign LUT_3[58044] = 32'b00000000000000010000001110001001;
assign LUT_3[58045] = 32'b00000000000000010110111001100110;
assign LUT_3[58046] = 32'b00000000000000010010010101101101;
assign LUT_3[58047] = 32'b00000000000000011001000001001010;
assign LUT_3[58048] = 32'b00000000000000001000111110010101;
assign LUT_3[58049] = 32'b00000000000000001111101001110010;
assign LUT_3[58050] = 32'b00000000000000001011000101111001;
assign LUT_3[58051] = 32'b00000000000000010001110001010110;
assign LUT_3[58052] = 32'b00000000000000000110001100001011;
assign LUT_3[58053] = 32'b00000000000000001100110111101000;
assign LUT_3[58054] = 32'b00000000000000001000010011101111;
assign LUT_3[58055] = 32'b00000000000000001110111111001100;
assign LUT_3[58056] = 32'b00000000000000001110010111011011;
assign LUT_3[58057] = 32'b00000000000000010101000010111000;
assign LUT_3[58058] = 32'b00000000000000010000011110111111;
assign LUT_3[58059] = 32'b00000000000000010111001010011100;
assign LUT_3[58060] = 32'b00000000000000001011100101010001;
assign LUT_3[58061] = 32'b00000000000000010010010000101110;
assign LUT_3[58062] = 32'b00000000000000001101101100110101;
assign LUT_3[58063] = 32'b00000000000000010100011000010010;
assign LUT_3[58064] = 32'b00000000000000001100010001011000;
assign LUT_3[58065] = 32'b00000000000000010010111100110101;
assign LUT_3[58066] = 32'b00000000000000001110011000111100;
assign LUT_3[58067] = 32'b00000000000000010101000100011001;
assign LUT_3[58068] = 32'b00000000000000001001011111001110;
assign LUT_3[58069] = 32'b00000000000000010000001010101011;
assign LUT_3[58070] = 32'b00000000000000001011100110110010;
assign LUT_3[58071] = 32'b00000000000000010010010010001111;
assign LUT_3[58072] = 32'b00000000000000010001101010011110;
assign LUT_3[58073] = 32'b00000000000000011000010101111011;
assign LUT_3[58074] = 32'b00000000000000010011110010000010;
assign LUT_3[58075] = 32'b00000000000000011010011101011111;
assign LUT_3[58076] = 32'b00000000000000001110111000010100;
assign LUT_3[58077] = 32'b00000000000000010101100011110001;
assign LUT_3[58078] = 32'b00000000000000010000111111111000;
assign LUT_3[58079] = 32'b00000000000000010111101011010101;
assign LUT_3[58080] = 32'b00000000000000001010001100110101;
assign LUT_3[58081] = 32'b00000000000000010000111000010010;
assign LUT_3[58082] = 32'b00000000000000001100010100011001;
assign LUT_3[58083] = 32'b00000000000000010010111111110110;
assign LUT_3[58084] = 32'b00000000000000000111011010101011;
assign LUT_3[58085] = 32'b00000000000000001110000110001000;
assign LUT_3[58086] = 32'b00000000000000001001100010001111;
assign LUT_3[58087] = 32'b00000000000000010000001101101100;
assign LUT_3[58088] = 32'b00000000000000001111100101111011;
assign LUT_3[58089] = 32'b00000000000000010110010001011000;
assign LUT_3[58090] = 32'b00000000000000010001101101011111;
assign LUT_3[58091] = 32'b00000000000000011000011000111100;
assign LUT_3[58092] = 32'b00000000000000001100110011110001;
assign LUT_3[58093] = 32'b00000000000000010011011111001110;
assign LUT_3[58094] = 32'b00000000000000001110111011010101;
assign LUT_3[58095] = 32'b00000000000000010101100110110010;
assign LUT_3[58096] = 32'b00000000000000001101011111111000;
assign LUT_3[58097] = 32'b00000000000000010100001011010101;
assign LUT_3[58098] = 32'b00000000000000001111100111011100;
assign LUT_3[58099] = 32'b00000000000000010110010010111001;
assign LUT_3[58100] = 32'b00000000000000001010101101101110;
assign LUT_3[58101] = 32'b00000000000000010001011001001011;
assign LUT_3[58102] = 32'b00000000000000001100110101010010;
assign LUT_3[58103] = 32'b00000000000000010011100000101111;
assign LUT_3[58104] = 32'b00000000000000010010111000111110;
assign LUT_3[58105] = 32'b00000000000000011001100100011011;
assign LUT_3[58106] = 32'b00000000000000010101000000100010;
assign LUT_3[58107] = 32'b00000000000000011011101011111111;
assign LUT_3[58108] = 32'b00000000000000010000000110110100;
assign LUT_3[58109] = 32'b00000000000000010110110010010001;
assign LUT_3[58110] = 32'b00000000000000010010001110011000;
assign LUT_3[58111] = 32'b00000000000000011000111001110101;
assign LUT_3[58112] = 32'b00000000000000000011001010001101;
assign LUT_3[58113] = 32'b00000000000000001001110101101010;
assign LUT_3[58114] = 32'b00000000000000000101010001110001;
assign LUT_3[58115] = 32'b00000000000000001011111101001110;
assign LUT_3[58116] = 32'b00000000000000000000011000000011;
assign LUT_3[58117] = 32'b00000000000000000111000011100000;
assign LUT_3[58118] = 32'b00000000000000000010011111100111;
assign LUT_3[58119] = 32'b00000000000000001001001011000100;
assign LUT_3[58120] = 32'b00000000000000001000100011010011;
assign LUT_3[58121] = 32'b00000000000000001111001110110000;
assign LUT_3[58122] = 32'b00000000000000001010101010110111;
assign LUT_3[58123] = 32'b00000000000000010001010110010100;
assign LUT_3[58124] = 32'b00000000000000000101110001001001;
assign LUT_3[58125] = 32'b00000000000000001100011100100110;
assign LUT_3[58126] = 32'b00000000000000000111111000101101;
assign LUT_3[58127] = 32'b00000000000000001110100100001010;
assign LUT_3[58128] = 32'b00000000000000000110011101010000;
assign LUT_3[58129] = 32'b00000000000000001101001000101101;
assign LUT_3[58130] = 32'b00000000000000001000100100110100;
assign LUT_3[58131] = 32'b00000000000000001111010000010001;
assign LUT_3[58132] = 32'b00000000000000000011101011000110;
assign LUT_3[58133] = 32'b00000000000000001010010110100011;
assign LUT_3[58134] = 32'b00000000000000000101110010101010;
assign LUT_3[58135] = 32'b00000000000000001100011110000111;
assign LUT_3[58136] = 32'b00000000000000001011110110010110;
assign LUT_3[58137] = 32'b00000000000000010010100001110011;
assign LUT_3[58138] = 32'b00000000000000001101111101111010;
assign LUT_3[58139] = 32'b00000000000000010100101001010111;
assign LUT_3[58140] = 32'b00000000000000001001000100001100;
assign LUT_3[58141] = 32'b00000000000000001111101111101001;
assign LUT_3[58142] = 32'b00000000000000001011001011110000;
assign LUT_3[58143] = 32'b00000000000000010001110111001101;
assign LUT_3[58144] = 32'b00000000000000000100011000101101;
assign LUT_3[58145] = 32'b00000000000000001011000100001010;
assign LUT_3[58146] = 32'b00000000000000000110100000010001;
assign LUT_3[58147] = 32'b00000000000000001101001011101110;
assign LUT_3[58148] = 32'b00000000000000000001100110100011;
assign LUT_3[58149] = 32'b00000000000000001000010010000000;
assign LUT_3[58150] = 32'b00000000000000000011101110000111;
assign LUT_3[58151] = 32'b00000000000000001010011001100100;
assign LUT_3[58152] = 32'b00000000000000001001110001110011;
assign LUT_3[58153] = 32'b00000000000000010000011101010000;
assign LUT_3[58154] = 32'b00000000000000001011111001010111;
assign LUT_3[58155] = 32'b00000000000000010010100100110100;
assign LUT_3[58156] = 32'b00000000000000000110111111101001;
assign LUT_3[58157] = 32'b00000000000000001101101011000110;
assign LUT_3[58158] = 32'b00000000000000001001000111001101;
assign LUT_3[58159] = 32'b00000000000000001111110010101010;
assign LUT_3[58160] = 32'b00000000000000000111101011110000;
assign LUT_3[58161] = 32'b00000000000000001110010111001101;
assign LUT_3[58162] = 32'b00000000000000001001110011010100;
assign LUT_3[58163] = 32'b00000000000000010000011110110001;
assign LUT_3[58164] = 32'b00000000000000000100111001100110;
assign LUT_3[58165] = 32'b00000000000000001011100101000011;
assign LUT_3[58166] = 32'b00000000000000000111000001001010;
assign LUT_3[58167] = 32'b00000000000000001101101100100111;
assign LUT_3[58168] = 32'b00000000000000001101000100110110;
assign LUT_3[58169] = 32'b00000000000000010011110000010011;
assign LUT_3[58170] = 32'b00000000000000001111001100011010;
assign LUT_3[58171] = 32'b00000000000000010101110111110111;
assign LUT_3[58172] = 32'b00000000000000001010010010101100;
assign LUT_3[58173] = 32'b00000000000000010000111110001001;
assign LUT_3[58174] = 32'b00000000000000001100011010010000;
assign LUT_3[58175] = 32'b00000000000000010011000101101101;
assign LUT_3[58176] = 32'b00000000000000000011000010111000;
assign LUT_3[58177] = 32'b00000000000000001001101110010101;
assign LUT_3[58178] = 32'b00000000000000000101001010011100;
assign LUT_3[58179] = 32'b00000000000000001011110101111001;
assign LUT_3[58180] = 32'b00000000000000000000010000101110;
assign LUT_3[58181] = 32'b00000000000000000110111100001011;
assign LUT_3[58182] = 32'b00000000000000000010011000010010;
assign LUT_3[58183] = 32'b00000000000000001001000011101111;
assign LUT_3[58184] = 32'b00000000000000001000011011111110;
assign LUT_3[58185] = 32'b00000000000000001111000111011011;
assign LUT_3[58186] = 32'b00000000000000001010100011100010;
assign LUT_3[58187] = 32'b00000000000000010001001110111111;
assign LUT_3[58188] = 32'b00000000000000000101101001110100;
assign LUT_3[58189] = 32'b00000000000000001100010101010001;
assign LUT_3[58190] = 32'b00000000000000000111110001011000;
assign LUT_3[58191] = 32'b00000000000000001110011100110101;
assign LUT_3[58192] = 32'b00000000000000000110010101111011;
assign LUT_3[58193] = 32'b00000000000000001101000001011000;
assign LUT_3[58194] = 32'b00000000000000001000011101011111;
assign LUT_3[58195] = 32'b00000000000000001111001000111100;
assign LUT_3[58196] = 32'b00000000000000000011100011110001;
assign LUT_3[58197] = 32'b00000000000000001010001111001110;
assign LUT_3[58198] = 32'b00000000000000000101101011010101;
assign LUT_3[58199] = 32'b00000000000000001100010110110010;
assign LUT_3[58200] = 32'b00000000000000001011101111000001;
assign LUT_3[58201] = 32'b00000000000000010010011010011110;
assign LUT_3[58202] = 32'b00000000000000001101110110100101;
assign LUT_3[58203] = 32'b00000000000000010100100010000010;
assign LUT_3[58204] = 32'b00000000000000001000111100110111;
assign LUT_3[58205] = 32'b00000000000000001111101000010100;
assign LUT_3[58206] = 32'b00000000000000001011000100011011;
assign LUT_3[58207] = 32'b00000000000000010001101111111000;
assign LUT_3[58208] = 32'b00000000000000000100010001011000;
assign LUT_3[58209] = 32'b00000000000000001010111100110101;
assign LUT_3[58210] = 32'b00000000000000000110011000111100;
assign LUT_3[58211] = 32'b00000000000000001101000100011001;
assign LUT_3[58212] = 32'b00000000000000000001011111001110;
assign LUT_3[58213] = 32'b00000000000000001000001010101011;
assign LUT_3[58214] = 32'b00000000000000000011100110110010;
assign LUT_3[58215] = 32'b00000000000000001010010010001111;
assign LUT_3[58216] = 32'b00000000000000001001101010011110;
assign LUT_3[58217] = 32'b00000000000000010000010101111011;
assign LUT_3[58218] = 32'b00000000000000001011110010000010;
assign LUT_3[58219] = 32'b00000000000000010010011101011111;
assign LUT_3[58220] = 32'b00000000000000000110111000010100;
assign LUT_3[58221] = 32'b00000000000000001101100011110001;
assign LUT_3[58222] = 32'b00000000000000001000111111111000;
assign LUT_3[58223] = 32'b00000000000000001111101011010101;
assign LUT_3[58224] = 32'b00000000000000000111100100011011;
assign LUT_3[58225] = 32'b00000000000000001110001111111000;
assign LUT_3[58226] = 32'b00000000000000001001101011111111;
assign LUT_3[58227] = 32'b00000000000000010000010111011100;
assign LUT_3[58228] = 32'b00000000000000000100110010010001;
assign LUT_3[58229] = 32'b00000000000000001011011101101110;
assign LUT_3[58230] = 32'b00000000000000000110111001110101;
assign LUT_3[58231] = 32'b00000000000000001101100101010010;
assign LUT_3[58232] = 32'b00000000000000001100111101100001;
assign LUT_3[58233] = 32'b00000000000000010011101000111110;
assign LUT_3[58234] = 32'b00000000000000001111000101000101;
assign LUT_3[58235] = 32'b00000000000000010101110000100010;
assign LUT_3[58236] = 32'b00000000000000001010001011010111;
assign LUT_3[58237] = 32'b00000000000000010000110110110100;
assign LUT_3[58238] = 32'b00000000000000001100010010111011;
assign LUT_3[58239] = 32'b00000000000000010010111110011000;
assign LUT_3[58240] = 32'b00000000000000000101010101001011;
assign LUT_3[58241] = 32'b00000000000000001100000000101000;
assign LUT_3[58242] = 32'b00000000000000000111011100101111;
assign LUT_3[58243] = 32'b00000000000000001110001000001100;
assign LUT_3[58244] = 32'b00000000000000000010100011000001;
assign LUT_3[58245] = 32'b00000000000000001001001110011110;
assign LUT_3[58246] = 32'b00000000000000000100101010100101;
assign LUT_3[58247] = 32'b00000000000000001011010110000010;
assign LUT_3[58248] = 32'b00000000000000001010101110010001;
assign LUT_3[58249] = 32'b00000000000000010001011001101110;
assign LUT_3[58250] = 32'b00000000000000001100110101110101;
assign LUT_3[58251] = 32'b00000000000000010011100001010010;
assign LUT_3[58252] = 32'b00000000000000000111111100000111;
assign LUT_3[58253] = 32'b00000000000000001110100111100100;
assign LUT_3[58254] = 32'b00000000000000001010000011101011;
assign LUT_3[58255] = 32'b00000000000000010000101111001000;
assign LUT_3[58256] = 32'b00000000000000001000101000001110;
assign LUT_3[58257] = 32'b00000000000000001111010011101011;
assign LUT_3[58258] = 32'b00000000000000001010101111110010;
assign LUT_3[58259] = 32'b00000000000000010001011011001111;
assign LUT_3[58260] = 32'b00000000000000000101110110000100;
assign LUT_3[58261] = 32'b00000000000000001100100001100001;
assign LUT_3[58262] = 32'b00000000000000000111111101101000;
assign LUT_3[58263] = 32'b00000000000000001110101001000101;
assign LUT_3[58264] = 32'b00000000000000001110000001010100;
assign LUT_3[58265] = 32'b00000000000000010100101100110001;
assign LUT_3[58266] = 32'b00000000000000010000001000111000;
assign LUT_3[58267] = 32'b00000000000000010110110100010101;
assign LUT_3[58268] = 32'b00000000000000001011001111001010;
assign LUT_3[58269] = 32'b00000000000000010001111010100111;
assign LUT_3[58270] = 32'b00000000000000001101010110101110;
assign LUT_3[58271] = 32'b00000000000000010100000010001011;
assign LUT_3[58272] = 32'b00000000000000000110100011101011;
assign LUT_3[58273] = 32'b00000000000000001101001111001000;
assign LUT_3[58274] = 32'b00000000000000001000101011001111;
assign LUT_3[58275] = 32'b00000000000000001111010110101100;
assign LUT_3[58276] = 32'b00000000000000000011110001100001;
assign LUT_3[58277] = 32'b00000000000000001010011100111110;
assign LUT_3[58278] = 32'b00000000000000000101111001000101;
assign LUT_3[58279] = 32'b00000000000000001100100100100010;
assign LUT_3[58280] = 32'b00000000000000001011111100110001;
assign LUT_3[58281] = 32'b00000000000000010010101000001110;
assign LUT_3[58282] = 32'b00000000000000001110000100010101;
assign LUT_3[58283] = 32'b00000000000000010100101111110010;
assign LUT_3[58284] = 32'b00000000000000001001001010100111;
assign LUT_3[58285] = 32'b00000000000000001111110110000100;
assign LUT_3[58286] = 32'b00000000000000001011010010001011;
assign LUT_3[58287] = 32'b00000000000000010001111101101000;
assign LUT_3[58288] = 32'b00000000000000001001110110101110;
assign LUT_3[58289] = 32'b00000000000000010000100010001011;
assign LUT_3[58290] = 32'b00000000000000001011111110010010;
assign LUT_3[58291] = 32'b00000000000000010010101001101111;
assign LUT_3[58292] = 32'b00000000000000000111000100100100;
assign LUT_3[58293] = 32'b00000000000000001101110000000001;
assign LUT_3[58294] = 32'b00000000000000001001001100001000;
assign LUT_3[58295] = 32'b00000000000000001111110111100101;
assign LUT_3[58296] = 32'b00000000000000001111001111110100;
assign LUT_3[58297] = 32'b00000000000000010101111011010001;
assign LUT_3[58298] = 32'b00000000000000010001010111011000;
assign LUT_3[58299] = 32'b00000000000000011000000010110101;
assign LUT_3[58300] = 32'b00000000000000001100011101101010;
assign LUT_3[58301] = 32'b00000000000000010011001001000111;
assign LUT_3[58302] = 32'b00000000000000001110100101001110;
assign LUT_3[58303] = 32'b00000000000000010101010000101011;
assign LUT_3[58304] = 32'b00000000000000000101001101110110;
assign LUT_3[58305] = 32'b00000000000000001011111001010011;
assign LUT_3[58306] = 32'b00000000000000000111010101011010;
assign LUT_3[58307] = 32'b00000000000000001110000000110111;
assign LUT_3[58308] = 32'b00000000000000000010011011101100;
assign LUT_3[58309] = 32'b00000000000000001001000111001001;
assign LUT_3[58310] = 32'b00000000000000000100100011010000;
assign LUT_3[58311] = 32'b00000000000000001011001110101101;
assign LUT_3[58312] = 32'b00000000000000001010100110111100;
assign LUT_3[58313] = 32'b00000000000000010001010010011001;
assign LUT_3[58314] = 32'b00000000000000001100101110100000;
assign LUT_3[58315] = 32'b00000000000000010011011001111101;
assign LUT_3[58316] = 32'b00000000000000000111110100110010;
assign LUT_3[58317] = 32'b00000000000000001110100000001111;
assign LUT_3[58318] = 32'b00000000000000001001111100010110;
assign LUT_3[58319] = 32'b00000000000000010000100111110011;
assign LUT_3[58320] = 32'b00000000000000001000100000111001;
assign LUT_3[58321] = 32'b00000000000000001111001100010110;
assign LUT_3[58322] = 32'b00000000000000001010101000011101;
assign LUT_3[58323] = 32'b00000000000000010001010011111010;
assign LUT_3[58324] = 32'b00000000000000000101101110101111;
assign LUT_3[58325] = 32'b00000000000000001100011010001100;
assign LUT_3[58326] = 32'b00000000000000000111110110010011;
assign LUT_3[58327] = 32'b00000000000000001110100001110000;
assign LUT_3[58328] = 32'b00000000000000001101111001111111;
assign LUT_3[58329] = 32'b00000000000000010100100101011100;
assign LUT_3[58330] = 32'b00000000000000010000000001100011;
assign LUT_3[58331] = 32'b00000000000000010110101101000000;
assign LUT_3[58332] = 32'b00000000000000001011000111110101;
assign LUT_3[58333] = 32'b00000000000000010001110011010010;
assign LUT_3[58334] = 32'b00000000000000001101001111011001;
assign LUT_3[58335] = 32'b00000000000000010011111010110110;
assign LUT_3[58336] = 32'b00000000000000000110011100010110;
assign LUT_3[58337] = 32'b00000000000000001101000111110011;
assign LUT_3[58338] = 32'b00000000000000001000100011111010;
assign LUT_3[58339] = 32'b00000000000000001111001111010111;
assign LUT_3[58340] = 32'b00000000000000000011101010001100;
assign LUT_3[58341] = 32'b00000000000000001010010101101001;
assign LUT_3[58342] = 32'b00000000000000000101110001110000;
assign LUT_3[58343] = 32'b00000000000000001100011101001101;
assign LUT_3[58344] = 32'b00000000000000001011110101011100;
assign LUT_3[58345] = 32'b00000000000000010010100000111001;
assign LUT_3[58346] = 32'b00000000000000001101111101000000;
assign LUT_3[58347] = 32'b00000000000000010100101000011101;
assign LUT_3[58348] = 32'b00000000000000001001000011010010;
assign LUT_3[58349] = 32'b00000000000000001111101110101111;
assign LUT_3[58350] = 32'b00000000000000001011001010110110;
assign LUT_3[58351] = 32'b00000000000000010001110110010011;
assign LUT_3[58352] = 32'b00000000000000001001101111011001;
assign LUT_3[58353] = 32'b00000000000000010000011010110110;
assign LUT_3[58354] = 32'b00000000000000001011110110111101;
assign LUT_3[58355] = 32'b00000000000000010010100010011010;
assign LUT_3[58356] = 32'b00000000000000000110111101001111;
assign LUT_3[58357] = 32'b00000000000000001101101000101100;
assign LUT_3[58358] = 32'b00000000000000001001000100110011;
assign LUT_3[58359] = 32'b00000000000000001111110000010000;
assign LUT_3[58360] = 32'b00000000000000001111001000011111;
assign LUT_3[58361] = 32'b00000000000000010101110011111100;
assign LUT_3[58362] = 32'b00000000000000010001010000000011;
assign LUT_3[58363] = 32'b00000000000000010111111011100000;
assign LUT_3[58364] = 32'b00000000000000001100010110010101;
assign LUT_3[58365] = 32'b00000000000000010011000001110010;
assign LUT_3[58366] = 32'b00000000000000001110011101111001;
assign LUT_3[58367] = 32'b00000000000000010101001001010110;
assign LUT_3[58368] = 32'b00000000000000001010001010011101;
assign LUT_3[58369] = 32'b00000000000000010000110101111010;
assign LUT_3[58370] = 32'b00000000000000001100010010000001;
assign LUT_3[58371] = 32'b00000000000000010010111101011110;
assign LUT_3[58372] = 32'b00000000000000000111011000010011;
assign LUT_3[58373] = 32'b00000000000000001110000011110000;
assign LUT_3[58374] = 32'b00000000000000001001011111110111;
assign LUT_3[58375] = 32'b00000000000000010000001011010100;
assign LUT_3[58376] = 32'b00000000000000001111100011100011;
assign LUT_3[58377] = 32'b00000000000000010110001111000000;
assign LUT_3[58378] = 32'b00000000000000010001101011000111;
assign LUT_3[58379] = 32'b00000000000000011000010110100100;
assign LUT_3[58380] = 32'b00000000000000001100110001011001;
assign LUT_3[58381] = 32'b00000000000000010011011100110110;
assign LUT_3[58382] = 32'b00000000000000001110111000111101;
assign LUT_3[58383] = 32'b00000000000000010101100100011010;
assign LUT_3[58384] = 32'b00000000000000001101011101100000;
assign LUT_3[58385] = 32'b00000000000000010100001000111101;
assign LUT_3[58386] = 32'b00000000000000001111100101000100;
assign LUT_3[58387] = 32'b00000000000000010110010000100001;
assign LUT_3[58388] = 32'b00000000000000001010101011010110;
assign LUT_3[58389] = 32'b00000000000000010001010110110011;
assign LUT_3[58390] = 32'b00000000000000001100110010111010;
assign LUT_3[58391] = 32'b00000000000000010011011110010111;
assign LUT_3[58392] = 32'b00000000000000010010110110100110;
assign LUT_3[58393] = 32'b00000000000000011001100010000011;
assign LUT_3[58394] = 32'b00000000000000010100111110001010;
assign LUT_3[58395] = 32'b00000000000000011011101001100111;
assign LUT_3[58396] = 32'b00000000000000010000000100011100;
assign LUT_3[58397] = 32'b00000000000000010110101111111001;
assign LUT_3[58398] = 32'b00000000000000010010001100000000;
assign LUT_3[58399] = 32'b00000000000000011000110111011101;
assign LUT_3[58400] = 32'b00000000000000001011011000111101;
assign LUT_3[58401] = 32'b00000000000000010010000100011010;
assign LUT_3[58402] = 32'b00000000000000001101100000100001;
assign LUT_3[58403] = 32'b00000000000000010100001011111110;
assign LUT_3[58404] = 32'b00000000000000001000100110110011;
assign LUT_3[58405] = 32'b00000000000000001111010010010000;
assign LUT_3[58406] = 32'b00000000000000001010101110010111;
assign LUT_3[58407] = 32'b00000000000000010001011001110100;
assign LUT_3[58408] = 32'b00000000000000010000110010000011;
assign LUT_3[58409] = 32'b00000000000000010111011101100000;
assign LUT_3[58410] = 32'b00000000000000010010111001100111;
assign LUT_3[58411] = 32'b00000000000000011001100101000100;
assign LUT_3[58412] = 32'b00000000000000001101111111111001;
assign LUT_3[58413] = 32'b00000000000000010100101011010110;
assign LUT_3[58414] = 32'b00000000000000010000000111011101;
assign LUT_3[58415] = 32'b00000000000000010110110010111010;
assign LUT_3[58416] = 32'b00000000000000001110101100000000;
assign LUT_3[58417] = 32'b00000000000000010101010111011101;
assign LUT_3[58418] = 32'b00000000000000010000110011100100;
assign LUT_3[58419] = 32'b00000000000000010111011111000001;
assign LUT_3[58420] = 32'b00000000000000001011111001110110;
assign LUT_3[58421] = 32'b00000000000000010010100101010011;
assign LUT_3[58422] = 32'b00000000000000001110000001011010;
assign LUT_3[58423] = 32'b00000000000000010100101100110111;
assign LUT_3[58424] = 32'b00000000000000010100000101000110;
assign LUT_3[58425] = 32'b00000000000000011010110000100011;
assign LUT_3[58426] = 32'b00000000000000010110001100101010;
assign LUT_3[58427] = 32'b00000000000000011100111000000111;
assign LUT_3[58428] = 32'b00000000000000010001010010111100;
assign LUT_3[58429] = 32'b00000000000000010111111110011001;
assign LUT_3[58430] = 32'b00000000000000010011011010100000;
assign LUT_3[58431] = 32'b00000000000000011010000101111101;
assign LUT_3[58432] = 32'b00000000000000001010000011001000;
assign LUT_3[58433] = 32'b00000000000000010000101110100101;
assign LUT_3[58434] = 32'b00000000000000001100001010101100;
assign LUT_3[58435] = 32'b00000000000000010010110110001001;
assign LUT_3[58436] = 32'b00000000000000000111010000111110;
assign LUT_3[58437] = 32'b00000000000000001101111100011011;
assign LUT_3[58438] = 32'b00000000000000001001011000100010;
assign LUT_3[58439] = 32'b00000000000000010000000011111111;
assign LUT_3[58440] = 32'b00000000000000001111011100001110;
assign LUT_3[58441] = 32'b00000000000000010110000111101011;
assign LUT_3[58442] = 32'b00000000000000010001100011110010;
assign LUT_3[58443] = 32'b00000000000000011000001111001111;
assign LUT_3[58444] = 32'b00000000000000001100101010000100;
assign LUT_3[58445] = 32'b00000000000000010011010101100001;
assign LUT_3[58446] = 32'b00000000000000001110110001101000;
assign LUT_3[58447] = 32'b00000000000000010101011101000101;
assign LUT_3[58448] = 32'b00000000000000001101010110001011;
assign LUT_3[58449] = 32'b00000000000000010100000001101000;
assign LUT_3[58450] = 32'b00000000000000001111011101101111;
assign LUT_3[58451] = 32'b00000000000000010110001001001100;
assign LUT_3[58452] = 32'b00000000000000001010100100000001;
assign LUT_3[58453] = 32'b00000000000000010001001111011110;
assign LUT_3[58454] = 32'b00000000000000001100101011100101;
assign LUT_3[58455] = 32'b00000000000000010011010111000010;
assign LUT_3[58456] = 32'b00000000000000010010101111010001;
assign LUT_3[58457] = 32'b00000000000000011001011010101110;
assign LUT_3[58458] = 32'b00000000000000010100110110110101;
assign LUT_3[58459] = 32'b00000000000000011011100010010010;
assign LUT_3[58460] = 32'b00000000000000001111111101000111;
assign LUT_3[58461] = 32'b00000000000000010110101000100100;
assign LUT_3[58462] = 32'b00000000000000010010000100101011;
assign LUT_3[58463] = 32'b00000000000000011000110000001000;
assign LUT_3[58464] = 32'b00000000000000001011010001101000;
assign LUT_3[58465] = 32'b00000000000000010001111101000101;
assign LUT_3[58466] = 32'b00000000000000001101011001001100;
assign LUT_3[58467] = 32'b00000000000000010100000100101001;
assign LUT_3[58468] = 32'b00000000000000001000011111011110;
assign LUT_3[58469] = 32'b00000000000000001111001010111011;
assign LUT_3[58470] = 32'b00000000000000001010100111000010;
assign LUT_3[58471] = 32'b00000000000000010001010010011111;
assign LUT_3[58472] = 32'b00000000000000010000101010101110;
assign LUT_3[58473] = 32'b00000000000000010111010110001011;
assign LUT_3[58474] = 32'b00000000000000010010110010010010;
assign LUT_3[58475] = 32'b00000000000000011001011101101111;
assign LUT_3[58476] = 32'b00000000000000001101111000100100;
assign LUT_3[58477] = 32'b00000000000000010100100100000001;
assign LUT_3[58478] = 32'b00000000000000010000000000001000;
assign LUT_3[58479] = 32'b00000000000000010110101011100101;
assign LUT_3[58480] = 32'b00000000000000001110100100101011;
assign LUT_3[58481] = 32'b00000000000000010101010000001000;
assign LUT_3[58482] = 32'b00000000000000010000101100001111;
assign LUT_3[58483] = 32'b00000000000000010111010111101100;
assign LUT_3[58484] = 32'b00000000000000001011110010100001;
assign LUT_3[58485] = 32'b00000000000000010010011101111110;
assign LUT_3[58486] = 32'b00000000000000001101111010000101;
assign LUT_3[58487] = 32'b00000000000000010100100101100010;
assign LUT_3[58488] = 32'b00000000000000010011111101110001;
assign LUT_3[58489] = 32'b00000000000000011010101001001110;
assign LUT_3[58490] = 32'b00000000000000010110000101010101;
assign LUT_3[58491] = 32'b00000000000000011100110000110010;
assign LUT_3[58492] = 32'b00000000000000010001001011100111;
assign LUT_3[58493] = 32'b00000000000000010111110111000100;
assign LUT_3[58494] = 32'b00000000000000010011010011001011;
assign LUT_3[58495] = 32'b00000000000000011001111110101000;
assign LUT_3[58496] = 32'b00000000000000001100010101011011;
assign LUT_3[58497] = 32'b00000000000000010011000000111000;
assign LUT_3[58498] = 32'b00000000000000001110011100111111;
assign LUT_3[58499] = 32'b00000000000000010101001000011100;
assign LUT_3[58500] = 32'b00000000000000001001100011010001;
assign LUT_3[58501] = 32'b00000000000000010000001110101110;
assign LUT_3[58502] = 32'b00000000000000001011101010110101;
assign LUT_3[58503] = 32'b00000000000000010010010110010010;
assign LUT_3[58504] = 32'b00000000000000010001101110100001;
assign LUT_3[58505] = 32'b00000000000000011000011001111110;
assign LUT_3[58506] = 32'b00000000000000010011110110000101;
assign LUT_3[58507] = 32'b00000000000000011010100001100010;
assign LUT_3[58508] = 32'b00000000000000001110111100010111;
assign LUT_3[58509] = 32'b00000000000000010101100111110100;
assign LUT_3[58510] = 32'b00000000000000010001000011111011;
assign LUT_3[58511] = 32'b00000000000000010111101111011000;
assign LUT_3[58512] = 32'b00000000000000001111101000011110;
assign LUT_3[58513] = 32'b00000000000000010110010011111011;
assign LUT_3[58514] = 32'b00000000000000010001110000000010;
assign LUT_3[58515] = 32'b00000000000000011000011011011111;
assign LUT_3[58516] = 32'b00000000000000001100110110010100;
assign LUT_3[58517] = 32'b00000000000000010011100001110001;
assign LUT_3[58518] = 32'b00000000000000001110111101111000;
assign LUT_3[58519] = 32'b00000000000000010101101001010101;
assign LUT_3[58520] = 32'b00000000000000010101000001100100;
assign LUT_3[58521] = 32'b00000000000000011011101101000001;
assign LUT_3[58522] = 32'b00000000000000010111001001001000;
assign LUT_3[58523] = 32'b00000000000000011101110100100101;
assign LUT_3[58524] = 32'b00000000000000010010001111011010;
assign LUT_3[58525] = 32'b00000000000000011000111010110111;
assign LUT_3[58526] = 32'b00000000000000010100010110111110;
assign LUT_3[58527] = 32'b00000000000000011011000010011011;
assign LUT_3[58528] = 32'b00000000000000001101100011111011;
assign LUT_3[58529] = 32'b00000000000000010100001111011000;
assign LUT_3[58530] = 32'b00000000000000001111101011011111;
assign LUT_3[58531] = 32'b00000000000000010110010110111100;
assign LUT_3[58532] = 32'b00000000000000001010110001110001;
assign LUT_3[58533] = 32'b00000000000000010001011101001110;
assign LUT_3[58534] = 32'b00000000000000001100111001010101;
assign LUT_3[58535] = 32'b00000000000000010011100100110010;
assign LUT_3[58536] = 32'b00000000000000010010111101000001;
assign LUT_3[58537] = 32'b00000000000000011001101000011110;
assign LUT_3[58538] = 32'b00000000000000010101000100100101;
assign LUT_3[58539] = 32'b00000000000000011011110000000010;
assign LUT_3[58540] = 32'b00000000000000010000001010110111;
assign LUT_3[58541] = 32'b00000000000000010110110110010100;
assign LUT_3[58542] = 32'b00000000000000010010010010011011;
assign LUT_3[58543] = 32'b00000000000000011000111101111000;
assign LUT_3[58544] = 32'b00000000000000010000110110111110;
assign LUT_3[58545] = 32'b00000000000000010111100010011011;
assign LUT_3[58546] = 32'b00000000000000010010111110100010;
assign LUT_3[58547] = 32'b00000000000000011001101001111111;
assign LUT_3[58548] = 32'b00000000000000001110000100110100;
assign LUT_3[58549] = 32'b00000000000000010100110000010001;
assign LUT_3[58550] = 32'b00000000000000010000001100011000;
assign LUT_3[58551] = 32'b00000000000000010110110111110101;
assign LUT_3[58552] = 32'b00000000000000010110010000000100;
assign LUT_3[58553] = 32'b00000000000000011100111011100001;
assign LUT_3[58554] = 32'b00000000000000011000010111101000;
assign LUT_3[58555] = 32'b00000000000000011111000011000101;
assign LUT_3[58556] = 32'b00000000000000010011011101111010;
assign LUT_3[58557] = 32'b00000000000000011010001001010111;
assign LUT_3[58558] = 32'b00000000000000010101100101011110;
assign LUT_3[58559] = 32'b00000000000000011100010000111011;
assign LUT_3[58560] = 32'b00000000000000001100001110000110;
assign LUT_3[58561] = 32'b00000000000000010010111001100011;
assign LUT_3[58562] = 32'b00000000000000001110010101101010;
assign LUT_3[58563] = 32'b00000000000000010101000001000111;
assign LUT_3[58564] = 32'b00000000000000001001011011111100;
assign LUT_3[58565] = 32'b00000000000000010000000111011001;
assign LUT_3[58566] = 32'b00000000000000001011100011100000;
assign LUT_3[58567] = 32'b00000000000000010010001110111101;
assign LUT_3[58568] = 32'b00000000000000010001100111001100;
assign LUT_3[58569] = 32'b00000000000000011000010010101001;
assign LUT_3[58570] = 32'b00000000000000010011101110110000;
assign LUT_3[58571] = 32'b00000000000000011010011010001101;
assign LUT_3[58572] = 32'b00000000000000001110110101000010;
assign LUT_3[58573] = 32'b00000000000000010101100000011111;
assign LUT_3[58574] = 32'b00000000000000010000111100100110;
assign LUT_3[58575] = 32'b00000000000000010111101000000011;
assign LUT_3[58576] = 32'b00000000000000001111100001001001;
assign LUT_3[58577] = 32'b00000000000000010110001100100110;
assign LUT_3[58578] = 32'b00000000000000010001101000101101;
assign LUT_3[58579] = 32'b00000000000000011000010100001010;
assign LUT_3[58580] = 32'b00000000000000001100101110111111;
assign LUT_3[58581] = 32'b00000000000000010011011010011100;
assign LUT_3[58582] = 32'b00000000000000001110110110100011;
assign LUT_3[58583] = 32'b00000000000000010101100010000000;
assign LUT_3[58584] = 32'b00000000000000010100111010001111;
assign LUT_3[58585] = 32'b00000000000000011011100101101100;
assign LUT_3[58586] = 32'b00000000000000010111000001110011;
assign LUT_3[58587] = 32'b00000000000000011101101101010000;
assign LUT_3[58588] = 32'b00000000000000010010001000000101;
assign LUT_3[58589] = 32'b00000000000000011000110011100010;
assign LUT_3[58590] = 32'b00000000000000010100001111101001;
assign LUT_3[58591] = 32'b00000000000000011010111011000110;
assign LUT_3[58592] = 32'b00000000000000001101011100100110;
assign LUT_3[58593] = 32'b00000000000000010100001000000011;
assign LUT_3[58594] = 32'b00000000000000001111100100001010;
assign LUT_3[58595] = 32'b00000000000000010110001111100111;
assign LUT_3[58596] = 32'b00000000000000001010101010011100;
assign LUT_3[58597] = 32'b00000000000000010001010101111001;
assign LUT_3[58598] = 32'b00000000000000001100110010000000;
assign LUT_3[58599] = 32'b00000000000000010011011101011101;
assign LUT_3[58600] = 32'b00000000000000010010110101101100;
assign LUT_3[58601] = 32'b00000000000000011001100001001001;
assign LUT_3[58602] = 32'b00000000000000010100111101010000;
assign LUT_3[58603] = 32'b00000000000000011011101000101101;
assign LUT_3[58604] = 32'b00000000000000010000000011100010;
assign LUT_3[58605] = 32'b00000000000000010110101110111111;
assign LUT_3[58606] = 32'b00000000000000010010001011000110;
assign LUT_3[58607] = 32'b00000000000000011000110110100011;
assign LUT_3[58608] = 32'b00000000000000010000101111101001;
assign LUT_3[58609] = 32'b00000000000000010111011011000110;
assign LUT_3[58610] = 32'b00000000000000010010110111001101;
assign LUT_3[58611] = 32'b00000000000000011001100010101010;
assign LUT_3[58612] = 32'b00000000000000001101111101011111;
assign LUT_3[58613] = 32'b00000000000000010100101000111100;
assign LUT_3[58614] = 32'b00000000000000010000000101000011;
assign LUT_3[58615] = 32'b00000000000000010110110000100000;
assign LUT_3[58616] = 32'b00000000000000010110001000101111;
assign LUT_3[58617] = 32'b00000000000000011100110100001100;
assign LUT_3[58618] = 32'b00000000000000011000010000010011;
assign LUT_3[58619] = 32'b00000000000000011110111011110000;
assign LUT_3[58620] = 32'b00000000000000010011010110100101;
assign LUT_3[58621] = 32'b00000000000000011010000010000010;
assign LUT_3[58622] = 32'b00000000000000010101011110001001;
assign LUT_3[58623] = 32'b00000000000000011100001001100110;
assign LUT_3[58624] = 32'b00000000000000000110011001111110;
assign LUT_3[58625] = 32'b00000000000000001101000101011011;
assign LUT_3[58626] = 32'b00000000000000001000100001100010;
assign LUT_3[58627] = 32'b00000000000000001111001100111111;
assign LUT_3[58628] = 32'b00000000000000000011100111110100;
assign LUT_3[58629] = 32'b00000000000000001010010011010001;
assign LUT_3[58630] = 32'b00000000000000000101101111011000;
assign LUT_3[58631] = 32'b00000000000000001100011010110101;
assign LUT_3[58632] = 32'b00000000000000001011110011000100;
assign LUT_3[58633] = 32'b00000000000000010010011110100001;
assign LUT_3[58634] = 32'b00000000000000001101111010101000;
assign LUT_3[58635] = 32'b00000000000000010100100110000101;
assign LUT_3[58636] = 32'b00000000000000001001000000111010;
assign LUT_3[58637] = 32'b00000000000000001111101100010111;
assign LUT_3[58638] = 32'b00000000000000001011001000011110;
assign LUT_3[58639] = 32'b00000000000000010001110011111011;
assign LUT_3[58640] = 32'b00000000000000001001101101000001;
assign LUT_3[58641] = 32'b00000000000000010000011000011110;
assign LUT_3[58642] = 32'b00000000000000001011110100100101;
assign LUT_3[58643] = 32'b00000000000000010010100000000010;
assign LUT_3[58644] = 32'b00000000000000000110111010110111;
assign LUT_3[58645] = 32'b00000000000000001101100110010100;
assign LUT_3[58646] = 32'b00000000000000001001000010011011;
assign LUT_3[58647] = 32'b00000000000000001111101101111000;
assign LUT_3[58648] = 32'b00000000000000001111000110000111;
assign LUT_3[58649] = 32'b00000000000000010101110001100100;
assign LUT_3[58650] = 32'b00000000000000010001001101101011;
assign LUT_3[58651] = 32'b00000000000000010111111001001000;
assign LUT_3[58652] = 32'b00000000000000001100010011111101;
assign LUT_3[58653] = 32'b00000000000000010010111111011010;
assign LUT_3[58654] = 32'b00000000000000001110011011100001;
assign LUT_3[58655] = 32'b00000000000000010101000110111110;
assign LUT_3[58656] = 32'b00000000000000000111101000011110;
assign LUT_3[58657] = 32'b00000000000000001110010011111011;
assign LUT_3[58658] = 32'b00000000000000001001110000000010;
assign LUT_3[58659] = 32'b00000000000000010000011011011111;
assign LUT_3[58660] = 32'b00000000000000000100110110010100;
assign LUT_3[58661] = 32'b00000000000000001011100001110001;
assign LUT_3[58662] = 32'b00000000000000000110111101111000;
assign LUT_3[58663] = 32'b00000000000000001101101001010101;
assign LUT_3[58664] = 32'b00000000000000001101000001100100;
assign LUT_3[58665] = 32'b00000000000000010011101101000001;
assign LUT_3[58666] = 32'b00000000000000001111001001001000;
assign LUT_3[58667] = 32'b00000000000000010101110100100101;
assign LUT_3[58668] = 32'b00000000000000001010001111011010;
assign LUT_3[58669] = 32'b00000000000000010000111010110111;
assign LUT_3[58670] = 32'b00000000000000001100010110111110;
assign LUT_3[58671] = 32'b00000000000000010011000010011011;
assign LUT_3[58672] = 32'b00000000000000001010111011100001;
assign LUT_3[58673] = 32'b00000000000000010001100110111110;
assign LUT_3[58674] = 32'b00000000000000001101000011000101;
assign LUT_3[58675] = 32'b00000000000000010011101110100010;
assign LUT_3[58676] = 32'b00000000000000001000001001010111;
assign LUT_3[58677] = 32'b00000000000000001110110100110100;
assign LUT_3[58678] = 32'b00000000000000001010010000111011;
assign LUT_3[58679] = 32'b00000000000000010000111100011000;
assign LUT_3[58680] = 32'b00000000000000010000010100100111;
assign LUT_3[58681] = 32'b00000000000000010111000000000100;
assign LUT_3[58682] = 32'b00000000000000010010011100001011;
assign LUT_3[58683] = 32'b00000000000000011001000111101000;
assign LUT_3[58684] = 32'b00000000000000001101100010011101;
assign LUT_3[58685] = 32'b00000000000000010100001101111010;
assign LUT_3[58686] = 32'b00000000000000001111101010000001;
assign LUT_3[58687] = 32'b00000000000000010110010101011110;
assign LUT_3[58688] = 32'b00000000000000000110010010101001;
assign LUT_3[58689] = 32'b00000000000000001100111110000110;
assign LUT_3[58690] = 32'b00000000000000001000011010001101;
assign LUT_3[58691] = 32'b00000000000000001111000101101010;
assign LUT_3[58692] = 32'b00000000000000000011100000011111;
assign LUT_3[58693] = 32'b00000000000000001010001011111100;
assign LUT_3[58694] = 32'b00000000000000000101101000000011;
assign LUT_3[58695] = 32'b00000000000000001100010011100000;
assign LUT_3[58696] = 32'b00000000000000001011101011101111;
assign LUT_3[58697] = 32'b00000000000000010010010111001100;
assign LUT_3[58698] = 32'b00000000000000001101110011010011;
assign LUT_3[58699] = 32'b00000000000000010100011110110000;
assign LUT_3[58700] = 32'b00000000000000001000111001100101;
assign LUT_3[58701] = 32'b00000000000000001111100101000010;
assign LUT_3[58702] = 32'b00000000000000001011000001001001;
assign LUT_3[58703] = 32'b00000000000000010001101100100110;
assign LUT_3[58704] = 32'b00000000000000001001100101101100;
assign LUT_3[58705] = 32'b00000000000000010000010001001001;
assign LUT_3[58706] = 32'b00000000000000001011101101010000;
assign LUT_3[58707] = 32'b00000000000000010010011000101101;
assign LUT_3[58708] = 32'b00000000000000000110110011100010;
assign LUT_3[58709] = 32'b00000000000000001101011110111111;
assign LUT_3[58710] = 32'b00000000000000001000111011000110;
assign LUT_3[58711] = 32'b00000000000000001111100110100011;
assign LUT_3[58712] = 32'b00000000000000001110111110110010;
assign LUT_3[58713] = 32'b00000000000000010101101010001111;
assign LUT_3[58714] = 32'b00000000000000010001000110010110;
assign LUT_3[58715] = 32'b00000000000000010111110001110011;
assign LUT_3[58716] = 32'b00000000000000001100001100101000;
assign LUT_3[58717] = 32'b00000000000000010010111000000101;
assign LUT_3[58718] = 32'b00000000000000001110010100001100;
assign LUT_3[58719] = 32'b00000000000000010100111111101001;
assign LUT_3[58720] = 32'b00000000000000000111100001001001;
assign LUT_3[58721] = 32'b00000000000000001110001100100110;
assign LUT_3[58722] = 32'b00000000000000001001101000101101;
assign LUT_3[58723] = 32'b00000000000000010000010100001010;
assign LUT_3[58724] = 32'b00000000000000000100101110111111;
assign LUT_3[58725] = 32'b00000000000000001011011010011100;
assign LUT_3[58726] = 32'b00000000000000000110110110100011;
assign LUT_3[58727] = 32'b00000000000000001101100010000000;
assign LUT_3[58728] = 32'b00000000000000001100111010001111;
assign LUT_3[58729] = 32'b00000000000000010011100101101100;
assign LUT_3[58730] = 32'b00000000000000001111000001110011;
assign LUT_3[58731] = 32'b00000000000000010101101101010000;
assign LUT_3[58732] = 32'b00000000000000001010001000000101;
assign LUT_3[58733] = 32'b00000000000000010000110011100010;
assign LUT_3[58734] = 32'b00000000000000001100001111101001;
assign LUT_3[58735] = 32'b00000000000000010010111011000110;
assign LUT_3[58736] = 32'b00000000000000001010110100001100;
assign LUT_3[58737] = 32'b00000000000000010001011111101001;
assign LUT_3[58738] = 32'b00000000000000001100111011110000;
assign LUT_3[58739] = 32'b00000000000000010011100111001101;
assign LUT_3[58740] = 32'b00000000000000001000000010000010;
assign LUT_3[58741] = 32'b00000000000000001110101101011111;
assign LUT_3[58742] = 32'b00000000000000001010001001100110;
assign LUT_3[58743] = 32'b00000000000000010000110101000011;
assign LUT_3[58744] = 32'b00000000000000010000001101010010;
assign LUT_3[58745] = 32'b00000000000000010110111000101111;
assign LUT_3[58746] = 32'b00000000000000010010010100110110;
assign LUT_3[58747] = 32'b00000000000000011001000000010011;
assign LUT_3[58748] = 32'b00000000000000001101011011001000;
assign LUT_3[58749] = 32'b00000000000000010100000110100101;
assign LUT_3[58750] = 32'b00000000000000001111100010101100;
assign LUT_3[58751] = 32'b00000000000000010110001110001001;
assign LUT_3[58752] = 32'b00000000000000001000100100111100;
assign LUT_3[58753] = 32'b00000000000000001111010000011001;
assign LUT_3[58754] = 32'b00000000000000001010101100100000;
assign LUT_3[58755] = 32'b00000000000000010001010111111101;
assign LUT_3[58756] = 32'b00000000000000000101110010110010;
assign LUT_3[58757] = 32'b00000000000000001100011110001111;
assign LUT_3[58758] = 32'b00000000000000000111111010010110;
assign LUT_3[58759] = 32'b00000000000000001110100101110011;
assign LUT_3[58760] = 32'b00000000000000001101111110000010;
assign LUT_3[58761] = 32'b00000000000000010100101001011111;
assign LUT_3[58762] = 32'b00000000000000010000000101100110;
assign LUT_3[58763] = 32'b00000000000000010110110001000011;
assign LUT_3[58764] = 32'b00000000000000001011001011111000;
assign LUT_3[58765] = 32'b00000000000000010001110111010101;
assign LUT_3[58766] = 32'b00000000000000001101010011011100;
assign LUT_3[58767] = 32'b00000000000000010011111110111001;
assign LUT_3[58768] = 32'b00000000000000001011110111111111;
assign LUT_3[58769] = 32'b00000000000000010010100011011100;
assign LUT_3[58770] = 32'b00000000000000001101111111100011;
assign LUT_3[58771] = 32'b00000000000000010100101011000000;
assign LUT_3[58772] = 32'b00000000000000001001000101110101;
assign LUT_3[58773] = 32'b00000000000000001111110001010010;
assign LUT_3[58774] = 32'b00000000000000001011001101011001;
assign LUT_3[58775] = 32'b00000000000000010001111000110110;
assign LUT_3[58776] = 32'b00000000000000010001010001000101;
assign LUT_3[58777] = 32'b00000000000000010111111100100010;
assign LUT_3[58778] = 32'b00000000000000010011011000101001;
assign LUT_3[58779] = 32'b00000000000000011010000100000110;
assign LUT_3[58780] = 32'b00000000000000001110011110111011;
assign LUT_3[58781] = 32'b00000000000000010101001010011000;
assign LUT_3[58782] = 32'b00000000000000010000100110011111;
assign LUT_3[58783] = 32'b00000000000000010111010001111100;
assign LUT_3[58784] = 32'b00000000000000001001110011011100;
assign LUT_3[58785] = 32'b00000000000000010000011110111001;
assign LUT_3[58786] = 32'b00000000000000001011111011000000;
assign LUT_3[58787] = 32'b00000000000000010010100110011101;
assign LUT_3[58788] = 32'b00000000000000000111000001010010;
assign LUT_3[58789] = 32'b00000000000000001101101100101111;
assign LUT_3[58790] = 32'b00000000000000001001001000110110;
assign LUT_3[58791] = 32'b00000000000000001111110100010011;
assign LUT_3[58792] = 32'b00000000000000001111001100100010;
assign LUT_3[58793] = 32'b00000000000000010101110111111111;
assign LUT_3[58794] = 32'b00000000000000010001010100000110;
assign LUT_3[58795] = 32'b00000000000000010111111111100011;
assign LUT_3[58796] = 32'b00000000000000001100011010011000;
assign LUT_3[58797] = 32'b00000000000000010011000101110101;
assign LUT_3[58798] = 32'b00000000000000001110100001111100;
assign LUT_3[58799] = 32'b00000000000000010101001101011001;
assign LUT_3[58800] = 32'b00000000000000001101000110011111;
assign LUT_3[58801] = 32'b00000000000000010011110001111100;
assign LUT_3[58802] = 32'b00000000000000001111001110000011;
assign LUT_3[58803] = 32'b00000000000000010101111001100000;
assign LUT_3[58804] = 32'b00000000000000001010010100010101;
assign LUT_3[58805] = 32'b00000000000000010000111111110010;
assign LUT_3[58806] = 32'b00000000000000001100011011111001;
assign LUT_3[58807] = 32'b00000000000000010011000111010110;
assign LUT_3[58808] = 32'b00000000000000010010011111100101;
assign LUT_3[58809] = 32'b00000000000000011001001011000010;
assign LUT_3[58810] = 32'b00000000000000010100100111001001;
assign LUT_3[58811] = 32'b00000000000000011011010010100110;
assign LUT_3[58812] = 32'b00000000000000001111101101011011;
assign LUT_3[58813] = 32'b00000000000000010110011000111000;
assign LUT_3[58814] = 32'b00000000000000010001110100111111;
assign LUT_3[58815] = 32'b00000000000000011000100000011100;
assign LUT_3[58816] = 32'b00000000000000001000011101100111;
assign LUT_3[58817] = 32'b00000000000000001111001001000100;
assign LUT_3[58818] = 32'b00000000000000001010100101001011;
assign LUT_3[58819] = 32'b00000000000000010001010000101000;
assign LUT_3[58820] = 32'b00000000000000000101101011011101;
assign LUT_3[58821] = 32'b00000000000000001100010110111010;
assign LUT_3[58822] = 32'b00000000000000000111110011000001;
assign LUT_3[58823] = 32'b00000000000000001110011110011110;
assign LUT_3[58824] = 32'b00000000000000001101110110101101;
assign LUT_3[58825] = 32'b00000000000000010100100010001010;
assign LUT_3[58826] = 32'b00000000000000001111111110010001;
assign LUT_3[58827] = 32'b00000000000000010110101001101110;
assign LUT_3[58828] = 32'b00000000000000001011000100100011;
assign LUT_3[58829] = 32'b00000000000000010001110000000000;
assign LUT_3[58830] = 32'b00000000000000001101001100000111;
assign LUT_3[58831] = 32'b00000000000000010011110111100100;
assign LUT_3[58832] = 32'b00000000000000001011110000101010;
assign LUT_3[58833] = 32'b00000000000000010010011100000111;
assign LUT_3[58834] = 32'b00000000000000001101111000001110;
assign LUT_3[58835] = 32'b00000000000000010100100011101011;
assign LUT_3[58836] = 32'b00000000000000001000111110100000;
assign LUT_3[58837] = 32'b00000000000000001111101001111101;
assign LUT_3[58838] = 32'b00000000000000001011000110000100;
assign LUT_3[58839] = 32'b00000000000000010001110001100001;
assign LUT_3[58840] = 32'b00000000000000010001001001110000;
assign LUT_3[58841] = 32'b00000000000000010111110101001101;
assign LUT_3[58842] = 32'b00000000000000010011010001010100;
assign LUT_3[58843] = 32'b00000000000000011001111100110001;
assign LUT_3[58844] = 32'b00000000000000001110010111100110;
assign LUT_3[58845] = 32'b00000000000000010101000011000011;
assign LUT_3[58846] = 32'b00000000000000010000011111001010;
assign LUT_3[58847] = 32'b00000000000000010111001010100111;
assign LUT_3[58848] = 32'b00000000000000001001101100000111;
assign LUT_3[58849] = 32'b00000000000000010000010111100100;
assign LUT_3[58850] = 32'b00000000000000001011110011101011;
assign LUT_3[58851] = 32'b00000000000000010010011111001000;
assign LUT_3[58852] = 32'b00000000000000000110111001111101;
assign LUT_3[58853] = 32'b00000000000000001101100101011010;
assign LUT_3[58854] = 32'b00000000000000001001000001100001;
assign LUT_3[58855] = 32'b00000000000000001111101100111110;
assign LUT_3[58856] = 32'b00000000000000001111000101001101;
assign LUT_3[58857] = 32'b00000000000000010101110000101010;
assign LUT_3[58858] = 32'b00000000000000010001001100110001;
assign LUT_3[58859] = 32'b00000000000000010111111000001110;
assign LUT_3[58860] = 32'b00000000000000001100010011000011;
assign LUT_3[58861] = 32'b00000000000000010010111110100000;
assign LUT_3[58862] = 32'b00000000000000001110011010100111;
assign LUT_3[58863] = 32'b00000000000000010101000110000100;
assign LUT_3[58864] = 32'b00000000000000001100111111001010;
assign LUT_3[58865] = 32'b00000000000000010011101010100111;
assign LUT_3[58866] = 32'b00000000000000001111000110101110;
assign LUT_3[58867] = 32'b00000000000000010101110010001011;
assign LUT_3[58868] = 32'b00000000000000001010001101000000;
assign LUT_3[58869] = 32'b00000000000000010000111000011101;
assign LUT_3[58870] = 32'b00000000000000001100010100100100;
assign LUT_3[58871] = 32'b00000000000000010011000000000001;
assign LUT_3[58872] = 32'b00000000000000010010011000010000;
assign LUT_3[58873] = 32'b00000000000000011001000011101101;
assign LUT_3[58874] = 32'b00000000000000010100011111110100;
assign LUT_3[58875] = 32'b00000000000000011011001011010001;
assign LUT_3[58876] = 32'b00000000000000001111100110000110;
assign LUT_3[58877] = 32'b00000000000000010110010001100011;
assign LUT_3[58878] = 32'b00000000000000010001101101101010;
assign LUT_3[58879] = 32'b00000000000000011000011001000111;
assign LUT_3[58880] = 32'b00000000000000001101011111101001;
assign LUT_3[58881] = 32'b00000000000000010100001011000110;
assign LUT_3[58882] = 32'b00000000000000001111100111001101;
assign LUT_3[58883] = 32'b00000000000000010110010010101010;
assign LUT_3[58884] = 32'b00000000000000001010101101011111;
assign LUT_3[58885] = 32'b00000000000000010001011000111100;
assign LUT_3[58886] = 32'b00000000000000001100110101000011;
assign LUT_3[58887] = 32'b00000000000000010011100000100000;
assign LUT_3[58888] = 32'b00000000000000010010111000101111;
assign LUT_3[58889] = 32'b00000000000000011001100100001100;
assign LUT_3[58890] = 32'b00000000000000010101000000010011;
assign LUT_3[58891] = 32'b00000000000000011011101011110000;
assign LUT_3[58892] = 32'b00000000000000010000000110100101;
assign LUT_3[58893] = 32'b00000000000000010110110010000010;
assign LUT_3[58894] = 32'b00000000000000010010001110001001;
assign LUT_3[58895] = 32'b00000000000000011000111001100110;
assign LUT_3[58896] = 32'b00000000000000010000110010101100;
assign LUT_3[58897] = 32'b00000000000000010111011110001001;
assign LUT_3[58898] = 32'b00000000000000010010111010010000;
assign LUT_3[58899] = 32'b00000000000000011001100101101101;
assign LUT_3[58900] = 32'b00000000000000001110000000100010;
assign LUT_3[58901] = 32'b00000000000000010100101011111111;
assign LUT_3[58902] = 32'b00000000000000010000001000000110;
assign LUT_3[58903] = 32'b00000000000000010110110011100011;
assign LUT_3[58904] = 32'b00000000000000010110001011110010;
assign LUT_3[58905] = 32'b00000000000000011100110111001111;
assign LUT_3[58906] = 32'b00000000000000011000010011010110;
assign LUT_3[58907] = 32'b00000000000000011110111110110011;
assign LUT_3[58908] = 32'b00000000000000010011011001101000;
assign LUT_3[58909] = 32'b00000000000000011010000101000101;
assign LUT_3[58910] = 32'b00000000000000010101100001001100;
assign LUT_3[58911] = 32'b00000000000000011100001100101001;
assign LUT_3[58912] = 32'b00000000000000001110101110001001;
assign LUT_3[58913] = 32'b00000000000000010101011001100110;
assign LUT_3[58914] = 32'b00000000000000010000110101101101;
assign LUT_3[58915] = 32'b00000000000000010111100001001010;
assign LUT_3[58916] = 32'b00000000000000001011111011111111;
assign LUT_3[58917] = 32'b00000000000000010010100111011100;
assign LUT_3[58918] = 32'b00000000000000001110000011100011;
assign LUT_3[58919] = 32'b00000000000000010100101111000000;
assign LUT_3[58920] = 32'b00000000000000010100000111001111;
assign LUT_3[58921] = 32'b00000000000000011010110010101100;
assign LUT_3[58922] = 32'b00000000000000010110001110110011;
assign LUT_3[58923] = 32'b00000000000000011100111010010000;
assign LUT_3[58924] = 32'b00000000000000010001010101000101;
assign LUT_3[58925] = 32'b00000000000000011000000000100010;
assign LUT_3[58926] = 32'b00000000000000010011011100101001;
assign LUT_3[58927] = 32'b00000000000000011010001000000110;
assign LUT_3[58928] = 32'b00000000000000010010000001001100;
assign LUT_3[58929] = 32'b00000000000000011000101100101001;
assign LUT_3[58930] = 32'b00000000000000010100001000110000;
assign LUT_3[58931] = 32'b00000000000000011010110100001101;
assign LUT_3[58932] = 32'b00000000000000001111001111000010;
assign LUT_3[58933] = 32'b00000000000000010101111010011111;
assign LUT_3[58934] = 32'b00000000000000010001010110100110;
assign LUT_3[58935] = 32'b00000000000000011000000010000011;
assign LUT_3[58936] = 32'b00000000000000010111011010010010;
assign LUT_3[58937] = 32'b00000000000000011110000101101111;
assign LUT_3[58938] = 32'b00000000000000011001100001110110;
assign LUT_3[58939] = 32'b00000000000000100000001101010011;
assign LUT_3[58940] = 32'b00000000000000010100101000001000;
assign LUT_3[58941] = 32'b00000000000000011011010011100101;
assign LUT_3[58942] = 32'b00000000000000010110101111101100;
assign LUT_3[58943] = 32'b00000000000000011101011011001001;
assign LUT_3[58944] = 32'b00000000000000001101011000010100;
assign LUT_3[58945] = 32'b00000000000000010100000011110001;
assign LUT_3[58946] = 32'b00000000000000001111011111111000;
assign LUT_3[58947] = 32'b00000000000000010110001011010101;
assign LUT_3[58948] = 32'b00000000000000001010100110001010;
assign LUT_3[58949] = 32'b00000000000000010001010001100111;
assign LUT_3[58950] = 32'b00000000000000001100101101101110;
assign LUT_3[58951] = 32'b00000000000000010011011001001011;
assign LUT_3[58952] = 32'b00000000000000010010110001011010;
assign LUT_3[58953] = 32'b00000000000000011001011100110111;
assign LUT_3[58954] = 32'b00000000000000010100111000111110;
assign LUT_3[58955] = 32'b00000000000000011011100100011011;
assign LUT_3[58956] = 32'b00000000000000001111111111010000;
assign LUT_3[58957] = 32'b00000000000000010110101010101101;
assign LUT_3[58958] = 32'b00000000000000010010000110110100;
assign LUT_3[58959] = 32'b00000000000000011000110010010001;
assign LUT_3[58960] = 32'b00000000000000010000101011010111;
assign LUT_3[58961] = 32'b00000000000000010111010110110100;
assign LUT_3[58962] = 32'b00000000000000010010110010111011;
assign LUT_3[58963] = 32'b00000000000000011001011110011000;
assign LUT_3[58964] = 32'b00000000000000001101111001001101;
assign LUT_3[58965] = 32'b00000000000000010100100100101010;
assign LUT_3[58966] = 32'b00000000000000010000000000110001;
assign LUT_3[58967] = 32'b00000000000000010110101100001110;
assign LUT_3[58968] = 32'b00000000000000010110000100011101;
assign LUT_3[58969] = 32'b00000000000000011100101111111010;
assign LUT_3[58970] = 32'b00000000000000011000001100000001;
assign LUT_3[58971] = 32'b00000000000000011110110111011110;
assign LUT_3[58972] = 32'b00000000000000010011010010010011;
assign LUT_3[58973] = 32'b00000000000000011001111101110000;
assign LUT_3[58974] = 32'b00000000000000010101011001110111;
assign LUT_3[58975] = 32'b00000000000000011100000101010100;
assign LUT_3[58976] = 32'b00000000000000001110100110110100;
assign LUT_3[58977] = 32'b00000000000000010101010010010001;
assign LUT_3[58978] = 32'b00000000000000010000101110011000;
assign LUT_3[58979] = 32'b00000000000000010111011001110101;
assign LUT_3[58980] = 32'b00000000000000001011110100101010;
assign LUT_3[58981] = 32'b00000000000000010010100000000111;
assign LUT_3[58982] = 32'b00000000000000001101111100001110;
assign LUT_3[58983] = 32'b00000000000000010100100111101011;
assign LUT_3[58984] = 32'b00000000000000010011111111111010;
assign LUT_3[58985] = 32'b00000000000000011010101011010111;
assign LUT_3[58986] = 32'b00000000000000010110000111011110;
assign LUT_3[58987] = 32'b00000000000000011100110010111011;
assign LUT_3[58988] = 32'b00000000000000010001001101110000;
assign LUT_3[58989] = 32'b00000000000000010111111001001101;
assign LUT_3[58990] = 32'b00000000000000010011010101010100;
assign LUT_3[58991] = 32'b00000000000000011010000000110001;
assign LUT_3[58992] = 32'b00000000000000010001111001110111;
assign LUT_3[58993] = 32'b00000000000000011000100101010100;
assign LUT_3[58994] = 32'b00000000000000010100000001011011;
assign LUT_3[58995] = 32'b00000000000000011010101100111000;
assign LUT_3[58996] = 32'b00000000000000001111000111101101;
assign LUT_3[58997] = 32'b00000000000000010101110011001010;
assign LUT_3[58998] = 32'b00000000000000010001001111010001;
assign LUT_3[58999] = 32'b00000000000000010111111010101110;
assign LUT_3[59000] = 32'b00000000000000010111010010111101;
assign LUT_3[59001] = 32'b00000000000000011101111110011010;
assign LUT_3[59002] = 32'b00000000000000011001011010100001;
assign LUT_3[59003] = 32'b00000000000000100000000101111110;
assign LUT_3[59004] = 32'b00000000000000010100100000110011;
assign LUT_3[59005] = 32'b00000000000000011011001100010000;
assign LUT_3[59006] = 32'b00000000000000010110101000010111;
assign LUT_3[59007] = 32'b00000000000000011101010011110100;
assign LUT_3[59008] = 32'b00000000000000001111101010100111;
assign LUT_3[59009] = 32'b00000000000000010110010110000100;
assign LUT_3[59010] = 32'b00000000000000010001110010001011;
assign LUT_3[59011] = 32'b00000000000000011000011101101000;
assign LUT_3[59012] = 32'b00000000000000001100111000011101;
assign LUT_3[59013] = 32'b00000000000000010011100011111010;
assign LUT_3[59014] = 32'b00000000000000001111000000000001;
assign LUT_3[59015] = 32'b00000000000000010101101011011110;
assign LUT_3[59016] = 32'b00000000000000010101000011101101;
assign LUT_3[59017] = 32'b00000000000000011011101111001010;
assign LUT_3[59018] = 32'b00000000000000010111001011010001;
assign LUT_3[59019] = 32'b00000000000000011101110110101110;
assign LUT_3[59020] = 32'b00000000000000010010010001100011;
assign LUT_3[59021] = 32'b00000000000000011000111101000000;
assign LUT_3[59022] = 32'b00000000000000010100011001000111;
assign LUT_3[59023] = 32'b00000000000000011011000100100100;
assign LUT_3[59024] = 32'b00000000000000010010111101101010;
assign LUT_3[59025] = 32'b00000000000000011001101001000111;
assign LUT_3[59026] = 32'b00000000000000010101000101001110;
assign LUT_3[59027] = 32'b00000000000000011011110000101011;
assign LUT_3[59028] = 32'b00000000000000010000001011100000;
assign LUT_3[59029] = 32'b00000000000000010110110110111101;
assign LUT_3[59030] = 32'b00000000000000010010010011000100;
assign LUT_3[59031] = 32'b00000000000000011000111110100001;
assign LUT_3[59032] = 32'b00000000000000011000010110110000;
assign LUT_3[59033] = 32'b00000000000000011111000010001101;
assign LUT_3[59034] = 32'b00000000000000011010011110010100;
assign LUT_3[59035] = 32'b00000000000000100001001001110001;
assign LUT_3[59036] = 32'b00000000000000010101100100100110;
assign LUT_3[59037] = 32'b00000000000000011100010000000011;
assign LUT_3[59038] = 32'b00000000000000010111101100001010;
assign LUT_3[59039] = 32'b00000000000000011110010111100111;
assign LUT_3[59040] = 32'b00000000000000010000111001000111;
assign LUT_3[59041] = 32'b00000000000000010111100100100100;
assign LUT_3[59042] = 32'b00000000000000010011000000101011;
assign LUT_3[59043] = 32'b00000000000000011001101100001000;
assign LUT_3[59044] = 32'b00000000000000001110000110111101;
assign LUT_3[59045] = 32'b00000000000000010100110010011010;
assign LUT_3[59046] = 32'b00000000000000010000001110100001;
assign LUT_3[59047] = 32'b00000000000000010110111001111110;
assign LUT_3[59048] = 32'b00000000000000010110010010001101;
assign LUT_3[59049] = 32'b00000000000000011100111101101010;
assign LUT_3[59050] = 32'b00000000000000011000011001110001;
assign LUT_3[59051] = 32'b00000000000000011111000101001110;
assign LUT_3[59052] = 32'b00000000000000010011100000000011;
assign LUT_3[59053] = 32'b00000000000000011010001011100000;
assign LUT_3[59054] = 32'b00000000000000010101100111100111;
assign LUT_3[59055] = 32'b00000000000000011100010011000100;
assign LUT_3[59056] = 32'b00000000000000010100001100001010;
assign LUT_3[59057] = 32'b00000000000000011010110111100111;
assign LUT_3[59058] = 32'b00000000000000010110010011101110;
assign LUT_3[59059] = 32'b00000000000000011100111111001011;
assign LUT_3[59060] = 32'b00000000000000010001011010000000;
assign LUT_3[59061] = 32'b00000000000000011000000101011101;
assign LUT_3[59062] = 32'b00000000000000010011100001100100;
assign LUT_3[59063] = 32'b00000000000000011010001101000001;
assign LUT_3[59064] = 32'b00000000000000011001100101010000;
assign LUT_3[59065] = 32'b00000000000000100000010000101101;
assign LUT_3[59066] = 32'b00000000000000011011101100110100;
assign LUT_3[59067] = 32'b00000000000000100010011000010001;
assign LUT_3[59068] = 32'b00000000000000010110110011000110;
assign LUT_3[59069] = 32'b00000000000000011101011110100011;
assign LUT_3[59070] = 32'b00000000000000011000111010101010;
assign LUT_3[59071] = 32'b00000000000000011111100110000111;
assign LUT_3[59072] = 32'b00000000000000001111100011010010;
assign LUT_3[59073] = 32'b00000000000000010110001110101111;
assign LUT_3[59074] = 32'b00000000000000010001101010110110;
assign LUT_3[59075] = 32'b00000000000000011000010110010011;
assign LUT_3[59076] = 32'b00000000000000001100110001001000;
assign LUT_3[59077] = 32'b00000000000000010011011100100101;
assign LUT_3[59078] = 32'b00000000000000001110111000101100;
assign LUT_3[59079] = 32'b00000000000000010101100100001001;
assign LUT_3[59080] = 32'b00000000000000010100111100011000;
assign LUT_3[59081] = 32'b00000000000000011011100111110101;
assign LUT_3[59082] = 32'b00000000000000010111000011111100;
assign LUT_3[59083] = 32'b00000000000000011101101111011001;
assign LUT_3[59084] = 32'b00000000000000010010001010001110;
assign LUT_3[59085] = 32'b00000000000000011000110101101011;
assign LUT_3[59086] = 32'b00000000000000010100010001110010;
assign LUT_3[59087] = 32'b00000000000000011010111101001111;
assign LUT_3[59088] = 32'b00000000000000010010110110010101;
assign LUT_3[59089] = 32'b00000000000000011001100001110010;
assign LUT_3[59090] = 32'b00000000000000010100111101111001;
assign LUT_3[59091] = 32'b00000000000000011011101001010110;
assign LUT_3[59092] = 32'b00000000000000010000000100001011;
assign LUT_3[59093] = 32'b00000000000000010110101111101000;
assign LUT_3[59094] = 32'b00000000000000010010001011101111;
assign LUT_3[59095] = 32'b00000000000000011000110111001100;
assign LUT_3[59096] = 32'b00000000000000011000001111011011;
assign LUT_3[59097] = 32'b00000000000000011110111010111000;
assign LUT_3[59098] = 32'b00000000000000011010010110111111;
assign LUT_3[59099] = 32'b00000000000000100001000010011100;
assign LUT_3[59100] = 32'b00000000000000010101011101010001;
assign LUT_3[59101] = 32'b00000000000000011100001000101110;
assign LUT_3[59102] = 32'b00000000000000010111100100110101;
assign LUT_3[59103] = 32'b00000000000000011110010000010010;
assign LUT_3[59104] = 32'b00000000000000010000110001110010;
assign LUT_3[59105] = 32'b00000000000000010111011101001111;
assign LUT_3[59106] = 32'b00000000000000010010111001010110;
assign LUT_3[59107] = 32'b00000000000000011001100100110011;
assign LUT_3[59108] = 32'b00000000000000001101111111101000;
assign LUT_3[59109] = 32'b00000000000000010100101011000101;
assign LUT_3[59110] = 32'b00000000000000010000000111001100;
assign LUT_3[59111] = 32'b00000000000000010110110010101001;
assign LUT_3[59112] = 32'b00000000000000010110001010111000;
assign LUT_3[59113] = 32'b00000000000000011100110110010101;
assign LUT_3[59114] = 32'b00000000000000011000010010011100;
assign LUT_3[59115] = 32'b00000000000000011110111101111001;
assign LUT_3[59116] = 32'b00000000000000010011011000101110;
assign LUT_3[59117] = 32'b00000000000000011010000100001011;
assign LUT_3[59118] = 32'b00000000000000010101100000010010;
assign LUT_3[59119] = 32'b00000000000000011100001011101111;
assign LUT_3[59120] = 32'b00000000000000010100000100110101;
assign LUT_3[59121] = 32'b00000000000000011010110000010010;
assign LUT_3[59122] = 32'b00000000000000010110001100011001;
assign LUT_3[59123] = 32'b00000000000000011100110111110110;
assign LUT_3[59124] = 32'b00000000000000010001010010101011;
assign LUT_3[59125] = 32'b00000000000000010111111110001000;
assign LUT_3[59126] = 32'b00000000000000010011011010001111;
assign LUT_3[59127] = 32'b00000000000000011010000101101100;
assign LUT_3[59128] = 32'b00000000000000011001011101111011;
assign LUT_3[59129] = 32'b00000000000000100000001001011000;
assign LUT_3[59130] = 32'b00000000000000011011100101011111;
assign LUT_3[59131] = 32'b00000000000000100010010000111100;
assign LUT_3[59132] = 32'b00000000000000010110101011110001;
assign LUT_3[59133] = 32'b00000000000000011101010111001110;
assign LUT_3[59134] = 32'b00000000000000011000110011010101;
assign LUT_3[59135] = 32'b00000000000000011111011110110010;
assign LUT_3[59136] = 32'b00000000000000001001101111001010;
assign LUT_3[59137] = 32'b00000000000000010000011010100111;
assign LUT_3[59138] = 32'b00000000000000001011110110101110;
assign LUT_3[59139] = 32'b00000000000000010010100010001011;
assign LUT_3[59140] = 32'b00000000000000000110111101000000;
assign LUT_3[59141] = 32'b00000000000000001101101000011101;
assign LUT_3[59142] = 32'b00000000000000001001000100100100;
assign LUT_3[59143] = 32'b00000000000000001111110000000001;
assign LUT_3[59144] = 32'b00000000000000001111001000010000;
assign LUT_3[59145] = 32'b00000000000000010101110011101101;
assign LUT_3[59146] = 32'b00000000000000010001001111110100;
assign LUT_3[59147] = 32'b00000000000000010111111011010001;
assign LUT_3[59148] = 32'b00000000000000001100010110000110;
assign LUT_3[59149] = 32'b00000000000000010011000001100011;
assign LUT_3[59150] = 32'b00000000000000001110011101101010;
assign LUT_3[59151] = 32'b00000000000000010101001001000111;
assign LUT_3[59152] = 32'b00000000000000001101000010001101;
assign LUT_3[59153] = 32'b00000000000000010011101101101010;
assign LUT_3[59154] = 32'b00000000000000001111001001110001;
assign LUT_3[59155] = 32'b00000000000000010101110101001110;
assign LUT_3[59156] = 32'b00000000000000001010010000000011;
assign LUT_3[59157] = 32'b00000000000000010000111011100000;
assign LUT_3[59158] = 32'b00000000000000001100010111100111;
assign LUT_3[59159] = 32'b00000000000000010011000011000100;
assign LUT_3[59160] = 32'b00000000000000010010011011010011;
assign LUT_3[59161] = 32'b00000000000000011001000110110000;
assign LUT_3[59162] = 32'b00000000000000010100100010110111;
assign LUT_3[59163] = 32'b00000000000000011011001110010100;
assign LUT_3[59164] = 32'b00000000000000001111101001001001;
assign LUT_3[59165] = 32'b00000000000000010110010100100110;
assign LUT_3[59166] = 32'b00000000000000010001110000101101;
assign LUT_3[59167] = 32'b00000000000000011000011100001010;
assign LUT_3[59168] = 32'b00000000000000001010111101101010;
assign LUT_3[59169] = 32'b00000000000000010001101001000111;
assign LUT_3[59170] = 32'b00000000000000001101000101001110;
assign LUT_3[59171] = 32'b00000000000000010011110000101011;
assign LUT_3[59172] = 32'b00000000000000001000001011100000;
assign LUT_3[59173] = 32'b00000000000000001110110110111101;
assign LUT_3[59174] = 32'b00000000000000001010010011000100;
assign LUT_3[59175] = 32'b00000000000000010000111110100001;
assign LUT_3[59176] = 32'b00000000000000010000010110110000;
assign LUT_3[59177] = 32'b00000000000000010111000010001101;
assign LUT_3[59178] = 32'b00000000000000010010011110010100;
assign LUT_3[59179] = 32'b00000000000000011001001001110001;
assign LUT_3[59180] = 32'b00000000000000001101100100100110;
assign LUT_3[59181] = 32'b00000000000000010100010000000011;
assign LUT_3[59182] = 32'b00000000000000001111101100001010;
assign LUT_3[59183] = 32'b00000000000000010110010111100111;
assign LUT_3[59184] = 32'b00000000000000001110010000101101;
assign LUT_3[59185] = 32'b00000000000000010100111100001010;
assign LUT_3[59186] = 32'b00000000000000010000011000010001;
assign LUT_3[59187] = 32'b00000000000000010111000011101110;
assign LUT_3[59188] = 32'b00000000000000001011011110100011;
assign LUT_3[59189] = 32'b00000000000000010010001010000000;
assign LUT_3[59190] = 32'b00000000000000001101100110000111;
assign LUT_3[59191] = 32'b00000000000000010100010001100100;
assign LUT_3[59192] = 32'b00000000000000010011101001110011;
assign LUT_3[59193] = 32'b00000000000000011010010101010000;
assign LUT_3[59194] = 32'b00000000000000010101110001010111;
assign LUT_3[59195] = 32'b00000000000000011100011100110100;
assign LUT_3[59196] = 32'b00000000000000010000110111101001;
assign LUT_3[59197] = 32'b00000000000000010111100011000110;
assign LUT_3[59198] = 32'b00000000000000010010111111001101;
assign LUT_3[59199] = 32'b00000000000000011001101010101010;
assign LUT_3[59200] = 32'b00000000000000001001100111110101;
assign LUT_3[59201] = 32'b00000000000000010000010011010010;
assign LUT_3[59202] = 32'b00000000000000001011101111011001;
assign LUT_3[59203] = 32'b00000000000000010010011010110110;
assign LUT_3[59204] = 32'b00000000000000000110110101101011;
assign LUT_3[59205] = 32'b00000000000000001101100001001000;
assign LUT_3[59206] = 32'b00000000000000001000111101001111;
assign LUT_3[59207] = 32'b00000000000000001111101000101100;
assign LUT_3[59208] = 32'b00000000000000001111000000111011;
assign LUT_3[59209] = 32'b00000000000000010101101100011000;
assign LUT_3[59210] = 32'b00000000000000010001001000011111;
assign LUT_3[59211] = 32'b00000000000000010111110011111100;
assign LUT_3[59212] = 32'b00000000000000001100001110110001;
assign LUT_3[59213] = 32'b00000000000000010010111010001110;
assign LUT_3[59214] = 32'b00000000000000001110010110010101;
assign LUT_3[59215] = 32'b00000000000000010101000001110010;
assign LUT_3[59216] = 32'b00000000000000001100111010111000;
assign LUT_3[59217] = 32'b00000000000000010011100110010101;
assign LUT_3[59218] = 32'b00000000000000001111000010011100;
assign LUT_3[59219] = 32'b00000000000000010101101101111001;
assign LUT_3[59220] = 32'b00000000000000001010001000101110;
assign LUT_3[59221] = 32'b00000000000000010000110100001011;
assign LUT_3[59222] = 32'b00000000000000001100010000010010;
assign LUT_3[59223] = 32'b00000000000000010010111011101111;
assign LUT_3[59224] = 32'b00000000000000010010010011111110;
assign LUT_3[59225] = 32'b00000000000000011000111111011011;
assign LUT_3[59226] = 32'b00000000000000010100011011100010;
assign LUT_3[59227] = 32'b00000000000000011011000110111111;
assign LUT_3[59228] = 32'b00000000000000001111100001110100;
assign LUT_3[59229] = 32'b00000000000000010110001101010001;
assign LUT_3[59230] = 32'b00000000000000010001101001011000;
assign LUT_3[59231] = 32'b00000000000000011000010100110101;
assign LUT_3[59232] = 32'b00000000000000001010110110010101;
assign LUT_3[59233] = 32'b00000000000000010001100001110010;
assign LUT_3[59234] = 32'b00000000000000001100111101111001;
assign LUT_3[59235] = 32'b00000000000000010011101001010110;
assign LUT_3[59236] = 32'b00000000000000001000000100001011;
assign LUT_3[59237] = 32'b00000000000000001110101111101000;
assign LUT_3[59238] = 32'b00000000000000001010001011101111;
assign LUT_3[59239] = 32'b00000000000000010000110111001100;
assign LUT_3[59240] = 32'b00000000000000010000001111011011;
assign LUT_3[59241] = 32'b00000000000000010110111010111000;
assign LUT_3[59242] = 32'b00000000000000010010010110111111;
assign LUT_3[59243] = 32'b00000000000000011001000010011100;
assign LUT_3[59244] = 32'b00000000000000001101011101010001;
assign LUT_3[59245] = 32'b00000000000000010100001000101110;
assign LUT_3[59246] = 32'b00000000000000001111100100110101;
assign LUT_3[59247] = 32'b00000000000000010110010000010010;
assign LUT_3[59248] = 32'b00000000000000001110001001011000;
assign LUT_3[59249] = 32'b00000000000000010100110100110101;
assign LUT_3[59250] = 32'b00000000000000010000010000111100;
assign LUT_3[59251] = 32'b00000000000000010110111100011001;
assign LUT_3[59252] = 32'b00000000000000001011010111001110;
assign LUT_3[59253] = 32'b00000000000000010010000010101011;
assign LUT_3[59254] = 32'b00000000000000001101011110110010;
assign LUT_3[59255] = 32'b00000000000000010100001010001111;
assign LUT_3[59256] = 32'b00000000000000010011100010011110;
assign LUT_3[59257] = 32'b00000000000000011010001101111011;
assign LUT_3[59258] = 32'b00000000000000010101101010000010;
assign LUT_3[59259] = 32'b00000000000000011100010101011111;
assign LUT_3[59260] = 32'b00000000000000010000110000010100;
assign LUT_3[59261] = 32'b00000000000000010111011011110001;
assign LUT_3[59262] = 32'b00000000000000010010110111111000;
assign LUT_3[59263] = 32'b00000000000000011001100011010101;
assign LUT_3[59264] = 32'b00000000000000001011111010001000;
assign LUT_3[59265] = 32'b00000000000000010010100101100101;
assign LUT_3[59266] = 32'b00000000000000001110000001101100;
assign LUT_3[59267] = 32'b00000000000000010100101101001001;
assign LUT_3[59268] = 32'b00000000000000001001000111111110;
assign LUT_3[59269] = 32'b00000000000000001111110011011011;
assign LUT_3[59270] = 32'b00000000000000001011001111100010;
assign LUT_3[59271] = 32'b00000000000000010001111010111111;
assign LUT_3[59272] = 32'b00000000000000010001010011001110;
assign LUT_3[59273] = 32'b00000000000000010111111110101011;
assign LUT_3[59274] = 32'b00000000000000010011011010110010;
assign LUT_3[59275] = 32'b00000000000000011010000110001111;
assign LUT_3[59276] = 32'b00000000000000001110100001000100;
assign LUT_3[59277] = 32'b00000000000000010101001100100001;
assign LUT_3[59278] = 32'b00000000000000010000101000101000;
assign LUT_3[59279] = 32'b00000000000000010111010100000101;
assign LUT_3[59280] = 32'b00000000000000001111001101001011;
assign LUT_3[59281] = 32'b00000000000000010101111000101000;
assign LUT_3[59282] = 32'b00000000000000010001010100101111;
assign LUT_3[59283] = 32'b00000000000000011000000000001100;
assign LUT_3[59284] = 32'b00000000000000001100011011000001;
assign LUT_3[59285] = 32'b00000000000000010011000110011110;
assign LUT_3[59286] = 32'b00000000000000001110100010100101;
assign LUT_3[59287] = 32'b00000000000000010101001110000010;
assign LUT_3[59288] = 32'b00000000000000010100100110010001;
assign LUT_3[59289] = 32'b00000000000000011011010001101110;
assign LUT_3[59290] = 32'b00000000000000010110101101110101;
assign LUT_3[59291] = 32'b00000000000000011101011001010010;
assign LUT_3[59292] = 32'b00000000000000010001110100000111;
assign LUT_3[59293] = 32'b00000000000000011000011111100100;
assign LUT_3[59294] = 32'b00000000000000010011111011101011;
assign LUT_3[59295] = 32'b00000000000000011010100111001000;
assign LUT_3[59296] = 32'b00000000000000001101001000101000;
assign LUT_3[59297] = 32'b00000000000000010011110100000101;
assign LUT_3[59298] = 32'b00000000000000001111010000001100;
assign LUT_3[59299] = 32'b00000000000000010101111011101001;
assign LUT_3[59300] = 32'b00000000000000001010010110011110;
assign LUT_3[59301] = 32'b00000000000000010001000001111011;
assign LUT_3[59302] = 32'b00000000000000001100011110000010;
assign LUT_3[59303] = 32'b00000000000000010011001001011111;
assign LUT_3[59304] = 32'b00000000000000010010100001101110;
assign LUT_3[59305] = 32'b00000000000000011001001101001011;
assign LUT_3[59306] = 32'b00000000000000010100101001010010;
assign LUT_3[59307] = 32'b00000000000000011011010100101111;
assign LUT_3[59308] = 32'b00000000000000001111101111100100;
assign LUT_3[59309] = 32'b00000000000000010110011011000001;
assign LUT_3[59310] = 32'b00000000000000010001110111001000;
assign LUT_3[59311] = 32'b00000000000000011000100010100101;
assign LUT_3[59312] = 32'b00000000000000010000011011101011;
assign LUT_3[59313] = 32'b00000000000000010111000111001000;
assign LUT_3[59314] = 32'b00000000000000010010100011001111;
assign LUT_3[59315] = 32'b00000000000000011001001110101100;
assign LUT_3[59316] = 32'b00000000000000001101101001100001;
assign LUT_3[59317] = 32'b00000000000000010100010100111110;
assign LUT_3[59318] = 32'b00000000000000001111110001000101;
assign LUT_3[59319] = 32'b00000000000000010110011100100010;
assign LUT_3[59320] = 32'b00000000000000010101110100110001;
assign LUT_3[59321] = 32'b00000000000000011100100000001110;
assign LUT_3[59322] = 32'b00000000000000010111111100010101;
assign LUT_3[59323] = 32'b00000000000000011110100111110010;
assign LUT_3[59324] = 32'b00000000000000010011000010100111;
assign LUT_3[59325] = 32'b00000000000000011001101110000100;
assign LUT_3[59326] = 32'b00000000000000010101001010001011;
assign LUT_3[59327] = 32'b00000000000000011011110101101000;
assign LUT_3[59328] = 32'b00000000000000001011110010110011;
assign LUT_3[59329] = 32'b00000000000000010010011110010000;
assign LUT_3[59330] = 32'b00000000000000001101111010010111;
assign LUT_3[59331] = 32'b00000000000000010100100101110100;
assign LUT_3[59332] = 32'b00000000000000001001000000101001;
assign LUT_3[59333] = 32'b00000000000000001111101100000110;
assign LUT_3[59334] = 32'b00000000000000001011001000001101;
assign LUT_3[59335] = 32'b00000000000000010001110011101010;
assign LUT_3[59336] = 32'b00000000000000010001001011111001;
assign LUT_3[59337] = 32'b00000000000000010111110111010110;
assign LUT_3[59338] = 32'b00000000000000010011010011011101;
assign LUT_3[59339] = 32'b00000000000000011001111110111010;
assign LUT_3[59340] = 32'b00000000000000001110011001101111;
assign LUT_3[59341] = 32'b00000000000000010101000101001100;
assign LUT_3[59342] = 32'b00000000000000010000100001010011;
assign LUT_3[59343] = 32'b00000000000000010111001100110000;
assign LUT_3[59344] = 32'b00000000000000001111000101110110;
assign LUT_3[59345] = 32'b00000000000000010101110001010011;
assign LUT_3[59346] = 32'b00000000000000010001001101011010;
assign LUT_3[59347] = 32'b00000000000000010111111000110111;
assign LUT_3[59348] = 32'b00000000000000001100010011101100;
assign LUT_3[59349] = 32'b00000000000000010010111111001001;
assign LUT_3[59350] = 32'b00000000000000001110011011010000;
assign LUT_3[59351] = 32'b00000000000000010101000110101101;
assign LUT_3[59352] = 32'b00000000000000010100011110111100;
assign LUT_3[59353] = 32'b00000000000000011011001010011001;
assign LUT_3[59354] = 32'b00000000000000010110100110100000;
assign LUT_3[59355] = 32'b00000000000000011101010001111101;
assign LUT_3[59356] = 32'b00000000000000010001101100110010;
assign LUT_3[59357] = 32'b00000000000000011000011000001111;
assign LUT_3[59358] = 32'b00000000000000010011110100010110;
assign LUT_3[59359] = 32'b00000000000000011010011111110011;
assign LUT_3[59360] = 32'b00000000000000001101000001010011;
assign LUT_3[59361] = 32'b00000000000000010011101100110000;
assign LUT_3[59362] = 32'b00000000000000001111001000110111;
assign LUT_3[59363] = 32'b00000000000000010101110100010100;
assign LUT_3[59364] = 32'b00000000000000001010001111001001;
assign LUT_3[59365] = 32'b00000000000000010000111010100110;
assign LUT_3[59366] = 32'b00000000000000001100010110101101;
assign LUT_3[59367] = 32'b00000000000000010011000010001010;
assign LUT_3[59368] = 32'b00000000000000010010011010011001;
assign LUT_3[59369] = 32'b00000000000000011001000101110110;
assign LUT_3[59370] = 32'b00000000000000010100100001111101;
assign LUT_3[59371] = 32'b00000000000000011011001101011010;
assign LUT_3[59372] = 32'b00000000000000001111101000001111;
assign LUT_3[59373] = 32'b00000000000000010110010011101100;
assign LUT_3[59374] = 32'b00000000000000010001101111110011;
assign LUT_3[59375] = 32'b00000000000000011000011011010000;
assign LUT_3[59376] = 32'b00000000000000010000010100010110;
assign LUT_3[59377] = 32'b00000000000000010110111111110011;
assign LUT_3[59378] = 32'b00000000000000010010011011111010;
assign LUT_3[59379] = 32'b00000000000000011001000111010111;
assign LUT_3[59380] = 32'b00000000000000001101100010001100;
assign LUT_3[59381] = 32'b00000000000000010100001101101001;
assign LUT_3[59382] = 32'b00000000000000001111101001110000;
assign LUT_3[59383] = 32'b00000000000000010110010101001101;
assign LUT_3[59384] = 32'b00000000000000010101101101011100;
assign LUT_3[59385] = 32'b00000000000000011100011000111001;
assign LUT_3[59386] = 32'b00000000000000010111110101000000;
assign LUT_3[59387] = 32'b00000000000000011110100000011101;
assign LUT_3[59388] = 32'b00000000000000010010111011010010;
assign LUT_3[59389] = 32'b00000000000000011001100110101111;
assign LUT_3[59390] = 32'b00000000000000010101000010110110;
assign LUT_3[59391] = 32'b00000000000000011011101110010011;
assign LUT_3[59392] = 32'b00000000000000000101011011101110;
assign LUT_3[59393] = 32'b00000000000000001100000111001011;
assign LUT_3[59394] = 32'b00000000000000000111100011010010;
assign LUT_3[59395] = 32'b00000000000000001110001110101111;
assign LUT_3[59396] = 32'b00000000000000000010101001100100;
assign LUT_3[59397] = 32'b00000000000000001001010101000001;
assign LUT_3[59398] = 32'b00000000000000000100110001001000;
assign LUT_3[59399] = 32'b00000000000000001011011100100101;
assign LUT_3[59400] = 32'b00000000000000001010110100110100;
assign LUT_3[59401] = 32'b00000000000000010001100000010001;
assign LUT_3[59402] = 32'b00000000000000001100111100011000;
assign LUT_3[59403] = 32'b00000000000000010011100111110101;
assign LUT_3[59404] = 32'b00000000000000001000000010101010;
assign LUT_3[59405] = 32'b00000000000000001110101110000111;
assign LUT_3[59406] = 32'b00000000000000001010001010001110;
assign LUT_3[59407] = 32'b00000000000000010000110101101011;
assign LUT_3[59408] = 32'b00000000000000001000101110110001;
assign LUT_3[59409] = 32'b00000000000000001111011010001110;
assign LUT_3[59410] = 32'b00000000000000001010110110010101;
assign LUT_3[59411] = 32'b00000000000000010001100001110010;
assign LUT_3[59412] = 32'b00000000000000000101111100100111;
assign LUT_3[59413] = 32'b00000000000000001100101000000100;
assign LUT_3[59414] = 32'b00000000000000001000000100001011;
assign LUT_3[59415] = 32'b00000000000000001110101111101000;
assign LUT_3[59416] = 32'b00000000000000001110000111110111;
assign LUT_3[59417] = 32'b00000000000000010100110011010100;
assign LUT_3[59418] = 32'b00000000000000010000001111011011;
assign LUT_3[59419] = 32'b00000000000000010110111010111000;
assign LUT_3[59420] = 32'b00000000000000001011010101101101;
assign LUT_3[59421] = 32'b00000000000000010010000001001010;
assign LUT_3[59422] = 32'b00000000000000001101011101010001;
assign LUT_3[59423] = 32'b00000000000000010100001000101110;
assign LUT_3[59424] = 32'b00000000000000000110101010001110;
assign LUT_3[59425] = 32'b00000000000000001101010101101011;
assign LUT_3[59426] = 32'b00000000000000001000110001110010;
assign LUT_3[59427] = 32'b00000000000000001111011101001111;
assign LUT_3[59428] = 32'b00000000000000000011111000000100;
assign LUT_3[59429] = 32'b00000000000000001010100011100001;
assign LUT_3[59430] = 32'b00000000000000000101111111101000;
assign LUT_3[59431] = 32'b00000000000000001100101011000101;
assign LUT_3[59432] = 32'b00000000000000001100000011010100;
assign LUT_3[59433] = 32'b00000000000000010010101110110001;
assign LUT_3[59434] = 32'b00000000000000001110001010111000;
assign LUT_3[59435] = 32'b00000000000000010100110110010101;
assign LUT_3[59436] = 32'b00000000000000001001010001001010;
assign LUT_3[59437] = 32'b00000000000000001111111100100111;
assign LUT_3[59438] = 32'b00000000000000001011011000101110;
assign LUT_3[59439] = 32'b00000000000000010010000100001011;
assign LUT_3[59440] = 32'b00000000000000001001111101010001;
assign LUT_3[59441] = 32'b00000000000000010000101000101110;
assign LUT_3[59442] = 32'b00000000000000001100000100110101;
assign LUT_3[59443] = 32'b00000000000000010010110000010010;
assign LUT_3[59444] = 32'b00000000000000000111001011000111;
assign LUT_3[59445] = 32'b00000000000000001101110110100100;
assign LUT_3[59446] = 32'b00000000000000001001010010101011;
assign LUT_3[59447] = 32'b00000000000000001111111110001000;
assign LUT_3[59448] = 32'b00000000000000001111010110010111;
assign LUT_3[59449] = 32'b00000000000000010110000001110100;
assign LUT_3[59450] = 32'b00000000000000010001011101111011;
assign LUT_3[59451] = 32'b00000000000000011000001001011000;
assign LUT_3[59452] = 32'b00000000000000001100100100001101;
assign LUT_3[59453] = 32'b00000000000000010011001111101010;
assign LUT_3[59454] = 32'b00000000000000001110101011110001;
assign LUT_3[59455] = 32'b00000000000000010101010111001110;
assign LUT_3[59456] = 32'b00000000000000000101010100011001;
assign LUT_3[59457] = 32'b00000000000000001011111111110110;
assign LUT_3[59458] = 32'b00000000000000000111011011111101;
assign LUT_3[59459] = 32'b00000000000000001110000111011010;
assign LUT_3[59460] = 32'b00000000000000000010100010001111;
assign LUT_3[59461] = 32'b00000000000000001001001101101100;
assign LUT_3[59462] = 32'b00000000000000000100101001110011;
assign LUT_3[59463] = 32'b00000000000000001011010101010000;
assign LUT_3[59464] = 32'b00000000000000001010101101011111;
assign LUT_3[59465] = 32'b00000000000000010001011000111100;
assign LUT_3[59466] = 32'b00000000000000001100110101000011;
assign LUT_3[59467] = 32'b00000000000000010011100000100000;
assign LUT_3[59468] = 32'b00000000000000000111111011010101;
assign LUT_3[59469] = 32'b00000000000000001110100110110010;
assign LUT_3[59470] = 32'b00000000000000001010000010111001;
assign LUT_3[59471] = 32'b00000000000000010000101110010110;
assign LUT_3[59472] = 32'b00000000000000001000100111011100;
assign LUT_3[59473] = 32'b00000000000000001111010010111001;
assign LUT_3[59474] = 32'b00000000000000001010101111000000;
assign LUT_3[59475] = 32'b00000000000000010001011010011101;
assign LUT_3[59476] = 32'b00000000000000000101110101010010;
assign LUT_3[59477] = 32'b00000000000000001100100000101111;
assign LUT_3[59478] = 32'b00000000000000000111111100110110;
assign LUT_3[59479] = 32'b00000000000000001110101000010011;
assign LUT_3[59480] = 32'b00000000000000001110000000100010;
assign LUT_3[59481] = 32'b00000000000000010100101011111111;
assign LUT_3[59482] = 32'b00000000000000010000001000000110;
assign LUT_3[59483] = 32'b00000000000000010110110011100011;
assign LUT_3[59484] = 32'b00000000000000001011001110011000;
assign LUT_3[59485] = 32'b00000000000000010001111001110101;
assign LUT_3[59486] = 32'b00000000000000001101010101111100;
assign LUT_3[59487] = 32'b00000000000000010100000001011001;
assign LUT_3[59488] = 32'b00000000000000000110100010111001;
assign LUT_3[59489] = 32'b00000000000000001101001110010110;
assign LUT_3[59490] = 32'b00000000000000001000101010011101;
assign LUT_3[59491] = 32'b00000000000000001111010101111010;
assign LUT_3[59492] = 32'b00000000000000000011110000101111;
assign LUT_3[59493] = 32'b00000000000000001010011100001100;
assign LUT_3[59494] = 32'b00000000000000000101111000010011;
assign LUT_3[59495] = 32'b00000000000000001100100011110000;
assign LUT_3[59496] = 32'b00000000000000001011111011111111;
assign LUT_3[59497] = 32'b00000000000000010010100111011100;
assign LUT_3[59498] = 32'b00000000000000001110000011100011;
assign LUT_3[59499] = 32'b00000000000000010100101111000000;
assign LUT_3[59500] = 32'b00000000000000001001001001110101;
assign LUT_3[59501] = 32'b00000000000000001111110101010010;
assign LUT_3[59502] = 32'b00000000000000001011010001011001;
assign LUT_3[59503] = 32'b00000000000000010001111100110110;
assign LUT_3[59504] = 32'b00000000000000001001110101111100;
assign LUT_3[59505] = 32'b00000000000000010000100001011001;
assign LUT_3[59506] = 32'b00000000000000001011111101100000;
assign LUT_3[59507] = 32'b00000000000000010010101000111101;
assign LUT_3[59508] = 32'b00000000000000000111000011110010;
assign LUT_3[59509] = 32'b00000000000000001101101111001111;
assign LUT_3[59510] = 32'b00000000000000001001001011010110;
assign LUT_3[59511] = 32'b00000000000000001111110110110011;
assign LUT_3[59512] = 32'b00000000000000001111001111000010;
assign LUT_3[59513] = 32'b00000000000000010101111010011111;
assign LUT_3[59514] = 32'b00000000000000010001010110100110;
assign LUT_3[59515] = 32'b00000000000000011000000010000011;
assign LUT_3[59516] = 32'b00000000000000001100011100111000;
assign LUT_3[59517] = 32'b00000000000000010011001000010101;
assign LUT_3[59518] = 32'b00000000000000001110100100011100;
assign LUT_3[59519] = 32'b00000000000000010101001111111001;
assign LUT_3[59520] = 32'b00000000000000000111100110101100;
assign LUT_3[59521] = 32'b00000000000000001110010010001001;
assign LUT_3[59522] = 32'b00000000000000001001101110010000;
assign LUT_3[59523] = 32'b00000000000000010000011001101101;
assign LUT_3[59524] = 32'b00000000000000000100110100100010;
assign LUT_3[59525] = 32'b00000000000000001011011111111111;
assign LUT_3[59526] = 32'b00000000000000000110111100000110;
assign LUT_3[59527] = 32'b00000000000000001101100111100011;
assign LUT_3[59528] = 32'b00000000000000001100111111110010;
assign LUT_3[59529] = 32'b00000000000000010011101011001111;
assign LUT_3[59530] = 32'b00000000000000001111000111010110;
assign LUT_3[59531] = 32'b00000000000000010101110010110011;
assign LUT_3[59532] = 32'b00000000000000001010001101101000;
assign LUT_3[59533] = 32'b00000000000000010000111001000101;
assign LUT_3[59534] = 32'b00000000000000001100010101001100;
assign LUT_3[59535] = 32'b00000000000000010011000000101001;
assign LUT_3[59536] = 32'b00000000000000001010111001101111;
assign LUT_3[59537] = 32'b00000000000000010001100101001100;
assign LUT_3[59538] = 32'b00000000000000001101000001010011;
assign LUT_3[59539] = 32'b00000000000000010011101100110000;
assign LUT_3[59540] = 32'b00000000000000001000000111100101;
assign LUT_3[59541] = 32'b00000000000000001110110011000010;
assign LUT_3[59542] = 32'b00000000000000001010001111001001;
assign LUT_3[59543] = 32'b00000000000000010000111010100110;
assign LUT_3[59544] = 32'b00000000000000010000010010110101;
assign LUT_3[59545] = 32'b00000000000000010110111110010010;
assign LUT_3[59546] = 32'b00000000000000010010011010011001;
assign LUT_3[59547] = 32'b00000000000000011001000101110110;
assign LUT_3[59548] = 32'b00000000000000001101100000101011;
assign LUT_3[59549] = 32'b00000000000000010100001100001000;
assign LUT_3[59550] = 32'b00000000000000001111101000001111;
assign LUT_3[59551] = 32'b00000000000000010110010011101100;
assign LUT_3[59552] = 32'b00000000000000001000110101001100;
assign LUT_3[59553] = 32'b00000000000000001111100000101001;
assign LUT_3[59554] = 32'b00000000000000001010111100110000;
assign LUT_3[59555] = 32'b00000000000000010001101000001101;
assign LUT_3[59556] = 32'b00000000000000000110000011000010;
assign LUT_3[59557] = 32'b00000000000000001100101110011111;
assign LUT_3[59558] = 32'b00000000000000001000001010100110;
assign LUT_3[59559] = 32'b00000000000000001110110110000011;
assign LUT_3[59560] = 32'b00000000000000001110001110010010;
assign LUT_3[59561] = 32'b00000000000000010100111001101111;
assign LUT_3[59562] = 32'b00000000000000010000010101110110;
assign LUT_3[59563] = 32'b00000000000000010111000001010011;
assign LUT_3[59564] = 32'b00000000000000001011011100001000;
assign LUT_3[59565] = 32'b00000000000000010010000111100101;
assign LUT_3[59566] = 32'b00000000000000001101100011101100;
assign LUT_3[59567] = 32'b00000000000000010100001111001001;
assign LUT_3[59568] = 32'b00000000000000001100001000001111;
assign LUT_3[59569] = 32'b00000000000000010010110011101100;
assign LUT_3[59570] = 32'b00000000000000001110001111110011;
assign LUT_3[59571] = 32'b00000000000000010100111011010000;
assign LUT_3[59572] = 32'b00000000000000001001010110000101;
assign LUT_3[59573] = 32'b00000000000000010000000001100010;
assign LUT_3[59574] = 32'b00000000000000001011011101101001;
assign LUT_3[59575] = 32'b00000000000000010010001001000110;
assign LUT_3[59576] = 32'b00000000000000010001100001010101;
assign LUT_3[59577] = 32'b00000000000000011000001100110010;
assign LUT_3[59578] = 32'b00000000000000010011101000111001;
assign LUT_3[59579] = 32'b00000000000000011010010100010110;
assign LUT_3[59580] = 32'b00000000000000001110101111001011;
assign LUT_3[59581] = 32'b00000000000000010101011010101000;
assign LUT_3[59582] = 32'b00000000000000010000110110101111;
assign LUT_3[59583] = 32'b00000000000000010111100010001100;
assign LUT_3[59584] = 32'b00000000000000000111011111010111;
assign LUT_3[59585] = 32'b00000000000000001110001010110100;
assign LUT_3[59586] = 32'b00000000000000001001100110111011;
assign LUT_3[59587] = 32'b00000000000000010000010010011000;
assign LUT_3[59588] = 32'b00000000000000000100101101001101;
assign LUT_3[59589] = 32'b00000000000000001011011000101010;
assign LUT_3[59590] = 32'b00000000000000000110110100110001;
assign LUT_3[59591] = 32'b00000000000000001101100000001110;
assign LUT_3[59592] = 32'b00000000000000001100111000011101;
assign LUT_3[59593] = 32'b00000000000000010011100011111010;
assign LUT_3[59594] = 32'b00000000000000001111000000000001;
assign LUT_3[59595] = 32'b00000000000000010101101011011110;
assign LUT_3[59596] = 32'b00000000000000001010000110010011;
assign LUT_3[59597] = 32'b00000000000000010000110001110000;
assign LUT_3[59598] = 32'b00000000000000001100001101110111;
assign LUT_3[59599] = 32'b00000000000000010010111001010100;
assign LUT_3[59600] = 32'b00000000000000001010110010011010;
assign LUT_3[59601] = 32'b00000000000000010001011101110111;
assign LUT_3[59602] = 32'b00000000000000001100111001111110;
assign LUT_3[59603] = 32'b00000000000000010011100101011011;
assign LUT_3[59604] = 32'b00000000000000001000000000010000;
assign LUT_3[59605] = 32'b00000000000000001110101011101101;
assign LUT_3[59606] = 32'b00000000000000001010000111110100;
assign LUT_3[59607] = 32'b00000000000000010000110011010001;
assign LUT_3[59608] = 32'b00000000000000010000001011100000;
assign LUT_3[59609] = 32'b00000000000000010110110110111101;
assign LUT_3[59610] = 32'b00000000000000010010010011000100;
assign LUT_3[59611] = 32'b00000000000000011000111110100001;
assign LUT_3[59612] = 32'b00000000000000001101011001010110;
assign LUT_3[59613] = 32'b00000000000000010100000100110011;
assign LUT_3[59614] = 32'b00000000000000001111100000111010;
assign LUT_3[59615] = 32'b00000000000000010110001100010111;
assign LUT_3[59616] = 32'b00000000000000001000101101110111;
assign LUT_3[59617] = 32'b00000000000000001111011001010100;
assign LUT_3[59618] = 32'b00000000000000001010110101011011;
assign LUT_3[59619] = 32'b00000000000000010001100000111000;
assign LUT_3[59620] = 32'b00000000000000000101111011101101;
assign LUT_3[59621] = 32'b00000000000000001100100111001010;
assign LUT_3[59622] = 32'b00000000000000001000000011010001;
assign LUT_3[59623] = 32'b00000000000000001110101110101110;
assign LUT_3[59624] = 32'b00000000000000001110000110111101;
assign LUT_3[59625] = 32'b00000000000000010100110010011010;
assign LUT_3[59626] = 32'b00000000000000010000001110100001;
assign LUT_3[59627] = 32'b00000000000000010110111001111110;
assign LUT_3[59628] = 32'b00000000000000001011010100110011;
assign LUT_3[59629] = 32'b00000000000000010010000000010000;
assign LUT_3[59630] = 32'b00000000000000001101011100010111;
assign LUT_3[59631] = 32'b00000000000000010100000111110100;
assign LUT_3[59632] = 32'b00000000000000001100000000111010;
assign LUT_3[59633] = 32'b00000000000000010010101100010111;
assign LUT_3[59634] = 32'b00000000000000001110001000011110;
assign LUT_3[59635] = 32'b00000000000000010100110011111011;
assign LUT_3[59636] = 32'b00000000000000001001001110110000;
assign LUT_3[59637] = 32'b00000000000000001111111010001101;
assign LUT_3[59638] = 32'b00000000000000001011010110010100;
assign LUT_3[59639] = 32'b00000000000000010010000001110001;
assign LUT_3[59640] = 32'b00000000000000010001011010000000;
assign LUT_3[59641] = 32'b00000000000000011000000101011101;
assign LUT_3[59642] = 32'b00000000000000010011100001100100;
assign LUT_3[59643] = 32'b00000000000000011010001101000001;
assign LUT_3[59644] = 32'b00000000000000001110100111110110;
assign LUT_3[59645] = 32'b00000000000000010101010011010011;
assign LUT_3[59646] = 32'b00000000000000010000101111011010;
assign LUT_3[59647] = 32'b00000000000000010111011010110111;
assign LUT_3[59648] = 32'b00000000000000000001101011001111;
assign LUT_3[59649] = 32'b00000000000000001000010110101100;
assign LUT_3[59650] = 32'b00000000000000000011110010110011;
assign LUT_3[59651] = 32'b00000000000000001010011110010000;
assign LUT_3[59652] = 32'b11111111111111111110111001000101;
assign LUT_3[59653] = 32'b00000000000000000101100100100010;
assign LUT_3[59654] = 32'b00000000000000000001000000101001;
assign LUT_3[59655] = 32'b00000000000000000111101100000110;
assign LUT_3[59656] = 32'b00000000000000000111000100010101;
assign LUT_3[59657] = 32'b00000000000000001101101111110010;
assign LUT_3[59658] = 32'b00000000000000001001001011111001;
assign LUT_3[59659] = 32'b00000000000000001111110111010110;
assign LUT_3[59660] = 32'b00000000000000000100010010001011;
assign LUT_3[59661] = 32'b00000000000000001010111101101000;
assign LUT_3[59662] = 32'b00000000000000000110011001101111;
assign LUT_3[59663] = 32'b00000000000000001101000101001100;
assign LUT_3[59664] = 32'b00000000000000000100111110010010;
assign LUT_3[59665] = 32'b00000000000000001011101001101111;
assign LUT_3[59666] = 32'b00000000000000000111000101110110;
assign LUT_3[59667] = 32'b00000000000000001101110001010011;
assign LUT_3[59668] = 32'b00000000000000000010001100001000;
assign LUT_3[59669] = 32'b00000000000000001000110111100101;
assign LUT_3[59670] = 32'b00000000000000000100010011101100;
assign LUT_3[59671] = 32'b00000000000000001010111111001001;
assign LUT_3[59672] = 32'b00000000000000001010010111011000;
assign LUT_3[59673] = 32'b00000000000000010001000010110101;
assign LUT_3[59674] = 32'b00000000000000001100011110111100;
assign LUT_3[59675] = 32'b00000000000000010011001010011001;
assign LUT_3[59676] = 32'b00000000000000000111100101001110;
assign LUT_3[59677] = 32'b00000000000000001110010000101011;
assign LUT_3[59678] = 32'b00000000000000001001101100110010;
assign LUT_3[59679] = 32'b00000000000000010000011000001111;
assign LUT_3[59680] = 32'b00000000000000000010111001101111;
assign LUT_3[59681] = 32'b00000000000000001001100101001100;
assign LUT_3[59682] = 32'b00000000000000000101000001010011;
assign LUT_3[59683] = 32'b00000000000000001011101100110000;
assign LUT_3[59684] = 32'b00000000000000000000000111100101;
assign LUT_3[59685] = 32'b00000000000000000110110011000010;
assign LUT_3[59686] = 32'b00000000000000000010001111001001;
assign LUT_3[59687] = 32'b00000000000000001000111010100110;
assign LUT_3[59688] = 32'b00000000000000001000010010110101;
assign LUT_3[59689] = 32'b00000000000000001110111110010010;
assign LUT_3[59690] = 32'b00000000000000001010011010011001;
assign LUT_3[59691] = 32'b00000000000000010001000101110110;
assign LUT_3[59692] = 32'b00000000000000000101100000101011;
assign LUT_3[59693] = 32'b00000000000000001100001100001000;
assign LUT_3[59694] = 32'b00000000000000000111101000001111;
assign LUT_3[59695] = 32'b00000000000000001110010011101100;
assign LUT_3[59696] = 32'b00000000000000000110001100110010;
assign LUT_3[59697] = 32'b00000000000000001100111000001111;
assign LUT_3[59698] = 32'b00000000000000001000010100010110;
assign LUT_3[59699] = 32'b00000000000000001110111111110011;
assign LUT_3[59700] = 32'b00000000000000000011011010101000;
assign LUT_3[59701] = 32'b00000000000000001010000110000101;
assign LUT_3[59702] = 32'b00000000000000000101100010001100;
assign LUT_3[59703] = 32'b00000000000000001100001101101001;
assign LUT_3[59704] = 32'b00000000000000001011100101111000;
assign LUT_3[59705] = 32'b00000000000000010010010001010101;
assign LUT_3[59706] = 32'b00000000000000001101101101011100;
assign LUT_3[59707] = 32'b00000000000000010100011000111001;
assign LUT_3[59708] = 32'b00000000000000001000110011101110;
assign LUT_3[59709] = 32'b00000000000000001111011111001011;
assign LUT_3[59710] = 32'b00000000000000001010111011010010;
assign LUT_3[59711] = 32'b00000000000000010001100110101111;
assign LUT_3[59712] = 32'b00000000000000000001100011111010;
assign LUT_3[59713] = 32'b00000000000000001000001111010111;
assign LUT_3[59714] = 32'b00000000000000000011101011011110;
assign LUT_3[59715] = 32'b00000000000000001010010110111011;
assign LUT_3[59716] = 32'b11111111111111111110110001110000;
assign LUT_3[59717] = 32'b00000000000000000101011101001101;
assign LUT_3[59718] = 32'b00000000000000000000111001010100;
assign LUT_3[59719] = 32'b00000000000000000111100100110001;
assign LUT_3[59720] = 32'b00000000000000000110111101000000;
assign LUT_3[59721] = 32'b00000000000000001101101000011101;
assign LUT_3[59722] = 32'b00000000000000001001000100100100;
assign LUT_3[59723] = 32'b00000000000000001111110000000001;
assign LUT_3[59724] = 32'b00000000000000000100001010110110;
assign LUT_3[59725] = 32'b00000000000000001010110110010011;
assign LUT_3[59726] = 32'b00000000000000000110010010011010;
assign LUT_3[59727] = 32'b00000000000000001100111101110111;
assign LUT_3[59728] = 32'b00000000000000000100110110111101;
assign LUT_3[59729] = 32'b00000000000000001011100010011010;
assign LUT_3[59730] = 32'b00000000000000000110111110100001;
assign LUT_3[59731] = 32'b00000000000000001101101001111110;
assign LUT_3[59732] = 32'b00000000000000000010000100110011;
assign LUT_3[59733] = 32'b00000000000000001000110000010000;
assign LUT_3[59734] = 32'b00000000000000000100001100010111;
assign LUT_3[59735] = 32'b00000000000000001010110111110100;
assign LUT_3[59736] = 32'b00000000000000001010010000000011;
assign LUT_3[59737] = 32'b00000000000000010000111011100000;
assign LUT_3[59738] = 32'b00000000000000001100010111100111;
assign LUT_3[59739] = 32'b00000000000000010011000011000100;
assign LUT_3[59740] = 32'b00000000000000000111011101111001;
assign LUT_3[59741] = 32'b00000000000000001110001001010110;
assign LUT_3[59742] = 32'b00000000000000001001100101011101;
assign LUT_3[59743] = 32'b00000000000000010000010000111010;
assign LUT_3[59744] = 32'b00000000000000000010110010011010;
assign LUT_3[59745] = 32'b00000000000000001001011101110111;
assign LUT_3[59746] = 32'b00000000000000000100111001111110;
assign LUT_3[59747] = 32'b00000000000000001011100101011011;
assign LUT_3[59748] = 32'b00000000000000000000000000010000;
assign LUT_3[59749] = 32'b00000000000000000110101011101101;
assign LUT_3[59750] = 32'b00000000000000000010000111110100;
assign LUT_3[59751] = 32'b00000000000000001000110011010001;
assign LUT_3[59752] = 32'b00000000000000001000001011100000;
assign LUT_3[59753] = 32'b00000000000000001110110110111101;
assign LUT_3[59754] = 32'b00000000000000001010010011000100;
assign LUT_3[59755] = 32'b00000000000000010000111110100001;
assign LUT_3[59756] = 32'b00000000000000000101011001010110;
assign LUT_3[59757] = 32'b00000000000000001100000100110011;
assign LUT_3[59758] = 32'b00000000000000000111100000111010;
assign LUT_3[59759] = 32'b00000000000000001110001100010111;
assign LUT_3[59760] = 32'b00000000000000000110000101011101;
assign LUT_3[59761] = 32'b00000000000000001100110000111010;
assign LUT_3[59762] = 32'b00000000000000001000001101000001;
assign LUT_3[59763] = 32'b00000000000000001110111000011110;
assign LUT_3[59764] = 32'b00000000000000000011010011010011;
assign LUT_3[59765] = 32'b00000000000000001001111110110000;
assign LUT_3[59766] = 32'b00000000000000000101011010110111;
assign LUT_3[59767] = 32'b00000000000000001100000110010100;
assign LUT_3[59768] = 32'b00000000000000001011011110100011;
assign LUT_3[59769] = 32'b00000000000000010010001010000000;
assign LUT_3[59770] = 32'b00000000000000001101100110000111;
assign LUT_3[59771] = 32'b00000000000000010100010001100100;
assign LUT_3[59772] = 32'b00000000000000001000101100011001;
assign LUT_3[59773] = 32'b00000000000000001111010111110110;
assign LUT_3[59774] = 32'b00000000000000001010110011111101;
assign LUT_3[59775] = 32'b00000000000000010001011111011010;
assign LUT_3[59776] = 32'b00000000000000000011110110001101;
assign LUT_3[59777] = 32'b00000000000000001010100001101010;
assign LUT_3[59778] = 32'b00000000000000000101111101110001;
assign LUT_3[59779] = 32'b00000000000000001100101001001110;
assign LUT_3[59780] = 32'b00000000000000000001000100000011;
assign LUT_3[59781] = 32'b00000000000000000111101111100000;
assign LUT_3[59782] = 32'b00000000000000000011001011100111;
assign LUT_3[59783] = 32'b00000000000000001001110111000100;
assign LUT_3[59784] = 32'b00000000000000001001001111010011;
assign LUT_3[59785] = 32'b00000000000000001111111010110000;
assign LUT_3[59786] = 32'b00000000000000001011010110110111;
assign LUT_3[59787] = 32'b00000000000000010010000010010100;
assign LUT_3[59788] = 32'b00000000000000000110011101001001;
assign LUT_3[59789] = 32'b00000000000000001101001000100110;
assign LUT_3[59790] = 32'b00000000000000001000100100101101;
assign LUT_3[59791] = 32'b00000000000000001111010000001010;
assign LUT_3[59792] = 32'b00000000000000000111001001010000;
assign LUT_3[59793] = 32'b00000000000000001101110100101101;
assign LUT_3[59794] = 32'b00000000000000001001010000110100;
assign LUT_3[59795] = 32'b00000000000000001111111100010001;
assign LUT_3[59796] = 32'b00000000000000000100010111000110;
assign LUT_3[59797] = 32'b00000000000000001011000010100011;
assign LUT_3[59798] = 32'b00000000000000000110011110101010;
assign LUT_3[59799] = 32'b00000000000000001101001010000111;
assign LUT_3[59800] = 32'b00000000000000001100100010010110;
assign LUT_3[59801] = 32'b00000000000000010011001101110011;
assign LUT_3[59802] = 32'b00000000000000001110101001111010;
assign LUT_3[59803] = 32'b00000000000000010101010101010111;
assign LUT_3[59804] = 32'b00000000000000001001110000001100;
assign LUT_3[59805] = 32'b00000000000000010000011011101001;
assign LUT_3[59806] = 32'b00000000000000001011110111110000;
assign LUT_3[59807] = 32'b00000000000000010010100011001101;
assign LUT_3[59808] = 32'b00000000000000000101000100101101;
assign LUT_3[59809] = 32'b00000000000000001011110000001010;
assign LUT_3[59810] = 32'b00000000000000000111001100010001;
assign LUT_3[59811] = 32'b00000000000000001101110111101110;
assign LUT_3[59812] = 32'b00000000000000000010010010100011;
assign LUT_3[59813] = 32'b00000000000000001000111110000000;
assign LUT_3[59814] = 32'b00000000000000000100011010000111;
assign LUT_3[59815] = 32'b00000000000000001011000101100100;
assign LUT_3[59816] = 32'b00000000000000001010011101110011;
assign LUT_3[59817] = 32'b00000000000000010001001001010000;
assign LUT_3[59818] = 32'b00000000000000001100100101010111;
assign LUT_3[59819] = 32'b00000000000000010011010000110100;
assign LUT_3[59820] = 32'b00000000000000000111101011101001;
assign LUT_3[59821] = 32'b00000000000000001110010111000110;
assign LUT_3[59822] = 32'b00000000000000001001110011001101;
assign LUT_3[59823] = 32'b00000000000000010000011110101010;
assign LUT_3[59824] = 32'b00000000000000001000010111110000;
assign LUT_3[59825] = 32'b00000000000000001111000011001101;
assign LUT_3[59826] = 32'b00000000000000001010011111010100;
assign LUT_3[59827] = 32'b00000000000000010001001010110001;
assign LUT_3[59828] = 32'b00000000000000000101100101100110;
assign LUT_3[59829] = 32'b00000000000000001100010001000011;
assign LUT_3[59830] = 32'b00000000000000000111101101001010;
assign LUT_3[59831] = 32'b00000000000000001110011000100111;
assign LUT_3[59832] = 32'b00000000000000001101110000110110;
assign LUT_3[59833] = 32'b00000000000000010100011100010011;
assign LUT_3[59834] = 32'b00000000000000001111111000011010;
assign LUT_3[59835] = 32'b00000000000000010110100011110111;
assign LUT_3[59836] = 32'b00000000000000001010111110101100;
assign LUT_3[59837] = 32'b00000000000000010001101010001001;
assign LUT_3[59838] = 32'b00000000000000001101000110010000;
assign LUT_3[59839] = 32'b00000000000000010011110001101101;
assign LUT_3[59840] = 32'b00000000000000000011101110111000;
assign LUT_3[59841] = 32'b00000000000000001010011010010101;
assign LUT_3[59842] = 32'b00000000000000000101110110011100;
assign LUT_3[59843] = 32'b00000000000000001100100001111001;
assign LUT_3[59844] = 32'b00000000000000000000111100101110;
assign LUT_3[59845] = 32'b00000000000000000111101000001011;
assign LUT_3[59846] = 32'b00000000000000000011000100010010;
assign LUT_3[59847] = 32'b00000000000000001001101111101111;
assign LUT_3[59848] = 32'b00000000000000001001000111111110;
assign LUT_3[59849] = 32'b00000000000000001111110011011011;
assign LUT_3[59850] = 32'b00000000000000001011001111100010;
assign LUT_3[59851] = 32'b00000000000000010001111010111111;
assign LUT_3[59852] = 32'b00000000000000000110010101110100;
assign LUT_3[59853] = 32'b00000000000000001101000001010001;
assign LUT_3[59854] = 32'b00000000000000001000011101011000;
assign LUT_3[59855] = 32'b00000000000000001111001000110101;
assign LUT_3[59856] = 32'b00000000000000000111000001111011;
assign LUT_3[59857] = 32'b00000000000000001101101101011000;
assign LUT_3[59858] = 32'b00000000000000001001001001011111;
assign LUT_3[59859] = 32'b00000000000000001111110100111100;
assign LUT_3[59860] = 32'b00000000000000000100001111110001;
assign LUT_3[59861] = 32'b00000000000000001010111011001110;
assign LUT_3[59862] = 32'b00000000000000000110010111010101;
assign LUT_3[59863] = 32'b00000000000000001101000010110010;
assign LUT_3[59864] = 32'b00000000000000001100011011000001;
assign LUT_3[59865] = 32'b00000000000000010011000110011110;
assign LUT_3[59866] = 32'b00000000000000001110100010100101;
assign LUT_3[59867] = 32'b00000000000000010101001110000010;
assign LUT_3[59868] = 32'b00000000000000001001101000110111;
assign LUT_3[59869] = 32'b00000000000000010000010100010100;
assign LUT_3[59870] = 32'b00000000000000001011110000011011;
assign LUT_3[59871] = 32'b00000000000000010010011011111000;
assign LUT_3[59872] = 32'b00000000000000000100111101011000;
assign LUT_3[59873] = 32'b00000000000000001011101000110101;
assign LUT_3[59874] = 32'b00000000000000000111000100111100;
assign LUT_3[59875] = 32'b00000000000000001101110000011001;
assign LUT_3[59876] = 32'b00000000000000000010001011001110;
assign LUT_3[59877] = 32'b00000000000000001000110110101011;
assign LUT_3[59878] = 32'b00000000000000000100010010110010;
assign LUT_3[59879] = 32'b00000000000000001010111110001111;
assign LUT_3[59880] = 32'b00000000000000001010010110011110;
assign LUT_3[59881] = 32'b00000000000000010001000001111011;
assign LUT_3[59882] = 32'b00000000000000001100011110000010;
assign LUT_3[59883] = 32'b00000000000000010011001001011111;
assign LUT_3[59884] = 32'b00000000000000000111100100010100;
assign LUT_3[59885] = 32'b00000000000000001110001111110001;
assign LUT_3[59886] = 32'b00000000000000001001101011111000;
assign LUT_3[59887] = 32'b00000000000000010000010111010101;
assign LUT_3[59888] = 32'b00000000000000001000010000011011;
assign LUT_3[59889] = 32'b00000000000000001110111011111000;
assign LUT_3[59890] = 32'b00000000000000001010010111111111;
assign LUT_3[59891] = 32'b00000000000000010001000011011100;
assign LUT_3[59892] = 32'b00000000000000000101011110010001;
assign LUT_3[59893] = 32'b00000000000000001100001001101110;
assign LUT_3[59894] = 32'b00000000000000000111100101110101;
assign LUT_3[59895] = 32'b00000000000000001110010001010010;
assign LUT_3[59896] = 32'b00000000000000001101101001100001;
assign LUT_3[59897] = 32'b00000000000000010100010100111110;
assign LUT_3[59898] = 32'b00000000000000001111110001000101;
assign LUT_3[59899] = 32'b00000000000000010110011100100010;
assign LUT_3[59900] = 32'b00000000000000001010110111010111;
assign LUT_3[59901] = 32'b00000000000000010001100010110100;
assign LUT_3[59902] = 32'b00000000000000001100111110111011;
assign LUT_3[59903] = 32'b00000000000000010011101010011000;
assign LUT_3[59904] = 32'b00000000000000001000110000111010;
assign LUT_3[59905] = 32'b00000000000000001111011100010111;
assign LUT_3[59906] = 32'b00000000000000001010111000011110;
assign LUT_3[59907] = 32'b00000000000000010001100011111011;
assign LUT_3[59908] = 32'b00000000000000000101111110110000;
assign LUT_3[59909] = 32'b00000000000000001100101010001101;
assign LUT_3[59910] = 32'b00000000000000001000000110010100;
assign LUT_3[59911] = 32'b00000000000000001110110001110001;
assign LUT_3[59912] = 32'b00000000000000001110001010000000;
assign LUT_3[59913] = 32'b00000000000000010100110101011101;
assign LUT_3[59914] = 32'b00000000000000010000010001100100;
assign LUT_3[59915] = 32'b00000000000000010110111101000001;
assign LUT_3[59916] = 32'b00000000000000001011010111110110;
assign LUT_3[59917] = 32'b00000000000000010010000011010011;
assign LUT_3[59918] = 32'b00000000000000001101011111011010;
assign LUT_3[59919] = 32'b00000000000000010100001010110111;
assign LUT_3[59920] = 32'b00000000000000001100000011111101;
assign LUT_3[59921] = 32'b00000000000000010010101111011010;
assign LUT_3[59922] = 32'b00000000000000001110001011100001;
assign LUT_3[59923] = 32'b00000000000000010100110110111110;
assign LUT_3[59924] = 32'b00000000000000001001010001110011;
assign LUT_3[59925] = 32'b00000000000000001111111101010000;
assign LUT_3[59926] = 32'b00000000000000001011011001010111;
assign LUT_3[59927] = 32'b00000000000000010010000100110100;
assign LUT_3[59928] = 32'b00000000000000010001011101000011;
assign LUT_3[59929] = 32'b00000000000000011000001000100000;
assign LUT_3[59930] = 32'b00000000000000010011100100100111;
assign LUT_3[59931] = 32'b00000000000000011010010000000100;
assign LUT_3[59932] = 32'b00000000000000001110101010111001;
assign LUT_3[59933] = 32'b00000000000000010101010110010110;
assign LUT_3[59934] = 32'b00000000000000010000110010011101;
assign LUT_3[59935] = 32'b00000000000000010111011101111010;
assign LUT_3[59936] = 32'b00000000000000001001111111011010;
assign LUT_3[59937] = 32'b00000000000000010000101010110111;
assign LUT_3[59938] = 32'b00000000000000001100000110111110;
assign LUT_3[59939] = 32'b00000000000000010010110010011011;
assign LUT_3[59940] = 32'b00000000000000000111001101010000;
assign LUT_3[59941] = 32'b00000000000000001101111000101101;
assign LUT_3[59942] = 32'b00000000000000001001010100110100;
assign LUT_3[59943] = 32'b00000000000000010000000000010001;
assign LUT_3[59944] = 32'b00000000000000001111011000100000;
assign LUT_3[59945] = 32'b00000000000000010110000011111101;
assign LUT_3[59946] = 32'b00000000000000010001100000000100;
assign LUT_3[59947] = 32'b00000000000000011000001011100001;
assign LUT_3[59948] = 32'b00000000000000001100100110010110;
assign LUT_3[59949] = 32'b00000000000000010011010001110011;
assign LUT_3[59950] = 32'b00000000000000001110101101111010;
assign LUT_3[59951] = 32'b00000000000000010101011001010111;
assign LUT_3[59952] = 32'b00000000000000001101010010011101;
assign LUT_3[59953] = 32'b00000000000000010011111101111010;
assign LUT_3[59954] = 32'b00000000000000001111011010000001;
assign LUT_3[59955] = 32'b00000000000000010110000101011110;
assign LUT_3[59956] = 32'b00000000000000001010100000010011;
assign LUT_3[59957] = 32'b00000000000000010001001011110000;
assign LUT_3[59958] = 32'b00000000000000001100100111110111;
assign LUT_3[59959] = 32'b00000000000000010011010011010100;
assign LUT_3[59960] = 32'b00000000000000010010101011100011;
assign LUT_3[59961] = 32'b00000000000000011001010111000000;
assign LUT_3[59962] = 32'b00000000000000010100110011000111;
assign LUT_3[59963] = 32'b00000000000000011011011110100100;
assign LUT_3[59964] = 32'b00000000000000001111111001011001;
assign LUT_3[59965] = 32'b00000000000000010110100100110110;
assign LUT_3[59966] = 32'b00000000000000010010000000111101;
assign LUT_3[59967] = 32'b00000000000000011000101100011010;
assign LUT_3[59968] = 32'b00000000000000001000101001100101;
assign LUT_3[59969] = 32'b00000000000000001111010101000010;
assign LUT_3[59970] = 32'b00000000000000001010110001001001;
assign LUT_3[59971] = 32'b00000000000000010001011100100110;
assign LUT_3[59972] = 32'b00000000000000000101110111011011;
assign LUT_3[59973] = 32'b00000000000000001100100010111000;
assign LUT_3[59974] = 32'b00000000000000000111111110111111;
assign LUT_3[59975] = 32'b00000000000000001110101010011100;
assign LUT_3[59976] = 32'b00000000000000001110000010101011;
assign LUT_3[59977] = 32'b00000000000000010100101110001000;
assign LUT_3[59978] = 32'b00000000000000010000001010001111;
assign LUT_3[59979] = 32'b00000000000000010110110101101100;
assign LUT_3[59980] = 32'b00000000000000001011010000100001;
assign LUT_3[59981] = 32'b00000000000000010001111011111110;
assign LUT_3[59982] = 32'b00000000000000001101011000000101;
assign LUT_3[59983] = 32'b00000000000000010100000011100010;
assign LUT_3[59984] = 32'b00000000000000001011111100101000;
assign LUT_3[59985] = 32'b00000000000000010010101000000101;
assign LUT_3[59986] = 32'b00000000000000001110000100001100;
assign LUT_3[59987] = 32'b00000000000000010100101111101001;
assign LUT_3[59988] = 32'b00000000000000001001001010011110;
assign LUT_3[59989] = 32'b00000000000000001111110101111011;
assign LUT_3[59990] = 32'b00000000000000001011010010000010;
assign LUT_3[59991] = 32'b00000000000000010001111101011111;
assign LUT_3[59992] = 32'b00000000000000010001010101101110;
assign LUT_3[59993] = 32'b00000000000000011000000001001011;
assign LUT_3[59994] = 32'b00000000000000010011011101010010;
assign LUT_3[59995] = 32'b00000000000000011010001000101111;
assign LUT_3[59996] = 32'b00000000000000001110100011100100;
assign LUT_3[59997] = 32'b00000000000000010101001111000001;
assign LUT_3[59998] = 32'b00000000000000010000101011001000;
assign LUT_3[59999] = 32'b00000000000000010111010110100101;
assign LUT_3[60000] = 32'b00000000000000001001111000000101;
assign LUT_3[60001] = 32'b00000000000000010000100011100010;
assign LUT_3[60002] = 32'b00000000000000001011111111101001;
assign LUT_3[60003] = 32'b00000000000000010010101011000110;
assign LUT_3[60004] = 32'b00000000000000000111000101111011;
assign LUT_3[60005] = 32'b00000000000000001101110001011000;
assign LUT_3[60006] = 32'b00000000000000001001001101011111;
assign LUT_3[60007] = 32'b00000000000000001111111000111100;
assign LUT_3[60008] = 32'b00000000000000001111010001001011;
assign LUT_3[60009] = 32'b00000000000000010101111100101000;
assign LUT_3[60010] = 32'b00000000000000010001011000101111;
assign LUT_3[60011] = 32'b00000000000000011000000100001100;
assign LUT_3[60012] = 32'b00000000000000001100011111000001;
assign LUT_3[60013] = 32'b00000000000000010011001010011110;
assign LUT_3[60014] = 32'b00000000000000001110100110100101;
assign LUT_3[60015] = 32'b00000000000000010101010010000010;
assign LUT_3[60016] = 32'b00000000000000001101001011001000;
assign LUT_3[60017] = 32'b00000000000000010011110110100101;
assign LUT_3[60018] = 32'b00000000000000001111010010101100;
assign LUT_3[60019] = 32'b00000000000000010101111110001001;
assign LUT_3[60020] = 32'b00000000000000001010011000111110;
assign LUT_3[60021] = 32'b00000000000000010001000100011011;
assign LUT_3[60022] = 32'b00000000000000001100100000100010;
assign LUT_3[60023] = 32'b00000000000000010011001011111111;
assign LUT_3[60024] = 32'b00000000000000010010100100001110;
assign LUT_3[60025] = 32'b00000000000000011001001111101011;
assign LUT_3[60026] = 32'b00000000000000010100101011110010;
assign LUT_3[60027] = 32'b00000000000000011011010111001111;
assign LUT_3[60028] = 32'b00000000000000001111110010000100;
assign LUT_3[60029] = 32'b00000000000000010110011101100001;
assign LUT_3[60030] = 32'b00000000000000010001111001101000;
assign LUT_3[60031] = 32'b00000000000000011000100101000101;
assign LUT_3[60032] = 32'b00000000000000001010111011111000;
assign LUT_3[60033] = 32'b00000000000000010001100111010101;
assign LUT_3[60034] = 32'b00000000000000001101000011011100;
assign LUT_3[60035] = 32'b00000000000000010011101110111001;
assign LUT_3[60036] = 32'b00000000000000001000001001101110;
assign LUT_3[60037] = 32'b00000000000000001110110101001011;
assign LUT_3[60038] = 32'b00000000000000001010010001010010;
assign LUT_3[60039] = 32'b00000000000000010000111100101111;
assign LUT_3[60040] = 32'b00000000000000010000010100111110;
assign LUT_3[60041] = 32'b00000000000000010111000000011011;
assign LUT_3[60042] = 32'b00000000000000010010011100100010;
assign LUT_3[60043] = 32'b00000000000000011001000111111111;
assign LUT_3[60044] = 32'b00000000000000001101100010110100;
assign LUT_3[60045] = 32'b00000000000000010100001110010001;
assign LUT_3[60046] = 32'b00000000000000001111101010011000;
assign LUT_3[60047] = 32'b00000000000000010110010101110101;
assign LUT_3[60048] = 32'b00000000000000001110001110111011;
assign LUT_3[60049] = 32'b00000000000000010100111010011000;
assign LUT_3[60050] = 32'b00000000000000010000010110011111;
assign LUT_3[60051] = 32'b00000000000000010111000001111100;
assign LUT_3[60052] = 32'b00000000000000001011011100110001;
assign LUT_3[60053] = 32'b00000000000000010010001000001110;
assign LUT_3[60054] = 32'b00000000000000001101100100010101;
assign LUT_3[60055] = 32'b00000000000000010100001111110010;
assign LUT_3[60056] = 32'b00000000000000010011101000000001;
assign LUT_3[60057] = 32'b00000000000000011010010011011110;
assign LUT_3[60058] = 32'b00000000000000010101101111100101;
assign LUT_3[60059] = 32'b00000000000000011100011011000010;
assign LUT_3[60060] = 32'b00000000000000010000110101110111;
assign LUT_3[60061] = 32'b00000000000000010111100001010100;
assign LUT_3[60062] = 32'b00000000000000010010111101011011;
assign LUT_3[60063] = 32'b00000000000000011001101000111000;
assign LUT_3[60064] = 32'b00000000000000001100001010011000;
assign LUT_3[60065] = 32'b00000000000000010010110101110101;
assign LUT_3[60066] = 32'b00000000000000001110010001111100;
assign LUT_3[60067] = 32'b00000000000000010100111101011001;
assign LUT_3[60068] = 32'b00000000000000001001011000001110;
assign LUT_3[60069] = 32'b00000000000000010000000011101011;
assign LUT_3[60070] = 32'b00000000000000001011011111110010;
assign LUT_3[60071] = 32'b00000000000000010010001011001111;
assign LUT_3[60072] = 32'b00000000000000010001100011011110;
assign LUT_3[60073] = 32'b00000000000000011000001110111011;
assign LUT_3[60074] = 32'b00000000000000010011101011000010;
assign LUT_3[60075] = 32'b00000000000000011010010110011111;
assign LUT_3[60076] = 32'b00000000000000001110110001010100;
assign LUT_3[60077] = 32'b00000000000000010101011100110001;
assign LUT_3[60078] = 32'b00000000000000010000111000111000;
assign LUT_3[60079] = 32'b00000000000000010111100100010101;
assign LUT_3[60080] = 32'b00000000000000001111011101011011;
assign LUT_3[60081] = 32'b00000000000000010110001000111000;
assign LUT_3[60082] = 32'b00000000000000010001100100111111;
assign LUT_3[60083] = 32'b00000000000000011000010000011100;
assign LUT_3[60084] = 32'b00000000000000001100101011010001;
assign LUT_3[60085] = 32'b00000000000000010011010110101110;
assign LUT_3[60086] = 32'b00000000000000001110110010110101;
assign LUT_3[60087] = 32'b00000000000000010101011110010010;
assign LUT_3[60088] = 32'b00000000000000010100110110100001;
assign LUT_3[60089] = 32'b00000000000000011011100001111110;
assign LUT_3[60090] = 32'b00000000000000010110111110000101;
assign LUT_3[60091] = 32'b00000000000000011101101001100010;
assign LUT_3[60092] = 32'b00000000000000010010000100010111;
assign LUT_3[60093] = 32'b00000000000000011000101111110100;
assign LUT_3[60094] = 32'b00000000000000010100001011111011;
assign LUT_3[60095] = 32'b00000000000000011010110111011000;
assign LUT_3[60096] = 32'b00000000000000001010110100100011;
assign LUT_3[60097] = 32'b00000000000000010001100000000000;
assign LUT_3[60098] = 32'b00000000000000001100111100000111;
assign LUT_3[60099] = 32'b00000000000000010011100111100100;
assign LUT_3[60100] = 32'b00000000000000001000000010011001;
assign LUT_3[60101] = 32'b00000000000000001110101101110110;
assign LUT_3[60102] = 32'b00000000000000001010001001111101;
assign LUT_3[60103] = 32'b00000000000000010000110101011010;
assign LUT_3[60104] = 32'b00000000000000010000001101101001;
assign LUT_3[60105] = 32'b00000000000000010110111001000110;
assign LUT_3[60106] = 32'b00000000000000010010010101001101;
assign LUT_3[60107] = 32'b00000000000000011001000000101010;
assign LUT_3[60108] = 32'b00000000000000001101011011011111;
assign LUT_3[60109] = 32'b00000000000000010100000110111100;
assign LUT_3[60110] = 32'b00000000000000001111100011000011;
assign LUT_3[60111] = 32'b00000000000000010110001110100000;
assign LUT_3[60112] = 32'b00000000000000001110000111100110;
assign LUT_3[60113] = 32'b00000000000000010100110011000011;
assign LUT_3[60114] = 32'b00000000000000010000001111001010;
assign LUT_3[60115] = 32'b00000000000000010110111010100111;
assign LUT_3[60116] = 32'b00000000000000001011010101011100;
assign LUT_3[60117] = 32'b00000000000000010010000000111001;
assign LUT_3[60118] = 32'b00000000000000001101011101000000;
assign LUT_3[60119] = 32'b00000000000000010100001000011101;
assign LUT_3[60120] = 32'b00000000000000010011100000101100;
assign LUT_3[60121] = 32'b00000000000000011010001100001001;
assign LUT_3[60122] = 32'b00000000000000010101101000010000;
assign LUT_3[60123] = 32'b00000000000000011100010011101101;
assign LUT_3[60124] = 32'b00000000000000010000101110100010;
assign LUT_3[60125] = 32'b00000000000000010111011001111111;
assign LUT_3[60126] = 32'b00000000000000010010110110000110;
assign LUT_3[60127] = 32'b00000000000000011001100001100011;
assign LUT_3[60128] = 32'b00000000000000001100000011000011;
assign LUT_3[60129] = 32'b00000000000000010010101110100000;
assign LUT_3[60130] = 32'b00000000000000001110001010100111;
assign LUT_3[60131] = 32'b00000000000000010100110110000100;
assign LUT_3[60132] = 32'b00000000000000001001010000111001;
assign LUT_3[60133] = 32'b00000000000000001111111100010110;
assign LUT_3[60134] = 32'b00000000000000001011011000011101;
assign LUT_3[60135] = 32'b00000000000000010010000011111010;
assign LUT_3[60136] = 32'b00000000000000010001011100001001;
assign LUT_3[60137] = 32'b00000000000000011000000111100110;
assign LUT_3[60138] = 32'b00000000000000010011100011101101;
assign LUT_3[60139] = 32'b00000000000000011010001111001010;
assign LUT_3[60140] = 32'b00000000000000001110101001111111;
assign LUT_3[60141] = 32'b00000000000000010101010101011100;
assign LUT_3[60142] = 32'b00000000000000010000110001100011;
assign LUT_3[60143] = 32'b00000000000000010111011101000000;
assign LUT_3[60144] = 32'b00000000000000001111010110000110;
assign LUT_3[60145] = 32'b00000000000000010110000001100011;
assign LUT_3[60146] = 32'b00000000000000010001011101101010;
assign LUT_3[60147] = 32'b00000000000000011000001001000111;
assign LUT_3[60148] = 32'b00000000000000001100100011111100;
assign LUT_3[60149] = 32'b00000000000000010011001111011001;
assign LUT_3[60150] = 32'b00000000000000001110101011100000;
assign LUT_3[60151] = 32'b00000000000000010101010110111101;
assign LUT_3[60152] = 32'b00000000000000010100101111001100;
assign LUT_3[60153] = 32'b00000000000000011011011010101001;
assign LUT_3[60154] = 32'b00000000000000010110110110110000;
assign LUT_3[60155] = 32'b00000000000000011101100010001101;
assign LUT_3[60156] = 32'b00000000000000010001111101000010;
assign LUT_3[60157] = 32'b00000000000000011000101000011111;
assign LUT_3[60158] = 32'b00000000000000010100000100100110;
assign LUT_3[60159] = 32'b00000000000000011010110000000011;
assign LUT_3[60160] = 32'b00000000000000000101000000011011;
assign LUT_3[60161] = 32'b00000000000000001011101011111000;
assign LUT_3[60162] = 32'b00000000000000000111000111111111;
assign LUT_3[60163] = 32'b00000000000000001101110011011100;
assign LUT_3[60164] = 32'b00000000000000000010001110010001;
assign LUT_3[60165] = 32'b00000000000000001000111001101110;
assign LUT_3[60166] = 32'b00000000000000000100010101110101;
assign LUT_3[60167] = 32'b00000000000000001011000001010010;
assign LUT_3[60168] = 32'b00000000000000001010011001100001;
assign LUT_3[60169] = 32'b00000000000000010001000100111110;
assign LUT_3[60170] = 32'b00000000000000001100100001000101;
assign LUT_3[60171] = 32'b00000000000000010011001100100010;
assign LUT_3[60172] = 32'b00000000000000000111100111010111;
assign LUT_3[60173] = 32'b00000000000000001110010010110100;
assign LUT_3[60174] = 32'b00000000000000001001101110111011;
assign LUT_3[60175] = 32'b00000000000000010000011010011000;
assign LUT_3[60176] = 32'b00000000000000001000010011011110;
assign LUT_3[60177] = 32'b00000000000000001110111110111011;
assign LUT_3[60178] = 32'b00000000000000001010011011000010;
assign LUT_3[60179] = 32'b00000000000000010001000110011111;
assign LUT_3[60180] = 32'b00000000000000000101100001010100;
assign LUT_3[60181] = 32'b00000000000000001100001100110001;
assign LUT_3[60182] = 32'b00000000000000000111101000111000;
assign LUT_3[60183] = 32'b00000000000000001110010100010101;
assign LUT_3[60184] = 32'b00000000000000001101101100100100;
assign LUT_3[60185] = 32'b00000000000000010100011000000001;
assign LUT_3[60186] = 32'b00000000000000001111110100001000;
assign LUT_3[60187] = 32'b00000000000000010110011111100101;
assign LUT_3[60188] = 32'b00000000000000001010111010011010;
assign LUT_3[60189] = 32'b00000000000000010001100101110111;
assign LUT_3[60190] = 32'b00000000000000001101000001111110;
assign LUT_3[60191] = 32'b00000000000000010011101101011011;
assign LUT_3[60192] = 32'b00000000000000000110001110111011;
assign LUT_3[60193] = 32'b00000000000000001100111010011000;
assign LUT_3[60194] = 32'b00000000000000001000010110011111;
assign LUT_3[60195] = 32'b00000000000000001111000001111100;
assign LUT_3[60196] = 32'b00000000000000000011011100110001;
assign LUT_3[60197] = 32'b00000000000000001010001000001110;
assign LUT_3[60198] = 32'b00000000000000000101100100010101;
assign LUT_3[60199] = 32'b00000000000000001100001111110010;
assign LUT_3[60200] = 32'b00000000000000001011101000000001;
assign LUT_3[60201] = 32'b00000000000000010010010011011110;
assign LUT_3[60202] = 32'b00000000000000001101101111100101;
assign LUT_3[60203] = 32'b00000000000000010100011011000010;
assign LUT_3[60204] = 32'b00000000000000001000110101110111;
assign LUT_3[60205] = 32'b00000000000000001111100001010100;
assign LUT_3[60206] = 32'b00000000000000001010111101011011;
assign LUT_3[60207] = 32'b00000000000000010001101000111000;
assign LUT_3[60208] = 32'b00000000000000001001100001111110;
assign LUT_3[60209] = 32'b00000000000000010000001101011011;
assign LUT_3[60210] = 32'b00000000000000001011101001100010;
assign LUT_3[60211] = 32'b00000000000000010010010100111111;
assign LUT_3[60212] = 32'b00000000000000000110101111110100;
assign LUT_3[60213] = 32'b00000000000000001101011011010001;
assign LUT_3[60214] = 32'b00000000000000001000110111011000;
assign LUT_3[60215] = 32'b00000000000000001111100010110101;
assign LUT_3[60216] = 32'b00000000000000001110111011000100;
assign LUT_3[60217] = 32'b00000000000000010101100110100001;
assign LUT_3[60218] = 32'b00000000000000010001000010101000;
assign LUT_3[60219] = 32'b00000000000000010111101110000101;
assign LUT_3[60220] = 32'b00000000000000001100001000111010;
assign LUT_3[60221] = 32'b00000000000000010010110100010111;
assign LUT_3[60222] = 32'b00000000000000001110010000011110;
assign LUT_3[60223] = 32'b00000000000000010100111011111011;
assign LUT_3[60224] = 32'b00000000000000000100111001000110;
assign LUT_3[60225] = 32'b00000000000000001011100100100011;
assign LUT_3[60226] = 32'b00000000000000000111000000101010;
assign LUT_3[60227] = 32'b00000000000000001101101100000111;
assign LUT_3[60228] = 32'b00000000000000000010000110111100;
assign LUT_3[60229] = 32'b00000000000000001000110010011001;
assign LUT_3[60230] = 32'b00000000000000000100001110100000;
assign LUT_3[60231] = 32'b00000000000000001010111001111101;
assign LUT_3[60232] = 32'b00000000000000001010010010001100;
assign LUT_3[60233] = 32'b00000000000000010000111101101001;
assign LUT_3[60234] = 32'b00000000000000001100011001110000;
assign LUT_3[60235] = 32'b00000000000000010011000101001101;
assign LUT_3[60236] = 32'b00000000000000000111100000000010;
assign LUT_3[60237] = 32'b00000000000000001110001011011111;
assign LUT_3[60238] = 32'b00000000000000001001100111100110;
assign LUT_3[60239] = 32'b00000000000000010000010011000011;
assign LUT_3[60240] = 32'b00000000000000001000001100001001;
assign LUT_3[60241] = 32'b00000000000000001110110111100110;
assign LUT_3[60242] = 32'b00000000000000001010010011101101;
assign LUT_3[60243] = 32'b00000000000000010000111111001010;
assign LUT_3[60244] = 32'b00000000000000000101011001111111;
assign LUT_3[60245] = 32'b00000000000000001100000101011100;
assign LUT_3[60246] = 32'b00000000000000000111100001100011;
assign LUT_3[60247] = 32'b00000000000000001110001101000000;
assign LUT_3[60248] = 32'b00000000000000001101100101001111;
assign LUT_3[60249] = 32'b00000000000000010100010000101100;
assign LUT_3[60250] = 32'b00000000000000001111101100110011;
assign LUT_3[60251] = 32'b00000000000000010110011000010000;
assign LUT_3[60252] = 32'b00000000000000001010110011000101;
assign LUT_3[60253] = 32'b00000000000000010001011110100010;
assign LUT_3[60254] = 32'b00000000000000001100111010101001;
assign LUT_3[60255] = 32'b00000000000000010011100110000110;
assign LUT_3[60256] = 32'b00000000000000000110000111100110;
assign LUT_3[60257] = 32'b00000000000000001100110011000011;
assign LUT_3[60258] = 32'b00000000000000001000001111001010;
assign LUT_3[60259] = 32'b00000000000000001110111010100111;
assign LUT_3[60260] = 32'b00000000000000000011010101011100;
assign LUT_3[60261] = 32'b00000000000000001010000000111001;
assign LUT_3[60262] = 32'b00000000000000000101011101000000;
assign LUT_3[60263] = 32'b00000000000000001100001000011101;
assign LUT_3[60264] = 32'b00000000000000001011100000101100;
assign LUT_3[60265] = 32'b00000000000000010010001100001001;
assign LUT_3[60266] = 32'b00000000000000001101101000010000;
assign LUT_3[60267] = 32'b00000000000000010100010011101101;
assign LUT_3[60268] = 32'b00000000000000001000101110100010;
assign LUT_3[60269] = 32'b00000000000000001111011001111111;
assign LUT_3[60270] = 32'b00000000000000001010110110000110;
assign LUT_3[60271] = 32'b00000000000000010001100001100011;
assign LUT_3[60272] = 32'b00000000000000001001011010101001;
assign LUT_3[60273] = 32'b00000000000000010000000110000110;
assign LUT_3[60274] = 32'b00000000000000001011100010001101;
assign LUT_3[60275] = 32'b00000000000000010010001101101010;
assign LUT_3[60276] = 32'b00000000000000000110101000011111;
assign LUT_3[60277] = 32'b00000000000000001101010011111100;
assign LUT_3[60278] = 32'b00000000000000001000110000000011;
assign LUT_3[60279] = 32'b00000000000000001111011011100000;
assign LUT_3[60280] = 32'b00000000000000001110110011101111;
assign LUT_3[60281] = 32'b00000000000000010101011111001100;
assign LUT_3[60282] = 32'b00000000000000010000111011010011;
assign LUT_3[60283] = 32'b00000000000000010111100110110000;
assign LUT_3[60284] = 32'b00000000000000001100000001100101;
assign LUT_3[60285] = 32'b00000000000000010010101101000010;
assign LUT_3[60286] = 32'b00000000000000001110001001001001;
assign LUT_3[60287] = 32'b00000000000000010100110100100110;
assign LUT_3[60288] = 32'b00000000000000000111001011011001;
assign LUT_3[60289] = 32'b00000000000000001101110110110110;
assign LUT_3[60290] = 32'b00000000000000001001010010111101;
assign LUT_3[60291] = 32'b00000000000000001111111110011010;
assign LUT_3[60292] = 32'b00000000000000000100011001001111;
assign LUT_3[60293] = 32'b00000000000000001011000100101100;
assign LUT_3[60294] = 32'b00000000000000000110100000110011;
assign LUT_3[60295] = 32'b00000000000000001101001100010000;
assign LUT_3[60296] = 32'b00000000000000001100100100011111;
assign LUT_3[60297] = 32'b00000000000000010011001111111100;
assign LUT_3[60298] = 32'b00000000000000001110101100000011;
assign LUT_3[60299] = 32'b00000000000000010101010111100000;
assign LUT_3[60300] = 32'b00000000000000001001110010010101;
assign LUT_3[60301] = 32'b00000000000000010000011101110010;
assign LUT_3[60302] = 32'b00000000000000001011111001111001;
assign LUT_3[60303] = 32'b00000000000000010010100101010110;
assign LUT_3[60304] = 32'b00000000000000001010011110011100;
assign LUT_3[60305] = 32'b00000000000000010001001001111001;
assign LUT_3[60306] = 32'b00000000000000001100100110000000;
assign LUT_3[60307] = 32'b00000000000000010011010001011101;
assign LUT_3[60308] = 32'b00000000000000000111101100010010;
assign LUT_3[60309] = 32'b00000000000000001110010111101111;
assign LUT_3[60310] = 32'b00000000000000001001110011110110;
assign LUT_3[60311] = 32'b00000000000000010000011111010011;
assign LUT_3[60312] = 32'b00000000000000001111110111100010;
assign LUT_3[60313] = 32'b00000000000000010110100010111111;
assign LUT_3[60314] = 32'b00000000000000010001111111000110;
assign LUT_3[60315] = 32'b00000000000000011000101010100011;
assign LUT_3[60316] = 32'b00000000000000001101000101011000;
assign LUT_3[60317] = 32'b00000000000000010011110000110101;
assign LUT_3[60318] = 32'b00000000000000001111001100111100;
assign LUT_3[60319] = 32'b00000000000000010101111000011001;
assign LUT_3[60320] = 32'b00000000000000001000011001111001;
assign LUT_3[60321] = 32'b00000000000000001111000101010110;
assign LUT_3[60322] = 32'b00000000000000001010100001011101;
assign LUT_3[60323] = 32'b00000000000000010001001100111010;
assign LUT_3[60324] = 32'b00000000000000000101100111101111;
assign LUT_3[60325] = 32'b00000000000000001100010011001100;
assign LUT_3[60326] = 32'b00000000000000000111101111010011;
assign LUT_3[60327] = 32'b00000000000000001110011010110000;
assign LUT_3[60328] = 32'b00000000000000001101110010111111;
assign LUT_3[60329] = 32'b00000000000000010100011110011100;
assign LUT_3[60330] = 32'b00000000000000001111111010100011;
assign LUT_3[60331] = 32'b00000000000000010110100110000000;
assign LUT_3[60332] = 32'b00000000000000001011000000110101;
assign LUT_3[60333] = 32'b00000000000000010001101100010010;
assign LUT_3[60334] = 32'b00000000000000001101001000011001;
assign LUT_3[60335] = 32'b00000000000000010011110011110110;
assign LUT_3[60336] = 32'b00000000000000001011101100111100;
assign LUT_3[60337] = 32'b00000000000000010010011000011001;
assign LUT_3[60338] = 32'b00000000000000001101110100100000;
assign LUT_3[60339] = 32'b00000000000000010100011111111101;
assign LUT_3[60340] = 32'b00000000000000001000111010110010;
assign LUT_3[60341] = 32'b00000000000000001111100110001111;
assign LUT_3[60342] = 32'b00000000000000001011000010010110;
assign LUT_3[60343] = 32'b00000000000000010001101101110011;
assign LUT_3[60344] = 32'b00000000000000010001000110000010;
assign LUT_3[60345] = 32'b00000000000000010111110001011111;
assign LUT_3[60346] = 32'b00000000000000010011001101100110;
assign LUT_3[60347] = 32'b00000000000000011001111001000011;
assign LUT_3[60348] = 32'b00000000000000001110010011111000;
assign LUT_3[60349] = 32'b00000000000000010100111111010101;
assign LUT_3[60350] = 32'b00000000000000010000011011011100;
assign LUT_3[60351] = 32'b00000000000000010111000110111001;
assign LUT_3[60352] = 32'b00000000000000000111000100000100;
assign LUT_3[60353] = 32'b00000000000000001101101111100001;
assign LUT_3[60354] = 32'b00000000000000001001001011101000;
assign LUT_3[60355] = 32'b00000000000000001111110111000101;
assign LUT_3[60356] = 32'b00000000000000000100010001111010;
assign LUT_3[60357] = 32'b00000000000000001010111101010111;
assign LUT_3[60358] = 32'b00000000000000000110011001011110;
assign LUT_3[60359] = 32'b00000000000000001101000100111011;
assign LUT_3[60360] = 32'b00000000000000001100011101001010;
assign LUT_3[60361] = 32'b00000000000000010011001000100111;
assign LUT_3[60362] = 32'b00000000000000001110100100101110;
assign LUT_3[60363] = 32'b00000000000000010101010000001011;
assign LUT_3[60364] = 32'b00000000000000001001101011000000;
assign LUT_3[60365] = 32'b00000000000000010000010110011101;
assign LUT_3[60366] = 32'b00000000000000001011110010100100;
assign LUT_3[60367] = 32'b00000000000000010010011110000001;
assign LUT_3[60368] = 32'b00000000000000001010010111000111;
assign LUT_3[60369] = 32'b00000000000000010001000010100100;
assign LUT_3[60370] = 32'b00000000000000001100011110101011;
assign LUT_3[60371] = 32'b00000000000000010011001010001000;
assign LUT_3[60372] = 32'b00000000000000000111100100111101;
assign LUT_3[60373] = 32'b00000000000000001110010000011010;
assign LUT_3[60374] = 32'b00000000000000001001101100100001;
assign LUT_3[60375] = 32'b00000000000000010000010111111110;
assign LUT_3[60376] = 32'b00000000000000001111110000001101;
assign LUT_3[60377] = 32'b00000000000000010110011011101010;
assign LUT_3[60378] = 32'b00000000000000010001110111110001;
assign LUT_3[60379] = 32'b00000000000000011000100011001110;
assign LUT_3[60380] = 32'b00000000000000001100111110000011;
assign LUT_3[60381] = 32'b00000000000000010011101001100000;
assign LUT_3[60382] = 32'b00000000000000001111000101100111;
assign LUT_3[60383] = 32'b00000000000000010101110001000100;
assign LUT_3[60384] = 32'b00000000000000001000010010100100;
assign LUT_3[60385] = 32'b00000000000000001110111110000001;
assign LUT_3[60386] = 32'b00000000000000001010011010001000;
assign LUT_3[60387] = 32'b00000000000000010001000101100101;
assign LUT_3[60388] = 32'b00000000000000000101100000011010;
assign LUT_3[60389] = 32'b00000000000000001100001011110111;
assign LUT_3[60390] = 32'b00000000000000000111100111111110;
assign LUT_3[60391] = 32'b00000000000000001110010011011011;
assign LUT_3[60392] = 32'b00000000000000001101101011101010;
assign LUT_3[60393] = 32'b00000000000000010100010111000111;
assign LUT_3[60394] = 32'b00000000000000001111110011001110;
assign LUT_3[60395] = 32'b00000000000000010110011110101011;
assign LUT_3[60396] = 32'b00000000000000001010111001100000;
assign LUT_3[60397] = 32'b00000000000000010001100100111101;
assign LUT_3[60398] = 32'b00000000000000001101000001000100;
assign LUT_3[60399] = 32'b00000000000000010011101100100001;
assign LUT_3[60400] = 32'b00000000000000001011100101100111;
assign LUT_3[60401] = 32'b00000000000000010010010001000100;
assign LUT_3[60402] = 32'b00000000000000001101101101001011;
assign LUT_3[60403] = 32'b00000000000000010100011000101000;
assign LUT_3[60404] = 32'b00000000000000001000110011011101;
assign LUT_3[60405] = 32'b00000000000000001111011110111010;
assign LUT_3[60406] = 32'b00000000000000001010111011000001;
assign LUT_3[60407] = 32'b00000000000000010001100110011110;
assign LUT_3[60408] = 32'b00000000000000010000111110101101;
assign LUT_3[60409] = 32'b00000000000000010111101010001010;
assign LUT_3[60410] = 32'b00000000000000010011000110010001;
assign LUT_3[60411] = 32'b00000000000000011001110001101110;
assign LUT_3[60412] = 32'b00000000000000001110001100100011;
assign LUT_3[60413] = 32'b00000000000000010100111000000000;
assign LUT_3[60414] = 32'b00000000000000010000010100000111;
assign LUT_3[60415] = 32'b00000000000000010110111111100100;
assign LUT_3[60416] = 32'b00000000000000001100000000101011;
assign LUT_3[60417] = 32'b00000000000000010010101100001000;
assign LUT_3[60418] = 32'b00000000000000001110001000001111;
assign LUT_3[60419] = 32'b00000000000000010100110011101100;
assign LUT_3[60420] = 32'b00000000000000001001001110100001;
assign LUT_3[60421] = 32'b00000000000000001111111001111110;
assign LUT_3[60422] = 32'b00000000000000001011010110000101;
assign LUT_3[60423] = 32'b00000000000000010010000001100010;
assign LUT_3[60424] = 32'b00000000000000010001011001110001;
assign LUT_3[60425] = 32'b00000000000000011000000101001110;
assign LUT_3[60426] = 32'b00000000000000010011100001010101;
assign LUT_3[60427] = 32'b00000000000000011010001100110010;
assign LUT_3[60428] = 32'b00000000000000001110100111100111;
assign LUT_3[60429] = 32'b00000000000000010101010011000100;
assign LUT_3[60430] = 32'b00000000000000010000101111001011;
assign LUT_3[60431] = 32'b00000000000000010111011010101000;
assign LUT_3[60432] = 32'b00000000000000001111010011101110;
assign LUT_3[60433] = 32'b00000000000000010101111111001011;
assign LUT_3[60434] = 32'b00000000000000010001011011010010;
assign LUT_3[60435] = 32'b00000000000000011000000110101111;
assign LUT_3[60436] = 32'b00000000000000001100100001100100;
assign LUT_3[60437] = 32'b00000000000000010011001101000001;
assign LUT_3[60438] = 32'b00000000000000001110101001001000;
assign LUT_3[60439] = 32'b00000000000000010101010100100101;
assign LUT_3[60440] = 32'b00000000000000010100101100110100;
assign LUT_3[60441] = 32'b00000000000000011011011000010001;
assign LUT_3[60442] = 32'b00000000000000010110110100011000;
assign LUT_3[60443] = 32'b00000000000000011101011111110101;
assign LUT_3[60444] = 32'b00000000000000010001111010101010;
assign LUT_3[60445] = 32'b00000000000000011000100110000111;
assign LUT_3[60446] = 32'b00000000000000010100000010001110;
assign LUT_3[60447] = 32'b00000000000000011010101101101011;
assign LUT_3[60448] = 32'b00000000000000001101001111001011;
assign LUT_3[60449] = 32'b00000000000000010011111010101000;
assign LUT_3[60450] = 32'b00000000000000001111010110101111;
assign LUT_3[60451] = 32'b00000000000000010110000010001100;
assign LUT_3[60452] = 32'b00000000000000001010011101000001;
assign LUT_3[60453] = 32'b00000000000000010001001000011110;
assign LUT_3[60454] = 32'b00000000000000001100100100100101;
assign LUT_3[60455] = 32'b00000000000000010011010000000010;
assign LUT_3[60456] = 32'b00000000000000010010101000010001;
assign LUT_3[60457] = 32'b00000000000000011001010011101110;
assign LUT_3[60458] = 32'b00000000000000010100101111110101;
assign LUT_3[60459] = 32'b00000000000000011011011011010010;
assign LUT_3[60460] = 32'b00000000000000001111110110000111;
assign LUT_3[60461] = 32'b00000000000000010110100001100100;
assign LUT_3[60462] = 32'b00000000000000010001111101101011;
assign LUT_3[60463] = 32'b00000000000000011000101001001000;
assign LUT_3[60464] = 32'b00000000000000010000100010001110;
assign LUT_3[60465] = 32'b00000000000000010111001101101011;
assign LUT_3[60466] = 32'b00000000000000010010101001110010;
assign LUT_3[60467] = 32'b00000000000000011001010101001111;
assign LUT_3[60468] = 32'b00000000000000001101110000000100;
assign LUT_3[60469] = 32'b00000000000000010100011011100001;
assign LUT_3[60470] = 32'b00000000000000001111110111101000;
assign LUT_3[60471] = 32'b00000000000000010110100011000101;
assign LUT_3[60472] = 32'b00000000000000010101111011010100;
assign LUT_3[60473] = 32'b00000000000000011100100110110001;
assign LUT_3[60474] = 32'b00000000000000011000000010111000;
assign LUT_3[60475] = 32'b00000000000000011110101110010101;
assign LUT_3[60476] = 32'b00000000000000010011001001001010;
assign LUT_3[60477] = 32'b00000000000000011001110100100111;
assign LUT_3[60478] = 32'b00000000000000010101010000101110;
assign LUT_3[60479] = 32'b00000000000000011011111100001011;
assign LUT_3[60480] = 32'b00000000000000001011111001010110;
assign LUT_3[60481] = 32'b00000000000000010010100100110011;
assign LUT_3[60482] = 32'b00000000000000001110000000111010;
assign LUT_3[60483] = 32'b00000000000000010100101100010111;
assign LUT_3[60484] = 32'b00000000000000001001000111001100;
assign LUT_3[60485] = 32'b00000000000000001111110010101001;
assign LUT_3[60486] = 32'b00000000000000001011001110110000;
assign LUT_3[60487] = 32'b00000000000000010001111010001101;
assign LUT_3[60488] = 32'b00000000000000010001010010011100;
assign LUT_3[60489] = 32'b00000000000000010111111101111001;
assign LUT_3[60490] = 32'b00000000000000010011011010000000;
assign LUT_3[60491] = 32'b00000000000000011010000101011101;
assign LUT_3[60492] = 32'b00000000000000001110100000010010;
assign LUT_3[60493] = 32'b00000000000000010101001011101111;
assign LUT_3[60494] = 32'b00000000000000010000100111110110;
assign LUT_3[60495] = 32'b00000000000000010111010011010011;
assign LUT_3[60496] = 32'b00000000000000001111001100011001;
assign LUT_3[60497] = 32'b00000000000000010101110111110110;
assign LUT_3[60498] = 32'b00000000000000010001010011111101;
assign LUT_3[60499] = 32'b00000000000000010111111111011010;
assign LUT_3[60500] = 32'b00000000000000001100011010001111;
assign LUT_3[60501] = 32'b00000000000000010011000101101100;
assign LUT_3[60502] = 32'b00000000000000001110100001110011;
assign LUT_3[60503] = 32'b00000000000000010101001101010000;
assign LUT_3[60504] = 32'b00000000000000010100100101011111;
assign LUT_3[60505] = 32'b00000000000000011011010000111100;
assign LUT_3[60506] = 32'b00000000000000010110101101000011;
assign LUT_3[60507] = 32'b00000000000000011101011000100000;
assign LUT_3[60508] = 32'b00000000000000010001110011010101;
assign LUT_3[60509] = 32'b00000000000000011000011110110010;
assign LUT_3[60510] = 32'b00000000000000010011111010111001;
assign LUT_3[60511] = 32'b00000000000000011010100110010110;
assign LUT_3[60512] = 32'b00000000000000001101000111110110;
assign LUT_3[60513] = 32'b00000000000000010011110011010011;
assign LUT_3[60514] = 32'b00000000000000001111001111011010;
assign LUT_3[60515] = 32'b00000000000000010101111010110111;
assign LUT_3[60516] = 32'b00000000000000001010010101101100;
assign LUT_3[60517] = 32'b00000000000000010001000001001001;
assign LUT_3[60518] = 32'b00000000000000001100011101010000;
assign LUT_3[60519] = 32'b00000000000000010011001000101101;
assign LUT_3[60520] = 32'b00000000000000010010100000111100;
assign LUT_3[60521] = 32'b00000000000000011001001100011001;
assign LUT_3[60522] = 32'b00000000000000010100101000100000;
assign LUT_3[60523] = 32'b00000000000000011011010011111101;
assign LUT_3[60524] = 32'b00000000000000001111101110110010;
assign LUT_3[60525] = 32'b00000000000000010110011010001111;
assign LUT_3[60526] = 32'b00000000000000010001110110010110;
assign LUT_3[60527] = 32'b00000000000000011000100001110011;
assign LUT_3[60528] = 32'b00000000000000010000011010111001;
assign LUT_3[60529] = 32'b00000000000000010111000110010110;
assign LUT_3[60530] = 32'b00000000000000010010100010011101;
assign LUT_3[60531] = 32'b00000000000000011001001101111010;
assign LUT_3[60532] = 32'b00000000000000001101101000101111;
assign LUT_3[60533] = 32'b00000000000000010100010100001100;
assign LUT_3[60534] = 32'b00000000000000001111110000010011;
assign LUT_3[60535] = 32'b00000000000000010110011011110000;
assign LUT_3[60536] = 32'b00000000000000010101110011111111;
assign LUT_3[60537] = 32'b00000000000000011100011111011100;
assign LUT_3[60538] = 32'b00000000000000010111111011100011;
assign LUT_3[60539] = 32'b00000000000000011110100111000000;
assign LUT_3[60540] = 32'b00000000000000010011000001110101;
assign LUT_3[60541] = 32'b00000000000000011001101101010010;
assign LUT_3[60542] = 32'b00000000000000010101001001011001;
assign LUT_3[60543] = 32'b00000000000000011011110100110110;
assign LUT_3[60544] = 32'b00000000000000001110001011101001;
assign LUT_3[60545] = 32'b00000000000000010100110111000110;
assign LUT_3[60546] = 32'b00000000000000010000010011001101;
assign LUT_3[60547] = 32'b00000000000000010110111110101010;
assign LUT_3[60548] = 32'b00000000000000001011011001011111;
assign LUT_3[60549] = 32'b00000000000000010010000100111100;
assign LUT_3[60550] = 32'b00000000000000001101100001000011;
assign LUT_3[60551] = 32'b00000000000000010100001100100000;
assign LUT_3[60552] = 32'b00000000000000010011100100101111;
assign LUT_3[60553] = 32'b00000000000000011010010000001100;
assign LUT_3[60554] = 32'b00000000000000010101101100010011;
assign LUT_3[60555] = 32'b00000000000000011100010111110000;
assign LUT_3[60556] = 32'b00000000000000010000110010100101;
assign LUT_3[60557] = 32'b00000000000000010111011110000010;
assign LUT_3[60558] = 32'b00000000000000010010111010001001;
assign LUT_3[60559] = 32'b00000000000000011001100101100110;
assign LUT_3[60560] = 32'b00000000000000010001011110101100;
assign LUT_3[60561] = 32'b00000000000000011000001010001001;
assign LUT_3[60562] = 32'b00000000000000010011100110010000;
assign LUT_3[60563] = 32'b00000000000000011010010001101101;
assign LUT_3[60564] = 32'b00000000000000001110101100100010;
assign LUT_3[60565] = 32'b00000000000000010101010111111111;
assign LUT_3[60566] = 32'b00000000000000010000110100000110;
assign LUT_3[60567] = 32'b00000000000000010111011111100011;
assign LUT_3[60568] = 32'b00000000000000010110110111110010;
assign LUT_3[60569] = 32'b00000000000000011101100011001111;
assign LUT_3[60570] = 32'b00000000000000011000111111010110;
assign LUT_3[60571] = 32'b00000000000000011111101010110011;
assign LUT_3[60572] = 32'b00000000000000010100000101101000;
assign LUT_3[60573] = 32'b00000000000000011010110001000101;
assign LUT_3[60574] = 32'b00000000000000010110001101001100;
assign LUT_3[60575] = 32'b00000000000000011100111000101001;
assign LUT_3[60576] = 32'b00000000000000001111011010001001;
assign LUT_3[60577] = 32'b00000000000000010110000101100110;
assign LUT_3[60578] = 32'b00000000000000010001100001101101;
assign LUT_3[60579] = 32'b00000000000000011000001101001010;
assign LUT_3[60580] = 32'b00000000000000001100100111111111;
assign LUT_3[60581] = 32'b00000000000000010011010011011100;
assign LUT_3[60582] = 32'b00000000000000001110101111100011;
assign LUT_3[60583] = 32'b00000000000000010101011011000000;
assign LUT_3[60584] = 32'b00000000000000010100110011001111;
assign LUT_3[60585] = 32'b00000000000000011011011110101100;
assign LUT_3[60586] = 32'b00000000000000010110111010110011;
assign LUT_3[60587] = 32'b00000000000000011101100110010000;
assign LUT_3[60588] = 32'b00000000000000010010000001000101;
assign LUT_3[60589] = 32'b00000000000000011000101100100010;
assign LUT_3[60590] = 32'b00000000000000010100001000101001;
assign LUT_3[60591] = 32'b00000000000000011010110100000110;
assign LUT_3[60592] = 32'b00000000000000010010101101001100;
assign LUT_3[60593] = 32'b00000000000000011001011000101001;
assign LUT_3[60594] = 32'b00000000000000010100110100110000;
assign LUT_3[60595] = 32'b00000000000000011011100000001101;
assign LUT_3[60596] = 32'b00000000000000001111111011000010;
assign LUT_3[60597] = 32'b00000000000000010110100110011111;
assign LUT_3[60598] = 32'b00000000000000010010000010100110;
assign LUT_3[60599] = 32'b00000000000000011000101110000011;
assign LUT_3[60600] = 32'b00000000000000011000000110010010;
assign LUT_3[60601] = 32'b00000000000000011110110001101111;
assign LUT_3[60602] = 32'b00000000000000011010001101110110;
assign LUT_3[60603] = 32'b00000000000000100000111001010011;
assign LUT_3[60604] = 32'b00000000000000010101010100001000;
assign LUT_3[60605] = 32'b00000000000000011011111111100101;
assign LUT_3[60606] = 32'b00000000000000010111011011101100;
assign LUT_3[60607] = 32'b00000000000000011110000111001001;
assign LUT_3[60608] = 32'b00000000000000001110000100010100;
assign LUT_3[60609] = 32'b00000000000000010100101111110001;
assign LUT_3[60610] = 32'b00000000000000010000001011111000;
assign LUT_3[60611] = 32'b00000000000000010110110111010101;
assign LUT_3[60612] = 32'b00000000000000001011010010001010;
assign LUT_3[60613] = 32'b00000000000000010001111101100111;
assign LUT_3[60614] = 32'b00000000000000001101011001101110;
assign LUT_3[60615] = 32'b00000000000000010100000101001011;
assign LUT_3[60616] = 32'b00000000000000010011011101011010;
assign LUT_3[60617] = 32'b00000000000000011010001000110111;
assign LUT_3[60618] = 32'b00000000000000010101100100111110;
assign LUT_3[60619] = 32'b00000000000000011100010000011011;
assign LUT_3[60620] = 32'b00000000000000010000101011010000;
assign LUT_3[60621] = 32'b00000000000000010111010110101101;
assign LUT_3[60622] = 32'b00000000000000010010110010110100;
assign LUT_3[60623] = 32'b00000000000000011001011110010001;
assign LUT_3[60624] = 32'b00000000000000010001010111010111;
assign LUT_3[60625] = 32'b00000000000000011000000010110100;
assign LUT_3[60626] = 32'b00000000000000010011011110111011;
assign LUT_3[60627] = 32'b00000000000000011010001010011000;
assign LUT_3[60628] = 32'b00000000000000001110100101001101;
assign LUT_3[60629] = 32'b00000000000000010101010000101010;
assign LUT_3[60630] = 32'b00000000000000010000101100110001;
assign LUT_3[60631] = 32'b00000000000000010111011000001110;
assign LUT_3[60632] = 32'b00000000000000010110110000011101;
assign LUT_3[60633] = 32'b00000000000000011101011011111010;
assign LUT_3[60634] = 32'b00000000000000011000111000000001;
assign LUT_3[60635] = 32'b00000000000000011111100011011110;
assign LUT_3[60636] = 32'b00000000000000010011111110010011;
assign LUT_3[60637] = 32'b00000000000000011010101001110000;
assign LUT_3[60638] = 32'b00000000000000010110000101110111;
assign LUT_3[60639] = 32'b00000000000000011100110001010100;
assign LUT_3[60640] = 32'b00000000000000001111010010110100;
assign LUT_3[60641] = 32'b00000000000000010101111110010001;
assign LUT_3[60642] = 32'b00000000000000010001011010011000;
assign LUT_3[60643] = 32'b00000000000000011000000101110101;
assign LUT_3[60644] = 32'b00000000000000001100100000101010;
assign LUT_3[60645] = 32'b00000000000000010011001100000111;
assign LUT_3[60646] = 32'b00000000000000001110101000001110;
assign LUT_3[60647] = 32'b00000000000000010101010011101011;
assign LUT_3[60648] = 32'b00000000000000010100101011111010;
assign LUT_3[60649] = 32'b00000000000000011011010111010111;
assign LUT_3[60650] = 32'b00000000000000010110110011011110;
assign LUT_3[60651] = 32'b00000000000000011101011110111011;
assign LUT_3[60652] = 32'b00000000000000010001111001110000;
assign LUT_3[60653] = 32'b00000000000000011000100101001101;
assign LUT_3[60654] = 32'b00000000000000010100000001010100;
assign LUT_3[60655] = 32'b00000000000000011010101100110001;
assign LUT_3[60656] = 32'b00000000000000010010100101110111;
assign LUT_3[60657] = 32'b00000000000000011001010001010100;
assign LUT_3[60658] = 32'b00000000000000010100101101011011;
assign LUT_3[60659] = 32'b00000000000000011011011000111000;
assign LUT_3[60660] = 32'b00000000000000001111110011101101;
assign LUT_3[60661] = 32'b00000000000000010110011111001010;
assign LUT_3[60662] = 32'b00000000000000010001111011010001;
assign LUT_3[60663] = 32'b00000000000000011000100110101110;
assign LUT_3[60664] = 32'b00000000000000010111111110111101;
assign LUT_3[60665] = 32'b00000000000000011110101010011010;
assign LUT_3[60666] = 32'b00000000000000011010000110100001;
assign LUT_3[60667] = 32'b00000000000000100000110001111110;
assign LUT_3[60668] = 32'b00000000000000010101001100110011;
assign LUT_3[60669] = 32'b00000000000000011011111000010000;
assign LUT_3[60670] = 32'b00000000000000010111010100010111;
assign LUT_3[60671] = 32'b00000000000000011101111111110100;
assign LUT_3[60672] = 32'b00000000000000001000010000001100;
assign LUT_3[60673] = 32'b00000000000000001110111011101001;
assign LUT_3[60674] = 32'b00000000000000001010010111110000;
assign LUT_3[60675] = 32'b00000000000000010001000011001101;
assign LUT_3[60676] = 32'b00000000000000000101011110000010;
assign LUT_3[60677] = 32'b00000000000000001100001001011111;
assign LUT_3[60678] = 32'b00000000000000000111100101100110;
assign LUT_3[60679] = 32'b00000000000000001110010001000011;
assign LUT_3[60680] = 32'b00000000000000001101101001010010;
assign LUT_3[60681] = 32'b00000000000000010100010100101111;
assign LUT_3[60682] = 32'b00000000000000001111110000110110;
assign LUT_3[60683] = 32'b00000000000000010110011100010011;
assign LUT_3[60684] = 32'b00000000000000001010110111001000;
assign LUT_3[60685] = 32'b00000000000000010001100010100101;
assign LUT_3[60686] = 32'b00000000000000001100111110101100;
assign LUT_3[60687] = 32'b00000000000000010011101010001001;
assign LUT_3[60688] = 32'b00000000000000001011100011001111;
assign LUT_3[60689] = 32'b00000000000000010010001110101100;
assign LUT_3[60690] = 32'b00000000000000001101101010110011;
assign LUT_3[60691] = 32'b00000000000000010100010110010000;
assign LUT_3[60692] = 32'b00000000000000001000110001000101;
assign LUT_3[60693] = 32'b00000000000000001111011100100010;
assign LUT_3[60694] = 32'b00000000000000001010111000101001;
assign LUT_3[60695] = 32'b00000000000000010001100100000110;
assign LUT_3[60696] = 32'b00000000000000010000111100010101;
assign LUT_3[60697] = 32'b00000000000000010111100111110010;
assign LUT_3[60698] = 32'b00000000000000010011000011111001;
assign LUT_3[60699] = 32'b00000000000000011001101111010110;
assign LUT_3[60700] = 32'b00000000000000001110001010001011;
assign LUT_3[60701] = 32'b00000000000000010100110101101000;
assign LUT_3[60702] = 32'b00000000000000010000010001101111;
assign LUT_3[60703] = 32'b00000000000000010110111101001100;
assign LUT_3[60704] = 32'b00000000000000001001011110101100;
assign LUT_3[60705] = 32'b00000000000000010000001010001001;
assign LUT_3[60706] = 32'b00000000000000001011100110010000;
assign LUT_3[60707] = 32'b00000000000000010010010001101101;
assign LUT_3[60708] = 32'b00000000000000000110101100100010;
assign LUT_3[60709] = 32'b00000000000000001101010111111111;
assign LUT_3[60710] = 32'b00000000000000001000110100000110;
assign LUT_3[60711] = 32'b00000000000000001111011111100011;
assign LUT_3[60712] = 32'b00000000000000001110110111110010;
assign LUT_3[60713] = 32'b00000000000000010101100011001111;
assign LUT_3[60714] = 32'b00000000000000010000111111010110;
assign LUT_3[60715] = 32'b00000000000000010111101010110011;
assign LUT_3[60716] = 32'b00000000000000001100000101101000;
assign LUT_3[60717] = 32'b00000000000000010010110001000101;
assign LUT_3[60718] = 32'b00000000000000001110001101001100;
assign LUT_3[60719] = 32'b00000000000000010100111000101001;
assign LUT_3[60720] = 32'b00000000000000001100110001101111;
assign LUT_3[60721] = 32'b00000000000000010011011101001100;
assign LUT_3[60722] = 32'b00000000000000001110111001010011;
assign LUT_3[60723] = 32'b00000000000000010101100100110000;
assign LUT_3[60724] = 32'b00000000000000001001111111100101;
assign LUT_3[60725] = 32'b00000000000000010000101011000010;
assign LUT_3[60726] = 32'b00000000000000001100000111001001;
assign LUT_3[60727] = 32'b00000000000000010010110010100110;
assign LUT_3[60728] = 32'b00000000000000010010001010110101;
assign LUT_3[60729] = 32'b00000000000000011000110110010010;
assign LUT_3[60730] = 32'b00000000000000010100010010011001;
assign LUT_3[60731] = 32'b00000000000000011010111101110110;
assign LUT_3[60732] = 32'b00000000000000001111011000101011;
assign LUT_3[60733] = 32'b00000000000000010110000100001000;
assign LUT_3[60734] = 32'b00000000000000010001100000001111;
assign LUT_3[60735] = 32'b00000000000000011000001011101100;
assign LUT_3[60736] = 32'b00000000000000001000001000110111;
assign LUT_3[60737] = 32'b00000000000000001110110100010100;
assign LUT_3[60738] = 32'b00000000000000001010010000011011;
assign LUT_3[60739] = 32'b00000000000000010000111011111000;
assign LUT_3[60740] = 32'b00000000000000000101010110101101;
assign LUT_3[60741] = 32'b00000000000000001100000010001010;
assign LUT_3[60742] = 32'b00000000000000000111011110010001;
assign LUT_3[60743] = 32'b00000000000000001110001001101110;
assign LUT_3[60744] = 32'b00000000000000001101100001111101;
assign LUT_3[60745] = 32'b00000000000000010100001101011010;
assign LUT_3[60746] = 32'b00000000000000001111101001100001;
assign LUT_3[60747] = 32'b00000000000000010110010100111110;
assign LUT_3[60748] = 32'b00000000000000001010101111110011;
assign LUT_3[60749] = 32'b00000000000000010001011011010000;
assign LUT_3[60750] = 32'b00000000000000001100110111010111;
assign LUT_3[60751] = 32'b00000000000000010011100010110100;
assign LUT_3[60752] = 32'b00000000000000001011011011111010;
assign LUT_3[60753] = 32'b00000000000000010010000111010111;
assign LUT_3[60754] = 32'b00000000000000001101100011011110;
assign LUT_3[60755] = 32'b00000000000000010100001110111011;
assign LUT_3[60756] = 32'b00000000000000001000101001110000;
assign LUT_3[60757] = 32'b00000000000000001111010101001101;
assign LUT_3[60758] = 32'b00000000000000001010110001010100;
assign LUT_3[60759] = 32'b00000000000000010001011100110001;
assign LUT_3[60760] = 32'b00000000000000010000110101000000;
assign LUT_3[60761] = 32'b00000000000000010111100000011101;
assign LUT_3[60762] = 32'b00000000000000010010111100100100;
assign LUT_3[60763] = 32'b00000000000000011001101000000001;
assign LUT_3[60764] = 32'b00000000000000001110000010110110;
assign LUT_3[60765] = 32'b00000000000000010100101110010011;
assign LUT_3[60766] = 32'b00000000000000010000001010011010;
assign LUT_3[60767] = 32'b00000000000000010110110101110111;
assign LUT_3[60768] = 32'b00000000000000001001010111010111;
assign LUT_3[60769] = 32'b00000000000000010000000010110100;
assign LUT_3[60770] = 32'b00000000000000001011011110111011;
assign LUT_3[60771] = 32'b00000000000000010010001010011000;
assign LUT_3[60772] = 32'b00000000000000000110100101001101;
assign LUT_3[60773] = 32'b00000000000000001101010000101010;
assign LUT_3[60774] = 32'b00000000000000001000101100110001;
assign LUT_3[60775] = 32'b00000000000000001111011000001110;
assign LUT_3[60776] = 32'b00000000000000001110110000011101;
assign LUT_3[60777] = 32'b00000000000000010101011011111010;
assign LUT_3[60778] = 32'b00000000000000010000111000000001;
assign LUT_3[60779] = 32'b00000000000000010111100011011110;
assign LUT_3[60780] = 32'b00000000000000001011111110010011;
assign LUT_3[60781] = 32'b00000000000000010010101001110000;
assign LUT_3[60782] = 32'b00000000000000001110000101110111;
assign LUT_3[60783] = 32'b00000000000000010100110001010100;
assign LUT_3[60784] = 32'b00000000000000001100101010011010;
assign LUT_3[60785] = 32'b00000000000000010011010101110111;
assign LUT_3[60786] = 32'b00000000000000001110110001111110;
assign LUT_3[60787] = 32'b00000000000000010101011101011011;
assign LUT_3[60788] = 32'b00000000000000001001111000010000;
assign LUT_3[60789] = 32'b00000000000000010000100011101101;
assign LUT_3[60790] = 32'b00000000000000001011111111110100;
assign LUT_3[60791] = 32'b00000000000000010010101011010001;
assign LUT_3[60792] = 32'b00000000000000010010000011100000;
assign LUT_3[60793] = 32'b00000000000000011000101110111101;
assign LUT_3[60794] = 32'b00000000000000010100001011000100;
assign LUT_3[60795] = 32'b00000000000000011010110110100001;
assign LUT_3[60796] = 32'b00000000000000001111010001010110;
assign LUT_3[60797] = 32'b00000000000000010101111100110011;
assign LUT_3[60798] = 32'b00000000000000010001011000111010;
assign LUT_3[60799] = 32'b00000000000000011000000100010111;
assign LUT_3[60800] = 32'b00000000000000001010011011001010;
assign LUT_3[60801] = 32'b00000000000000010001000110100111;
assign LUT_3[60802] = 32'b00000000000000001100100010101110;
assign LUT_3[60803] = 32'b00000000000000010011001110001011;
assign LUT_3[60804] = 32'b00000000000000000111101001000000;
assign LUT_3[60805] = 32'b00000000000000001110010100011101;
assign LUT_3[60806] = 32'b00000000000000001001110000100100;
assign LUT_3[60807] = 32'b00000000000000010000011100000001;
assign LUT_3[60808] = 32'b00000000000000001111110100010000;
assign LUT_3[60809] = 32'b00000000000000010110011111101101;
assign LUT_3[60810] = 32'b00000000000000010001111011110100;
assign LUT_3[60811] = 32'b00000000000000011000100111010001;
assign LUT_3[60812] = 32'b00000000000000001101000010000110;
assign LUT_3[60813] = 32'b00000000000000010011101101100011;
assign LUT_3[60814] = 32'b00000000000000001111001001101010;
assign LUT_3[60815] = 32'b00000000000000010101110101000111;
assign LUT_3[60816] = 32'b00000000000000001101101110001101;
assign LUT_3[60817] = 32'b00000000000000010100011001101010;
assign LUT_3[60818] = 32'b00000000000000001111110101110001;
assign LUT_3[60819] = 32'b00000000000000010110100001001110;
assign LUT_3[60820] = 32'b00000000000000001010111100000011;
assign LUT_3[60821] = 32'b00000000000000010001100111100000;
assign LUT_3[60822] = 32'b00000000000000001101000011100111;
assign LUT_3[60823] = 32'b00000000000000010011101111000100;
assign LUT_3[60824] = 32'b00000000000000010011000111010011;
assign LUT_3[60825] = 32'b00000000000000011001110010110000;
assign LUT_3[60826] = 32'b00000000000000010101001110110111;
assign LUT_3[60827] = 32'b00000000000000011011111010010100;
assign LUT_3[60828] = 32'b00000000000000010000010101001001;
assign LUT_3[60829] = 32'b00000000000000010111000000100110;
assign LUT_3[60830] = 32'b00000000000000010010011100101101;
assign LUT_3[60831] = 32'b00000000000000011001001000001010;
assign LUT_3[60832] = 32'b00000000000000001011101001101010;
assign LUT_3[60833] = 32'b00000000000000010010010101000111;
assign LUT_3[60834] = 32'b00000000000000001101110001001110;
assign LUT_3[60835] = 32'b00000000000000010100011100101011;
assign LUT_3[60836] = 32'b00000000000000001000110111100000;
assign LUT_3[60837] = 32'b00000000000000001111100010111101;
assign LUT_3[60838] = 32'b00000000000000001010111111000100;
assign LUT_3[60839] = 32'b00000000000000010001101010100001;
assign LUT_3[60840] = 32'b00000000000000010001000010110000;
assign LUT_3[60841] = 32'b00000000000000010111101110001101;
assign LUT_3[60842] = 32'b00000000000000010011001010010100;
assign LUT_3[60843] = 32'b00000000000000011001110101110001;
assign LUT_3[60844] = 32'b00000000000000001110010000100110;
assign LUT_3[60845] = 32'b00000000000000010100111100000011;
assign LUT_3[60846] = 32'b00000000000000010000011000001010;
assign LUT_3[60847] = 32'b00000000000000010111000011100111;
assign LUT_3[60848] = 32'b00000000000000001110111100101101;
assign LUT_3[60849] = 32'b00000000000000010101101000001010;
assign LUT_3[60850] = 32'b00000000000000010001000100010001;
assign LUT_3[60851] = 32'b00000000000000010111101111101110;
assign LUT_3[60852] = 32'b00000000000000001100001010100011;
assign LUT_3[60853] = 32'b00000000000000010010110110000000;
assign LUT_3[60854] = 32'b00000000000000001110010010000111;
assign LUT_3[60855] = 32'b00000000000000010100111101100100;
assign LUT_3[60856] = 32'b00000000000000010100010101110011;
assign LUT_3[60857] = 32'b00000000000000011011000001010000;
assign LUT_3[60858] = 32'b00000000000000010110011101010111;
assign LUT_3[60859] = 32'b00000000000000011101001000110100;
assign LUT_3[60860] = 32'b00000000000000010001100011101001;
assign LUT_3[60861] = 32'b00000000000000011000001111000110;
assign LUT_3[60862] = 32'b00000000000000010011101011001101;
assign LUT_3[60863] = 32'b00000000000000011010010110101010;
assign LUT_3[60864] = 32'b00000000000000001010010011110101;
assign LUT_3[60865] = 32'b00000000000000010000111111010010;
assign LUT_3[60866] = 32'b00000000000000001100011011011001;
assign LUT_3[60867] = 32'b00000000000000010011000110110110;
assign LUT_3[60868] = 32'b00000000000000000111100001101011;
assign LUT_3[60869] = 32'b00000000000000001110001101001000;
assign LUT_3[60870] = 32'b00000000000000001001101001001111;
assign LUT_3[60871] = 32'b00000000000000010000010100101100;
assign LUT_3[60872] = 32'b00000000000000001111101100111011;
assign LUT_3[60873] = 32'b00000000000000010110011000011000;
assign LUT_3[60874] = 32'b00000000000000010001110100011111;
assign LUT_3[60875] = 32'b00000000000000011000011111111100;
assign LUT_3[60876] = 32'b00000000000000001100111010110001;
assign LUT_3[60877] = 32'b00000000000000010011100110001110;
assign LUT_3[60878] = 32'b00000000000000001111000010010101;
assign LUT_3[60879] = 32'b00000000000000010101101101110010;
assign LUT_3[60880] = 32'b00000000000000001101100110111000;
assign LUT_3[60881] = 32'b00000000000000010100010010010101;
assign LUT_3[60882] = 32'b00000000000000001111101110011100;
assign LUT_3[60883] = 32'b00000000000000010110011001111001;
assign LUT_3[60884] = 32'b00000000000000001010110100101110;
assign LUT_3[60885] = 32'b00000000000000010001100000001011;
assign LUT_3[60886] = 32'b00000000000000001100111100010010;
assign LUT_3[60887] = 32'b00000000000000010011100111101111;
assign LUT_3[60888] = 32'b00000000000000010010111111111110;
assign LUT_3[60889] = 32'b00000000000000011001101011011011;
assign LUT_3[60890] = 32'b00000000000000010101000111100010;
assign LUT_3[60891] = 32'b00000000000000011011110010111111;
assign LUT_3[60892] = 32'b00000000000000010000001101110100;
assign LUT_3[60893] = 32'b00000000000000010110111001010001;
assign LUT_3[60894] = 32'b00000000000000010010010101011000;
assign LUT_3[60895] = 32'b00000000000000011001000000110101;
assign LUT_3[60896] = 32'b00000000000000001011100010010101;
assign LUT_3[60897] = 32'b00000000000000010010001101110010;
assign LUT_3[60898] = 32'b00000000000000001101101001111001;
assign LUT_3[60899] = 32'b00000000000000010100010101010110;
assign LUT_3[60900] = 32'b00000000000000001000110000001011;
assign LUT_3[60901] = 32'b00000000000000001111011011101000;
assign LUT_3[60902] = 32'b00000000000000001010110111101111;
assign LUT_3[60903] = 32'b00000000000000010001100011001100;
assign LUT_3[60904] = 32'b00000000000000010000111011011011;
assign LUT_3[60905] = 32'b00000000000000010111100110111000;
assign LUT_3[60906] = 32'b00000000000000010011000010111111;
assign LUT_3[60907] = 32'b00000000000000011001101110011100;
assign LUT_3[60908] = 32'b00000000000000001110001001010001;
assign LUT_3[60909] = 32'b00000000000000010100110100101110;
assign LUT_3[60910] = 32'b00000000000000010000010000110101;
assign LUT_3[60911] = 32'b00000000000000010110111100010010;
assign LUT_3[60912] = 32'b00000000000000001110110101011000;
assign LUT_3[60913] = 32'b00000000000000010101100000110101;
assign LUT_3[60914] = 32'b00000000000000010000111100111100;
assign LUT_3[60915] = 32'b00000000000000010111101000011001;
assign LUT_3[60916] = 32'b00000000000000001100000011001110;
assign LUT_3[60917] = 32'b00000000000000010010101110101011;
assign LUT_3[60918] = 32'b00000000000000001110001010110010;
assign LUT_3[60919] = 32'b00000000000000010100110110001111;
assign LUT_3[60920] = 32'b00000000000000010100001110011110;
assign LUT_3[60921] = 32'b00000000000000011010111001111011;
assign LUT_3[60922] = 32'b00000000000000010110010110000010;
assign LUT_3[60923] = 32'b00000000000000011101000001011111;
assign LUT_3[60924] = 32'b00000000000000010001011100010100;
assign LUT_3[60925] = 32'b00000000000000011000000111110001;
assign LUT_3[60926] = 32'b00000000000000010011100011111000;
assign LUT_3[60927] = 32'b00000000000000011010001111010101;
assign LUT_3[60928] = 32'b00000000000000001111010101110111;
assign LUT_3[60929] = 32'b00000000000000010110000001010100;
assign LUT_3[60930] = 32'b00000000000000010001011101011011;
assign LUT_3[60931] = 32'b00000000000000011000001000111000;
assign LUT_3[60932] = 32'b00000000000000001100100011101101;
assign LUT_3[60933] = 32'b00000000000000010011001111001010;
assign LUT_3[60934] = 32'b00000000000000001110101011010001;
assign LUT_3[60935] = 32'b00000000000000010101010110101110;
assign LUT_3[60936] = 32'b00000000000000010100101110111101;
assign LUT_3[60937] = 32'b00000000000000011011011010011010;
assign LUT_3[60938] = 32'b00000000000000010110110110100001;
assign LUT_3[60939] = 32'b00000000000000011101100001111110;
assign LUT_3[60940] = 32'b00000000000000010001111100110011;
assign LUT_3[60941] = 32'b00000000000000011000101000010000;
assign LUT_3[60942] = 32'b00000000000000010100000100010111;
assign LUT_3[60943] = 32'b00000000000000011010101111110100;
assign LUT_3[60944] = 32'b00000000000000010010101000111010;
assign LUT_3[60945] = 32'b00000000000000011001010100010111;
assign LUT_3[60946] = 32'b00000000000000010100110000011110;
assign LUT_3[60947] = 32'b00000000000000011011011011111011;
assign LUT_3[60948] = 32'b00000000000000001111110110110000;
assign LUT_3[60949] = 32'b00000000000000010110100010001101;
assign LUT_3[60950] = 32'b00000000000000010001111110010100;
assign LUT_3[60951] = 32'b00000000000000011000101001110001;
assign LUT_3[60952] = 32'b00000000000000011000000010000000;
assign LUT_3[60953] = 32'b00000000000000011110101101011101;
assign LUT_3[60954] = 32'b00000000000000011010001001100100;
assign LUT_3[60955] = 32'b00000000000000100000110101000001;
assign LUT_3[60956] = 32'b00000000000000010101001111110110;
assign LUT_3[60957] = 32'b00000000000000011011111011010011;
assign LUT_3[60958] = 32'b00000000000000010111010111011010;
assign LUT_3[60959] = 32'b00000000000000011110000010110111;
assign LUT_3[60960] = 32'b00000000000000010000100100010111;
assign LUT_3[60961] = 32'b00000000000000010111001111110100;
assign LUT_3[60962] = 32'b00000000000000010010101011111011;
assign LUT_3[60963] = 32'b00000000000000011001010111011000;
assign LUT_3[60964] = 32'b00000000000000001101110010001101;
assign LUT_3[60965] = 32'b00000000000000010100011101101010;
assign LUT_3[60966] = 32'b00000000000000001111111001110001;
assign LUT_3[60967] = 32'b00000000000000010110100101001110;
assign LUT_3[60968] = 32'b00000000000000010101111101011101;
assign LUT_3[60969] = 32'b00000000000000011100101000111010;
assign LUT_3[60970] = 32'b00000000000000011000000101000001;
assign LUT_3[60971] = 32'b00000000000000011110110000011110;
assign LUT_3[60972] = 32'b00000000000000010011001011010011;
assign LUT_3[60973] = 32'b00000000000000011001110110110000;
assign LUT_3[60974] = 32'b00000000000000010101010010110111;
assign LUT_3[60975] = 32'b00000000000000011011111110010100;
assign LUT_3[60976] = 32'b00000000000000010011110111011010;
assign LUT_3[60977] = 32'b00000000000000011010100010110111;
assign LUT_3[60978] = 32'b00000000000000010101111110111110;
assign LUT_3[60979] = 32'b00000000000000011100101010011011;
assign LUT_3[60980] = 32'b00000000000000010001000101010000;
assign LUT_3[60981] = 32'b00000000000000010111110000101101;
assign LUT_3[60982] = 32'b00000000000000010011001100110100;
assign LUT_3[60983] = 32'b00000000000000011001111000010001;
assign LUT_3[60984] = 32'b00000000000000011001010000100000;
assign LUT_3[60985] = 32'b00000000000000011111111011111101;
assign LUT_3[60986] = 32'b00000000000000011011011000000100;
assign LUT_3[60987] = 32'b00000000000000100010000011100001;
assign LUT_3[60988] = 32'b00000000000000010110011110010110;
assign LUT_3[60989] = 32'b00000000000000011101001001110011;
assign LUT_3[60990] = 32'b00000000000000011000100101111010;
assign LUT_3[60991] = 32'b00000000000000011111010001010111;
assign LUT_3[60992] = 32'b00000000000000001111001110100010;
assign LUT_3[60993] = 32'b00000000000000010101111001111111;
assign LUT_3[60994] = 32'b00000000000000010001010110000110;
assign LUT_3[60995] = 32'b00000000000000011000000001100011;
assign LUT_3[60996] = 32'b00000000000000001100011100011000;
assign LUT_3[60997] = 32'b00000000000000010011000111110101;
assign LUT_3[60998] = 32'b00000000000000001110100011111100;
assign LUT_3[60999] = 32'b00000000000000010101001111011001;
assign LUT_3[61000] = 32'b00000000000000010100100111101000;
assign LUT_3[61001] = 32'b00000000000000011011010011000101;
assign LUT_3[61002] = 32'b00000000000000010110101111001100;
assign LUT_3[61003] = 32'b00000000000000011101011010101001;
assign LUT_3[61004] = 32'b00000000000000010001110101011110;
assign LUT_3[61005] = 32'b00000000000000011000100000111011;
assign LUT_3[61006] = 32'b00000000000000010011111101000010;
assign LUT_3[61007] = 32'b00000000000000011010101000011111;
assign LUT_3[61008] = 32'b00000000000000010010100001100101;
assign LUT_3[61009] = 32'b00000000000000011001001101000010;
assign LUT_3[61010] = 32'b00000000000000010100101001001001;
assign LUT_3[61011] = 32'b00000000000000011011010100100110;
assign LUT_3[61012] = 32'b00000000000000001111101111011011;
assign LUT_3[61013] = 32'b00000000000000010110011010111000;
assign LUT_3[61014] = 32'b00000000000000010001110110111111;
assign LUT_3[61015] = 32'b00000000000000011000100010011100;
assign LUT_3[61016] = 32'b00000000000000010111111010101011;
assign LUT_3[61017] = 32'b00000000000000011110100110001000;
assign LUT_3[61018] = 32'b00000000000000011010000010001111;
assign LUT_3[61019] = 32'b00000000000000100000101101101100;
assign LUT_3[61020] = 32'b00000000000000010101001000100001;
assign LUT_3[61021] = 32'b00000000000000011011110011111110;
assign LUT_3[61022] = 32'b00000000000000010111010000000101;
assign LUT_3[61023] = 32'b00000000000000011101111011100010;
assign LUT_3[61024] = 32'b00000000000000010000011101000010;
assign LUT_3[61025] = 32'b00000000000000010111001000011111;
assign LUT_3[61026] = 32'b00000000000000010010100100100110;
assign LUT_3[61027] = 32'b00000000000000011001010000000011;
assign LUT_3[61028] = 32'b00000000000000001101101010111000;
assign LUT_3[61029] = 32'b00000000000000010100010110010101;
assign LUT_3[61030] = 32'b00000000000000001111110010011100;
assign LUT_3[61031] = 32'b00000000000000010110011101111001;
assign LUT_3[61032] = 32'b00000000000000010101110110001000;
assign LUT_3[61033] = 32'b00000000000000011100100001100101;
assign LUT_3[61034] = 32'b00000000000000010111111101101100;
assign LUT_3[61035] = 32'b00000000000000011110101001001001;
assign LUT_3[61036] = 32'b00000000000000010011000011111110;
assign LUT_3[61037] = 32'b00000000000000011001101111011011;
assign LUT_3[61038] = 32'b00000000000000010101001011100010;
assign LUT_3[61039] = 32'b00000000000000011011110110111111;
assign LUT_3[61040] = 32'b00000000000000010011110000000101;
assign LUT_3[61041] = 32'b00000000000000011010011011100010;
assign LUT_3[61042] = 32'b00000000000000010101110111101001;
assign LUT_3[61043] = 32'b00000000000000011100100011000110;
assign LUT_3[61044] = 32'b00000000000000010000111101111011;
assign LUT_3[61045] = 32'b00000000000000010111101001011000;
assign LUT_3[61046] = 32'b00000000000000010011000101011111;
assign LUT_3[61047] = 32'b00000000000000011001110000111100;
assign LUT_3[61048] = 32'b00000000000000011001001001001011;
assign LUT_3[61049] = 32'b00000000000000011111110100101000;
assign LUT_3[61050] = 32'b00000000000000011011010000101111;
assign LUT_3[61051] = 32'b00000000000000100001111100001100;
assign LUT_3[61052] = 32'b00000000000000010110010111000001;
assign LUT_3[61053] = 32'b00000000000000011101000010011110;
assign LUT_3[61054] = 32'b00000000000000011000011110100101;
assign LUT_3[61055] = 32'b00000000000000011111001010000010;
assign LUT_3[61056] = 32'b00000000000000010001100000110101;
assign LUT_3[61057] = 32'b00000000000000011000001100010010;
assign LUT_3[61058] = 32'b00000000000000010011101000011001;
assign LUT_3[61059] = 32'b00000000000000011010010011110110;
assign LUT_3[61060] = 32'b00000000000000001110101110101011;
assign LUT_3[61061] = 32'b00000000000000010101011010001000;
assign LUT_3[61062] = 32'b00000000000000010000110110001111;
assign LUT_3[61063] = 32'b00000000000000010111100001101100;
assign LUT_3[61064] = 32'b00000000000000010110111001111011;
assign LUT_3[61065] = 32'b00000000000000011101100101011000;
assign LUT_3[61066] = 32'b00000000000000011001000001011111;
assign LUT_3[61067] = 32'b00000000000000011111101100111100;
assign LUT_3[61068] = 32'b00000000000000010100000111110001;
assign LUT_3[61069] = 32'b00000000000000011010110011001110;
assign LUT_3[61070] = 32'b00000000000000010110001111010101;
assign LUT_3[61071] = 32'b00000000000000011100111010110010;
assign LUT_3[61072] = 32'b00000000000000010100110011111000;
assign LUT_3[61073] = 32'b00000000000000011011011111010101;
assign LUT_3[61074] = 32'b00000000000000010110111011011100;
assign LUT_3[61075] = 32'b00000000000000011101100110111001;
assign LUT_3[61076] = 32'b00000000000000010010000001101110;
assign LUT_3[61077] = 32'b00000000000000011000101101001011;
assign LUT_3[61078] = 32'b00000000000000010100001001010010;
assign LUT_3[61079] = 32'b00000000000000011010110100101111;
assign LUT_3[61080] = 32'b00000000000000011010001100111110;
assign LUT_3[61081] = 32'b00000000000000100000111000011011;
assign LUT_3[61082] = 32'b00000000000000011100010100100010;
assign LUT_3[61083] = 32'b00000000000000100010111111111111;
assign LUT_3[61084] = 32'b00000000000000010111011010110100;
assign LUT_3[61085] = 32'b00000000000000011110000110010001;
assign LUT_3[61086] = 32'b00000000000000011001100010011000;
assign LUT_3[61087] = 32'b00000000000000100000001101110101;
assign LUT_3[61088] = 32'b00000000000000010010101111010101;
assign LUT_3[61089] = 32'b00000000000000011001011010110010;
assign LUT_3[61090] = 32'b00000000000000010100110110111001;
assign LUT_3[61091] = 32'b00000000000000011011100010010110;
assign LUT_3[61092] = 32'b00000000000000001111111101001011;
assign LUT_3[61093] = 32'b00000000000000010110101000101000;
assign LUT_3[61094] = 32'b00000000000000010010000100101111;
assign LUT_3[61095] = 32'b00000000000000011000110000001100;
assign LUT_3[61096] = 32'b00000000000000011000001000011011;
assign LUT_3[61097] = 32'b00000000000000011110110011111000;
assign LUT_3[61098] = 32'b00000000000000011010001111111111;
assign LUT_3[61099] = 32'b00000000000000100000111011011100;
assign LUT_3[61100] = 32'b00000000000000010101010110010001;
assign LUT_3[61101] = 32'b00000000000000011100000001101110;
assign LUT_3[61102] = 32'b00000000000000010111011101110101;
assign LUT_3[61103] = 32'b00000000000000011110001001010010;
assign LUT_3[61104] = 32'b00000000000000010110000010011000;
assign LUT_3[61105] = 32'b00000000000000011100101101110101;
assign LUT_3[61106] = 32'b00000000000000011000001001111100;
assign LUT_3[61107] = 32'b00000000000000011110110101011001;
assign LUT_3[61108] = 32'b00000000000000010011010000001110;
assign LUT_3[61109] = 32'b00000000000000011001111011101011;
assign LUT_3[61110] = 32'b00000000000000010101010111110010;
assign LUT_3[61111] = 32'b00000000000000011100000011001111;
assign LUT_3[61112] = 32'b00000000000000011011011011011110;
assign LUT_3[61113] = 32'b00000000000000100010000110111011;
assign LUT_3[61114] = 32'b00000000000000011101100011000010;
assign LUT_3[61115] = 32'b00000000000000100100001110011111;
assign LUT_3[61116] = 32'b00000000000000011000101001010100;
assign LUT_3[61117] = 32'b00000000000000011111010100110001;
assign LUT_3[61118] = 32'b00000000000000011010110000111000;
assign LUT_3[61119] = 32'b00000000000000100001011100010101;
assign LUT_3[61120] = 32'b00000000000000010001011001100000;
assign LUT_3[61121] = 32'b00000000000000011000000100111101;
assign LUT_3[61122] = 32'b00000000000000010011100001000100;
assign LUT_3[61123] = 32'b00000000000000011010001100100001;
assign LUT_3[61124] = 32'b00000000000000001110100111010110;
assign LUT_3[61125] = 32'b00000000000000010101010010110011;
assign LUT_3[61126] = 32'b00000000000000010000101110111010;
assign LUT_3[61127] = 32'b00000000000000010111011010010111;
assign LUT_3[61128] = 32'b00000000000000010110110010100110;
assign LUT_3[61129] = 32'b00000000000000011101011110000011;
assign LUT_3[61130] = 32'b00000000000000011000111010001010;
assign LUT_3[61131] = 32'b00000000000000011111100101100111;
assign LUT_3[61132] = 32'b00000000000000010100000000011100;
assign LUT_3[61133] = 32'b00000000000000011010101011111001;
assign LUT_3[61134] = 32'b00000000000000010110001000000000;
assign LUT_3[61135] = 32'b00000000000000011100110011011101;
assign LUT_3[61136] = 32'b00000000000000010100101100100011;
assign LUT_3[61137] = 32'b00000000000000011011011000000000;
assign LUT_3[61138] = 32'b00000000000000010110110100000111;
assign LUT_3[61139] = 32'b00000000000000011101011111100100;
assign LUT_3[61140] = 32'b00000000000000010001111010011001;
assign LUT_3[61141] = 32'b00000000000000011000100101110110;
assign LUT_3[61142] = 32'b00000000000000010100000001111101;
assign LUT_3[61143] = 32'b00000000000000011010101101011010;
assign LUT_3[61144] = 32'b00000000000000011010000101101001;
assign LUT_3[61145] = 32'b00000000000000100000110001000110;
assign LUT_3[61146] = 32'b00000000000000011100001101001101;
assign LUT_3[61147] = 32'b00000000000000100010111000101010;
assign LUT_3[61148] = 32'b00000000000000010111010011011111;
assign LUT_3[61149] = 32'b00000000000000011101111110111100;
assign LUT_3[61150] = 32'b00000000000000011001011011000011;
assign LUT_3[61151] = 32'b00000000000000100000000110100000;
assign LUT_3[61152] = 32'b00000000000000010010101000000000;
assign LUT_3[61153] = 32'b00000000000000011001010011011101;
assign LUT_3[61154] = 32'b00000000000000010100101111100100;
assign LUT_3[61155] = 32'b00000000000000011011011011000001;
assign LUT_3[61156] = 32'b00000000000000001111110101110110;
assign LUT_3[61157] = 32'b00000000000000010110100001010011;
assign LUT_3[61158] = 32'b00000000000000010001111101011010;
assign LUT_3[61159] = 32'b00000000000000011000101000110111;
assign LUT_3[61160] = 32'b00000000000000011000000001000110;
assign LUT_3[61161] = 32'b00000000000000011110101100100011;
assign LUT_3[61162] = 32'b00000000000000011010001000101010;
assign LUT_3[61163] = 32'b00000000000000100000110100000111;
assign LUT_3[61164] = 32'b00000000000000010101001110111100;
assign LUT_3[61165] = 32'b00000000000000011011111010011001;
assign LUT_3[61166] = 32'b00000000000000010111010110100000;
assign LUT_3[61167] = 32'b00000000000000011110000001111101;
assign LUT_3[61168] = 32'b00000000000000010101111011000011;
assign LUT_3[61169] = 32'b00000000000000011100100110100000;
assign LUT_3[61170] = 32'b00000000000000011000000010100111;
assign LUT_3[61171] = 32'b00000000000000011110101110000100;
assign LUT_3[61172] = 32'b00000000000000010011001000111001;
assign LUT_3[61173] = 32'b00000000000000011001110100010110;
assign LUT_3[61174] = 32'b00000000000000010101010000011101;
assign LUT_3[61175] = 32'b00000000000000011011111011111010;
assign LUT_3[61176] = 32'b00000000000000011011010100001001;
assign LUT_3[61177] = 32'b00000000000000100001111111100110;
assign LUT_3[61178] = 32'b00000000000000011101011011101101;
assign LUT_3[61179] = 32'b00000000000000100100000111001010;
assign LUT_3[61180] = 32'b00000000000000011000100001111111;
assign LUT_3[61181] = 32'b00000000000000011111001101011100;
assign LUT_3[61182] = 32'b00000000000000011010101001100011;
assign LUT_3[61183] = 32'b00000000000000100001010101000000;
assign LUT_3[61184] = 32'b00000000000000001011100101011000;
assign LUT_3[61185] = 32'b00000000000000010010010000110101;
assign LUT_3[61186] = 32'b00000000000000001101101100111100;
assign LUT_3[61187] = 32'b00000000000000010100011000011001;
assign LUT_3[61188] = 32'b00000000000000001000110011001110;
assign LUT_3[61189] = 32'b00000000000000001111011110101011;
assign LUT_3[61190] = 32'b00000000000000001010111010110010;
assign LUT_3[61191] = 32'b00000000000000010001100110001111;
assign LUT_3[61192] = 32'b00000000000000010000111110011110;
assign LUT_3[61193] = 32'b00000000000000010111101001111011;
assign LUT_3[61194] = 32'b00000000000000010011000110000010;
assign LUT_3[61195] = 32'b00000000000000011001110001011111;
assign LUT_3[61196] = 32'b00000000000000001110001100010100;
assign LUT_3[61197] = 32'b00000000000000010100110111110001;
assign LUT_3[61198] = 32'b00000000000000010000010011111000;
assign LUT_3[61199] = 32'b00000000000000010110111111010101;
assign LUT_3[61200] = 32'b00000000000000001110111000011011;
assign LUT_3[61201] = 32'b00000000000000010101100011111000;
assign LUT_3[61202] = 32'b00000000000000010000111111111111;
assign LUT_3[61203] = 32'b00000000000000010111101011011100;
assign LUT_3[61204] = 32'b00000000000000001100000110010001;
assign LUT_3[61205] = 32'b00000000000000010010110001101110;
assign LUT_3[61206] = 32'b00000000000000001110001101110101;
assign LUT_3[61207] = 32'b00000000000000010100111001010010;
assign LUT_3[61208] = 32'b00000000000000010100010001100001;
assign LUT_3[61209] = 32'b00000000000000011010111100111110;
assign LUT_3[61210] = 32'b00000000000000010110011001000101;
assign LUT_3[61211] = 32'b00000000000000011101000100100010;
assign LUT_3[61212] = 32'b00000000000000010001011111010111;
assign LUT_3[61213] = 32'b00000000000000011000001010110100;
assign LUT_3[61214] = 32'b00000000000000010011100110111011;
assign LUT_3[61215] = 32'b00000000000000011010010010011000;
assign LUT_3[61216] = 32'b00000000000000001100110011111000;
assign LUT_3[61217] = 32'b00000000000000010011011111010101;
assign LUT_3[61218] = 32'b00000000000000001110111011011100;
assign LUT_3[61219] = 32'b00000000000000010101100110111001;
assign LUT_3[61220] = 32'b00000000000000001010000001101110;
assign LUT_3[61221] = 32'b00000000000000010000101101001011;
assign LUT_3[61222] = 32'b00000000000000001100001001010010;
assign LUT_3[61223] = 32'b00000000000000010010110100101111;
assign LUT_3[61224] = 32'b00000000000000010010001100111110;
assign LUT_3[61225] = 32'b00000000000000011000111000011011;
assign LUT_3[61226] = 32'b00000000000000010100010100100010;
assign LUT_3[61227] = 32'b00000000000000011010111111111111;
assign LUT_3[61228] = 32'b00000000000000001111011010110100;
assign LUT_3[61229] = 32'b00000000000000010110000110010001;
assign LUT_3[61230] = 32'b00000000000000010001100010011000;
assign LUT_3[61231] = 32'b00000000000000011000001101110101;
assign LUT_3[61232] = 32'b00000000000000010000000110111011;
assign LUT_3[61233] = 32'b00000000000000010110110010011000;
assign LUT_3[61234] = 32'b00000000000000010010001110011111;
assign LUT_3[61235] = 32'b00000000000000011000111001111100;
assign LUT_3[61236] = 32'b00000000000000001101010100110001;
assign LUT_3[61237] = 32'b00000000000000010100000000001110;
assign LUT_3[61238] = 32'b00000000000000001111011100010101;
assign LUT_3[61239] = 32'b00000000000000010110000111110010;
assign LUT_3[61240] = 32'b00000000000000010101100000000001;
assign LUT_3[61241] = 32'b00000000000000011100001011011110;
assign LUT_3[61242] = 32'b00000000000000010111100111100101;
assign LUT_3[61243] = 32'b00000000000000011110010011000010;
assign LUT_3[61244] = 32'b00000000000000010010101101110111;
assign LUT_3[61245] = 32'b00000000000000011001011001010100;
assign LUT_3[61246] = 32'b00000000000000010100110101011011;
assign LUT_3[61247] = 32'b00000000000000011011100000111000;
assign LUT_3[61248] = 32'b00000000000000001011011110000011;
assign LUT_3[61249] = 32'b00000000000000010010001001100000;
assign LUT_3[61250] = 32'b00000000000000001101100101100111;
assign LUT_3[61251] = 32'b00000000000000010100010001000100;
assign LUT_3[61252] = 32'b00000000000000001000101011111001;
assign LUT_3[61253] = 32'b00000000000000001111010111010110;
assign LUT_3[61254] = 32'b00000000000000001010110011011101;
assign LUT_3[61255] = 32'b00000000000000010001011110111010;
assign LUT_3[61256] = 32'b00000000000000010000110111001001;
assign LUT_3[61257] = 32'b00000000000000010111100010100110;
assign LUT_3[61258] = 32'b00000000000000010010111110101101;
assign LUT_3[61259] = 32'b00000000000000011001101010001010;
assign LUT_3[61260] = 32'b00000000000000001110000100111111;
assign LUT_3[61261] = 32'b00000000000000010100110000011100;
assign LUT_3[61262] = 32'b00000000000000010000001100100011;
assign LUT_3[61263] = 32'b00000000000000010110111000000000;
assign LUT_3[61264] = 32'b00000000000000001110110001000110;
assign LUT_3[61265] = 32'b00000000000000010101011100100011;
assign LUT_3[61266] = 32'b00000000000000010000111000101010;
assign LUT_3[61267] = 32'b00000000000000010111100100000111;
assign LUT_3[61268] = 32'b00000000000000001011111110111100;
assign LUT_3[61269] = 32'b00000000000000010010101010011001;
assign LUT_3[61270] = 32'b00000000000000001110000110100000;
assign LUT_3[61271] = 32'b00000000000000010100110001111101;
assign LUT_3[61272] = 32'b00000000000000010100001010001100;
assign LUT_3[61273] = 32'b00000000000000011010110101101001;
assign LUT_3[61274] = 32'b00000000000000010110010001110000;
assign LUT_3[61275] = 32'b00000000000000011100111101001101;
assign LUT_3[61276] = 32'b00000000000000010001011000000010;
assign LUT_3[61277] = 32'b00000000000000011000000011011111;
assign LUT_3[61278] = 32'b00000000000000010011011111100110;
assign LUT_3[61279] = 32'b00000000000000011010001011000011;
assign LUT_3[61280] = 32'b00000000000000001100101100100011;
assign LUT_3[61281] = 32'b00000000000000010011011000000000;
assign LUT_3[61282] = 32'b00000000000000001110110100000111;
assign LUT_3[61283] = 32'b00000000000000010101011111100100;
assign LUT_3[61284] = 32'b00000000000000001001111010011001;
assign LUT_3[61285] = 32'b00000000000000010000100101110110;
assign LUT_3[61286] = 32'b00000000000000001100000001111101;
assign LUT_3[61287] = 32'b00000000000000010010101101011010;
assign LUT_3[61288] = 32'b00000000000000010010000101101001;
assign LUT_3[61289] = 32'b00000000000000011000110001000110;
assign LUT_3[61290] = 32'b00000000000000010100001101001101;
assign LUT_3[61291] = 32'b00000000000000011010111000101010;
assign LUT_3[61292] = 32'b00000000000000001111010011011111;
assign LUT_3[61293] = 32'b00000000000000010101111110111100;
assign LUT_3[61294] = 32'b00000000000000010001011011000011;
assign LUT_3[61295] = 32'b00000000000000011000000110100000;
assign LUT_3[61296] = 32'b00000000000000001111111111100110;
assign LUT_3[61297] = 32'b00000000000000010110101011000011;
assign LUT_3[61298] = 32'b00000000000000010010000111001010;
assign LUT_3[61299] = 32'b00000000000000011000110010100111;
assign LUT_3[61300] = 32'b00000000000000001101001101011100;
assign LUT_3[61301] = 32'b00000000000000010011111000111001;
assign LUT_3[61302] = 32'b00000000000000001111010101000000;
assign LUT_3[61303] = 32'b00000000000000010110000000011101;
assign LUT_3[61304] = 32'b00000000000000010101011000101100;
assign LUT_3[61305] = 32'b00000000000000011100000100001001;
assign LUT_3[61306] = 32'b00000000000000010111100000010000;
assign LUT_3[61307] = 32'b00000000000000011110001011101101;
assign LUT_3[61308] = 32'b00000000000000010010100110100010;
assign LUT_3[61309] = 32'b00000000000000011001010001111111;
assign LUT_3[61310] = 32'b00000000000000010100101110000110;
assign LUT_3[61311] = 32'b00000000000000011011011001100011;
assign LUT_3[61312] = 32'b00000000000000001101110000010110;
assign LUT_3[61313] = 32'b00000000000000010100011011110011;
assign LUT_3[61314] = 32'b00000000000000001111110111111010;
assign LUT_3[61315] = 32'b00000000000000010110100011010111;
assign LUT_3[61316] = 32'b00000000000000001010111110001100;
assign LUT_3[61317] = 32'b00000000000000010001101001101001;
assign LUT_3[61318] = 32'b00000000000000001101000101110000;
assign LUT_3[61319] = 32'b00000000000000010011110001001101;
assign LUT_3[61320] = 32'b00000000000000010011001001011100;
assign LUT_3[61321] = 32'b00000000000000011001110100111001;
assign LUT_3[61322] = 32'b00000000000000010101010001000000;
assign LUT_3[61323] = 32'b00000000000000011011111100011101;
assign LUT_3[61324] = 32'b00000000000000010000010111010010;
assign LUT_3[61325] = 32'b00000000000000010111000010101111;
assign LUT_3[61326] = 32'b00000000000000010010011110110110;
assign LUT_3[61327] = 32'b00000000000000011001001010010011;
assign LUT_3[61328] = 32'b00000000000000010001000011011001;
assign LUT_3[61329] = 32'b00000000000000010111101110110110;
assign LUT_3[61330] = 32'b00000000000000010011001010111101;
assign LUT_3[61331] = 32'b00000000000000011001110110011010;
assign LUT_3[61332] = 32'b00000000000000001110010001001111;
assign LUT_3[61333] = 32'b00000000000000010100111100101100;
assign LUT_3[61334] = 32'b00000000000000010000011000110011;
assign LUT_3[61335] = 32'b00000000000000010111000100010000;
assign LUT_3[61336] = 32'b00000000000000010110011100011111;
assign LUT_3[61337] = 32'b00000000000000011101000111111100;
assign LUT_3[61338] = 32'b00000000000000011000100100000011;
assign LUT_3[61339] = 32'b00000000000000011111001111100000;
assign LUT_3[61340] = 32'b00000000000000010011101010010101;
assign LUT_3[61341] = 32'b00000000000000011010010101110010;
assign LUT_3[61342] = 32'b00000000000000010101110001111001;
assign LUT_3[61343] = 32'b00000000000000011100011101010110;
assign LUT_3[61344] = 32'b00000000000000001110111110110110;
assign LUT_3[61345] = 32'b00000000000000010101101010010011;
assign LUT_3[61346] = 32'b00000000000000010001000110011010;
assign LUT_3[61347] = 32'b00000000000000010111110001110111;
assign LUT_3[61348] = 32'b00000000000000001100001100101100;
assign LUT_3[61349] = 32'b00000000000000010010111000001001;
assign LUT_3[61350] = 32'b00000000000000001110010100010000;
assign LUT_3[61351] = 32'b00000000000000010100111111101101;
assign LUT_3[61352] = 32'b00000000000000010100010111111100;
assign LUT_3[61353] = 32'b00000000000000011011000011011001;
assign LUT_3[61354] = 32'b00000000000000010110011111100000;
assign LUT_3[61355] = 32'b00000000000000011101001010111101;
assign LUT_3[61356] = 32'b00000000000000010001100101110010;
assign LUT_3[61357] = 32'b00000000000000011000010001001111;
assign LUT_3[61358] = 32'b00000000000000010011101101010110;
assign LUT_3[61359] = 32'b00000000000000011010011000110011;
assign LUT_3[61360] = 32'b00000000000000010010010001111001;
assign LUT_3[61361] = 32'b00000000000000011000111101010110;
assign LUT_3[61362] = 32'b00000000000000010100011001011101;
assign LUT_3[61363] = 32'b00000000000000011011000100111010;
assign LUT_3[61364] = 32'b00000000000000001111011111101111;
assign LUT_3[61365] = 32'b00000000000000010110001011001100;
assign LUT_3[61366] = 32'b00000000000000010001100111010011;
assign LUT_3[61367] = 32'b00000000000000011000010010110000;
assign LUT_3[61368] = 32'b00000000000000010111101010111111;
assign LUT_3[61369] = 32'b00000000000000011110010110011100;
assign LUT_3[61370] = 32'b00000000000000011001110010100011;
assign LUT_3[61371] = 32'b00000000000000100000011110000000;
assign LUT_3[61372] = 32'b00000000000000010100111000110101;
assign LUT_3[61373] = 32'b00000000000000011011100100010010;
assign LUT_3[61374] = 32'b00000000000000010111000000011001;
assign LUT_3[61375] = 32'b00000000000000011101101011110110;
assign LUT_3[61376] = 32'b00000000000000001101101001000001;
assign LUT_3[61377] = 32'b00000000000000010100010100011110;
assign LUT_3[61378] = 32'b00000000000000001111110000100101;
assign LUT_3[61379] = 32'b00000000000000010110011100000010;
assign LUT_3[61380] = 32'b00000000000000001010110110110111;
assign LUT_3[61381] = 32'b00000000000000010001100010010100;
assign LUT_3[61382] = 32'b00000000000000001100111110011011;
assign LUT_3[61383] = 32'b00000000000000010011101001111000;
assign LUT_3[61384] = 32'b00000000000000010011000010000111;
assign LUT_3[61385] = 32'b00000000000000011001101101100100;
assign LUT_3[61386] = 32'b00000000000000010101001001101011;
assign LUT_3[61387] = 32'b00000000000000011011110101001000;
assign LUT_3[61388] = 32'b00000000000000010000001111111101;
assign LUT_3[61389] = 32'b00000000000000010110111011011010;
assign LUT_3[61390] = 32'b00000000000000010010010111100001;
assign LUT_3[61391] = 32'b00000000000000011001000010111110;
assign LUT_3[61392] = 32'b00000000000000010000111100000100;
assign LUT_3[61393] = 32'b00000000000000010111100111100001;
assign LUT_3[61394] = 32'b00000000000000010011000011101000;
assign LUT_3[61395] = 32'b00000000000000011001101111000101;
assign LUT_3[61396] = 32'b00000000000000001110001001111010;
assign LUT_3[61397] = 32'b00000000000000010100110101010111;
assign LUT_3[61398] = 32'b00000000000000010000010001011110;
assign LUT_3[61399] = 32'b00000000000000010110111100111011;
assign LUT_3[61400] = 32'b00000000000000010110010101001010;
assign LUT_3[61401] = 32'b00000000000000011101000000100111;
assign LUT_3[61402] = 32'b00000000000000011000011100101110;
assign LUT_3[61403] = 32'b00000000000000011111001000001011;
assign LUT_3[61404] = 32'b00000000000000010011100011000000;
assign LUT_3[61405] = 32'b00000000000000011010001110011101;
assign LUT_3[61406] = 32'b00000000000000010101101010100100;
assign LUT_3[61407] = 32'b00000000000000011100010110000001;
assign LUT_3[61408] = 32'b00000000000000001110110111100001;
assign LUT_3[61409] = 32'b00000000000000010101100010111110;
assign LUT_3[61410] = 32'b00000000000000010000111111000101;
assign LUT_3[61411] = 32'b00000000000000010111101010100010;
assign LUT_3[61412] = 32'b00000000000000001100000101010111;
assign LUT_3[61413] = 32'b00000000000000010010110000110100;
assign LUT_3[61414] = 32'b00000000000000001110001100111011;
assign LUT_3[61415] = 32'b00000000000000010100111000011000;
assign LUT_3[61416] = 32'b00000000000000010100010000100111;
assign LUT_3[61417] = 32'b00000000000000011010111100000100;
assign LUT_3[61418] = 32'b00000000000000010110011000001011;
assign LUT_3[61419] = 32'b00000000000000011101000011101000;
assign LUT_3[61420] = 32'b00000000000000010001011110011101;
assign LUT_3[61421] = 32'b00000000000000011000001001111010;
assign LUT_3[61422] = 32'b00000000000000010011100110000001;
assign LUT_3[61423] = 32'b00000000000000011010010001011110;
assign LUT_3[61424] = 32'b00000000000000010010001010100100;
assign LUT_3[61425] = 32'b00000000000000011000110110000001;
assign LUT_3[61426] = 32'b00000000000000010100010010001000;
assign LUT_3[61427] = 32'b00000000000000011010111101100101;
assign LUT_3[61428] = 32'b00000000000000001111011000011010;
assign LUT_3[61429] = 32'b00000000000000010110000011110111;
assign LUT_3[61430] = 32'b00000000000000010001011111111110;
assign LUT_3[61431] = 32'b00000000000000011000001011011011;
assign LUT_3[61432] = 32'b00000000000000010111100011101010;
assign LUT_3[61433] = 32'b00000000000000011110001111000111;
assign LUT_3[61434] = 32'b00000000000000011001101011001110;
assign LUT_3[61435] = 32'b00000000000000100000010110101011;
assign LUT_3[61436] = 32'b00000000000000010100110001100000;
assign LUT_3[61437] = 32'b00000000000000011011011100111101;
assign LUT_3[61438] = 32'b00000000000000010110111001000100;
assign LUT_3[61439] = 32'b00000000000000011101100100100001;
assign LUT_3[61440] = 32'b00000000000000000111110110111011;
assign LUT_3[61441] = 32'b00000000000000001110100010011000;
assign LUT_3[61442] = 32'b00000000000000001001111110011111;
assign LUT_3[61443] = 32'b00000000000000010000101001111100;
assign LUT_3[61444] = 32'b00000000000000000101000100110001;
assign LUT_3[61445] = 32'b00000000000000001011110000001110;
assign LUT_3[61446] = 32'b00000000000000000111001100010101;
assign LUT_3[61447] = 32'b00000000000000001101110111110010;
assign LUT_3[61448] = 32'b00000000000000001101010000000001;
assign LUT_3[61449] = 32'b00000000000000010011111011011110;
assign LUT_3[61450] = 32'b00000000000000001111010111100101;
assign LUT_3[61451] = 32'b00000000000000010110000011000010;
assign LUT_3[61452] = 32'b00000000000000001010011101110111;
assign LUT_3[61453] = 32'b00000000000000010001001001010100;
assign LUT_3[61454] = 32'b00000000000000001100100101011011;
assign LUT_3[61455] = 32'b00000000000000010011010000111000;
assign LUT_3[61456] = 32'b00000000000000001011001001111110;
assign LUT_3[61457] = 32'b00000000000000010001110101011011;
assign LUT_3[61458] = 32'b00000000000000001101010001100010;
assign LUT_3[61459] = 32'b00000000000000010011111100111111;
assign LUT_3[61460] = 32'b00000000000000001000010111110100;
assign LUT_3[61461] = 32'b00000000000000001111000011010001;
assign LUT_3[61462] = 32'b00000000000000001010011111011000;
assign LUT_3[61463] = 32'b00000000000000010001001010110101;
assign LUT_3[61464] = 32'b00000000000000010000100011000100;
assign LUT_3[61465] = 32'b00000000000000010111001110100001;
assign LUT_3[61466] = 32'b00000000000000010010101010101000;
assign LUT_3[61467] = 32'b00000000000000011001010110000101;
assign LUT_3[61468] = 32'b00000000000000001101110000111010;
assign LUT_3[61469] = 32'b00000000000000010100011100010111;
assign LUT_3[61470] = 32'b00000000000000001111111000011110;
assign LUT_3[61471] = 32'b00000000000000010110100011111011;
assign LUT_3[61472] = 32'b00000000000000001001000101011011;
assign LUT_3[61473] = 32'b00000000000000001111110000111000;
assign LUT_3[61474] = 32'b00000000000000001011001100111111;
assign LUT_3[61475] = 32'b00000000000000010001111000011100;
assign LUT_3[61476] = 32'b00000000000000000110010011010001;
assign LUT_3[61477] = 32'b00000000000000001100111110101110;
assign LUT_3[61478] = 32'b00000000000000001000011010110101;
assign LUT_3[61479] = 32'b00000000000000001111000110010010;
assign LUT_3[61480] = 32'b00000000000000001110011110100001;
assign LUT_3[61481] = 32'b00000000000000010101001001111110;
assign LUT_3[61482] = 32'b00000000000000010000100110000101;
assign LUT_3[61483] = 32'b00000000000000010111010001100010;
assign LUT_3[61484] = 32'b00000000000000001011101100010111;
assign LUT_3[61485] = 32'b00000000000000010010010111110100;
assign LUT_3[61486] = 32'b00000000000000001101110011111011;
assign LUT_3[61487] = 32'b00000000000000010100011111011000;
assign LUT_3[61488] = 32'b00000000000000001100011000011110;
assign LUT_3[61489] = 32'b00000000000000010011000011111011;
assign LUT_3[61490] = 32'b00000000000000001110100000000010;
assign LUT_3[61491] = 32'b00000000000000010101001011011111;
assign LUT_3[61492] = 32'b00000000000000001001100110010100;
assign LUT_3[61493] = 32'b00000000000000010000010001110001;
assign LUT_3[61494] = 32'b00000000000000001011101101111000;
assign LUT_3[61495] = 32'b00000000000000010010011001010101;
assign LUT_3[61496] = 32'b00000000000000010001110001100100;
assign LUT_3[61497] = 32'b00000000000000011000011101000001;
assign LUT_3[61498] = 32'b00000000000000010011111001001000;
assign LUT_3[61499] = 32'b00000000000000011010100100100101;
assign LUT_3[61500] = 32'b00000000000000001110111111011010;
assign LUT_3[61501] = 32'b00000000000000010101101010110111;
assign LUT_3[61502] = 32'b00000000000000010001000110111110;
assign LUT_3[61503] = 32'b00000000000000010111110010011011;
assign LUT_3[61504] = 32'b00000000000000000111101111100110;
assign LUT_3[61505] = 32'b00000000000000001110011011000011;
assign LUT_3[61506] = 32'b00000000000000001001110111001010;
assign LUT_3[61507] = 32'b00000000000000010000100010100111;
assign LUT_3[61508] = 32'b00000000000000000100111101011100;
assign LUT_3[61509] = 32'b00000000000000001011101000111001;
assign LUT_3[61510] = 32'b00000000000000000111000101000000;
assign LUT_3[61511] = 32'b00000000000000001101110000011101;
assign LUT_3[61512] = 32'b00000000000000001101001000101100;
assign LUT_3[61513] = 32'b00000000000000010011110100001001;
assign LUT_3[61514] = 32'b00000000000000001111010000010000;
assign LUT_3[61515] = 32'b00000000000000010101111011101101;
assign LUT_3[61516] = 32'b00000000000000001010010110100010;
assign LUT_3[61517] = 32'b00000000000000010001000001111111;
assign LUT_3[61518] = 32'b00000000000000001100011110000110;
assign LUT_3[61519] = 32'b00000000000000010011001001100011;
assign LUT_3[61520] = 32'b00000000000000001011000010101001;
assign LUT_3[61521] = 32'b00000000000000010001101110000110;
assign LUT_3[61522] = 32'b00000000000000001101001010001101;
assign LUT_3[61523] = 32'b00000000000000010011110101101010;
assign LUT_3[61524] = 32'b00000000000000001000010000011111;
assign LUT_3[61525] = 32'b00000000000000001110111011111100;
assign LUT_3[61526] = 32'b00000000000000001010011000000011;
assign LUT_3[61527] = 32'b00000000000000010001000011100000;
assign LUT_3[61528] = 32'b00000000000000010000011011101111;
assign LUT_3[61529] = 32'b00000000000000010111000111001100;
assign LUT_3[61530] = 32'b00000000000000010010100011010011;
assign LUT_3[61531] = 32'b00000000000000011001001110110000;
assign LUT_3[61532] = 32'b00000000000000001101101001100101;
assign LUT_3[61533] = 32'b00000000000000010100010101000010;
assign LUT_3[61534] = 32'b00000000000000001111110001001001;
assign LUT_3[61535] = 32'b00000000000000010110011100100110;
assign LUT_3[61536] = 32'b00000000000000001000111110000110;
assign LUT_3[61537] = 32'b00000000000000001111101001100011;
assign LUT_3[61538] = 32'b00000000000000001011000101101010;
assign LUT_3[61539] = 32'b00000000000000010001110001000111;
assign LUT_3[61540] = 32'b00000000000000000110001011111100;
assign LUT_3[61541] = 32'b00000000000000001100110111011001;
assign LUT_3[61542] = 32'b00000000000000001000010011100000;
assign LUT_3[61543] = 32'b00000000000000001110111110111101;
assign LUT_3[61544] = 32'b00000000000000001110010111001100;
assign LUT_3[61545] = 32'b00000000000000010101000010101001;
assign LUT_3[61546] = 32'b00000000000000010000011110110000;
assign LUT_3[61547] = 32'b00000000000000010111001010001101;
assign LUT_3[61548] = 32'b00000000000000001011100101000010;
assign LUT_3[61549] = 32'b00000000000000010010010000011111;
assign LUT_3[61550] = 32'b00000000000000001101101100100110;
assign LUT_3[61551] = 32'b00000000000000010100011000000011;
assign LUT_3[61552] = 32'b00000000000000001100010001001001;
assign LUT_3[61553] = 32'b00000000000000010010111100100110;
assign LUT_3[61554] = 32'b00000000000000001110011000101101;
assign LUT_3[61555] = 32'b00000000000000010101000100001010;
assign LUT_3[61556] = 32'b00000000000000001001011110111111;
assign LUT_3[61557] = 32'b00000000000000010000001010011100;
assign LUT_3[61558] = 32'b00000000000000001011100110100011;
assign LUT_3[61559] = 32'b00000000000000010010010010000000;
assign LUT_3[61560] = 32'b00000000000000010001101010001111;
assign LUT_3[61561] = 32'b00000000000000011000010101101100;
assign LUT_3[61562] = 32'b00000000000000010011110001110011;
assign LUT_3[61563] = 32'b00000000000000011010011101010000;
assign LUT_3[61564] = 32'b00000000000000001110111000000101;
assign LUT_3[61565] = 32'b00000000000000010101100011100010;
assign LUT_3[61566] = 32'b00000000000000010000111111101001;
assign LUT_3[61567] = 32'b00000000000000010111101011000110;
assign LUT_3[61568] = 32'b00000000000000001010000001111001;
assign LUT_3[61569] = 32'b00000000000000010000101101010110;
assign LUT_3[61570] = 32'b00000000000000001100001001011101;
assign LUT_3[61571] = 32'b00000000000000010010110100111010;
assign LUT_3[61572] = 32'b00000000000000000111001111101111;
assign LUT_3[61573] = 32'b00000000000000001101111011001100;
assign LUT_3[61574] = 32'b00000000000000001001010111010011;
assign LUT_3[61575] = 32'b00000000000000010000000010110000;
assign LUT_3[61576] = 32'b00000000000000001111011010111111;
assign LUT_3[61577] = 32'b00000000000000010110000110011100;
assign LUT_3[61578] = 32'b00000000000000010001100010100011;
assign LUT_3[61579] = 32'b00000000000000011000001110000000;
assign LUT_3[61580] = 32'b00000000000000001100101000110101;
assign LUT_3[61581] = 32'b00000000000000010011010100010010;
assign LUT_3[61582] = 32'b00000000000000001110110000011001;
assign LUT_3[61583] = 32'b00000000000000010101011011110110;
assign LUT_3[61584] = 32'b00000000000000001101010100111100;
assign LUT_3[61585] = 32'b00000000000000010100000000011001;
assign LUT_3[61586] = 32'b00000000000000001111011100100000;
assign LUT_3[61587] = 32'b00000000000000010110000111111101;
assign LUT_3[61588] = 32'b00000000000000001010100010110010;
assign LUT_3[61589] = 32'b00000000000000010001001110001111;
assign LUT_3[61590] = 32'b00000000000000001100101010010110;
assign LUT_3[61591] = 32'b00000000000000010011010101110011;
assign LUT_3[61592] = 32'b00000000000000010010101110000010;
assign LUT_3[61593] = 32'b00000000000000011001011001011111;
assign LUT_3[61594] = 32'b00000000000000010100110101100110;
assign LUT_3[61595] = 32'b00000000000000011011100001000011;
assign LUT_3[61596] = 32'b00000000000000001111111011111000;
assign LUT_3[61597] = 32'b00000000000000010110100111010101;
assign LUT_3[61598] = 32'b00000000000000010010000011011100;
assign LUT_3[61599] = 32'b00000000000000011000101110111001;
assign LUT_3[61600] = 32'b00000000000000001011010000011001;
assign LUT_3[61601] = 32'b00000000000000010001111011110110;
assign LUT_3[61602] = 32'b00000000000000001101010111111101;
assign LUT_3[61603] = 32'b00000000000000010100000011011010;
assign LUT_3[61604] = 32'b00000000000000001000011110001111;
assign LUT_3[61605] = 32'b00000000000000001111001001101100;
assign LUT_3[61606] = 32'b00000000000000001010100101110011;
assign LUT_3[61607] = 32'b00000000000000010001010001010000;
assign LUT_3[61608] = 32'b00000000000000010000101001011111;
assign LUT_3[61609] = 32'b00000000000000010111010100111100;
assign LUT_3[61610] = 32'b00000000000000010010110001000011;
assign LUT_3[61611] = 32'b00000000000000011001011100100000;
assign LUT_3[61612] = 32'b00000000000000001101110111010101;
assign LUT_3[61613] = 32'b00000000000000010100100010110010;
assign LUT_3[61614] = 32'b00000000000000001111111110111001;
assign LUT_3[61615] = 32'b00000000000000010110101010010110;
assign LUT_3[61616] = 32'b00000000000000001110100011011100;
assign LUT_3[61617] = 32'b00000000000000010101001110111001;
assign LUT_3[61618] = 32'b00000000000000010000101011000000;
assign LUT_3[61619] = 32'b00000000000000010111010110011101;
assign LUT_3[61620] = 32'b00000000000000001011110001010010;
assign LUT_3[61621] = 32'b00000000000000010010011100101111;
assign LUT_3[61622] = 32'b00000000000000001101111000110110;
assign LUT_3[61623] = 32'b00000000000000010100100100010011;
assign LUT_3[61624] = 32'b00000000000000010011111100100010;
assign LUT_3[61625] = 32'b00000000000000011010100111111111;
assign LUT_3[61626] = 32'b00000000000000010110000100000110;
assign LUT_3[61627] = 32'b00000000000000011100101111100011;
assign LUT_3[61628] = 32'b00000000000000010001001010011000;
assign LUT_3[61629] = 32'b00000000000000010111110101110101;
assign LUT_3[61630] = 32'b00000000000000010011010001111100;
assign LUT_3[61631] = 32'b00000000000000011001111101011001;
assign LUT_3[61632] = 32'b00000000000000001001111010100100;
assign LUT_3[61633] = 32'b00000000000000010000100110000001;
assign LUT_3[61634] = 32'b00000000000000001100000010001000;
assign LUT_3[61635] = 32'b00000000000000010010101101100101;
assign LUT_3[61636] = 32'b00000000000000000111001000011010;
assign LUT_3[61637] = 32'b00000000000000001101110011110111;
assign LUT_3[61638] = 32'b00000000000000001001001111111110;
assign LUT_3[61639] = 32'b00000000000000001111111011011011;
assign LUT_3[61640] = 32'b00000000000000001111010011101010;
assign LUT_3[61641] = 32'b00000000000000010101111111000111;
assign LUT_3[61642] = 32'b00000000000000010001011011001110;
assign LUT_3[61643] = 32'b00000000000000011000000110101011;
assign LUT_3[61644] = 32'b00000000000000001100100001100000;
assign LUT_3[61645] = 32'b00000000000000010011001100111101;
assign LUT_3[61646] = 32'b00000000000000001110101001000100;
assign LUT_3[61647] = 32'b00000000000000010101010100100001;
assign LUT_3[61648] = 32'b00000000000000001101001101100111;
assign LUT_3[61649] = 32'b00000000000000010011111001000100;
assign LUT_3[61650] = 32'b00000000000000001111010101001011;
assign LUT_3[61651] = 32'b00000000000000010110000000101000;
assign LUT_3[61652] = 32'b00000000000000001010011011011101;
assign LUT_3[61653] = 32'b00000000000000010001000110111010;
assign LUT_3[61654] = 32'b00000000000000001100100011000001;
assign LUT_3[61655] = 32'b00000000000000010011001110011110;
assign LUT_3[61656] = 32'b00000000000000010010100110101101;
assign LUT_3[61657] = 32'b00000000000000011001010010001010;
assign LUT_3[61658] = 32'b00000000000000010100101110010001;
assign LUT_3[61659] = 32'b00000000000000011011011001101110;
assign LUT_3[61660] = 32'b00000000000000001111110100100011;
assign LUT_3[61661] = 32'b00000000000000010110100000000000;
assign LUT_3[61662] = 32'b00000000000000010001111100000111;
assign LUT_3[61663] = 32'b00000000000000011000100111100100;
assign LUT_3[61664] = 32'b00000000000000001011001001000100;
assign LUT_3[61665] = 32'b00000000000000010001110100100001;
assign LUT_3[61666] = 32'b00000000000000001101010000101000;
assign LUT_3[61667] = 32'b00000000000000010011111100000101;
assign LUT_3[61668] = 32'b00000000000000001000010110111010;
assign LUT_3[61669] = 32'b00000000000000001111000010010111;
assign LUT_3[61670] = 32'b00000000000000001010011110011110;
assign LUT_3[61671] = 32'b00000000000000010001001001111011;
assign LUT_3[61672] = 32'b00000000000000010000100010001010;
assign LUT_3[61673] = 32'b00000000000000010111001101100111;
assign LUT_3[61674] = 32'b00000000000000010010101001101110;
assign LUT_3[61675] = 32'b00000000000000011001010101001011;
assign LUT_3[61676] = 32'b00000000000000001101110000000000;
assign LUT_3[61677] = 32'b00000000000000010100011011011101;
assign LUT_3[61678] = 32'b00000000000000001111110111100100;
assign LUT_3[61679] = 32'b00000000000000010110100011000001;
assign LUT_3[61680] = 32'b00000000000000001110011100000111;
assign LUT_3[61681] = 32'b00000000000000010101000111100100;
assign LUT_3[61682] = 32'b00000000000000010000100011101011;
assign LUT_3[61683] = 32'b00000000000000010111001111001000;
assign LUT_3[61684] = 32'b00000000000000001011101001111101;
assign LUT_3[61685] = 32'b00000000000000010010010101011010;
assign LUT_3[61686] = 32'b00000000000000001101110001100001;
assign LUT_3[61687] = 32'b00000000000000010100011100111110;
assign LUT_3[61688] = 32'b00000000000000010011110101001101;
assign LUT_3[61689] = 32'b00000000000000011010100000101010;
assign LUT_3[61690] = 32'b00000000000000010101111100110001;
assign LUT_3[61691] = 32'b00000000000000011100101000001110;
assign LUT_3[61692] = 32'b00000000000000010001000011000011;
assign LUT_3[61693] = 32'b00000000000000010111101110100000;
assign LUT_3[61694] = 32'b00000000000000010011001010100111;
assign LUT_3[61695] = 32'b00000000000000011001110110000100;
assign LUT_3[61696] = 32'b00000000000000000100000110011100;
assign LUT_3[61697] = 32'b00000000000000001010110001111001;
assign LUT_3[61698] = 32'b00000000000000000110001110000000;
assign LUT_3[61699] = 32'b00000000000000001100111001011101;
assign LUT_3[61700] = 32'b00000000000000000001010100010010;
assign LUT_3[61701] = 32'b00000000000000000111111111101111;
assign LUT_3[61702] = 32'b00000000000000000011011011110110;
assign LUT_3[61703] = 32'b00000000000000001010000111010011;
assign LUT_3[61704] = 32'b00000000000000001001011111100010;
assign LUT_3[61705] = 32'b00000000000000010000001010111111;
assign LUT_3[61706] = 32'b00000000000000001011100111000110;
assign LUT_3[61707] = 32'b00000000000000010010010010100011;
assign LUT_3[61708] = 32'b00000000000000000110101101011000;
assign LUT_3[61709] = 32'b00000000000000001101011000110101;
assign LUT_3[61710] = 32'b00000000000000001000110100111100;
assign LUT_3[61711] = 32'b00000000000000001111100000011001;
assign LUT_3[61712] = 32'b00000000000000000111011001011111;
assign LUT_3[61713] = 32'b00000000000000001110000100111100;
assign LUT_3[61714] = 32'b00000000000000001001100001000011;
assign LUT_3[61715] = 32'b00000000000000010000001100100000;
assign LUT_3[61716] = 32'b00000000000000000100100111010101;
assign LUT_3[61717] = 32'b00000000000000001011010010110010;
assign LUT_3[61718] = 32'b00000000000000000110101110111001;
assign LUT_3[61719] = 32'b00000000000000001101011010010110;
assign LUT_3[61720] = 32'b00000000000000001100110010100101;
assign LUT_3[61721] = 32'b00000000000000010011011110000010;
assign LUT_3[61722] = 32'b00000000000000001110111010001001;
assign LUT_3[61723] = 32'b00000000000000010101100101100110;
assign LUT_3[61724] = 32'b00000000000000001010000000011011;
assign LUT_3[61725] = 32'b00000000000000010000101011111000;
assign LUT_3[61726] = 32'b00000000000000001100000111111111;
assign LUT_3[61727] = 32'b00000000000000010010110011011100;
assign LUT_3[61728] = 32'b00000000000000000101010100111100;
assign LUT_3[61729] = 32'b00000000000000001100000000011001;
assign LUT_3[61730] = 32'b00000000000000000111011100100000;
assign LUT_3[61731] = 32'b00000000000000001110000111111101;
assign LUT_3[61732] = 32'b00000000000000000010100010110010;
assign LUT_3[61733] = 32'b00000000000000001001001110001111;
assign LUT_3[61734] = 32'b00000000000000000100101010010110;
assign LUT_3[61735] = 32'b00000000000000001011010101110011;
assign LUT_3[61736] = 32'b00000000000000001010101110000010;
assign LUT_3[61737] = 32'b00000000000000010001011001011111;
assign LUT_3[61738] = 32'b00000000000000001100110101100110;
assign LUT_3[61739] = 32'b00000000000000010011100001000011;
assign LUT_3[61740] = 32'b00000000000000000111111011111000;
assign LUT_3[61741] = 32'b00000000000000001110100111010101;
assign LUT_3[61742] = 32'b00000000000000001010000011011100;
assign LUT_3[61743] = 32'b00000000000000010000101110111001;
assign LUT_3[61744] = 32'b00000000000000001000100111111111;
assign LUT_3[61745] = 32'b00000000000000001111010011011100;
assign LUT_3[61746] = 32'b00000000000000001010101111100011;
assign LUT_3[61747] = 32'b00000000000000010001011011000000;
assign LUT_3[61748] = 32'b00000000000000000101110101110101;
assign LUT_3[61749] = 32'b00000000000000001100100001010010;
assign LUT_3[61750] = 32'b00000000000000000111111101011001;
assign LUT_3[61751] = 32'b00000000000000001110101000110110;
assign LUT_3[61752] = 32'b00000000000000001110000001000101;
assign LUT_3[61753] = 32'b00000000000000010100101100100010;
assign LUT_3[61754] = 32'b00000000000000010000001000101001;
assign LUT_3[61755] = 32'b00000000000000010110110100000110;
assign LUT_3[61756] = 32'b00000000000000001011001110111011;
assign LUT_3[61757] = 32'b00000000000000010001111010011000;
assign LUT_3[61758] = 32'b00000000000000001101010110011111;
assign LUT_3[61759] = 32'b00000000000000010100000001111100;
assign LUT_3[61760] = 32'b00000000000000000011111111000111;
assign LUT_3[61761] = 32'b00000000000000001010101010100100;
assign LUT_3[61762] = 32'b00000000000000000110000110101011;
assign LUT_3[61763] = 32'b00000000000000001100110010001000;
assign LUT_3[61764] = 32'b00000000000000000001001100111101;
assign LUT_3[61765] = 32'b00000000000000000111111000011010;
assign LUT_3[61766] = 32'b00000000000000000011010100100001;
assign LUT_3[61767] = 32'b00000000000000001001111111111110;
assign LUT_3[61768] = 32'b00000000000000001001011000001101;
assign LUT_3[61769] = 32'b00000000000000010000000011101010;
assign LUT_3[61770] = 32'b00000000000000001011011111110001;
assign LUT_3[61771] = 32'b00000000000000010010001011001110;
assign LUT_3[61772] = 32'b00000000000000000110100110000011;
assign LUT_3[61773] = 32'b00000000000000001101010001100000;
assign LUT_3[61774] = 32'b00000000000000001000101101100111;
assign LUT_3[61775] = 32'b00000000000000001111011001000100;
assign LUT_3[61776] = 32'b00000000000000000111010010001010;
assign LUT_3[61777] = 32'b00000000000000001101111101100111;
assign LUT_3[61778] = 32'b00000000000000001001011001101110;
assign LUT_3[61779] = 32'b00000000000000010000000101001011;
assign LUT_3[61780] = 32'b00000000000000000100100000000000;
assign LUT_3[61781] = 32'b00000000000000001011001011011101;
assign LUT_3[61782] = 32'b00000000000000000110100111100100;
assign LUT_3[61783] = 32'b00000000000000001101010011000001;
assign LUT_3[61784] = 32'b00000000000000001100101011010000;
assign LUT_3[61785] = 32'b00000000000000010011010110101101;
assign LUT_3[61786] = 32'b00000000000000001110110010110100;
assign LUT_3[61787] = 32'b00000000000000010101011110010001;
assign LUT_3[61788] = 32'b00000000000000001001111001000110;
assign LUT_3[61789] = 32'b00000000000000010000100100100011;
assign LUT_3[61790] = 32'b00000000000000001100000000101010;
assign LUT_3[61791] = 32'b00000000000000010010101100000111;
assign LUT_3[61792] = 32'b00000000000000000101001101100111;
assign LUT_3[61793] = 32'b00000000000000001011111001000100;
assign LUT_3[61794] = 32'b00000000000000000111010101001011;
assign LUT_3[61795] = 32'b00000000000000001110000000101000;
assign LUT_3[61796] = 32'b00000000000000000010011011011101;
assign LUT_3[61797] = 32'b00000000000000001001000110111010;
assign LUT_3[61798] = 32'b00000000000000000100100011000001;
assign LUT_3[61799] = 32'b00000000000000001011001110011110;
assign LUT_3[61800] = 32'b00000000000000001010100110101101;
assign LUT_3[61801] = 32'b00000000000000010001010010001010;
assign LUT_3[61802] = 32'b00000000000000001100101110010001;
assign LUT_3[61803] = 32'b00000000000000010011011001101110;
assign LUT_3[61804] = 32'b00000000000000000111110100100011;
assign LUT_3[61805] = 32'b00000000000000001110100000000000;
assign LUT_3[61806] = 32'b00000000000000001001111100000111;
assign LUT_3[61807] = 32'b00000000000000010000100111100100;
assign LUT_3[61808] = 32'b00000000000000001000100000101010;
assign LUT_3[61809] = 32'b00000000000000001111001100000111;
assign LUT_3[61810] = 32'b00000000000000001010101000001110;
assign LUT_3[61811] = 32'b00000000000000010001010011101011;
assign LUT_3[61812] = 32'b00000000000000000101101110100000;
assign LUT_3[61813] = 32'b00000000000000001100011001111101;
assign LUT_3[61814] = 32'b00000000000000000111110110000100;
assign LUT_3[61815] = 32'b00000000000000001110100001100001;
assign LUT_3[61816] = 32'b00000000000000001101111001110000;
assign LUT_3[61817] = 32'b00000000000000010100100101001101;
assign LUT_3[61818] = 32'b00000000000000010000000001010100;
assign LUT_3[61819] = 32'b00000000000000010110101100110001;
assign LUT_3[61820] = 32'b00000000000000001011000111100110;
assign LUT_3[61821] = 32'b00000000000000010001110011000011;
assign LUT_3[61822] = 32'b00000000000000001101001111001010;
assign LUT_3[61823] = 32'b00000000000000010011111010100111;
assign LUT_3[61824] = 32'b00000000000000000110010001011010;
assign LUT_3[61825] = 32'b00000000000000001100111100110111;
assign LUT_3[61826] = 32'b00000000000000001000011000111110;
assign LUT_3[61827] = 32'b00000000000000001111000100011011;
assign LUT_3[61828] = 32'b00000000000000000011011111010000;
assign LUT_3[61829] = 32'b00000000000000001010001010101101;
assign LUT_3[61830] = 32'b00000000000000000101100110110100;
assign LUT_3[61831] = 32'b00000000000000001100010010010001;
assign LUT_3[61832] = 32'b00000000000000001011101010100000;
assign LUT_3[61833] = 32'b00000000000000010010010101111101;
assign LUT_3[61834] = 32'b00000000000000001101110010000100;
assign LUT_3[61835] = 32'b00000000000000010100011101100001;
assign LUT_3[61836] = 32'b00000000000000001000111000010110;
assign LUT_3[61837] = 32'b00000000000000001111100011110011;
assign LUT_3[61838] = 32'b00000000000000001010111111111010;
assign LUT_3[61839] = 32'b00000000000000010001101011010111;
assign LUT_3[61840] = 32'b00000000000000001001100100011101;
assign LUT_3[61841] = 32'b00000000000000010000001111111010;
assign LUT_3[61842] = 32'b00000000000000001011101100000001;
assign LUT_3[61843] = 32'b00000000000000010010010111011110;
assign LUT_3[61844] = 32'b00000000000000000110110010010011;
assign LUT_3[61845] = 32'b00000000000000001101011101110000;
assign LUT_3[61846] = 32'b00000000000000001000111001110111;
assign LUT_3[61847] = 32'b00000000000000001111100101010100;
assign LUT_3[61848] = 32'b00000000000000001110111101100011;
assign LUT_3[61849] = 32'b00000000000000010101101001000000;
assign LUT_3[61850] = 32'b00000000000000010001000101000111;
assign LUT_3[61851] = 32'b00000000000000010111110000100100;
assign LUT_3[61852] = 32'b00000000000000001100001011011001;
assign LUT_3[61853] = 32'b00000000000000010010110110110110;
assign LUT_3[61854] = 32'b00000000000000001110010010111101;
assign LUT_3[61855] = 32'b00000000000000010100111110011010;
assign LUT_3[61856] = 32'b00000000000000000111011111111010;
assign LUT_3[61857] = 32'b00000000000000001110001011010111;
assign LUT_3[61858] = 32'b00000000000000001001100111011110;
assign LUT_3[61859] = 32'b00000000000000010000010010111011;
assign LUT_3[61860] = 32'b00000000000000000100101101110000;
assign LUT_3[61861] = 32'b00000000000000001011011001001101;
assign LUT_3[61862] = 32'b00000000000000000110110101010100;
assign LUT_3[61863] = 32'b00000000000000001101100000110001;
assign LUT_3[61864] = 32'b00000000000000001100111001000000;
assign LUT_3[61865] = 32'b00000000000000010011100100011101;
assign LUT_3[61866] = 32'b00000000000000001111000000100100;
assign LUT_3[61867] = 32'b00000000000000010101101100000001;
assign LUT_3[61868] = 32'b00000000000000001010000110110110;
assign LUT_3[61869] = 32'b00000000000000010000110010010011;
assign LUT_3[61870] = 32'b00000000000000001100001110011010;
assign LUT_3[61871] = 32'b00000000000000010010111001110111;
assign LUT_3[61872] = 32'b00000000000000001010110010111101;
assign LUT_3[61873] = 32'b00000000000000010001011110011010;
assign LUT_3[61874] = 32'b00000000000000001100111010100001;
assign LUT_3[61875] = 32'b00000000000000010011100101111110;
assign LUT_3[61876] = 32'b00000000000000001000000000110011;
assign LUT_3[61877] = 32'b00000000000000001110101100010000;
assign LUT_3[61878] = 32'b00000000000000001010001000010111;
assign LUT_3[61879] = 32'b00000000000000010000110011110100;
assign LUT_3[61880] = 32'b00000000000000010000001100000011;
assign LUT_3[61881] = 32'b00000000000000010110110111100000;
assign LUT_3[61882] = 32'b00000000000000010010010011100111;
assign LUT_3[61883] = 32'b00000000000000011000111111000100;
assign LUT_3[61884] = 32'b00000000000000001101011001111001;
assign LUT_3[61885] = 32'b00000000000000010100000101010110;
assign LUT_3[61886] = 32'b00000000000000001111100001011101;
assign LUT_3[61887] = 32'b00000000000000010110001100111010;
assign LUT_3[61888] = 32'b00000000000000000110001010000101;
assign LUT_3[61889] = 32'b00000000000000001100110101100010;
assign LUT_3[61890] = 32'b00000000000000001000010001101001;
assign LUT_3[61891] = 32'b00000000000000001110111101000110;
assign LUT_3[61892] = 32'b00000000000000000011010111111011;
assign LUT_3[61893] = 32'b00000000000000001010000011011000;
assign LUT_3[61894] = 32'b00000000000000000101011111011111;
assign LUT_3[61895] = 32'b00000000000000001100001010111100;
assign LUT_3[61896] = 32'b00000000000000001011100011001011;
assign LUT_3[61897] = 32'b00000000000000010010001110101000;
assign LUT_3[61898] = 32'b00000000000000001101101010101111;
assign LUT_3[61899] = 32'b00000000000000010100010110001100;
assign LUT_3[61900] = 32'b00000000000000001000110001000001;
assign LUT_3[61901] = 32'b00000000000000001111011100011110;
assign LUT_3[61902] = 32'b00000000000000001010111000100101;
assign LUT_3[61903] = 32'b00000000000000010001100100000010;
assign LUT_3[61904] = 32'b00000000000000001001011101001000;
assign LUT_3[61905] = 32'b00000000000000010000001000100101;
assign LUT_3[61906] = 32'b00000000000000001011100100101100;
assign LUT_3[61907] = 32'b00000000000000010010010000001001;
assign LUT_3[61908] = 32'b00000000000000000110101010111110;
assign LUT_3[61909] = 32'b00000000000000001101010110011011;
assign LUT_3[61910] = 32'b00000000000000001000110010100010;
assign LUT_3[61911] = 32'b00000000000000001111011101111111;
assign LUT_3[61912] = 32'b00000000000000001110110110001110;
assign LUT_3[61913] = 32'b00000000000000010101100001101011;
assign LUT_3[61914] = 32'b00000000000000010000111101110010;
assign LUT_3[61915] = 32'b00000000000000010111101001001111;
assign LUT_3[61916] = 32'b00000000000000001100000100000100;
assign LUT_3[61917] = 32'b00000000000000010010101111100001;
assign LUT_3[61918] = 32'b00000000000000001110001011101000;
assign LUT_3[61919] = 32'b00000000000000010100110111000101;
assign LUT_3[61920] = 32'b00000000000000000111011000100101;
assign LUT_3[61921] = 32'b00000000000000001110000100000010;
assign LUT_3[61922] = 32'b00000000000000001001100000001001;
assign LUT_3[61923] = 32'b00000000000000010000001011100110;
assign LUT_3[61924] = 32'b00000000000000000100100110011011;
assign LUT_3[61925] = 32'b00000000000000001011010001111000;
assign LUT_3[61926] = 32'b00000000000000000110101101111111;
assign LUT_3[61927] = 32'b00000000000000001101011001011100;
assign LUT_3[61928] = 32'b00000000000000001100110001101011;
assign LUT_3[61929] = 32'b00000000000000010011011101001000;
assign LUT_3[61930] = 32'b00000000000000001110111001001111;
assign LUT_3[61931] = 32'b00000000000000010101100100101100;
assign LUT_3[61932] = 32'b00000000000000001001111111100001;
assign LUT_3[61933] = 32'b00000000000000010000101010111110;
assign LUT_3[61934] = 32'b00000000000000001100000111000101;
assign LUT_3[61935] = 32'b00000000000000010010110010100010;
assign LUT_3[61936] = 32'b00000000000000001010101011101000;
assign LUT_3[61937] = 32'b00000000000000010001010111000101;
assign LUT_3[61938] = 32'b00000000000000001100110011001100;
assign LUT_3[61939] = 32'b00000000000000010011011110101001;
assign LUT_3[61940] = 32'b00000000000000000111111001011110;
assign LUT_3[61941] = 32'b00000000000000001110100100111011;
assign LUT_3[61942] = 32'b00000000000000001010000001000010;
assign LUT_3[61943] = 32'b00000000000000010000101100011111;
assign LUT_3[61944] = 32'b00000000000000010000000100101110;
assign LUT_3[61945] = 32'b00000000000000010110110000001011;
assign LUT_3[61946] = 32'b00000000000000010010001100010010;
assign LUT_3[61947] = 32'b00000000000000011000110111101111;
assign LUT_3[61948] = 32'b00000000000000001101010010100100;
assign LUT_3[61949] = 32'b00000000000000010011111110000001;
assign LUT_3[61950] = 32'b00000000000000001111011010001000;
assign LUT_3[61951] = 32'b00000000000000010110000101100101;
assign LUT_3[61952] = 32'b00000000000000001011001100000111;
assign LUT_3[61953] = 32'b00000000000000010001110111100100;
assign LUT_3[61954] = 32'b00000000000000001101010011101011;
assign LUT_3[61955] = 32'b00000000000000010011111111001000;
assign LUT_3[61956] = 32'b00000000000000001000011001111101;
assign LUT_3[61957] = 32'b00000000000000001111000101011010;
assign LUT_3[61958] = 32'b00000000000000001010100001100001;
assign LUT_3[61959] = 32'b00000000000000010001001100111110;
assign LUT_3[61960] = 32'b00000000000000010000100101001101;
assign LUT_3[61961] = 32'b00000000000000010111010000101010;
assign LUT_3[61962] = 32'b00000000000000010010101100110001;
assign LUT_3[61963] = 32'b00000000000000011001011000001110;
assign LUT_3[61964] = 32'b00000000000000001101110011000011;
assign LUT_3[61965] = 32'b00000000000000010100011110100000;
assign LUT_3[61966] = 32'b00000000000000001111111010100111;
assign LUT_3[61967] = 32'b00000000000000010110100110000100;
assign LUT_3[61968] = 32'b00000000000000001110011111001010;
assign LUT_3[61969] = 32'b00000000000000010101001010100111;
assign LUT_3[61970] = 32'b00000000000000010000100110101110;
assign LUT_3[61971] = 32'b00000000000000010111010010001011;
assign LUT_3[61972] = 32'b00000000000000001011101101000000;
assign LUT_3[61973] = 32'b00000000000000010010011000011101;
assign LUT_3[61974] = 32'b00000000000000001101110100100100;
assign LUT_3[61975] = 32'b00000000000000010100100000000001;
assign LUT_3[61976] = 32'b00000000000000010011111000010000;
assign LUT_3[61977] = 32'b00000000000000011010100011101101;
assign LUT_3[61978] = 32'b00000000000000010101111111110100;
assign LUT_3[61979] = 32'b00000000000000011100101011010001;
assign LUT_3[61980] = 32'b00000000000000010001000110000110;
assign LUT_3[61981] = 32'b00000000000000010111110001100011;
assign LUT_3[61982] = 32'b00000000000000010011001101101010;
assign LUT_3[61983] = 32'b00000000000000011001111001000111;
assign LUT_3[61984] = 32'b00000000000000001100011010100111;
assign LUT_3[61985] = 32'b00000000000000010011000110000100;
assign LUT_3[61986] = 32'b00000000000000001110100010001011;
assign LUT_3[61987] = 32'b00000000000000010101001101101000;
assign LUT_3[61988] = 32'b00000000000000001001101000011101;
assign LUT_3[61989] = 32'b00000000000000010000010011111010;
assign LUT_3[61990] = 32'b00000000000000001011110000000001;
assign LUT_3[61991] = 32'b00000000000000010010011011011110;
assign LUT_3[61992] = 32'b00000000000000010001110011101101;
assign LUT_3[61993] = 32'b00000000000000011000011111001010;
assign LUT_3[61994] = 32'b00000000000000010011111011010001;
assign LUT_3[61995] = 32'b00000000000000011010100110101110;
assign LUT_3[61996] = 32'b00000000000000001111000001100011;
assign LUT_3[61997] = 32'b00000000000000010101101101000000;
assign LUT_3[61998] = 32'b00000000000000010001001001000111;
assign LUT_3[61999] = 32'b00000000000000010111110100100100;
assign LUT_3[62000] = 32'b00000000000000001111101101101010;
assign LUT_3[62001] = 32'b00000000000000010110011001000111;
assign LUT_3[62002] = 32'b00000000000000010001110101001110;
assign LUT_3[62003] = 32'b00000000000000011000100000101011;
assign LUT_3[62004] = 32'b00000000000000001100111011100000;
assign LUT_3[62005] = 32'b00000000000000010011100110111101;
assign LUT_3[62006] = 32'b00000000000000001111000011000100;
assign LUT_3[62007] = 32'b00000000000000010101101110100001;
assign LUT_3[62008] = 32'b00000000000000010101000110110000;
assign LUT_3[62009] = 32'b00000000000000011011110010001101;
assign LUT_3[62010] = 32'b00000000000000010111001110010100;
assign LUT_3[62011] = 32'b00000000000000011101111001110001;
assign LUT_3[62012] = 32'b00000000000000010010010100100110;
assign LUT_3[62013] = 32'b00000000000000011001000000000011;
assign LUT_3[62014] = 32'b00000000000000010100011100001010;
assign LUT_3[62015] = 32'b00000000000000011011000111100111;
assign LUT_3[62016] = 32'b00000000000000001011000100110010;
assign LUT_3[62017] = 32'b00000000000000010001110000001111;
assign LUT_3[62018] = 32'b00000000000000001101001100010110;
assign LUT_3[62019] = 32'b00000000000000010011110111110011;
assign LUT_3[62020] = 32'b00000000000000001000010010101000;
assign LUT_3[62021] = 32'b00000000000000001110111110000101;
assign LUT_3[62022] = 32'b00000000000000001010011010001100;
assign LUT_3[62023] = 32'b00000000000000010001000101101001;
assign LUT_3[62024] = 32'b00000000000000010000011101111000;
assign LUT_3[62025] = 32'b00000000000000010111001001010101;
assign LUT_3[62026] = 32'b00000000000000010010100101011100;
assign LUT_3[62027] = 32'b00000000000000011001010000111001;
assign LUT_3[62028] = 32'b00000000000000001101101011101110;
assign LUT_3[62029] = 32'b00000000000000010100010111001011;
assign LUT_3[62030] = 32'b00000000000000001111110011010010;
assign LUT_3[62031] = 32'b00000000000000010110011110101111;
assign LUT_3[62032] = 32'b00000000000000001110010111110101;
assign LUT_3[62033] = 32'b00000000000000010101000011010010;
assign LUT_3[62034] = 32'b00000000000000010000011111011001;
assign LUT_3[62035] = 32'b00000000000000010111001010110110;
assign LUT_3[62036] = 32'b00000000000000001011100101101011;
assign LUT_3[62037] = 32'b00000000000000010010010001001000;
assign LUT_3[62038] = 32'b00000000000000001101101101001111;
assign LUT_3[62039] = 32'b00000000000000010100011000101100;
assign LUT_3[62040] = 32'b00000000000000010011110000111011;
assign LUT_3[62041] = 32'b00000000000000011010011100011000;
assign LUT_3[62042] = 32'b00000000000000010101111000011111;
assign LUT_3[62043] = 32'b00000000000000011100100011111100;
assign LUT_3[62044] = 32'b00000000000000010000111110110001;
assign LUT_3[62045] = 32'b00000000000000010111101010001110;
assign LUT_3[62046] = 32'b00000000000000010011000110010101;
assign LUT_3[62047] = 32'b00000000000000011001110001110010;
assign LUT_3[62048] = 32'b00000000000000001100010011010010;
assign LUT_3[62049] = 32'b00000000000000010010111110101111;
assign LUT_3[62050] = 32'b00000000000000001110011010110110;
assign LUT_3[62051] = 32'b00000000000000010101000110010011;
assign LUT_3[62052] = 32'b00000000000000001001100001001000;
assign LUT_3[62053] = 32'b00000000000000010000001100100101;
assign LUT_3[62054] = 32'b00000000000000001011101000101100;
assign LUT_3[62055] = 32'b00000000000000010010010100001001;
assign LUT_3[62056] = 32'b00000000000000010001101100011000;
assign LUT_3[62057] = 32'b00000000000000011000010111110101;
assign LUT_3[62058] = 32'b00000000000000010011110011111100;
assign LUT_3[62059] = 32'b00000000000000011010011111011001;
assign LUT_3[62060] = 32'b00000000000000001110111010001110;
assign LUT_3[62061] = 32'b00000000000000010101100101101011;
assign LUT_3[62062] = 32'b00000000000000010001000001110010;
assign LUT_3[62063] = 32'b00000000000000010111101101001111;
assign LUT_3[62064] = 32'b00000000000000001111100110010101;
assign LUT_3[62065] = 32'b00000000000000010110010001110010;
assign LUT_3[62066] = 32'b00000000000000010001101101111001;
assign LUT_3[62067] = 32'b00000000000000011000011001010110;
assign LUT_3[62068] = 32'b00000000000000001100110100001011;
assign LUT_3[62069] = 32'b00000000000000010011011111101000;
assign LUT_3[62070] = 32'b00000000000000001110111011101111;
assign LUT_3[62071] = 32'b00000000000000010101100111001100;
assign LUT_3[62072] = 32'b00000000000000010100111111011011;
assign LUT_3[62073] = 32'b00000000000000011011101010111000;
assign LUT_3[62074] = 32'b00000000000000010111000110111111;
assign LUT_3[62075] = 32'b00000000000000011101110010011100;
assign LUT_3[62076] = 32'b00000000000000010010001101010001;
assign LUT_3[62077] = 32'b00000000000000011000111000101110;
assign LUT_3[62078] = 32'b00000000000000010100010100110101;
assign LUT_3[62079] = 32'b00000000000000011011000000010010;
assign LUT_3[62080] = 32'b00000000000000001101010111000101;
assign LUT_3[62081] = 32'b00000000000000010100000010100010;
assign LUT_3[62082] = 32'b00000000000000001111011110101001;
assign LUT_3[62083] = 32'b00000000000000010110001010000110;
assign LUT_3[62084] = 32'b00000000000000001010100100111011;
assign LUT_3[62085] = 32'b00000000000000010001010000011000;
assign LUT_3[62086] = 32'b00000000000000001100101100011111;
assign LUT_3[62087] = 32'b00000000000000010011010111111100;
assign LUT_3[62088] = 32'b00000000000000010010110000001011;
assign LUT_3[62089] = 32'b00000000000000011001011011101000;
assign LUT_3[62090] = 32'b00000000000000010100110111101111;
assign LUT_3[62091] = 32'b00000000000000011011100011001100;
assign LUT_3[62092] = 32'b00000000000000001111111110000001;
assign LUT_3[62093] = 32'b00000000000000010110101001011110;
assign LUT_3[62094] = 32'b00000000000000010010000101100101;
assign LUT_3[62095] = 32'b00000000000000011000110001000010;
assign LUT_3[62096] = 32'b00000000000000010000101010001000;
assign LUT_3[62097] = 32'b00000000000000010111010101100101;
assign LUT_3[62098] = 32'b00000000000000010010110001101100;
assign LUT_3[62099] = 32'b00000000000000011001011101001001;
assign LUT_3[62100] = 32'b00000000000000001101110111111110;
assign LUT_3[62101] = 32'b00000000000000010100100011011011;
assign LUT_3[62102] = 32'b00000000000000001111111111100010;
assign LUT_3[62103] = 32'b00000000000000010110101010111111;
assign LUT_3[62104] = 32'b00000000000000010110000011001110;
assign LUT_3[62105] = 32'b00000000000000011100101110101011;
assign LUT_3[62106] = 32'b00000000000000011000001010110010;
assign LUT_3[62107] = 32'b00000000000000011110110110001111;
assign LUT_3[62108] = 32'b00000000000000010011010001000100;
assign LUT_3[62109] = 32'b00000000000000011001111100100001;
assign LUT_3[62110] = 32'b00000000000000010101011000101000;
assign LUT_3[62111] = 32'b00000000000000011100000100000101;
assign LUT_3[62112] = 32'b00000000000000001110100101100101;
assign LUT_3[62113] = 32'b00000000000000010101010001000010;
assign LUT_3[62114] = 32'b00000000000000010000101101001001;
assign LUT_3[62115] = 32'b00000000000000010111011000100110;
assign LUT_3[62116] = 32'b00000000000000001011110011011011;
assign LUT_3[62117] = 32'b00000000000000010010011110111000;
assign LUT_3[62118] = 32'b00000000000000001101111010111111;
assign LUT_3[62119] = 32'b00000000000000010100100110011100;
assign LUT_3[62120] = 32'b00000000000000010011111110101011;
assign LUT_3[62121] = 32'b00000000000000011010101010001000;
assign LUT_3[62122] = 32'b00000000000000010110000110001111;
assign LUT_3[62123] = 32'b00000000000000011100110001101100;
assign LUT_3[62124] = 32'b00000000000000010001001100100001;
assign LUT_3[62125] = 32'b00000000000000010111110111111110;
assign LUT_3[62126] = 32'b00000000000000010011010100000101;
assign LUT_3[62127] = 32'b00000000000000011001111111100010;
assign LUT_3[62128] = 32'b00000000000000010001111000101000;
assign LUT_3[62129] = 32'b00000000000000011000100100000101;
assign LUT_3[62130] = 32'b00000000000000010100000000001100;
assign LUT_3[62131] = 32'b00000000000000011010101011101001;
assign LUT_3[62132] = 32'b00000000000000001111000110011110;
assign LUT_3[62133] = 32'b00000000000000010101110001111011;
assign LUT_3[62134] = 32'b00000000000000010001001110000010;
assign LUT_3[62135] = 32'b00000000000000010111111001011111;
assign LUT_3[62136] = 32'b00000000000000010111010001101110;
assign LUT_3[62137] = 32'b00000000000000011101111101001011;
assign LUT_3[62138] = 32'b00000000000000011001011001010010;
assign LUT_3[62139] = 32'b00000000000000100000000100101111;
assign LUT_3[62140] = 32'b00000000000000010100011111100100;
assign LUT_3[62141] = 32'b00000000000000011011001011000001;
assign LUT_3[62142] = 32'b00000000000000010110100111001000;
assign LUT_3[62143] = 32'b00000000000000011101010010100101;
assign LUT_3[62144] = 32'b00000000000000001101001111110000;
assign LUT_3[62145] = 32'b00000000000000010011111011001101;
assign LUT_3[62146] = 32'b00000000000000001111010111010100;
assign LUT_3[62147] = 32'b00000000000000010110000010110001;
assign LUT_3[62148] = 32'b00000000000000001010011101100110;
assign LUT_3[62149] = 32'b00000000000000010001001001000011;
assign LUT_3[62150] = 32'b00000000000000001100100101001010;
assign LUT_3[62151] = 32'b00000000000000010011010000100111;
assign LUT_3[62152] = 32'b00000000000000010010101000110110;
assign LUT_3[62153] = 32'b00000000000000011001010100010011;
assign LUT_3[62154] = 32'b00000000000000010100110000011010;
assign LUT_3[62155] = 32'b00000000000000011011011011110111;
assign LUT_3[62156] = 32'b00000000000000001111110110101100;
assign LUT_3[62157] = 32'b00000000000000010110100010001001;
assign LUT_3[62158] = 32'b00000000000000010001111110010000;
assign LUT_3[62159] = 32'b00000000000000011000101001101101;
assign LUT_3[62160] = 32'b00000000000000010000100010110011;
assign LUT_3[62161] = 32'b00000000000000010111001110010000;
assign LUT_3[62162] = 32'b00000000000000010010101010010111;
assign LUT_3[62163] = 32'b00000000000000011001010101110100;
assign LUT_3[62164] = 32'b00000000000000001101110000101001;
assign LUT_3[62165] = 32'b00000000000000010100011100000110;
assign LUT_3[62166] = 32'b00000000000000001111111000001101;
assign LUT_3[62167] = 32'b00000000000000010110100011101010;
assign LUT_3[62168] = 32'b00000000000000010101111011111001;
assign LUT_3[62169] = 32'b00000000000000011100100111010110;
assign LUT_3[62170] = 32'b00000000000000011000000011011101;
assign LUT_3[62171] = 32'b00000000000000011110101110111010;
assign LUT_3[62172] = 32'b00000000000000010011001001101111;
assign LUT_3[62173] = 32'b00000000000000011001110101001100;
assign LUT_3[62174] = 32'b00000000000000010101010001010011;
assign LUT_3[62175] = 32'b00000000000000011011111100110000;
assign LUT_3[62176] = 32'b00000000000000001110011110010000;
assign LUT_3[62177] = 32'b00000000000000010101001001101101;
assign LUT_3[62178] = 32'b00000000000000010000100101110100;
assign LUT_3[62179] = 32'b00000000000000010111010001010001;
assign LUT_3[62180] = 32'b00000000000000001011101100000110;
assign LUT_3[62181] = 32'b00000000000000010010010111100011;
assign LUT_3[62182] = 32'b00000000000000001101110011101010;
assign LUT_3[62183] = 32'b00000000000000010100011111000111;
assign LUT_3[62184] = 32'b00000000000000010011110111010110;
assign LUT_3[62185] = 32'b00000000000000011010100010110011;
assign LUT_3[62186] = 32'b00000000000000010101111110111010;
assign LUT_3[62187] = 32'b00000000000000011100101010010111;
assign LUT_3[62188] = 32'b00000000000000010001000101001100;
assign LUT_3[62189] = 32'b00000000000000010111110000101001;
assign LUT_3[62190] = 32'b00000000000000010011001100110000;
assign LUT_3[62191] = 32'b00000000000000011001111000001101;
assign LUT_3[62192] = 32'b00000000000000010001110001010011;
assign LUT_3[62193] = 32'b00000000000000011000011100110000;
assign LUT_3[62194] = 32'b00000000000000010011111000110111;
assign LUT_3[62195] = 32'b00000000000000011010100100010100;
assign LUT_3[62196] = 32'b00000000000000001110111111001001;
assign LUT_3[62197] = 32'b00000000000000010101101010100110;
assign LUT_3[62198] = 32'b00000000000000010001000110101101;
assign LUT_3[62199] = 32'b00000000000000010111110010001010;
assign LUT_3[62200] = 32'b00000000000000010111001010011001;
assign LUT_3[62201] = 32'b00000000000000011101110101110110;
assign LUT_3[62202] = 32'b00000000000000011001010001111101;
assign LUT_3[62203] = 32'b00000000000000011111111101011010;
assign LUT_3[62204] = 32'b00000000000000010100011000001111;
assign LUT_3[62205] = 32'b00000000000000011011000011101100;
assign LUT_3[62206] = 32'b00000000000000010110011111110011;
assign LUT_3[62207] = 32'b00000000000000011101001011010000;
assign LUT_3[62208] = 32'b00000000000000000111011011101000;
assign LUT_3[62209] = 32'b00000000000000001110000111000101;
assign LUT_3[62210] = 32'b00000000000000001001100011001100;
assign LUT_3[62211] = 32'b00000000000000010000001110101001;
assign LUT_3[62212] = 32'b00000000000000000100101001011110;
assign LUT_3[62213] = 32'b00000000000000001011010100111011;
assign LUT_3[62214] = 32'b00000000000000000110110001000010;
assign LUT_3[62215] = 32'b00000000000000001101011100011111;
assign LUT_3[62216] = 32'b00000000000000001100110100101110;
assign LUT_3[62217] = 32'b00000000000000010011100000001011;
assign LUT_3[62218] = 32'b00000000000000001110111100010010;
assign LUT_3[62219] = 32'b00000000000000010101100111101111;
assign LUT_3[62220] = 32'b00000000000000001010000010100100;
assign LUT_3[62221] = 32'b00000000000000010000101110000001;
assign LUT_3[62222] = 32'b00000000000000001100001010001000;
assign LUT_3[62223] = 32'b00000000000000010010110101100101;
assign LUT_3[62224] = 32'b00000000000000001010101110101011;
assign LUT_3[62225] = 32'b00000000000000010001011010001000;
assign LUT_3[62226] = 32'b00000000000000001100110110001111;
assign LUT_3[62227] = 32'b00000000000000010011100001101100;
assign LUT_3[62228] = 32'b00000000000000000111111100100001;
assign LUT_3[62229] = 32'b00000000000000001110100111111110;
assign LUT_3[62230] = 32'b00000000000000001010000100000101;
assign LUT_3[62231] = 32'b00000000000000010000101111100010;
assign LUT_3[62232] = 32'b00000000000000010000000111110001;
assign LUT_3[62233] = 32'b00000000000000010110110011001110;
assign LUT_3[62234] = 32'b00000000000000010010001111010101;
assign LUT_3[62235] = 32'b00000000000000011000111010110010;
assign LUT_3[62236] = 32'b00000000000000001101010101100111;
assign LUT_3[62237] = 32'b00000000000000010100000001000100;
assign LUT_3[62238] = 32'b00000000000000001111011101001011;
assign LUT_3[62239] = 32'b00000000000000010110001000101000;
assign LUT_3[62240] = 32'b00000000000000001000101010001000;
assign LUT_3[62241] = 32'b00000000000000001111010101100101;
assign LUT_3[62242] = 32'b00000000000000001010110001101100;
assign LUT_3[62243] = 32'b00000000000000010001011101001001;
assign LUT_3[62244] = 32'b00000000000000000101110111111110;
assign LUT_3[62245] = 32'b00000000000000001100100011011011;
assign LUT_3[62246] = 32'b00000000000000000111111111100010;
assign LUT_3[62247] = 32'b00000000000000001110101010111111;
assign LUT_3[62248] = 32'b00000000000000001110000011001110;
assign LUT_3[62249] = 32'b00000000000000010100101110101011;
assign LUT_3[62250] = 32'b00000000000000010000001010110010;
assign LUT_3[62251] = 32'b00000000000000010110110110001111;
assign LUT_3[62252] = 32'b00000000000000001011010001000100;
assign LUT_3[62253] = 32'b00000000000000010001111100100001;
assign LUT_3[62254] = 32'b00000000000000001101011000101000;
assign LUT_3[62255] = 32'b00000000000000010100000100000101;
assign LUT_3[62256] = 32'b00000000000000001011111101001011;
assign LUT_3[62257] = 32'b00000000000000010010101000101000;
assign LUT_3[62258] = 32'b00000000000000001110000100101111;
assign LUT_3[62259] = 32'b00000000000000010100110000001100;
assign LUT_3[62260] = 32'b00000000000000001001001011000001;
assign LUT_3[62261] = 32'b00000000000000001111110110011110;
assign LUT_3[62262] = 32'b00000000000000001011010010100101;
assign LUT_3[62263] = 32'b00000000000000010001111110000010;
assign LUT_3[62264] = 32'b00000000000000010001010110010001;
assign LUT_3[62265] = 32'b00000000000000011000000001101110;
assign LUT_3[62266] = 32'b00000000000000010011011101110101;
assign LUT_3[62267] = 32'b00000000000000011010001001010010;
assign LUT_3[62268] = 32'b00000000000000001110100100000111;
assign LUT_3[62269] = 32'b00000000000000010101001111100100;
assign LUT_3[62270] = 32'b00000000000000010000101011101011;
assign LUT_3[62271] = 32'b00000000000000010111010111001000;
assign LUT_3[62272] = 32'b00000000000000000111010100010011;
assign LUT_3[62273] = 32'b00000000000000001101111111110000;
assign LUT_3[62274] = 32'b00000000000000001001011011110111;
assign LUT_3[62275] = 32'b00000000000000010000000111010100;
assign LUT_3[62276] = 32'b00000000000000000100100010001001;
assign LUT_3[62277] = 32'b00000000000000001011001101100110;
assign LUT_3[62278] = 32'b00000000000000000110101001101101;
assign LUT_3[62279] = 32'b00000000000000001101010101001010;
assign LUT_3[62280] = 32'b00000000000000001100101101011001;
assign LUT_3[62281] = 32'b00000000000000010011011000110110;
assign LUT_3[62282] = 32'b00000000000000001110110100111101;
assign LUT_3[62283] = 32'b00000000000000010101100000011010;
assign LUT_3[62284] = 32'b00000000000000001001111011001111;
assign LUT_3[62285] = 32'b00000000000000010000100110101100;
assign LUT_3[62286] = 32'b00000000000000001100000010110011;
assign LUT_3[62287] = 32'b00000000000000010010101110010000;
assign LUT_3[62288] = 32'b00000000000000001010100111010110;
assign LUT_3[62289] = 32'b00000000000000010001010010110011;
assign LUT_3[62290] = 32'b00000000000000001100101110111010;
assign LUT_3[62291] = 32'b00000000000000010011011010010111;
assign LUT_3[62292] = 32'b00000000000000000111110101001100;
assign LUT_3[62293] = 32'b00000000000000001110100000101001;
assign LUT_3[62294] = 32'b00000000000000001001111100110000;
assign LUT_3[62295] = 32'b00000000000000010000101000001101;
assign LUT_3[62296] = 32'b00000000000000010000000000011100;
assign LUT_3[62297] = 32'b00000000000000010110101011111001;
assign LUT_3[62298] = 32'b00000000000000010010001000000000;
assign LUT_3[62299] = 32'b00000000000000011000110011011101;
assign LUT_3[62300] = 32'b00000000000000001101001110010010;
assign LUT_3[62301] = 32'b00000000000000010011111001101111;
assign LUT_3[62302] = 32'b00000000000000001111010101110110;
assign LUT_3[62303] = 32'b00000000000000010110000001010011;
assign LUT_3[62304] = 32'b00000000000000001000100010110011;
assign LUT_3[62305] = 32'b00000000000000001111001110010000;
assign LUT_3[62306] = 32'b00000000000000001010101010010111;
assign LUT_3[62307] = 32'b00000000000000010001010101110100;
assign LUT_3[62308] = 32'b00000000000000000101110000101001;
assign LUT_3[62309] = 32'b00000000000000001100011100000110;
assign LUT_3[62310] = 32'b00000000000000000111111000001101;
assign LUT_3[62311] = 32'b00000000000000001110100011101010;
assign LUT_3[62312] = 32'b00000000000000001101111011111001;
assign LUT_3[62313] = 32'b00000000000000010100100111010110;
assign LUT_3[62314] = 32'b00000000000000010000000011011101;
assign LUT_3[62315] = 32'b00000000000000010110101110111010;
assign LUT_3[62316] = 32'b00000000000000001011001001101111;
assign LUT_3[62317] = 32'b00000000000000010001110101001100;
assign LUT_3[62318] = 32'b00000000000000001101010001010011;
assign LUT_3[62319] = 32'b00000000000000010011111100110000;
assign LUT_3[62320] = 32'b00000000000000001011110101110110;
assign LUT_3[62321] = 32'b00000000000000010010100001010011;
assign LUT_3[62322] = 32'b00000000000000001101111101011010;
assign LUT_3[62323] = 32'b00000000000000010100101000110111;
assign LUT_3[62324] = 32'b00000000000000001001000011101100;
assign LUT_3[62325] = 32'b00000000000000001111101111001001;
assign LUT_3[62326] = 32'b00000000000000001011001011010000;
assign LUT_3[62327] = 32'b00000000000000010001110110101101;
assign LUT_3[62328] = 32'b00000000000000010001001110111100;
assign LUT_3[62329] = 32'b00000000000000010111111010011001;
assign LUT_3[62330] = 32'b00000000000000010011010110100000;
assign LUT_3[62331] = 32'b00000000000000011010000001111101;
assign LUT_3[62332] = 32'b00000000000000001110011100110010;
assign LUT_3[62333] = 32'b00000000000000010101001000001111;
assign LUT_3[62334] = 32'b00000000000000010000100100010110;
assign LUT_3[62335] = 32'b00000000000000010111001111110011;
assign LUT_3[62336] = 32'b00000000000000001001100110100110;
assign LUT_3[62337] = 32'b00000000000000010000010010000011;
assign LUT_3[62338] = 32'b00000000000000001011101110001010;
assign LUT_3[62339] = 32'b00000000000000010010011001100111;
assign LUT_3[62340] = 32'b00000000000000000110110100011100;
assign LUT_3[62341] = 32'b00000000000000001101011111111001;
assign LUT_3[62342] = 32'b00000000000000001000111100000000;
assign LUT_3[62343] = 32'b00000000000000001111100111011101;
assign LUT_3[62344] = 32'b00000000000000001110111111101100;
assign LUT_3[62345] = 32'b00000000000000010101101011001001;
assign LUT_3[62346] = 32'b00000000000000010001000111010000;
assign LUT_3[62347] = 32'b00000000000000010111110010101101;
assign LUT_3[62348] = 32'b00000000000000001100001101100010;
assign LUT_3[62349] = 32'b00000000000000010010111000111111;
assign LUT_3[62350] = 32'b00000000000000001110010101000110;
assign LUT_3[62351] = 32'b00000000000000010101000000100011;
assign LUT_3[62352] = 32'b00000000000000001100111001101001;
assign LUT_3[62353] = 32'b00000000000000010011100101000110;
assign LUT_3[62354] = 32'b00000000000000001111000001001101;
assign LUT_3[62355] = 32'b00000000000000010101101100101010;
assign LUT_3[62356] = 32'b00000000000000001010000111011111;
assign LUT_3[62357] = 32'b00000000000000010000110010111100;
assign LUT_3[62358] = 32'b00000000000000001100001111000011;
assign LUT_3[62359] = 32'b00000000000000010010111010100000;
assign LUT_3[62360] = 32'b00000000000000010010010010101111;
assign LUT_3[62361] = 32'b00000000000000011000111110001100;
assign LUT_3[62362] = 32'b00000000000000010100011010010011;
assign LUT_3[62363] = 32'b00000000000000011011000101110000;
assign LUT_3[62364] = 32'b00000000000000001111100000100101;
assign LUT_3[62365] = 32'b00000000000000010110001100000010;
assign LUT_3[62366] = 32'b00000000000000010001101000001001;
assign LUT_3[62367] = 32'b00000000000000011000010011100110;
assign LUT_3[62368] = 32'b00000000000000001010110101000110;
assign LUT_3[62369] = 32'b00000000000000010001100000100011;
assign LUT_3[62370] = 32'b00000000000000001100111100101010;
assign LUT_3[62371] = 32'b00000000000000010011101000000111;
assign LUT_3[62372] = 32'b00000000000000001000000010111100;
assign LUT_3[62373] = 32'b00000000000000001110101110011001;
assign LUT_3[62374] = 32'b00000000000000001010001010100000;
assign LUT_3[62375] = 32'b00000000000000010000110101111101;
assign LUT_3[62376] = 32'b00000000000000010000001110001100;
assign LUT_3[62377] = 32'b00000000000000010110111001101001;
assign LUT_3[62378] = 32'b00000000000000010010010101110000;
assign LUT_3[62379] = 32'b00000000000000011001000001001101;
assign LUT_3[62380] = 32'b00000000000000001101011100000010;
assign LUT_3[62381] = 32'b00000000000000010100000111011111;
assign LUT_3[62382] = 32'b00000000000000001111100011100110;
assign LUT_3[62383] = 32'b00000000000000010110001111000011;
assign LUT_3[62384] = 32'b00000000000000001110001000001001;
assign LUT_3[62385] = 32'b00000000000000010100110011100110;
assign LUT_3[62386] = 32'b00000000000000010000001111101101;
assign LUT_3[62387] = 32'b00000000000000010110111011001010;
assign LUT_3[62388] = 32'b00000000000000001011010101111111;
assign LUT_3[62389] = 32'b00000000000000010010000001011100;
assign LUT_3[62390] = 32'b00000000000000001101011101100011;
assign LUT_3[62391] = 32'b00000000000000010100001001000000;
assign LUT_3[62392] = 32'b00000000000000010011100001001111;
assign LUT_3[62393] = 32'b00000000000000011010001100101100;
assign LUT_3[62394] = 32'b00000000000000010101101000110011;
assign LUT_3[62395] = 32'b00000000000000011100010100010000;
assign LUT_3[62396] = 32'b00000000000000010000101111000101;
assign LUT_3[62397] = 32'b00000000000000010111011010100010;
assign LUT_3[62398] = 32'b00000000000000010010110110101001;
assign LUT_3[62399] = 32'b00000000000000011001100010000110;
assign LUT_3[62400] = 32'b00000000000000001001011111010001;
assign LUT_3[62401] = 32'b00000000000000010000001010101110;
assign LUT_3[62402] = 32'b00000000000000001011100110110101;
assign LUT_3[62403] = 32'b00000000000000010010010010010010;
assign LUT_3[62404] = 32'b00000000000000000110101101000111;
assign LUT_3[62405] = 32'b00000000000000001101011000100100;
assign LUT_3[62406] = 32'b00000000000000001000110100101011;
assign LUT_3[62407] = 32'b00000000000000001111100000001000;
assign LUT_3[62408] = 32'b00000000000000001110111000010111;
assign LUT_3[62409] = 32'b00000000000000010101100011110100;
assign LUT_3[62410] = 32'b00000000000000010000111111111011;
assign LUT_3[62411] = 32'b00000000000000010111101011011000;
assign LUT_3[62412] = 32'b00000000000000001100000110001101;
assign LUT_3[62413] = 32'b00000000000000010010110001101010;
assign LUT_3[62414] = 32'b00000000000000001110001101110001;
assign LUT_3[62415] = 32'b00000000000000010100111001001110;
assign LUT_3[62416] = 32'b00000000000000001100110010010100;
assign LUT_3[62417] = 32'b00000000000000010011011101110001;
assign LUT_3[62418] = 32'b00000000000000001110111001111000;
assign LUT_3[62419] = 32'b00000000000000010101100101010101;
assign LUT_3[62420] = 32'b00000000000000001010000000001010;
assign LUT_3[62421] = 32'b00000000000000010000101011100111;
assign LUT_3[62422] = 32'b00000000000000001100000111101110;
assign LUT_3[62423] = 32'b00000000000000010010110011001011;
assign LUT_3[62424] = 32'b00000000000000010010001011011010;
assign LUT_3[62425] = 32'b00000000000000011000110110110111;
assign LUT_3[62426] = 32'b00000000000000010100010010111110;
assign LUT_3[62427] = 32'b00000000000000011010111110011011;
assign LUT_3[62428] = 32'b00000000000000001111011001010000;
assign LUT_3[62429] = 32'b00000000000000010110000100101101;
assign LUT_3[62430] = 32'b00000000000000010001100000110100;
assign LUT_3[62431] = 32'b00000000000000011000001100010001;
assign LUT_3[62432] = 32'b00000000000000001010101101110001;
assign LUT_3[62433] = 32'b00000000000000010001011001001110;
assign LUT_3[62434] = 32'b00000000000000001100110101010101;
assign LUT_3[62435] = 32'b00000000000000010011100000110010;
assign LUT_3[62436] = 32'b00000000000000000111111011100111;
assign LUT_3[62437] = 32'b00000000000000001110100111000100;
assign LUT_3[62438] = 32'b00000000000000001010000011001011;
assign LUT_3[62439] = 32'b00000000000000010000101110101000;
assign LUT_3[62440] = 32'b00000000000000010000000110110111;
assign LUT_3[62441] = 32'b00000000000000010110110010010100;
assign LUT_3[62442] = 32'b00000000000000010010001110011011;
assign LUT_3[62443] = 32'b00000000000000011000111001111000;
assign LUT_3[62444] = 32'b00000000000000001101010100101101;
assign LUT_3[62445] = 32'b00000000000000010100000000001010;
assign LUT_3[62446] = 32'b00000000000000001111011100010001;
assign LUT_3[62447] = 32'b00000000000000010110000111101110;
assign LUT_3[62448] = 32'b00000000000000001110000000110100;
assign LUT_3[62449] = 32'b00000000000000010100101100010001;
assign LUT_3[62450] = 32'b00000000000000010000001000011000;
assign LUT_3[62451] = 32'b00000000000000010110110011110101;
assign LUT_3[62452] = 32'b00000000000000001011001110101010;
assign LUT_3[62453] = 32'b00000000000000010001111010000111;
assign LUT_3[62454] = 32'b00000000000000001101010110001110;
assign LUT_3[62455] = 32'b00000000000000010100000001101011;
assign LUT_3[62456] = 32'b00000000000000010011011001111010;
assign LUT_3[62457] = 32'b00000000000000011010000101010111;
assign LUT_3[62458] = 32'b00000000000000010101100001011110;
assign LUT_3[62459] = 32'b00000000000000011100001100111011;
assign LUT_3[62460] = 32'b00000000000000010000100111110000;
assign LUT_3[62461] = 32'b00000000000000010111010011001101;
assign LUT_3[62462] = 32'b00000000000000010010101111010100;
assign LUT_3[62463] = 32'b00000000000000011001011010110001;
assign LUT_3[62464] = 32'b00000000000000001110011011111000;
assign LUT_3[62465] = 32'b00000000000000010101000111010101;
assign LUT_3[62466] = 32'b00000000000000010000100011011100;
assign LUT_3[62467] = 32'b00000000000000010111001110111001;
assign LUT_3[62468] = 32'b00000000000000001011101001101110;
assign LUT_3[62469] = 32'b00000000000000010010010101001011;
assign LUT_3[62470] = 32'b00000000000000001101110001010010;
assign LUT_3[62471] = 32'b00000000000000010100011100101111;
assign LUT_3[62472] = 32'b00000000000000010011110100111110;
assign LUT_3[62473] = 32'b00000000000000011010100000011011;
assign LUT_3[62474] = 32'b00000000000000010101111100100010;
assign LUT_3[62475] = 32'b00000000000000011100100111111111;
assign LUT_3[62476] = 32'b00000000000000010001000010110100;
assign LUT_3[62477] = 32'b00000000000000010111101110010001;
assign LUT_3[62478] = 32'b00000000000000010011001010011000;
assign LUT_3[62479] = 32'b00000000000000011001110101110101;
assign LUT_3[62480] = 32'b00000000000000010001101110111011;
assign LUT_3[62481] = 32'b00000000000000011000011010011000;
assign LUT_3[62482] = 32'b00000000000000010011110110011111;
assign LUT_3[62483] = 32'b00000000000000011010100001111100;
assign LUT_3[62484] = 32'b00000000000000001110111100110001;
assign LUT_3[62485] = 32'b00000000000000010101101000001110;
assign LUT_3[62486] = 32'b00000000000000010001000100010101;
assign LUT_3[62487] = 32'b00000000000000010111101111110010;
assign LUT_3[62488] = 32'b00000000000000010111001000000001;
assign LUT_3[62489] = 32'b00000000000000011101110011011110;
assign LUT_3[62490] = 32'b00000000000000011001001111100101;
assign LUT_3[62491] = 32'b00000000000000011111111011000010;
assign LUT_3[62492] = 32'b00000000000000010100010101110111;
assign LUT_3[62493] = 32'b00000000000000011011000001010100;
assign LUT_3[62494] = 32'b00000000000000010110011101011011;
assign LUT_3[62495] = 32'b00000000000000011101001000111000;
assign LUT_3[62496] = 32'b00000000000000001111101010011000;
assign LUT_3[62497] = 32'b00000000000000010110010101110101;
assign LUT_3[62498] = 32'b00000000000000010001110001111100;
assign LUT_3[62499] = 32'b00000000000000011000011101011001;
assign LUT_3[62500] = 32'b00000000000000001100111000001110;
assign LUT_3[62501] = 32'b00000000000000010011100011101011;
assign LUT_3[62502] = 32'b00000000000000001110111111110010;
assign LUT_3[62503] = 32'b00000000000000010101101011001111;
assign LUT_3[62504] = 32'b00000000000000010101000011011110;
assign LUT_3[62505] = 32'b00000000000000011011101110111011;
assign LUT_3[62506] = 32'b00000000000000010111001011000010;
assign LUT_3[62507] = 32'b00000000000000011101110110011111;
assign LUT_3[62508] = 32'b00000000000000010010010001010100;
assign LUT_3[62509] = 32'b00000000000000011000111100110001;
assign LUT_3[62510] = 32'b00000000000000010100011000111000;
assign LUT_3[62511] = 32'b00000000000000011011000100010101;
assign LUT_3[62512] = 32'b00000000000000010010111101011011;
assign LUT_3[62513] = 32'b00000000000000011001101000111000;
assign LUT_3[62514] = 32'b00000000000000010101000100111111;
assign LUT_3[62515] = 32'b00000000000000011011110000011100;
assign LUT_3[62516] = 32'b00000000000000010000001011010001;
assign LUT_3[62517] = 32'b00000000000000010110110110101110;
assign LUT_3[62518] = 32'b00000000000000010010010010110101;
assign LUT_3[62519] = 32'b00000000000000011000111110010010;
assign LUT_3[62520] = 32'b00000000000000011000010110100001;
assign LUT_3[62521] = 32'b00000000000000011111000001111110;
assign LUT_3[62522] = 32'b00000000000000011010011110000101;
assign LUT_3[62523] = 32'b00000000000000100001001001100010;
assign LUT_3[62524] = 32'b00000000000000010101100100010111;
assign LUT_3[62525] = 32'b00000000000000011100001111110100;
assign LUT_3[62526] = 32'b00000000000000010111101011111011;
assign LUT_3[62527] = 32'b00000000000000011110010111011000;
assign LUT_3[62528] = 32'b00000000000000001110010100100011;
assign LUT_3[62529] = 32'b00000000000000010101000000000000;
assign LUT_3[62530] = 32'b00000000000000010000011100000111;
assign LUT_3[62531] = 32'b00000000000000010111000111100100;
assign LUT_3[62532] = 32'b00000000000000001011100010011001;
assign LUT_3[62533] = 32'b00000000000000010010001101110110;
assign LUT_3[62534] = 32'b00000000000000001101101001111101;
assign LUT_3[62535] = 32'b00000000000000010100010101011010;
assign LUT_3[62536] = 32'b00000000000000010011101101101001;
assign LUT_3[62537] = 32'b00000000000000011010011001000110;
assign LUT_3[62538] = 32'b00000000000000010101110101001101;
assign LUT_3[62539] = 32'b00000000000000011100100000101010;
assign LUT_3[62540] = 32'b00000000000000010000111011011111;
assign LUT_3[62541] = 32'b00000000000000010111100110111100;
assign LUT_3[62542] = 32'b00000000000000010011000011000011;
assign LUT_3[62543] = 32'b00000000000000011001101110100000;
assign LUT_3[62544] = 32'b00000000000000010001100111100110;
assign LUT_3[62545] = 32'b00000000000000011000010011000011;
assign LUT_3[62546] = 32'b00000000000000010011101111001010;
assign LUT_3[62547] = 32'b00000000000000011010011010100111;
assign LUT_3[62548] = 32'b00000000000000001110110101011100;
assign LUT_3[62549] = 32'b00000000000000010101100000111001;
assign LUT_3[62550] = 32'b00000000000000010000111101000000;
assign LUT_3[62551] = 32'b00000000000000010111101000011101;
assign LUT_3[62552] = 32'b00000000000000010111000000101100;
assign LUT_3[62553] = 32'b00000000000000011101101100001001;
assign LUT_3[62554] = 32'b00000000000000011001001000010000;
assign LUT_3[62555] = 32'b00000000000000011111110011101101;
assign LUT_3[62556] = 32'b00000000000000010100001110100010;
assign LUT_3[62557] = 32'b00000000000000011010111001111111;
assign LUT_3[62558] = 32'b00000000000000010110010110000110;
assign LUT_3[62559] = 32'b00000000000000011101000001100011;
assign LUT_3[62560] = 32'b00000000000000001111100011000011;
assign LUT_3[62561] = 32'b00000000000000010110001110100000;
assign LUT_3[62562] = 32'b00000000000000010001101010100111;
assign LUT_3[62563] = 32'b00000000000000011000010110000100;
assign LUT_3[62564] = 32'b00000000000000001100110000111001;
assign LUT_3[62565] = 32'b00000000000000010011011100010110;
assign LUT_3[62566] = 32'b00000000000000001110111000011101;
assign LUT_3[62567] = 32'b00000000000000010101100011111010;
assign LUT_3[62568] = 32'b00000000000000010100111100001001;
assign LUT_3[62569] = 32'b00000000000000011011100111100110;
assign LUT_3[62570] = 32'b00000000000000010111000011101101;
assign LUT_3[62571] = 32'b00000000000000011101101111001010;
assign LUT_3[62572] = 32'b00000000000000010010001001111111;
assign LUT_3[62573] = 32'b00000000000000011000110101011100;
assign LUT_3[62574] = 32'b00000000000000010100010001100011;
assign LUT_3[62575] = 32'b00000000000000011010111101000000;
assign LUT_3[62576] = 32'b00000000000000010010110110000110;
assign LUT_3[62577] = 32'b00000000000000011001100001100011;
assign LUT_3[62578] = 32'b00000000000000010100111101101010;
assign LUT_3[62579] = 32'b00000000000000011011101001000111;
assign LUT_3[62580] = 32'b00000000000000010000000011111100;
assign LUT_3[62581] = 32'b00000000000000010110101111011001;
assign LUT_3[62582] = 32'b00000000000000010010001011100000;
assign LUT_3[62583] = 32'b00000000000000011000110110111101;
assign LUT_3[62584] = 32'b00000000000000011000001111001100;
assign LUT_3[62585] = 32'b00000000000000011110111010101001;
assign LUT_3[62586] = 32'b00000000000000011010010110110000;
assign LUT_3[62587] = 32'b00000000000000100001000010001101;
assign LUT_3[62588] = 32'b00000000000000010101011101000010;
assign LUT_3[62589] = 32'b00000000000000011100001000011111;
assign LUT_3[62590] = 32'b00000000000000010111100100100110;
assign LUT_3[62591] = 32'b00000000000000011110010000000011;
assign LUT_3[62592] = 32'b00000000000000010000100110110110;
assign LUT_3[62593] = 32'b00000000000000010111010010010011;
assign LUT_3[62594] = 32'b00000000000000010010101110011010;
assign LUT_3[62595] = 32'b00000000000000011001011001110111;
assign LUT_3[62596] = 32'b00000000000000001101110100101100;
assign LUT_3[62597] = 32'b00000000000000010100100000001001;
assign LUT_3[62598] = 32'b00000000000000001111111100010000;
assign LUT_3[62599] = 32'b00000000000000010110100111101101;
assign LUT_3[62600] = 32'b00000000000000010101111111111100;
assign LUT_3[62601] = 32'b00000000000000011100101011011001;
assign LUT_3[62602] = 32'b00000000000000011000000111100000;
assign LUT_3[62603] = 32'b00000000000000011110110010111101;
assign LUT_3[62604] = 32'b00000000000000010011001101110010;
assign LUT_3[62605] = 32'b00000000000000011001111001001111;
assign LUT_3[62606] = 32'b00000000000000010101010101010110;
assign LUT_3[62607] = 32'b00000000000000011100000000110011;
assign LUT_3[62608] = 32'b00000000000000010011111001111001;
assign LUT_3[62609] = 32'b00000000000000011010100101010110;
assign LUT_3[62610] = 32'b00000000000000010110000001011101;
assign LUT_3[62611] = 32'b00000000000000011100101100111010;
assign LUT_3[62612] = 32'b00000000000000010001000111101111;
assign LUT_3[62613] = 32'b00000000000000010111110011001100;
assign LUT_3[62614] = 32'b00000000000000010011001111010011;
assign LUT_3[62615] = 32'b00000000000000011001111010110000;
assign LUT_3[62616] = 32'b00000000000000011001010010111111;
assign LUT_3[62617] = 32'b00000000000000011111111110011100;
assign LUT_3[62618] = 32'b00000000000000011011011010100011;
assign LUT_3[62619] = 32'b00000000000000100010000110000000;
assign LUT_3[62620] = 32'b00000000000000010110100000110101;
assign LUT_3[62621] = 32'b00000000000000011101001100010010;
assign LUT_3[62622] = 32'b00000000000000011000101000011001;
assign LUT_3[62623] = 32'b00000000000000011111010011110110;
assign LUT_3[62624] = 32'b00000000000000010001110101010110;
assign LUT_3[62625] = 32'b00000000000000011000100000110011;
assign LUT_3[62626] = 32'b00000000000000010011111100111010;
assign LUT_3[62627] = 32'b00000000000000011010101000010111;
assign LUT_3[62628] = 32'b00000000000000001111000011001100;
assign LUT_3[62629] = 32'b00000000000000010101101110101001;
assign LUT_3[62630] = 32'b00000000000000010001001010110000;
assign LUT_3[62631] = 32'b00000000000000010111110110001101;
assign LUT_3[62632] = 32'b00000000000000010111001110011100;
assign LUT_3[62633] = 32'b00000000000000011101111001111001;
assign LUT_3[62634] = 32'b00000000000000011001010110000000;
assign LUT_3[62635] = 32'b00000000000000100000000001011101;
assign LUT_3[62636] = 32'b00000000000000010100011100010010;
assign LUT_3[62637] = 32'b00000000000000011011000111101111;
assign LUT_3[62638] = 32'b00000000000000010110100011110110;
assign LUT_3[62639] = 32'b00000000000000011101001111010011;
assign LUT_3[62640] = 32'b00000000000000010101001000011001;
assign LUT_3[62641] = 32'b00000000000000011011110011110110;
assign LUT_3[62642] = 32'b00000000000000010111001111111101;
assign LUT_3[62643] = 32'b00000000000000011101111011011010;
assign LUT_3[62644] = 32'b00000000000000010010010110001111;
assign LUT_3[62645] = 32'b00000000000000011001000001101100;
assign LUT_3[62646] = 32'b00000000000000010100011101110011;
assign LUT_3[62647] = 32'b00000000000000011011001001010000;
assign LUT_3[62648] = 32'b00000000000000011010100001011111;
assign LUT_3[62649] = 32'b00000000000000100001001100111100;
assign LUT_3[62650] = 32'b00000000000000011100101001000011;
assign LUT_3[62651] = 32'b00000000000000100011010100100000;
assign LUT_3[62652] = 32'b00000000000000010111101111010101;
assign LUT_3[62653] = 32'b00000000000000011110011010110010;
assign LUT_3[62654] = 32'b00000000000000011001110110111001;
assign LUT_3[62655] = 32'b00000000000000100000100010010110;
assign LUT_3[62656] = 32'b00000000000000010000011111100001;
assign LUT_3[62657] = 32'b00000000000000010111001010111110;
assign LUT_3[62658] = 32'b00000000000000010010100111000101;
assign LUT_3[62659] = 32'b00000000000000011001010010100010;
assign LUT_3[62660] = 32'b00000000000000001101101101010111;
assign LUT_3[62661] = 32'b00000000000000010100011000110100;
assign LUT_3[62662] = 32'b00000000000000001111110100111011;
assign LUT_3[62663] = 32'b00000000000000010110100000011000;
assign LUT_3[62664] = 32'b00000000000000010101111000100111;
assign LUT_3[62665] = 32'b00000000000000011100100100000100;
assign LUT_3[62666] = 32'b00000000000000011000000000001011;
assign LUT_3[62667] = 32'b00000000000000011110101011101000;
assign LUT_3[62668] = 32'b00000000000000010011000110011101;
assign LUT_3[62669] = 32'b00000000000000011001110001111010;
assign LUT_3[62670] = 32'b00000000000000010101001110000001;
assign LUT_3[62671] = 32'b00000000000000011011111001011110;
assign LUT_3[62672] = 32'b00000000000000010011110010100100;
assign LUT_3[62673] = 32'b00000000000000011010011110000001;
assign LUT_3[62674] = 32'b00000000000000010101111010001000;
assign LUT_3[62675] = 32'b00000000000000011100100101100101;
assign LUT_3[62676] = 32'b00000000000000010001000000011010;
assign LUT_3[62677] = 32'b00000000000000010111101011110111;
assign LUT_3[62678] = 32'b00000000000000010011000111111110;
assign LUT_3[62679] = 32'b00000000000000011001110011011011;
assign LUT_3[62680] = 32'b00000000000000011001001011101010;
assign LUT_3[62681] = 32'b00000000000000011111110111000111;
assign LUT_3[62682] = 32'b00000000000000011011010011001110;
assign LUT_3[62683] = 32'b00000000000000100001111110101011;
assign LUT_3[62684] = 32'b00000000000000010110011001100000;
assign LUT_3[62685] = 32'b00000000000000011101000100111101;
assign LUT_3[62686] = 32'b00000000000000011000100001000100;
assign LUT_3[62687] = 32'b00000000000000011111001100100001;
assign LUT_3[62688] = 32'b00000000000000010001101110000001;
assign LUT_3[62689] = 32'b00000000000000011000011001011110;
assign LUT_3[62690] = 32'b00000000000000010011110101100101;
assign LUT_3[62691] = 32'b00000000000000011010100001000010;
assign LUT_3[62692] = 32'b00000000000000001110111011110111;
assign LUT_3[62693] = 32'b00000000000000010101100111010100;
assign LUT_3[62694] = 32'b00000000000000010001000011011011;
assign LUT_3[62695] = 32'b00000000000000010111101110111000;
assign LUT_3[62696] = 32'b00000000000000010111000111000111;
assign LUT_3[62697] = 32'b00000000000000011101110010100100;
assign LUT_3[62698] = 32'b00000000000000011001001110101011;
assign LUT_3[62699] = 32'b00000000000000011111111010001000;
assign LUT_3[62700] = 32'b00000000000000010100010100111101;
assign LUT_3[62701] = 32'b00000000000000011011000000011010;
assign LUT_3[62702] = 32'b00000000000000010110011100100001;
assign LUT_3[62703] = 32'b00000000000000011101000111111110;
assign LUT_3[62704] = 32'b00000000000000010101000001000100;
assign LUT_3[62705] = 32'b00000000000000011011101100100001;
assign LUT_3[62706] = 32'b00000000000000010111001000101000;
assign LUT_3[62707] = 32'b00000000000000011101110100000101;
assign LUT_3[62708] = 32'b00000000000000010010001110111010;
assign LUT_3[62709] = 32'b00000000000000011000111010010111;
assign LUT_3[62710] = 32'b00000000000000010100010110011110;
assign LUT_3[62711] = 32'b00000000000000011011000001111011;
assign LUT_3[62712] = 32'b00000000000000011010011010001010;
assign LUT_3[62713] = 32'b00000000000000100001000101100111;
assign LUT_3[62714] = 32'b00000000000000011100100001101110;
assign LUT_3[62715] = 32'b00000000000000100011001101001011;
assign LUT_3[62716] = 32'b00000000000000010111101000000000;
assign LUT_3[62717] = 32'b00000000000000011110010011011101;
assign LUT_3[62718] = 32'b00000000000000011001101111100100;
assign LUT_3[62719] = 32'b00000000000000100000011011000001;
assign LUT_3[62720] = 32'b00000000000000001010101011011001;
assign LUT_3[62721] = 32'b00000000000000010001010110110110;
assign LUT_3[62722] = 32'b00000000000000001100110010111101;
assign LUT_3[62723] = 32'b00000000000000010011011110011010;
assign LUT_3[62724] = 32'b00000000000000000111111001001111;
assign LUT_3[62725] = 32'b00000000000000001110100100101100;
assign LUT_3[62726] = 32'b00000000000000001010000000110011;
assign LUT_3[62727] = 32'b00000000000000010000101100010000;
assign LUT_3[62728] = 32'b00000000000000010000000100011111;
assign LUT_3[62729] = 32'b00000000000000010110101111111100;
assign LUT_3[62730] = 32'b00000000000000010010001100000011;
assign LUT_3[62731] = 32'b00000000000000011000110111100000;
assign LUT_3[62732] = 32'b00000000000000001101010010010101;
assign LUT_3[62733] = 32'b00000000000000010011111101110010;
assign LUT_3[62734] = 32'b00000000000000001111011001111001;
assign LUT_3[62735] = 32'b00000000000000010110000101010110;
assign LUT_3[62736] = 32'b00000000000000001101111110011100;
assign LUT_3[62737] = 32'b00000000000000010100101001111001;
assign LUT_3[62738] = 32'b00000000000000010000000110000000;
assign LUT_3[62739] = 32'b00000000000000010110110001011101;
assign LUT_3[62740] = 32'b00000000000000001011001100010010;
assign LUT_3[62741] = 32'b00000000000000010001110111101111;
assign LUT_3[62742] = 32'b00000000000000001101010011110110;
assign LUT_3[62743] = 32'b00000000000000010011111111010011;
assign LUT_3[62744] = 32'b00000000000000010011010111100010;
assign LUT_3[62745] = 32'b00000000000000011010000010111111;
assign LUT_3[62746] = 32'b00000000000000010101011111000110;
assign LUT_3[62747] = 32'b00000000000000011100001010100011;
assign LUT_3[62748] = 32'b00000000000000010000100101011000;
assign LUT_3[62749] = 32'b00000000000000010111010000110101;
assign LUT_3[62750] = 32'b00000000000000010010101100111100;
assign LUT_3[62751] = 32'b00000000000000011001011000011001;
assign LUT_3[62752] = 32'b00000000000000001011111001111001;
assign LUT_3[62753] = 32'b00000000000000010010100101010110;
assign LUT_3[62754] = 32'b00000000000000001110000001011101;
assign LUT_3[62755] = 32'b00000000000000010100101100111010;
assign LUT_3[62756] = 32'b00000000000000001001000111101111;
assign LUT_3[62757] = 32'b00000000000000001111110011001100;
assign LUT_3[62758] = 32'b00000000000000001011001111010011;
assign LUT_3[62759] = 32'b00000000000000010001111010110000;
assign LUT_3[62760] = 32'b00000000000000010001010010111111;
assign LUT_3[62761] = 32'b00000000000000010111111110011100;
assign LUT_3[62762] = 32'b00000000000000010011011010100011;
assign LUT_3[62763] = 32'b00000000000000011010000110000000;
assign LUT_3[62764] = 32'b00000000000000001110100000110101;
assign LUT_3[62765] = 32'b00000000000000010101001100010010;
assign LUT_3[62766] = 32'b00000000000000010000101000011001;
assign LUT_3[62767] = 32'b00000000000000010111010011110110;
assign LUT_3[62768] = 32'b00000000000000001111001100111100;
assign LUT_3[62769] = 32'b00000000000000010101111000011001;
assign LUT_3[62770] = 32'b00000000000000010001010100100000;
assign LUT_3[62771] = 32'b00000000000000010111111111111101;
assign LUT_3[62772] = 32'b00000000000000001100011010110010;
assign LUT_3[62773] = 32'b00000000000000010011000110001111;
assign LUT_3[62774] = 32'b00000000000000001110100010010110;
assign LUT_3[62775] = 32'b00000000000000010101001101110011;
assign LUT_3[62776] = 32'b00000000000000010100100110000010;
assign LUT_3[62777] = 32'b00000000000000011011010001011111;
assign LUT_3[62778] = 32'b00000000000000010110101101100110;
assign LUT_3[62779] = 32'b00000000000000011101011001000011;
assign LUT_3[62780] = 32'b00000000000000010001110011111000;
assign LUT_3[62781] = 32'b00000000000000011000011111010101;
assign LUT_3[62782] = 32'b00000000000000010011111011011100;
assign LUT_3[62783] = 32'b00000000000000011010100110111001;
assign LUT_3[62784] = 32'b00000000000000001010100100000100;
assign LUT_3[62785] = 32'b00000000000000010001001111100001;
assign LUT_3[62786] = 32'b00000000000000001100101011101000;
assign LUT_3[62787] = 32'b00000000000000010011010111000101;
assign LUT_3[62788] = 32'b00000000000000000111110001111010;
assign LUT_3[62789] = 32'b00000000000000001110011101010111;
assign LUT_3[62790] = 32'b00000000000000001001111001011110;
assign LUT_3[62791] = 32'b00000000000000010000100100111011;
assign LUT_3[62792] = 32'b00000000000000001111111101001010;
assign LUT_3[62793] = 32'b00000000000000010110101000100111;
assign LUT_3[62794] = 32'b00000000000000010010000100101110;
assign LUT_3[62795] = 32'b00000000000000011000110000001011;
assign LUT_3[62796] = 32'b00000000000000001101001011000000;
assign LUT_3[62797] = 32'b00000000000000010011110110011101;
assign LUT_3[62798] = 32'b00000000000000001111010010100100;
assign LUT_3[62799] = 32'b00000000000000010101111110000001;
assign LUT_3[62800] = 32'b00000000000000001101110111000111;
assign LUT_3[62801] = 32'b00000000000000010100100010100100;
assign LUT_3[62802] = 32'b00000000000000001111111110101011;
assign LUT_3[62803] = 32'b00000000000000010110101010001000;
assign LUT_3[62804] = 32'b00000000000000001011000100111101;
assign LUT_3[62805] = 32'b00000000000000010001110000011010;
assign LUT_3[62806] = 32'b00000000000000001101001100100001;
assign LUT_3[62807] = 32'b00000000000000010011110111111110;
assign LUT_3[62808] = 32'b00000000000000010011010000001101;
assign LUT_3[62809] = 32'b00000000000000011001111011101010;
assign LUT_3[62810] = 32'b00000000000000010101010111110001;
assign LUT_3[62811] = 32'b00000000000000011100000011001110;
assign LUT_3[62812] = 32'b00000000000000010000011110000011;
assign LUT_3[62813] = 32'b00000000000000010111001001100000;
assign LUT_3[62814] = 32'b00000000000000010010100101100111;
assign LUT_3[62815] = 32'b00000000000000011001010001000100;
assign LUT_3[62816] = 32'b00000000000000001011110010100100;
assign LUT_3[62817] = 32'b00000000000000010010011110000001;
assign LUT_3[62818] = 32'b00000000000000001101111010001000;
assign LUT_3[62819] = 32'b00000000000000010100100101100101;
assign LUT_3[62820] = 32'b00000000000000001001000000011010;
assign LUT_3[62821] = 32'b00000000000000001111101011110111;
assign LUT_3[62822] = 32'b00000000000000001011000111111110;
assign LUT_3[62823] = 32'b00000000000000010001110011011011;
assign LUT_3[62824] = 32'b00000000000000010001001011101010;
assign LUT_3[62825] = 32'b00000000000000010111110111000111;
assign LUT_3[62826] = 32'b00000000000000010011010011001110;
assign LUT_3[62827] = 32'b00000000000000011001111110101011;
assign LUT_3[62828] = 32'b00000000000000001110011001100000;
assign LUT_3[62829] = 32'b00000000000000010101000100111101;
assign LUT_3[62830] = 32'b00000000000000010000100001000100;
assign LUT_3[62831] = 32'b00000000000000010111001100100001;
assign LUT_3[62832] = 32'b00000000000000001111000101100111;
assign LUT_3[62833] = 32'b00000000000000010101110001000100;
assign LUT_3[62834] = 32'b00000000000000010001001101001011;
assign LUT_3[62835] = 32'b00000000000000010111111000101000;
assign LUT_3[62836] = 32'b00000000000000001100010011011101;
assign LUT_3[62837] = 32'b00000000000000010010111110111010;
assign LUT_3[62838] = 32'b00000000000000001110011011000001;
assign LUT_3[62839] = 32'b00000000000000010101000110011110;
assign LUT_3[62840] = 32'b00000000000000010100011110101101;
assign LUT_3[62841] = 32'b00000000000000011011001010001010;
assign LUT_3[62842] = 32'b00000000000000010110100110010001;
assign LUT_3[62843] = 32'b00000000000000011101010001101110;
assign LUT_3[62844] = 32'b00000000000000010001101100100011;
assign LUT_3[62845] = 32'b00000000000000011000011000000000;
assign LUT_3[62846] = 32'b00000000000000010011110100000111;
assign LUT_3[62847] = 32'b00000000000000011010011111100100;
assign LUT_3[62848] = 32'b00000000000000001100110110010111;
assign LUT_3[62849] = 32'b00000000000000010011100001110100;
assign LUT_3[62850] = 32'b00000000000000001110111101111011;
assign LUT_3[62851] = 32'b00000000000000010101101001011000;
assign LUT_3[62852] = 32'b00000000000000001010000100001101;
assign LUT_3[62853] = 32'b00000000000000010000101111101010;
assign LUT_3[62854] = 32'b00000000000000001100001011110001;
assign LUT_3[62855] = 32'b00000000000000010010110111001110;
assign LUT_3[62856] = 32'b00000000000000010010001111011101;
assign LUT_3[62857] = 32'b00000000000000011000111010111010;
assign LUT_3[62858] = 32'b00000000000000010100010111000001;
assign LUT_3[62859] = 32'b00000000000000011011000010011110;
assign LUT_3[62860] = 32'b00000000000000001111011101010011;
assign LUT_3[62861] = 32'b00000000000000010110001000110000;
assign LUT_3[62862] = 32'b00000000000000010001100100110111;
assign LUT_3[62863] = 32'b00000000000000011000010000010100;
assign LUT_3[62864] = 32'b00000000000000010000001001011010;
assign LUT_3[62865] = 32'b00000000000000010110110100110111;
assign LUT_3[62866] = 32'b00000000000000010010010000111110;
assign LUT_3[62867] = 32'b00000000000000011000111100011011;
assign LUT_3[62868] = 32'b00000000000000001101010111010000;
assign LUT_3[62869] = 32'b00000000000000010100000010101101;
assign LUT_3[62870] = 32'b00000000000000001111011110110100;
assign LUT_3[62871] = 32'b00000000000000010110001010010001;
assign LUT_3[62872] = 32'b00000000000000010101100010100000;
assign LUT_3[62873] = 32'b00000000000000011100001101111101;
assign LUT_3[62874] = 32'b00000000000000010111101010000100;
assign LUT_3[62875] = 32'b00000000000000011110010101100001;
assign LUT_3[62876] = 32'b00000000000000010010110000010110;
assign LUT_3[62877] = 32'b00000000000000011001011011110011;
assign LUT_3[62878] = 32'b00000000000000010100110111111010;
assign LUT_3[62879] = 32'b00000000000000011011100011010111;
assign LUT_3[62880] = 32'b00000000000000001110000100110111;
assign LUT_3[62881] = 32'b00000000000000010100110000010100;
assign LUT_3[62882] = 32'b00000000000000010000001100011011;
assign LUT_3[62883] = 32'b00000000000000010110110111111000;
assign LUT_3[62884] = 32'b00000000000000001011010010101101;
assign LUT_3[62885] = 32'b00000000000000010001111110001010;
assign LUT_3[62886] = 32'b00000000000000001101011010010001;
assign LUT_3[62887] = 32'b00000000000000010100000101101110;
assign LUT_3[62888] = 32'b00000000000000010011011101111101;
assign LUT_3[62889] = 32'b00000000000000011010001001011010;
assign LUT_3[62890] = 32'b00000000000000010101100101100001;
assign LUT_3[62891] = 32'b00000000000000011100010000111110;
assign LUT_3[62892] = 32'b00000000000000010000101011110011;
assign LUT_3[62893] = 32'b00000000000000010111010111010000;
assign LUT_3[62894] = 32'b00000000000000010010110011010111;
assign LUT_3[62895] = 32'b00000000000000011001011110110100;
assign LUT_3[62896] = 32'b00000000000000010001010111111010;
assign LUT_3[62897] = 32'b00000000000000011000000011010111;
assign LUT_3[62898] = 32'b00000000000000010011011111011110;
assign LUT_3[62899] = 32'b00000000000000011010001010111011;
assign LUT_3[62900] = 32'b00000000000000001110100101110000;
assign LUT_3[62901] = 32'b00000000000000010101010001001101;
assign LUT_3[62902] = 32'b00000000000000010000101101010100;
assign LUT_3[62903] = 32'b00000000000000010111011000110001;
assign LUT_3[62904] = 32'b00000000000000010110110001000000;
assign LUT_3[62905] = 32'b00000000000000011101011100011101;
assign LUT_3[62906] = 32'b00000000000000011000111000100100;
assign LUT_3[62907] = 32'b00000000000000011111100100000001;
assign LUT_3[62908] = 32'b00000000000000010011111110110110;
assign LUT_3[62909] = 32'b00000000000000011010101010010011;
assign LUT_3[62910] = 32'b00000000000000010110000110011010;
assign LUT_3[62911] = 32'b00000000000000011100110001110111;
assign LUT_3[62912] = 32'b00000000000000001100101111000010;
assign LUT_3[62913] = 32'b00000000000000010011011010011111;
assign LUT_3[62914] = 32'b00000000000000001110110110100110;
assign LUT_3[62915] = 32'b00000000000000010101100010000011;
assign LUT_3[62916] = 32'b00000000000000001001111100111000;
assign LUT_3[62917] = 32'b00000000000000010000101000010101;
assign LUT_3[62918] = 32'b00000000000000001100000100011100;
assign LUT_3[62919] = 32'b00000000000000010010101111111001;
assign LUT_3[62920] = 32'b00000000000000010010001000001000;
assign LUT_3[62921] = 32'b00000000000000011000110011100101;
assign LUT_3[62922] = 32'b00000000000000010100001111101100;
assign LUT_3[62923] = 32'b00000000000000011010111011001001;
assign LUT_3[62924] = 32'b00000000000000001111010101111110;
assign LUT_3[62925] = 32'b00000000000000010110000001011011;
assign LUT_3[62926] = 32'b00000000000000010001011101100010;
assign LUT_3[62927] = 32'b00000000000000011000001000111111;
assign LUT_3[62928] = 32'b00000000000000010000000010000101;
assign LUT_3[62929] = 32'b00000000000000010110101101100010;
assign LUT_3[62930] = 32'b00000000000000010010001001101001;
assign LUT_3[62931] = 32'b00000000000000011000110101000110;
assign LUT_3[62932] = 32'b00000000000000001101001111111011;
assign LUT_3[62933] = 32'b00000000000000010011111011011000;
assign LUT_3[62934] = 32'b00000000000000001111010111011111;
assign LUT_3[62935] = 32'b00000000000000010110000010111100;
assign LUT_3[62936] = 32'b00000000000000010101011011001011;
assign LUT_3[62937] = 32'b00000000000000011100000110101000;
assign LUT_3[62938] = 32'b00000000000000010111100010101111;
assign LUT_3[62939] = 32'b00000000000000011110001110001100;
assign LUT_3[62940] = 32'b00000000000000010010101001000001;
assign LUT_3[62941] = 32'b00000000000000011001010100011110;
assign LUT_3[62942] = 32'b00000000000000010100110000100101;
assign LUT_3[62943] = 32'b00000000000000011011011100000010;
assign LUT_3[62944] = 32'b00000000000000001101111101100010;
assign LUT_3[62945] = 32'b00000000000000010100101000111111;
assign LUT_3[62946] = 32'b00000000000000010000000101000110;
assign LUT_3[62947] = 32'b00000000000000010110110000100011;
assign LUT_3[62948] = 32'b00000000000000001011001011011000;
assign LUT_3[62949] = 32'b00000000000000010001110110110101;
assign LUT_3[62950] = 32'b00000000000000001101010010111100;
assign LUT_3[62951] = 32'b00000000000000010011111110011001;
assign LUT_3[62952] = 32'b00000000000000010011010110101000;
assign LUT_3[62953] = 32'b00000000000000011010000010000101;
assign LUT_3[62954] = 32'b00000000000000010101011110001100;
assign LUT_3[62955] = 32'b00000000000000011100001001101001;
assign LUT_3[62956] = 32'b00000000000000010000100100011110;
assign LUT_3[62957] = 32'b00000000000000010111001111111011;
assign LUT_3[62958] = 32'b00000000000000010010101100000010;
assign LUT_3[62959] = 32'b00000000000000011001010111011111;
assign LUT_3[62960] = 32'b00000000000000010001010000100101;
assign LUT_3[62961] = 32'b00000000000000010111111100000010;
assign LUT_3[62962] = 32'b00000000000000010011011000001001;
assign LUT_3[62963] = 32'b00000000000000011010000011100110;
assign LUT_3[62964] = 32'b00000000000000001110011110011011;
assign LUT_3[62965] = 32'b00000000000000010101001001111000;
assign LUT_3[62966] = 32'b00000000000000010000100101111111;
assign LUT_3[62967] = 32'b00000000000000010111010001011100;
assign LUT_3[62968] = 32'b00000000000000010110101001101011;
assign LUT_3[62969] = 32'b00000000000000011101010101001000;
assign LUT_3[62970] = 32'b00000000000000011000110001001111;
assign LUT_3[62971] = 32'b00000000000000011111011100101100;
assign LUT_3[62972] = 32'b00000000000000010011110111100001;
assign LUT_3[62973] = 32'b00000000000000011010100010111110;
assign LUT_3[62974] = 32'b00000000000000010101111111000101;
assign LUT_3[62975] = 32'b00000000000000011100101010100010;
assign LUT_3[62976] = 32'b00000000000000010001110001000100;
assign LUT_3[62977] = 32'b00000000000000011000011100100001;
assign LUT_3[62978] = 32'b00000000000000010011111000101000;
assign LUT_3[62979] = 32'b00000000000000011010100100000101;
assign LUT_3[62980] = 32'b00000000000000001110111110111010;
assign LUT_3[62981] = 32'b00000000000000010101101010010111;
assign LUT_3[62982] = 32'b00000000000000010001000110011110;
assign LUT_3[62983] = 32'b00000000000000010111110001111011;
assign LUT_3[62984] = 32'b00000000000000010111001010001010;
assign LUT_3[62985] = 32'b00000000000000011101110101100111;
assign LUT_3[62986] = 32'b00000000000000011001010001101110;
assign LUT_3[62987] = 32'b00000000000000011111111101001011;
assign LUT_3[62988] = 32'b00000000000000010100011000000000;
assign LUT_3[62989] = 32'b00000000000000011011000011011101;
assign LUT_3[62990] = 32'b00000000000000010110011111100100;
assign LUT_3[62991] = 32'b00000000000000011101001011000001;
assign LUT_3[62992] = 32'b00000000000000010101000100000111;
assign LUT_3[62993] = 32'b00000000000000011011101111100100;
assign LUT_3[62994] = 32'b00000000000000010111001011101011;
assign LUT_3[62995] = 32'b00000000000000011101110111001000;
assign LUT_3[62996] = 32'b00000000000000010010010001111101;
assign LUT_3[62997] = 32'b00000000000000011000111101011010;
assign LUT_3[62998] = 32'b00000000000000010100011001100001;
assign LUT_3[62999] = 32'b00000000000000011011000100111110;
assign LUT_3[63000] = 32'b00000000000000011010011101001101;
assign LUT_3[63001] = 32'b00000000000000100001001000101010;
assign LUT_3[63002] = 32'b00000000000000011100100100110001;
assign LUT_3[63003] = 32'b00000000000000100011010000001110;
assign LUT_3[63004] = 32'b00000000000000010111101011000011;
assign LUT_3[63005] = 32'b00000000000000011110010110100000;
assign LUT_3[63006] = 32'b00000000000000011001110010100111;
assign LUT_3[63007] = 32'b00000000000000100000011110000100;
assign LUT_3[63008] = 32'b00000000000000010010111111100100;
assign LUT_3[63009] = 32'b00000000000000011001101011000001;
assign LUT_3[63010] = 32'b00000000000000010101000111001000;
assign LUT_3[63011] = 32'b00000000000000011011110010100101;
assign LUT_3[63012] = 32'b00000000000000010000001101011010;
assign LUT_3[63013] = 32'b00000000000000010110111000110111;
assign LUT_3[63014] = 32'b00000000000000010010010100111110;
assign LUT_3[63015] = 32'b00000000000000011001000000011011;
assign LUT_3[63016] = 32'b00000000000000011000011000101010;
assign LUT_3[63017] = 32'b00000000000000011111000100000111;
assign LUT_3[63018] = 32'b00000000000000011010100000001110;
assign LUT_3[63019] = 32'b00000000000000100001001011101011;
assign LUT_3[63020] = 32'b00000000000000010101100110100000;
assign LUT_3[63021] = 32'b00000000000000011100010001111101;
assign LUT_3[63022] = 32'b00000000000000010111101110000100;
assign LUT_3[63023] = 32'b00000000000000011110011001100001;
assign LUT_3[63024] = 32'b00000000000000010110010010100111;
assign LUT_3[63025] = 32'b00000000000000011100111110000100;
assign LUT_3[63026] = 32'b00000000000000011000011010001011;
assign LUT_3[63027] = 32'b00000000000000011111000101101000;
assign LUT_3[63028] = 32'b00000000000000010011100000011101;
assign LUT_3[63029] = 32'b00000000000000011010001011111010;
assign LUT_3[63030] = 32'b00000000000000010101101000000001;
assign LUT_3[63031] = 32'b00000000000000011100010011011110;
assign LUT_3[63032] = 32'b00000000000000011011101011101101;
assign LUT_3[63033] = 32'b00000000000000100010010111001010;
assign LUT_3[63034] = 32'b00000000000000011101110011010001;
assign LUT_3[63035] = 32'b00000000000000100100011110101110;
assign LUT_3[63036] = 32'b00000000000000011000111001100011;
assign LUT_3[63037] = 32'b00000000000000011111100101000000;
assign LUT_3[63038] = 32'b00000000000000011011000001000111;
assign LUT_3[63039] = 32'b00000000000000100001101100100100;
assign LUT_3[63040] = 32'b00000000000000010001101001101111;
assign LUT_3[63041] = 32'b00000000000000011000010101001100;
assign LUT_3[63042] = 32'b00000000000000010011110001010011;
assign LUT_3[63043] = 32'b00000000000000011010011100110000;
assign LUT_3[63044] = 32'b00000000000000001110110111100101;
assign LUT_3[63045] = 32'b00000000000000010101100011000010;
assign LUT_3[63046] = 32'b00000000000000010000111111001001;
assign LUT_3[63047] = 32'b00000000000000010111101010100110;
assign LUT_3[63048] = 32'b00000000000000010111000010110101;
assign LUT_3[63049] = 32'b00000000000000011101101110010010;
assign LUT_3[63050] = 32'b00000000000000011001001010011001;
assign LUT_3[63051] = 32'b00000000000000011111110101110110;
assign LUT_3[63052] = 32'b00000000000000010100010000101011;
assign LUT_3[63053] = 32'b00000000000000011010111100001000;
assign LUT_3[63054] = 32'b00000000000000010110011000001111;
assign LUT_3[63055] = 32'b00000000000000011101000011101100;
assign LUT_3[63056] = 32'b00000000000000010100111100110010;
assign LUT_3[63057] = 32'b00000000000000011011101000001111;
assign LUT_3[63058] = 32'b00000000000000010111000100010110;
assign LUT_3[63059] = 32'b00000000000000011101101111110011;
assign LUT_3[63060] = 32'b00000000000000010010001010101000;
assign LUT_3[63061] = 32'b00000000000000011000110110000101;
assign LUT_3[63062] = 32'b00000000000000010100010010001100;
assign LUT_3[63063] = 32'b00000000000000011010111101101001;
assign LUT_3[63064] = 32'b00000000000000011010010101111000;
assign LUT_3[63065] = 32'b00000000000000100001000001010101;
assign LUT_3[63066] = 32'b00000000000000011100011101011100;
assign LUT_3[63067] = 32'b00000000000000100011001000111001;
assign LUT_3[63068] = 32'b00000000000000010111100011101110;
assign LUT_3[63069] = 32'b00000000000000011110001111001011;
assign LUT_3[63070] = 32'b00000000000000011001101011010010;
assign LUT_3[63071] = 32'b00000000000000100000010110101111;
assign LUT_3[63072] = 32'b00000000000000010010111000001111;
assign LUT_3[63073] = 32'b00000000000000011001100011101100;
assign LUT_3[63074] = 32'b00000000000000010100111111110011;
assign LUT_3[63075] = 32'b00000000000000011011101011010000;
assign LUT_3[63076] = 32'b00000000000000010000000110000101;
assign LUT_3[63077] = 32'b00000000000000010110110001100010;
assign LUT_3[63078] = 32'b00000000000000010010001101101001;
assign LUT_3[63079] = 32'b00000000000000011000111001000110;
assign LUT_3[63080] = 32'b00000000000000011000010001010101;
assign LUT_3[63081] = 32'b00000000000000011110111100110010;
assign LUT_3[63082] = 32'b00000000000000011010011000111001;
assign LUT_3[63083] = 32'b00000000000000100001000100010110;
assign LUT_3[63084] = 32'b00000000000000010101011111001011;
assign LUT_3[63085] = 32'b00000000000000011100001010101000;
assign LUT_3[63086] = 32'b00000000000000010111100110101111;
assign LUT_3[63087] = 32'b00000000000000011110010010001100;
assign LUT_3[63088] = 32'b00000000000000010110001011010010;
assign LUT_3[63089] = 32'b00000000000000011100110110101111;
assign LUT_3[63090] = 32'b00000000000000011000010010110110;
assign LUT_3[63091] = 32'b00000000000000011110111110010011;
assign LUT_3[63092] = 32'b00000000000000010011011001001000;
assign LUT_3[63093] = 32'b00000000000000011010000100100101;
assign LUT_3[63094] = 32'b00000000000000010101100000101100;
assign LUT_3[63095] = 32'b00000000000000011100001100001001;
assign LUT_3[63096] = 32'b00000000000000011011100100011000;
assign LUT_3[63097] = 32'b00000000000000100010001111110101;
assign LUT_3[63098] = 32'b00000000000000011101101011111100;
assign LUT_3[63099] = 32'b00000000000000100100010111011001;
assign LUT_3[63100] = 32'b00000000000000011000110010001110;
assign LUT_3[63101] = 32'b00000000000000011111011101101011;
assign LUT_3[63102] = 32'b00000000000000011010111001110010;
assign LUT_3[63103] = 32'b00000000000000100001100101001111;
assign LUT_3[63104] = 32'b00000000000000010011111100000010;
assign LUT_3[63105] = 32'b00000000000000011010100111011111;
assign LUT_3[63106] = 32'b00000000000000010110000011100110;
assign LUT_3[63107] = 32'b00000000000000011100101111000011;
assign LUT_3[63108] = 32'b00000000000000010001001001111000;
assign LUT_3[63109] = 32'b00000000000000010111110101010101;
assign LUT_3[63110] = 32'b00000000000000010011010001011100;
assign LUT_3[63111] = 32'b00000000000000011001111100111001;
assign LUT_3[63112] = 32'b00000000000000011001010101001000;
assign LUT_3[63113] = 32'b00000000000000100000000000100101;
assign LUT_3[63114] = 32'b00000000000000011011011100101100;
assign LUT_3[63115] = 32'b00000000000000100010001000001001;
assign LUT_3[63116] = 32'b00000000000000010110100010111110;
assign LUT_3[63117] = 32'b00000000000000011101001110011011;
assign LUT_3[63118] = 32'b00000000000000011000101010100010;
assign LUT_3[63119] = 32'b00000000000000011111010101111111;
assign LUT_3[63120] = 32'b00000000000000010111001111000101;
assign LUT_3[63121] = 32'b00000000000000011101111010100010;
assign LUT_3[63122] = 32'b00000000000000011001010110101001;
assign LUT_3[63123] = 32'b00000000000000100000000010000110;
assign LUT_3[63124] = 32'b00000000000000010100011100111011;
assign LUT_3[63125] = 32'b00000000000000011011001000011000;
assign LUT_3[63126] = 32'b00000000000000010110100100011111;
assign LUT_3[63127] = 32'b00000000000000011101001111111100;
assign LUT_3[63128] = 32'b00000000000000011100101000001011;
assign LUT_3[63129] = 32'b00000000000000100011010011101000;
assign LUT_3[63130] = 32'b00000000000000011110101111101111;
assign LUT_3[63131] = 32'b00000000000000100101011011001100;
assign LUT_3[63132] = 32'b00000000000000011001110110000001;
assign LUT_3[63133] = 32'b00000000000000100000100001011110;
assign LUT_3[63134] = 32'b00000000000000011011111101100101;
assign LUT_3[63135] = 32'b00000000000000100010101001000010;
assign LUT_3[63136] = 32'b00000000000000010101001010100010;
assign LUT_3[63137] = 32'b00000000000000011011110101111111;
assign LUT_3[63138] = 32'b00000000000000010111010010000110;
assign LUT_3[63139] = 32'b00000000000000011101111101100011;
assign LUT_3[63140] = 32'b00000000000000010010011000011000;
assign LUT_3[63141] = 32'b00000000000000011001000011110101;
assign LUT_3[63142] = 32'b00000000000000010100011111111100;
assign LUT_3[63143] = 32'b00000000000000011011001011011001;
assign LUT_3[63144] = 32'b00000000000000011010100011101000;
assign LUT_3[63145] = 32'b00000000000000100001001111000101;
assign LUT_3[63146] = 32'b00000000000000011100101011001100;
assign LUT_3[63147] = 32'b00000000000000100011010110101001;
assign LUT_3[63148] = 32'b00000000000000010111110001011110;
assign LUT_3[63149] = 32'b00000000000000011110011100111011;
assign LUT_3[63150] = 32'b00000000000000011001111001000010;
assign LUT_3[63151] = 32'b00000000000000100000100100011111;
assign LUT_3[63152] = 32'b00000000000000011000011101100101;
assign LUT_3[63153] = 32'b00000000000000011111001001000010;
assign LUT_3[63154] = 32'b00000000000000011010100101001001;
assign LUT_3[63155] = 32'b00000000000000100001010000100110;
assign LUT_3[63156] = 32'b00000000000000010101101011011011;
assign LUT_3[63157] = 32'b00000000000000011100010110111000;
assign LUT_3[63158] = 32'b00000000000000010111110010111111;
assign LUT_3[63159] = 32'b00000000000000011110011110011100;
assign LUT_3[63160] = 32'b00000000000000011101110110101011;
assign LUT_3[63161] = 32'b00000000000000100100100010001000;
assign LUT_3[63162] = 32'b00000000000000011111111110001111;
assign LUT_3[63163] = 32'b00000000000000100110101001101100;
assign LUT_3[63164] = 32'b00000000000000011011000100100001;
assign LUT_3[63165] = 32'b00000000000000100001101111111110;
assign LUT_3[63166] = 32'b00000000000000011101001100000101;
assign LUT_3[63167] = 32'b00000000000000100011110111100010;
assign LUT_3[63168] = 32'b00000000000000010011110100101101;
assign LUT_3[63169] = 32'b00000000000000011010100000001010;
assign LUT_3[63170] = 32'b00000000000000010101111100010001;
assign LUT_3[63171] = 32'b00000000000000011100100111101110;
assign LUT_3[63172] = 32'b00000000000000010001000010100011;
assign LUT_3[63173] = 32'b00000000000000010111101110000000;
assign LUT_3[63174] = 32'b00000000000000010011001010000111;
assign LUT_3[63175] = 32'b00000000000000011001110101100100;
assign LUT_3[63176] = 32'b00000000000000011001001101110011;
assign LUT_3[63177] = 32'b00000000000000011111111001010000;
assign LUT_3[63178] = 32'b00000000000000011011010101010111;
assign LUT_3[63179] = 32'b00000000000000100010000000110100;
assign LUT_3[63180] = 32'b00000000000000010110011011101001;
assign LUT_3[63181] = 32'b00000000000000011101000111000110;
assign LUT_3[63182] = 32'b00000000000000011000100011001101;
assign LUT_3[63183] = 32'b00000000000000011111001110101010;
assign LUT_3[63184] = 32'b00000000000000010111000111110000;
assign LUT_3[63185] = 32'b00000000000000011101110011001101;
assign LUT_3[63186] = 32'b00000000000000011001001111010100;
assign LUT_3[63187] = 32'b00000000000000011111111010110001;
assign LUT_3[63188] = 32'b00000000000000010100010101100110;
assign LUT_3[63189] = 32'b00000000000000011011000001000011;
assign LUT_3[63190] = 32'b00000000000000010110011101001010;
assign LUT_3[63191] = 32'b00000000000000011101001000100111;
assign LUT_3[63192] = 32'b00000000000000011100100000110110;
assign LUT_3[63193] = 32'b00000000000000100011001100010011;
assign LUT_3[63194] = 32'b00000000000000011110101000011010;
assign LUT_3[63195] = 32'b00000000000000100101010011110111;
assign LUT_3[63196] = 32'b00000000000000011001101110101100;
assign LUT_3[63197] = 32'b00000000000000100000011010001001;
assign LUT_3[63198] = 32'b00000000000000011011110110010000;
assign LUT_3[63199] = 32'b00000000000000100010100001101101;
assign LUT_3[63200] = 32'b00000000000000010101000011001101;
assign LUT_3[63201] = 32'b00000000000000011011101110101010;
assign LUT_3[63202] = 32'b00000000000000010111001010110001;
assign LUT_3[63203] = 32'b00000000000000011101110110001110;
assign LUT_3[63204] = 32'b00000000000000010010010001000011;
assign LUT_3[63205] = 32'b00000000000000011000111100100000;
assign LUT_3[63206] = 32'b00000000000000010100011000100111;
assign LUT_3[63207] = 32'b00000000000000011011000100000100;
assign LUT_3[63208] = 32'b00000000000000011010011100010011;
assign LUT_3[63209] = 32'b00000000000000100001000111110000;
assign LUT_3[63210] = 32'b00000000000000011100100011110111;
assign LUT_3[63211] = 32'b00000000000000100011001111010100;
assign LUT_3[63212] = 32'b00000000000000010111101010001001;
assign LUT_3[63213] = 32'b00000000000000011110010101100110;
assign LUT_3[63214] = 32'b00000000000000011001110001101101;
assign LUT_3[63215] = 32'b00000000000000100000011101001010;
assign LUT_3[63216] = 32'b00000000000000011000010110010000;
assign LUT_3[63217] = 32'b00000000000000011111000001101101;
assign LUT_3[63218] = 32'b00000000000000011010011101110100;
assign LUT_3[63219] = 32'b00000000000000100001001001010001;
assign LUT_3[63220] = 32'b00000000000000010101100100000110;
assign LUT_3[63221] = 32'b00000000000000011100001111100011;
assign LUT_3[63222] = 32'b00000000000000010111101011101010;
assign LUT_3[63223] = 32'b00000000000000011110010111000111;
assign LUT_3[63224] = 32'b00000000000000011101101111010110;
assign LUT_3[63225] = 32'b00000000000000100100011010110011;
assign LUT_3[63226] = 32'b00000000000000011111110110111010;
assign LUT_3[63227] = 32'b00000000000000100110100010010111;
assign LUT_3[63228] = 32'b00000000000000011010111101001100;
assign LUT_3[63229] = 32'b00000000000000100001101000101001;
assign LUT_3[63230] = 32'b00000000000000011101000100110000;
assign LUT_3[63231] = 32'b00000000000000100011110000001101;
assign LUT_3[63232] = 32'b00000000000000001110000000100101;
assign LUT_3[63233] = 32'b00000000000000010100101100000010;
assign LUT_3[63234] = 32'b00000000000000010000001000001001;
assign LUT_3[63235] = 32'b00000000000000010110110011100110;
assign LUT_3[63236] = 32'b00000000000000001011001110011011;
assign LUT_3[63237] = 32'b00000000000000010001111001111000;
assign LUT_3[63238] = 32'b00000000000000001101010101111111;
assign LUT_3[63239] = 32'b00000000000000010100000001011100;
assign LUT_3[63240] = 32'b00000000000000010011011001101011;
assign LUT_3[63241] = 32'b00000000000000011010000101001000;
assign LUT_3[63242] = 32'b00000000000000010101100001001111;
assign LUT_3[63243] = 32'b00000000000000011100001100101100;
assign LUT_3[63244] = 32'b00000000000000010000100111100001;
assign LUT_3[63245] = 32'b00000000000000010111010010111110;
assign LUT_3[63246] = 32'b00000000000000010010101111000101;
assign LUT_3[63247] = 32'b00000000000000011001011010100010;
assign LUT_3[63248] = 32'b00000000000000010001010011101000;
assign LUT_3[63249] = 32'b00000000000000010111111111000101;
assign LUT_3[63250] = 32'b00000000000000010011011011001100;
assign LUT_3[63251] = 32'b00000000000000011010000110101001;
assign LUT_3[63252] = 32'b00000000000000001110100001011110;
assign LUT_3[63253] = 32'b00000000000000010101001100111011;
assign LUT_3[63254] = 32'b00000000000000010000101001000010;
assign LUT_3[63255] = 32'b00000000000000010111010100011111;
assign LUT_3[63256] = 32'b00000000000000010110101100101110;
assign LUT_3[63257] = 32'b00000000000000011101011000001011;
assign LUT_3[63258] = 32'b00000000000000011000110100010010;
assign LUT_3[63259] = 32'b00000000000000011111011111101111;
assign LUT_3[63260] = 32'b00000000000000010011111010100100;
assign LUT_3[63261] = 32'b00000000000000011010100110000001;
assign LUT_3[63262] = 32'b00000000000000010110000010001000;
assign LUT_3[63263] = 32'b00000000000000011100101101100101;
assign LUT_3[63264] = 32'b00000000000000001111001111000101;
assign LUT_3[63265] = 32'b00000000000000010101111010100010;
assign LUT_3[63266] = 32'b00000000000000010001010110101001;
assign LUT_3[63267] = 32'b00000000000000011000000010000110;
assign LUT_3[63268] = 32'b00000000000000001100011100111011;
assign LUT_3[63269] = 32'b00000000000000010011001000011000;
assign LUT_3[63270] = 32'b00000000000000001110100100011111;
assign LUT_3[63271] = 32'b00000000000000010101001111111100;
assign LUT_3[63272] = 32'b00000000000000010100101000001011;
assign LUT_3[63273] = 32'b00000000000000011011010011101000;
assign LUT_3[63274] = 32'b00000000000000010110101111101111;
assign LUT_3[63275] = 32'b00000000000000011101011011001100;
assign LUT_3[63276] = 32'b00000000000000010001110110000001;
assign LUT_3[63277] = 32'b00000000000000011000100001011110;
assign LUT_3[63278] = 32'b00000000000000010011111101100101;
assign LUT_3[63279] = 32'b00000000000000011010101001000010;
assign LUT_3[63280] = 32'b00000000000000010010100010001000;
assign LUT_3[63281] = 32'b00000000000000011001001101100101;
assign LUT_3[63282] = 32'b00000000000000010100101001101100;
assign LUT_3[63283] = 32'b00000000000000011011010101001001;
assign LUT_3[63284] = 32'b00000000000000001111101111111110;
assign LUT_3[63285] = 32'b00000000000000010110011011011011;
assign LUT_3[63286] = 32'b00000000000000010001110111100010;
assign LUT_3[63287] = 32'b00000000000000011000100010111111;
assign LUT_3[63288] = 32'b00000000000000010111111011001110;
assign LUT_3[63289] = 32'b00000000000000011110100110101011;
assign LUT_3[63290] = 32'b00000000000000011010000010110010;
assign LUT_3[63291] = 32'b00000000000000100000101110001111;
assign LUT_3[63292] = 32'b00000000000000010101001001000100;
assign LUT_3[63293] = 32'b00000000000000011011110100100001;
assign LUT_3[63294] = 32'b00000000000000010111010000101000;
assign LUT_3[63295] = 32'b00000000000000011101111100000101;
assign LUT_3[63296] = 32'b00000000000000001101111001010000;
assign LUT_3[63297] = 32'b00000000000000010100100100101101;
assign LUT_3[63298] = 32'b00000000000000010000000000110100;
assign LUT_3[63299] = 32'b00000000000000010110101100010001;
assign LUT_3[63300] = 32'b00000000000000001011000111000110;
assign LUT_3[63301] = 32'b00000000000000010001110010100011;
assign LUT_3[63302] = 32'b00000000000000001101001110101010;
assign LUT_3[63303] = 32'b00000000000000010011111010000111;
assign LUT_3[63304] = 32'b00000000000000010011010010010110;
assign LUT_3[63305] = 32'b00000000000000011001111101110011;
assign LUT_3[63306] = 32'b00000000000000010101011001111010;
assign LUT_3[63307] = 32'b00000000000000011100000101010111;
assign LUT_3[63308] = 32'b00000000000000010000100000001100;
assign LUT_3[63309] = 32'b00000000000000010111001011101001;
assign LUT_3[63310] = 32'b00000000000000010010100111110000;
assign LUT_3[63311] = 32'b00000000000000011001010011001101;
assign LUT_3[63312] = 32'b00000000000000010001001100010011;
assign LUT_3[63313] = 32'b00000000000000010111110111110000;
assign LUT_3[63314] = 32'b00000000000000010011010011110111;
assign LUT_3[63315] = 32'b00000000000000011001111111010100;
assign LUT_3[63316] = 32'b00000000000000001110011010001001;
assign LUT_3[63317] = 32'b00000000000000010101000101100110;
assign LUT_3[63318] = 32'b00000000000000010000100001101101;
assign LUT_3[63319] = 32'b00000000000000010111001101001010;
assign LUT_3[63320] = 32'b00000000000000010110100101011001;
assign LUT_3[63321] = 32'b00000000000000011101010000110110;
assign LUT_3[63322] = 32'b00000000000000011000101100111101;
assign LUT_3[63323] = 32'b00000000000000011111011000011010;
assign LUT_3[63324] = 32'b00000000000000010011110011001111;
assign LUT_3[63325] = 32'b00000000000000011010011110101100;
assign LUT_3[63326] = 32'b00000000000000010101111010110011;
assign LUT_3[63327] = 32'b00000000000000011100100110010000;
assign LUT_3[63328] = 32'b00000000000000001111000111110000;
assign LUT_3[63329] = 32'b00000000000000010101110011001101;
assign LUT_3[63330] = 32'b00000000000000010001001111010100;
assign LUT_3[63331] = 32'b00000000000000010111111010110001;
assign LUT_3[63332] = 32'b00000000000000001100010101100110;
assign LUT_3[63333] = 32'b00000000000000010011000001000011;
assign LUT_3[63334] = 32'b00000000000000001110011101001010;
assign LUT_3[63335] = 32'b00000000000000010101001000100111;
assign LUT_3[63336] = 32'b00000000000000010100100000110110;
assign LUT_3[63337] = 32'b00000000000000011011001100010011;
assign LUT_3[63338] = 32'b00000000000000010110101000011010;
assign LUT_3[63339] = 32'b00000000000000011101010011110111;
assign LUT_3[63340] = 32'b00000000000000010001101110101100;
assign LUT_3[63341] = 32'b00000000000000011000011010001001;
assign LUT_3[63342] = 32'b00000000000000010011110110010000;
assign LUT_3[63343] = 32'b00000000000000011010100001101101;
assign LUT_3[63344] = 32'b00000000000000010010011010110011;
assign LUT_3[63345] = 32'b00000000000000011001000110010000;
assign LUT_3[63346] = 32'b00000000000000010100100010010111;
assign LUT_3[63347] = 32'b00000000000000011011001101110100;
assign LUT_3[63348] = 32'b00000000000000001111101000101001;
assign LUT_3[63349] = 32'b00000000000000010110010100000110;
assign LUT_3[63350] = 32'b00000000000000010001110000001101;
assign LUT_3[63351] = 32'b00000000000000011000011011101010;
assign LUT_3[63352] = 32'b00000000000000010111110011111001;
assign LUT_3[63353] = 32'b00000000000000011110011111010110;
assign LUT_3[63354] = 32'b00000000000000011001111011011101;
assign LUT_3[63355] = 32'b00000000000000100000100110111010;
assign LUT_3[63356] = 32'b00000000000000010101000001101111;
assign LUT_3[63357] = 32'b00000000000000011011101101001100;
assign LUT_3[63358] = 32'b00000000000000010111001001010011;
assign LUT_3[63359] = 32'b00000000000000011101110100110000;
assign LUT_3[63360] = 32'b00000000000000010000001011100011;
assign LUT_3[63361] = 32'b00000000000000010110110111000000;
assign LUT_3[63362] = 32'b00000000000000010010010011000111;
assign LUT_3[63363] = 32'b00000000000000011000111110100100;
assign LUT_3[63364] = 32'b00000000000000001101011001011001;
assign LUT_3[63365] = 32'b00000000000000010100000100110110;
assign LUT_3[63366] = 32'b00000000000000001111100000111101;
assign LUT_3[63367] = 32'b00000000000000010110001100011010;
assign LUT_3[63368] = 32'b00000000000000010101100100101001;
assign LUT_3[63369] = 32'b00000000000000011100010000000110;
assign LUT_3[63370] = 32'b00000000000000010111101100001101;
assign LUT_3[63371] = 32'b00000000000000011110010111101010;
assign LUT_3[63372] = 32'b00000000000000010010110010011111;
assign LUT_3[63373] = 32'b00000000000000011001011101111100;
assign LUT_3[63374] = 32'b00000000000000010100111010000011;
assign LUT_3[63375] = 32'b00000000000000011011100101100000;
assign LUT_3[63376] = 32'b00000000000000010011011110100110;
assign LUT_3[63377] = 32'b00000000000000011010001010000011;
assign LUT_3[63378] = 32'b00000000000000010101100110001010;
assign LUT_3[63379] = 32'b00000000000000011100010001100111;
assign LUT_3[63380] = 32'b00000000000000010000101100011100;
assign LUT_3[63381] = 32'b00000000000000010111010111111001;
assign LUT_3[63382] = 32'b00000000000000010010110100000000;
assign LUT_3[63383] = 32'b00000000000000011001011111011101;
assign LUT_3[63384] = 32'b00000000000000011000110111101100;
assign LUT_3[63385] = 32'b00000000000000011111100011001001;
assign LUT_3[63386] = 32'b00000000000000011010111111010000;
assign LUT_3[63387] = 32'b00000000000000100001101010101101;
assign LUT_3[63388] = 32'b00000000000000010110000101100010;
assign LUT_3[63389] = 32'b00000000000000011100110000111111;
assign LUT_3[63390] = 32'b00000000000000011000001101000110;
assign LUT_3[63391] = 32'b00000000000000011110111000100011;
assign LUT_3[63392] = 32'b00000000000000010001011010000011;
assign LUT_3[63393] = 32'b00000000000000011000000101100000;
assign LUT_3[63394] = 32'b00000000000000010011100001100111;
assign LUT_3[63395] = 32'b00000000000000011010001101000100;
assign LUT_3[63396] = 32'b00000000000000001110100111111001;
assign LUT_3[63397] = 32'b00000000000000010101010011010110;
assign LUT_3[63398] = 32'b00000000000000010000101111011101;
assign LUT_3[63399] = 32'b00000000000000010111011010111010;
assign LUT_3[63400] = 32'b00000000000000010110110011001001;
assign LUT_3[63401] = 32'b00000000000000011101011110100110;
assign LUT_3[63402] = 32'b00000000000000011000111010101101;
assign LUT_3[63403] = 32'b00000000000000011111100110001010;
assign LUT_3[63404] = 32'b00000000000000010100000000111111;
assign LUT_3[63405] = 32'b00000000000000011010101100011100;
assign LUT_3[63406] = 32'b00000000000000010110001000100011;
assign LUT_3[63407] = 32'b00000000000000011100110100000000;
assign LUT_3[63408] = 32'b00000000000000010100101101000110;
assign LUT_3[63409] = 32'b00000000000000011011011000100011;
assign LUT_3[63410] = 32'b00000000000000010110110100101010;
assign LUT_3[63411] = 32'b00000000000000011101100000000111;
assign LUT_3[63412] = 32'b00000000000000010001111010111100;
assign LUT_3[63413] = 32'b00000000000000011000100110011001;
assign LUT_3[63414] = 32'b00000000000000010100000010100000;
assign LUT_3[63415] = 32'b00000000000000011010101101111101;
assign LUT_3[63416] = 32'b00000000000000011010000110001100;
assign LUT_3[63417] = 32'b00000000000000100000110001101001;
assign LUT_3[63418] = 32'b00000000000000011100001101110000;
assign LUT_3[63419] = 32'b00000000000000100010111001001101;
assign LUT_3[63420] = 32'b00000000000000010111010100000010;
assign LUT_3[63421] = 32'b00000000000000011101111111011111;
assign LUT_3[63422] = 32'b00000000000000011001011011100110;
assign LUT_3[63423] = 32'b00000000000000100000000111000011;
assign LUT_3[63424] = 32'b00000000000000010000000100001110;
assign LUT_3[63425] = 32'b00000000000000010110101111101011;
assign LUT_3[63426] = 32'b00000000000000010010001011110010;
assign LUT_3[63427] = 32'b00000000000000011000110111001111;
assign LUT_3[63428] = 32'b00000000000000001101010010000100;
assign LUT_3[63429] = 32'b00000000000000010011111101100001;
assign LUT_3[63430] = 32'b00000000000000001111011001101000;
assign LUT_3[63431] = 32'b00000000000000010110000101000101;
assign LUT_3[63432] = 32'b00000000000000010101011101010100;
assign LUT_3[63433] = 32'b00000000000000011100001000110001;
assign LUT_3[63434] = 32'b00000000000000010111100100111000;
assign LUT_3[63435] = 32'b00000000000000011110010000010101;
assign LUT_3[63436] = 32'b00000000000000010010101011001010;
assign LUT_3[63437] = 32'b00000000000000011001010110100111;
assign LUT_3[63438] = 32'b00000000000000010100110010101110;
assign LUT_3[63439] = 32'b00000000000000011011011110001011;
assign LUT_3[63440] = 32'b00000000000000010011010111010001;
assign LUT_3[63441] = 32'b00000000000000011010000010101110;
assign LUT_3[63442] = 32'b00000000000000010101011110110101;
assign LUT_3[63443] = 32'b00000000000000011100001010010010;
assign LUT_3[63444] = 32'b00000000000000010000100101000111;
assign LUT_3[63445] = 32'b00000000000000010111010000100100;
assign LUT_3[63446] = 32'b00000000000000010010101100101011;
assign LUT_3[63447] = 32'b00000000000000011001011000001000;
assign LUT_3[63448] = 32'b00000000000000011000110000010111;
assign LUT_3[63449] = 32'b00000000000000011111011011110100;
assign LUT_3[63450] = 32'b00000000000000011010110111111011;
assign LUT_3[63451] = 32'b00000000000000100001100011011000;
assign LUT_3[63452] = 32'b00000000000000010101111110001101;
assign LUT_3[63453] = 32'b00000000000000011100101001101010;
assign LUT_3[63454] = 32'b00000000000000011000000101110001;
assign LUT_3[63455] = 32'b00000000000000011110110001001110;
assign LUT_3[63456] = 32'b00000000000000010001010010101110;
assign LUT_3[63457] = 32'b00000000000000010111111110001011;
assign LUT_3[63458] = 32'b00000000000000010011011010010010;
assign LUT_3[63459] = 32'b00000000000000011010000101101111;
assign LUT_3[63460] = 32'b00000000000000001110100000100100;
assign LUT_3[63461] = 32'b00000000000000010101001100000001;
assign LUT_3[63462] = 32'b00000000000000010000101000001000;
assign LUT_3[63463] = 32'b00000000000000010111010011100101;
assign LUT_3[63464] = 32'b00000000000000010110101011110100;
assign LUT_3[63465] = 32'b00000000000000011101010111010001;
assign LUT_3[63466] = 32'b00000000000000011000110011011000;
assign LUT_3[63467] = 32'b00000000000000011111011110110101;
assign LUT_3[63468] = 32'b00000000000000010011111001101010;
assign LUT_3[63469] = 32'b00000000000000011010100101000111;
assign LUT_3[63470] = 32'b00000000000000010110000001001110;
assign LUT_3[63471] = 32'b00000000000000011100101100101011;
assign LUT_3[63472] = 32'b00000000000000010100100101110001;
assign LUT_3[63473] = 32'b00000000000000011011010001001110;
assign LUT_3[63474] = 32'b00000000000000010110101101010101;
assign LUT_3[63475] = 32'b00000000000000011101011000110010;
assign LUT_3[63476] = 32'b00000000000000010001110011100111;
assign LUT_3[63477] = 32'b00000000000000011000011111000100;
assign LUT_3[63478] = 32'b00000000000000010011111011001011;
assign LUT_3[63479] = 32'b00000000000000011010100110101000;
assign LUT_3[63480] = 32'b00000000000000011001111110110111;
assign LUT_3[63481] = 32'b00000000000000100000101010010100;
assign LUT_3[63482] = 32'b00000000000000011100000110011011;
assign LUT_3[63483] = 32'b00000000000000100010110001111000;
assign LUT_3[63484] = 32'b00000000000000010111001100101101;
assign LUT_3[63485] = 32'b00000000000000011101111000001010;
assign LUT_3[63486] = 32'b00000000000000011001010100010001;
assign LUT_3[63487] = 32'b00000000000000011111111111101110;
assign LUT_3[63488] = 32'b00000000000000001001101101001001;
assign LUT_3[63489] = 32'b00000000000000010000011000100110;
assign LUT_3[63490] = 32'b00000000000000001011110100101101;
assign LUT_3[63491] = 32'b00000000000000010010100000001010;
assign LUT_3[63492] = 32'b00000000000000000110111010111111;
assign LUT_3[63493] = 32'b00000000000000001101100110011100;
assign LUT_3[63494] = 32'b00000000000000001001000010100011;
assign LUT_3[63495] = 32'b00000000000000001111101110000000;
assign LUT_3[63496] = 32'b00000000000000001111000110001111;
assign LUT_3[63497] = 32'b00000000000000010101110001101100;
assign LUT_3[63498] = 32'b00000000000000010001001101110011;
assign LUT_3[63499] = 32'b00000000000000010111111001010000;
assign LUT_3[63500] = 32'b00000000000000001100010100000101;
assign LUT_3[63501] = 32'b00000000000000010010111111100010;
assign LUT_3[63502] = 32'b00000000000000001110011011101001;
assign LUT_3[63503] = 32'b00000000000000010101000111000110;
assign LUT_3[63504] = 32'b00000000000000001101000000001100;
assign LUT_3[63505] = 32'b00000000000000010011101011101001;
assign LUT_3[63506] = 32'b00000000000000001111000111110000;
assign LUT_3[63507] = 32'b00000000000000010101110011001101;
assign LUT_3[63508] = 32'b00000000000000001010001110000010;
assign LUT_3[63509] = 32'b00000000000000010000111001011111;
assign LUT_3[63510] = 32'b00000000000000001100010101100110;
assign LUT_3[63511] = 32'b00000000000000010011000001000011;
assign LUT_3[63512] = 32'b00000000000000010010011001010010;
assign LUT_3[63513] = 32'b00000000000000011001000100101111;
assign LUT_3[63514] = 32'b00000000000000010100100000110110;
assign LUT_3[63515] = 32'b00000000000000011011001100010011;
assign LUT_3[63516] = 32'b00000000000000001111100111001000;
assign LUT_3[63517] = 32'b00000000000000010110010010100101;
assign LUT_3[63518] = 32'b00000000000000010001101110101100;
assign LUT_3[63519] = 32'b00000000000000011000011010001001;
assign LUT_3[63520] = 32'b00000000000000001010111011101001;
assign LUT_3[63521] = 32'b00000000000000010001100111000110;
assign LUT_3[63522] = 32'b00000000000000001101000011001101;
assign LUT_3[63523] = 32'b00000000000000010011101110101010;
assign LUT_3[63524] = 32'b00000000000000001000001001011111;
assign LUT_3[63525] = 32'b00000000000000001110110100111100;
assign LUT_3[63526] = 32'b00000000000000001010010001000011;
assign LUT_3[63527] = 32'b00000000000000010000111100100000;
assign LUT_3[63528] = 32'b00000000000000010000010100101111;
assign LUT_3[63529] = 32'b00000000000000010111000000001100;
assign LUT_3[63530] = 32'b00000000000000010010011100010011;
assign LUT_3[63531] = 32'b00000000000000011001000111110000;
assign LUT_3[63532] = 32'b00000000000000001101100010100101;
assign LUT_3[63533] = 32'b00000000000000010100001110000010;
assign LUT_3[63534] = 32'b00000000000000001111101010001001;
assign LUT_3[63535] = 32'b00000000000000010110010101100110;
assign LUT_3[63536] = 32'b00000000000000001110001110101100;
assign LUT_3[63537] = 32'b00000000000000010100111010001001;
assign LUT_3[63538] = 32'b00000000000000010000010110010000;
assign LUT_3[63539] = 32'b00000000000000010111000001101101;
assign LUT_3[63540] = 32'b00000000000000001011011100100010;
assign LUT_3[63541] = 32'b00000000000000010010000111111111;
assign LUT_3[63542] = 32'b00000000000000001101100100000110;
assign LUT_3[63543] = 32'b00000000000000010100001111100011;
assign LUT_3[63544] = 32'b00000000000000010011100111110010;
assign LUT_3[63545] = 32'b00000000000000011010010011001111;
assign LUT_3[63546] = 32'b00000000000000010101101111010110;
assign LUT_3[63547] = 32'b00000000000000011100011010110011;
assign LUT_3[63548] = 32'b00000000000000010000110101101000;
assign LUT_3[63549] = 32'b00000000000000010111100001000101;
assign LUT_3[63550] = 32'b00000000000000010010111101001100;
assign LUT_3[63551] = 32'b00000000000000011001101000101001;
assign LUT_3[63552] = 32'b00000000000000001001100101110100;
assign LUT_3[63553] = 32'b00000000000000010000010001010001;
assign LUT_3[63554] = 32'b00000000000000001011101101011000;
assign LUT_3[63555] = 32'b00000000000000010010011000110101;
assign LUT_3[63556] = 32'b00000000000000000110110011101010;
assign LUT_3[63557] = 32'b00000000000000001101011111000111;
assign LUT_3[63558] = 32'b00000000000000001000111011001110;
assign LUT_3[63559] = 32'b00000000000000001111100110101011;
assign LUT_3[63560] = 32'b00000000000000001110111110111010;
assign LUT_3[63561] = 32'b00000000000000010101101010010111;
assign LUT_3[63562] = 32'b00000000000000010001000110011110;
assign LUT_3[63563] = 32'b00000000000000010111110001111011;
assign LUT_3[63564] = 32'b00000000000000001100001100110000;
assign LUT_3[63565] = 32'b00000000000000010010111000001101;
assign LUT_3[63566] = 32'b00000000000000001110010100010100;
assign LUT_3[63567] = 32'b00000000000000010100111111110001;
assign LUT_3[63568] = 32'b00000000000000001100111000110111;
assign LUT_3[63569] = 32'b00000000000000010011100100010100;
assign LUT_3[63570] = 32'b00000000000000001111000000011011;
assign LUT_3[63571] = 32'b00000000000000010101101011111000;
assign LUT_3[63572] = 32'b00000000000000001010000110101101;
assign LUT_3[63573] = 32'b00000000000000010000110010001010;
assign LUT_3[63574] = 32'b00000000000000001100001110010001;
assign LUT_3[63575] = 32'b00000000000000010010111001101110;
assign LUT_3[63576] = 32'b00000000000000010010010001111101;
assign LUT_3[63577] = 32'b00000000000000011000111101011010;
assign LUT_3[63578] = 32'b00000000000000010100011001100001;
assign LUT_3[63579] = 32'b00000000000000011011000100111110;
assign LUT_3[63580] = 32'b00000000000000001111011111110011;
assign LUT_3[63581] = 32'b00000000000000010110001011010000;
assign LUT_3[63582] = 32'b00000000000000010001100111010111;
assign LUT_3[63583] = 32'b00000000000000011000010010110100;
assign LUT_3[63584] = 32'b00000000000000001010110100010100;
assign LUT_3[63585] = 32'b00000000000000010001011111110001;
assign LUT_3[63586] = 32'b00000000000000001100111011111000;
assign LUT_3[63587] = 32'b00000000000000010011100111010101;
assign LUT_3[63588] = 32'b00000000000000001000000010001010;
assign LUT_3[63589] = 32'b00000000000000001110101101100111;
assign LUT_3[63590] = 32'b00000000000000001010001001101110;
assign LUT_3[63591] = 32'b00000000000000010000110101001011;
assign LUT_3[63592] = 32'b00000000000000010000001101011010;
assign LUT_3[63593] = 32'b00000000000000010110111000110111;
assign LUT_3[63594] = 32'b00000000000000010010010100111110;
assign LUT_3[63595] = 32'b00000000000000011001000000011011;
assign LUT_3[63596] = 32'b00000000000000001101011011010000;
assign LUT_3[63597] = 32'b00000000000000010100000110101101;
assign LUT_3[63598] = 32'b00000000000000001111100010110100;
assign LUT_3[63599] = 32'b00000000000000010110001110010001;
assign LUT_3[63600] = 32'b00000000000000001110000111010111;
assign LUT_3[63601] = 32'b00000000000000010100110010110100;
assign LUT_3[63602] = 32'b00000000000000010000001110111011;
assign LUT_3[63603] = 32'b00000000000000010110111010011000;
assign LUT_3[63604] = 32'b00000000000000001011010101001101;
assign LUT_3[63605] = 32'b00000000000000010010000000101010;
assign LUT_3[63606] = 32'b00000000000000001101011100110001;
assign LUT_3[63607] = 32'b00000000000000010100001000001110;
assign LUT_3[63608] = 32'b00000000000000010011100000011101;
assign LUT_3[63609] = 32'b00000000000000011010001011111010;
assign LUT_3[63610] = 32'b00000000000000010101101000000001;
assign LUT_3[63611] = 32'b00000000000000011100010011011110;
assign LUT_3[63612] = 32'b00000000000000010000101110010011;
assign LUT_3[63613] = 32'b00000000000000010111011001110000;
assign LUT_3[63614] = 32'b00000000000000010010110101110111;
assign LUT_3[63615] = 32'b00000000000000011001100001010100;
assign LUT_3[63616] = 32'b00000000000000001011111000000111;
assign LUT_3[63617] = 32'b00000000000000010010100011100100;
assign LUT_3[63618] = 32'b00000000000000001101111111101011;
assign LUT_3[63619] = 32'b00000000000000010100101011001000;
assign LUT_3[63620] = 32'b00000000000000001001000101111101;
assign LUT_3[63621] = 32'b00000000000000001111110001011010;
assign LUT_3[63622] = 32'b00000000000000001011001101100001;
assign LUT_3[63623] = 32'b00000000000000010001111000111110;
assign LUT_3[63624] = 32'b00000000000000010001010001001101;
assign LUT_3[63625] = 32'b00000000000000010111111100101010;
assign LUT_3[63626] = 32'b00000000000000010011011000110001;
assign LUT_3[63627] = 32'b00000000000000011010000100001110;
assign LUT_3[63628] = 32'b00000000000000001110011111000011;
assign LUT_3[63629] = 32'b00000000000000010101001010100000;
assign LUT_3[63630] = 32'b00000000000000010000100110100111;
assign LUT_3[63631] = 32'b00000000000000010111010010000100;
assign LUT_3[63632] = 32'b00000000000000001111001011001010;
assign LUT_3[63633] = 32'b00000000000000010101110110100111;
assign LUT_3[63634] = 32'b00000000000000010001010010101110;
assign LUT_3[63635] = 32'b00000000000000010111111110001011;
assign LUT_3[63636] = 32'b00000000000000001100011001000000;
assign LUT_3[63637] = 32'b00000000000000010011000100011101;
assign LUT_3[63638] = 32'b00000000000000001110100000100100;
assign LUT_3[63639] = 32'b00000000000000010101001100000001;
assign LUT_3[63640] = 32'b00000000000000010100100100010000;
assign LUT_3[63641] = 32'b00000000000000011011001111101101;
assign LUT_3[63642] = 32'b00000000000000010110101011110100;
assign LUT_3[63643] = 32'b00000000000000011101010111010001;
assign LUT_3[63644] = 32'b00000000000000010001110010000110;
assign LUT_3[63645] = 32'b00000000000000011000011101100011;
assign LUT_3[63646] = 32'b00000000000000010011111001101010;
assign LUT_3[63647] = 32'b00000000000000011010100101000111;
assign LUT_3[63648] = 32'b00000000000000001101000110100111;
assign LUT_3[63649] = 32'b00000000000000010011110010000100;
assign LUT_3[63650] = 32'b00000000000000001111001110001011;
assign LUT_3[63651] = 32'b00000000000000010101111001101000;
assign LUT_3[63652] = 32'b00000000000000001010010100011101;
assign LUT_3[63653] = 32'b00000000000000010000111111111010;
assign LUT_3[63654] = 32'b00000000000000001100011100000001;
assign LUT_3[63655] = 32'b00000000000000010011000111011110;
assign LUT_3[63656] = 32'b00000000000000010010011111101101;
assign LUT_3[63657] = 32'b00000000000000011001001011001010;
assign LUT_3[63658] = 32'b00000000000000010100100111010001;
assign LUT_3[63659] = 32'b00000000000000011011010010101110;
assign LUT_3[63660] = 32'b00000000000000001111101101100011;
assign LUT_3[63661] = 32'b00000000000000010110011001000000;
assign LUT_3[63662] = 32'b00000000000000010001110101000111;
assign LUT_3[63663] = 32'b00000000000000011000100000100100;
assign LUT_3[63664] = 32'b00000000000000010000011001101010;
assign LUT_3[63665] = 32'b00000000000000010111000101000111;
assign LUT_3[63666] = 32'b00000000000000010010100001001110;
assign LUT_3[63667] = 32'b00000000000000011001001100101011;
assign LUT_3[63668] = 32'b00000000000000001101100111100000;
assign LUT_3[63669] = 32'b00000000000000010100010010111101;
assign LUT_3[63670] = 32'b00000000000000001111101111000100;
assign LUT_3[63671] = 32'b00000000000000010110011010100001;
assign LUT_3[63672] = 32'b00000000000000010101110010110000;
assign LUT_3[63673] = 32'b00000000000000011100011110001101;
assign LUT_3[63674] = 32'b00000000000000010111111010010100;
assign LUT_3[63675] = 32'b00000000000000011110100101110001;
assign LUT_3[63676] = 32'b00000000000000010011000000100110;
assign LUT_3[63677] = 32'b00000000000000011001101100000011;
assign LUT_3[63678] = 32'b00000000000000010101001000001010;
assign LUT_3[63679] = 32'b00000000000000011011110011100111;
assign LUT_3[63680] = 32'b00000000000000001011110000110010;
assign LUT_3[63681] = 32'b00000000000000010010011100001111;
assign LUT_3[63682] = 32'b00000000000000001101111000010110;
assign LUT_3[63683] = 32'b00000000000000010100100011110011;
assign LUT_3[63684] = 32'b00000000000000001000111110101000;
assign LUT_3[63685] = 32'b00000000000000001111101010000101;
assign LUT_3[63686] = 32'b00000000000000001011000110001100;
assign LUT_3[63687] = 32'b00000000000000010001110001101001;
assign LUT_3[63688] = 32'b00000000000000010001001001111000;
assign LUT_3[63689] = 32'b00000000000000010111110101010101;
assign LUT_3[63690] = 32'b00000000000000010011010001011100;
assign LUT_3[63691] = 32'b00000000000000011001111100111001;
assign LUT_3[63692] = 32'b00000000000000001110010111101110;
assign LUT_3[63693] = 32'b00000000000000010101000011001011;
assign LUT_3[63694] = 32'b00000000000000010000011111010010;
assign LUT_3[63695] = 32'b00000000000000010111001010101111;
assign LUT_3[63696] = 32'b00000000000000001111000011110101;
assign LUT_3[63697] = 32'b00000000000000010101101111010010;
assign LUT_3[63698] = 32'b00000000000000010001001011011001;
assign LUT_3[63699] = 32'b00000000000000010111110110110110;
assign LUT_3[63700] = 32'b00000000000000001100010001101011;
assign LUT_3[63701] = 32'b00000000000000010010111101001000;
assign LUT_3[63702] = 32'b00000000000000001110011001001111;
assign LUT_3[63703] = 32'b00000000000000010101000100101100;
assign LUT_3[63704] = 32'b00000000000000010100011100111011;
assign LUT_3[63705] = 32'b00000000000000011011001000011000;
assign LUT_3[63706] = 32'b00000000000000010110100100011111;
assign LUT_3[63707] = 32'b00000000000000011101001111111100;
assign LUT_3[63708] = 32'b00000000000000010001101010110001;
assign LUT_3[63709] = 32'b00000000000000011000010110001110;
assign LUT_3[63710] = 32'b00000000000000010011110010010101;
assign LUT_3[63711] = 32'b00000000000000011010011101110010;
assign LUT_3[63712] = 32'b00000000000000001100111111010010;
assign LUT_3[63713] = 32'b00000000000000010011101010101111;
assign LUT_3[63714] = 32'b00000000000000001111000110110110;
assign LUT_3[63715] = 32'b00000000000000010101110010010011;
assign LUT_3[63716] = 32'b00000000000000001010001101001000;
assign LUT_3[63717] = 32'b00000000000000010000111000100101;
assign LUT_3[63718] = 32'b00000000000000001100010100101100;
assign LUT_3[63719] = 32'b00000000000000010011000000001001;
assign LUT_3[63720] = 32'b00000000000000010010011000011000;
assign LUT_3[63721] = 32'b00000000000000011001000011110101;
assign LUT_3[63722] = 32'b00000000000000010100011111111100;
assign LUT_3[63723] = 32'b00000000000000011011001011011001;
assign LUT_3[63724] = 32'b00000000000000001111100110001110;
assign LUT_3[63725] = 32'b00000000000000010110010001101011;
assign LUT_3[63726] = 32'b00000000000000010001101101110010;
assign LUT_3[63727] = 32'b00000000000000011000011001001111;
assign LUT_3[63728] = 32'b00000000000000010000010010010101;
assign LUT_3[63729] = 32'b00000000000000010110111101110010;
assign LUT_3[63730] = 32'b00000000000000010010011001111001;
assign LUT_3[63731] = 32'b00000000000000011001000101010110;
assign LUT_3[63732] = 32'b00000000000000001101100000001011;
assign LUT_3[63733] = 32'b00000000000000010100001011101000;
assign LUT_3[63734] = 32'b00000000000000001111100111101111;
assign LUT_3[63735] = 32'b00000000000000010110010011001100;
assign LUT_3[63736] = 32'b00000000000000010101101011011011;
assign LUT_3[63737] = 32'b00000000000000011100010110111000;
assign LUT_3[63738] = 32'b00000000000000010111110010111111;
assign LUT_3[63739] = 32'b00000000000000011110011110011100;
assign LUT_3[63740] = 32'b00000000000000010010111001010001;
assign LUT_3[63741] = 32'b00000000000000011001100100101110;
assign LUT_3[63742] = 32'b00000000000000010101000000110101;
assign LUT_3[63743] = 32'b00000000000000011011101100010010;
assign LUT_3[63744] = 32'b00000000000000000101111100101010;
assign LUT_3[63745] = 32'b00000000000000001100101000000111;
assign LUT_3[63746] = 32'b00000000000000001000000100001110;
assign LUT_3[63747] = 32'b00000000000000001110101111101011;
assign LUT_3[63748] = 32'b00000000000000000011001010100000;
assign LUT_3[63749] = 32'b00000000000000001001110101111101;
assign LUT_3[63750] = 32'b00000000000000000101010010000100;
assign LUT_3[63751] = 32'b00000000000000001011111101100001;
assign LUT_3[63752] = 32'b00000000000000001011010101110000;
assign LUT_3[63753] = 32'b00000000000000010010000001001101;
assign LUT_3[63754] = 32'b00000000000000001101011101010100;
assign LUT_3[63755] = 32'b00000000000000010100001000110001;
assign LUT_3[63756] = 32'b00000000000000001000100011100110;
assign LUT_3[63757] = 32'b00000000000000001111001111000011;
assign LUT_3[63758] = 32'b00000000000000001010101011001010;
assign LUT_3[63759] = 32'b00000000000000010001010110100111;
assign LUT_3[63760] = 32'b00000000000000001001001111101101;
assign LUT_3[63761] = 32'b00000000000000001111111011001010;
assign LUT_3[63762] = 32'b00000000000000001011010111010001;
assign LUT_3[63763] = 32'b00000000000000010010000010101110;
assign LUT_3[63764] = 32'b00000000000000000110011101100011;
assign LUT_3[63765] = 32'b00000000000000001101001001000000;
assign LUT_3[63766] = 32'b00000000000000001000100101000111;
assign LUT_3[63767] = 32'b00000000000000001111010000100100;
assign LUT_3[63768] = 32'b00000000000000001110101000110011;
assign LUT_3[63769] = 32'b00000000000000010101010100010000;
assign LUT_3[63770] = 32'b00000000000000010000110000010111;
assign LUT_3[63771] = 32'b00000000000000010111011011110100;
assign LUT_3[63772] = 32'b00000000000000001011110110101001;
assign LUT_3[63773] = 32'b00000000000000010010100010000110;
assign LUT_3[63774] = 32'b00000000000000001101111110001101;
assign LUT_3[63775] = 32'b00000000000000010100101001101010;
assign LUT_3[63776] = 32'b00000000000000000111001011001010;
assign LUT_3[63777] = 32'b00000000000000001101110110100111;
assign LUT_3[63778] = 32'b00000000000000001001010010101110;
assign LUT_3[63779] = 32'b00000000000000001111111110001011;
assign LUT_3[63780] = 32'b00000000000000000100011001000000;
assign LUT_3[63781] = 32'b00000000000000001011000100011101;
assign LUT_3[63782] = 32'b00000000000000000110100000100100;
assign LUT_3[63783] = 32'b00000000000000001101001100000001;
assign LUT_3[63784] = 32'b00000000000000001100100100010000;
assign LUT_3[63785] = 32'b00000000000000010011001111101101;
assign LUT_3[63786] = 32'b00000000000000001110101011110100;
assign LUT_3[63787] = 32'b00000000000000010101010111010001;
assign LUT_3[63788] = 32'b00000000000000001001110010000110;
assign LUT_3[63789] = 32'b00000000000000010000011101100011;
assign LUT_3[63790] = 32'b00000000000000001011111001101010;
assign LUT_3[63791] = 32'b00000000000000010010100101000111;
assign LUT_3[63792] = 32'b00000000000000001010011110001101;
assign LUT_3[63793] = 32'b00000000000000010001001001101010;
assign LUT_3[63794] = 32'b00000000000000001100100101110001;
assign LUT_3[63795] = 32'b00000000000000010011010001001110;
assign LUT_3[63796] = 32'b00000000000000000111101100000011;
assign LUT_3[63797] = 32'b00000000000000001110010111100000;
assign LUT_3[63798] = 32'b00000000000000001001110011100111;
assign LUT_3[63799] = 32'b00000000000000010000011111000100;
assign LUT_3[63800] = 32'b00000000000000001111110111010011;
assign LUT_3[63801] = 32'b00000000000000010110100010110000;
assign LUT_3[63802] = 32'b00000000000000010001111110110111;
assign LUT_3[63803] = 32'b00000000000000011000101010010100;
assign LUT_3[63804] = 32'b00000000000000001101000101001001;
assign LUT_3[63805] = 32'b00000000000000010011110000100110;
assign LUT_3[63806] = 32'b00000000000000001111001100101101;
assign LUT_3[63807] = 32'b00000000000000010101111000001010;
assign LUT_3[63808] = 32'b00000000000000000101110101010101;
assign LUT_3[63809] = 32'b00000000000000001100100000110010;
assign LUT_3[63810] = 32'b00000000000000000111111100111001;
assign LUT_3[63811] = 32'b00000000000000001110101000010110;
assign LUT_3[63812] = 32'b00000000000000000011000011001011;
assign LUT_3[63813] = 32'b00000000000000001001101110101000;
assign LUT_3[63814] = 32'b00000000000000000101001010101111;
assign LUT_3[63815] = 32'b00000000000000001011110110001100;
assign LUT_3[63816] = 32'b00000000000000001011001110011011;
assign LUT_3[63817] = 32'b00000000000000010001111001111000;
assign LUT_3[63818] = 32'b00000000000000001101010101111111;
assign LUT_3[63819] = 32'b00000000000000010100000001011100;
assign LUT_3[63820] = 32'b00000000000000001000011100010001;
assign LUT_3[63821] = 32'b00000000000000001111000111101110;
assign LUT_3[63822] = 32'b00000000000000001010100011110101;
assign LUT_3[63823] = 32'b00000000000000010001001111010010;
assign LUT_3[63824] = 32'b00000000000000001001001000011000;
assign LUT_3[63825] = 32'b00000000000000001111110011110101;
assign LUT_3[63826] = 32'b00000000000000001011001111111100;
assign LUT_3[63827] = 32'b00000000000000010001111011011001;
assign LUT_3[63828] = 32'b00000000000000000110010110001110;
assign LUT_3[63829] = 32'b00000000000000001101000001101011;
assign LUT_3[63830] = 32'b00000000000000001000011101110010;
assign LUT_3[63831] = 32'b00000000000000001111001001001111;
assign LUT_3[63832] = 32'b00000000000000001110100001011110;
assign LUT_3[63833] = 32'b00000000000000010101001100111011;
assign LUT_3[63834] = 32'b00000000000000010000101001000010;
assign LUT_3[63835] = 32'b00000000000000010111010100011111;
assign LUT_3[63836] = 32'b00000000000000001011101111010100;
assign LUT_3[63837] = 32'b00000000000000010010011010110001;
assign LUT_3[63838] = 32'b00000000000000001101110110111000;
assign LUT_3[63839] = 32'b00000000000000010100100010010101;
assign LUT_3[63840] = 32'b00000000000000000111000011110101;
assign LUT_3[63841] = 32'b00000000000000001101101111010010;
assign LUT_3[63842] = 32'b00000000000000001001001011011001;
assign LUT_3[63843] = 32'b00000000000000001111110110110110;
assign LUT_3[63844] = 32'b00000000000000000100010001101011;
assign LUT_3[63845] = 32'b00000000000000001010111101001000;
assign LUT_3[63846] = 32'b00000000000000000110011001001111;
assign LUT_3[63847] = 32'b00000000000000001101000100101100;
assign LUT_3[63848] = 32'b00000000000000001100011100111011;
assign LUT_3[63849] = 32'b00000000000000010011001000011000;
assign LUT_3[63850] = 32'b00000000000000001110100100011111;
assign LUT_3[63851] = 32'b00000000000000010101001111111100;
assign LUT_3[63852] = 32'b00000000000000001001101010110001;
assign LUT_3[63853] = 32'b00000000000000010000010110001110;
assign LUT_3[63854] = 32'b00000000000000001011110010010101;
assign LUT_3[63855] = 32'b00000000000000010010011101110010;
assign LUT_3[63856] = 32'b00000000000000001010010110111000;
assign LUT_3[63857] = 32'b00000000000000010001000010010101;
assign LUT_3[63858] = 32'b00000000000000001100011110011100;
assign LUT_3[63859] = 32'b00000000000000010011001001111001;
assign LUT_3[63860] = 32'b00000000000000000111100100101110;
assign LUT_3[63861] = 32'b00000000000000001110010000001011;
assign LUT_3[63862] = 32'b00000000000000001001101100010010;
assign LUT_3[63863] = 32'b00000000000000010000010111101111;
assign LUT_3[63864] = 32'b00000000000000001111101111111110;
assign LUT_3[63865] = 32'b00000000000000010110011011011011;
assign LUT_3[63866] = 32'b00000000000000010001110111100010;
assign LUT_3[63867] = 32'b00000000000000011000100010111111;
assign LUT_3[63868] = 32'b00000000000000001100111101110100;
assign LUT_3[63869] = 32'b00000000000000010011101001010001;
assign LUT_3[63870] = 32'b00000000000000001111000101011000;
assign LUT_3[63871] = 32'b00000000000000010101110000110101;
assign LUT_3[63872] = 32'b00000000000000001000000111101000;
assign LUT_3[63873] = 32'b00000000000000001110110011000101;
assign LUT_3[63874] = 32'b00000000000000001010001111001100;
assign LUT_3[63875] = 32'b00000000000000010000111010101001;
assign LUT_3[63876] = 32'b00000000000000000101010101011110;
assign LUT_3[63877] = 32'b00000000000000001100000000111011;
assign LUT_3[63878] = 32'b00000000000000000111011101000010;
assign LUT_3[63879] = 32'b00000000000000001110001000011111;
assign LUT_3[63880] = 32'b00000000000000001101100000101110;
assign LUT_3[63881] = 32'b00000000000000010100001100001011;
assign LUT_3[63882] = 32'b00000000000000001111101000010010;
assign LUT_3[63883] = 32'b00000000000000010110010011101111;
assign LUT_3[63884] = 32'b00000000000000001010101110100100;
assign LUT_3[63885] = 32'b00000000000000010001011010000001;
assign LUT_3[63886] = 32'b00000000000000001100110110001000;
assign LUT_3[63887] = 32'b00000000000000010011100001100101;
assign LUT_3[63888] = 32'b00000000000000001011011010101011;
assign LUT_3[63889] = 32'b00000000000000010010000110001000;
assign LUT_3[63890] = 32'b00000000000000001101100010001111;
assign LUT_3[63891] = 32'b00000000000000010100001101101100;
assign LUT_3[63892] = 32'b00000000000000001000101000100001;
assign LUT_3[63893] = 32'b00000000000000001111010011111110;
assign LUT_3[63894] = 32'b00000000000000001010110000000101;
assign LUT_3[63895] = 32'b00000000000000010001011011100010;
assign LUT_3[63896] = 32'b00000000000000010000110011110001;
assign LUT_3[63897] = 32'b00000000000000010111011111001110;
assign LUT_3[63898] = 32'b00000000000000010010111011010101;
assign LUT_3[63899] = 32'b00000000000000011001100110110010;
assign LUT_3[63900] = 32'b00000000000000001110000001100111;
assign LUT_3[63901] = 32'b00000000000000010100101101000100;
assign LUT_3[63902] = 32'b00000000000000010000001001001011;
assign LUT_3[63903] = 32'b00000000000000010110110100101000;
assign LUT_3[63904] = 32'b00000000000000001001010110001000;
assign LUT_3[63905] = 32'b00000000000000010000000001100101;
assign LUT_3[63906] = 32'b00000000000000001011011101101100;
assign LUT_3[63907] = 32'b00000000000000010010001001001001;
assign LUT_3[63908] = 32'b00000000000000000110100011111110;
assign LUT_3[63909] = 32'b00000000000000001101001111011011;
assign LUT_3[63910] = 32'b00000000000000001000101011100010;
assign LUT_3[63911] = 32'b00000000000000001111010110111111;
assign LUT_3[63912] = 32'b00000000000000001110101111001110;
assign LUT_3[63913] = 32'b00000000000000010101011010101011;
assign LUT_3[63914] = 32'b00000000000000010000110110110010;
assign LUT_3[63915] = 32'b00000000000000010111100010001111;
assign LUT_3[63916] = 32'b00000000000000001011111101000100;
assign LUT_3[63917] = 32'b00000000000000010010101000100001;
assign LUT_3[63918] = 32'b00000000000000001110000100101000;
assign LUT_3[63919] = 32'b00000000000000010100110000000101;
assign LUT_3[63920] = 32'b00000000000000001100101001001011;
assign LUT_3[63921] = 32'b00000000000000010011010100101000;
assign LUT_3[63922] = 32'b00000000000000001110110000101111;
assign LUT_3[63923] = 32'b00000000000000010101011100001100;
assign LUT_3[63924] = 32'b00000000000000001001110111000001;
assign LUT_3[63925] = 32'b00000000000000010000100010011110;
assign LUT_3[63926] = 32'b00000000000000001011111110100101;
assign LUT_3[63927] = 32'b00000000000000010010101010000010;
assign LUT_3[63928] = 32'b00000000000000010010000010010001;
assign LUT_3[63929] = 32'b00000000000000011000101101101110;
assign LUT_3[63930] = 32'b00000000000000010100001001110101;
assign LUT_3[63931] = 32'b00000000000000011010110101010010;
assign LUT_3[63932] = 32'b00000000000000001111010000000111;
assign LUT_3[63933] = 32'b00000000000000010101111011100100;
assign LUT_3[63934] = 32'b00000000000000010001010111101011;
assign LUT_3[63935] = 32'b00000000000000011000000011001000;
assign LUT_3[63936] = 32'b00000000000000001000000000010011;
assign LUT_3[63937] = 32'b00000000000000001110101011110000;
assign LUT_3[63938] = 32'b00000000000000001010000111110111;
assign LUT_3[63939] = 32'b00000000000000010000110011010100;
assign LUT_3[63940] = 32'b00000000000000000101001110001001;
assign LUT_3[63941] = 32'b00000000000000001011111001100110;
assign LUT_3[63942] = 32'b00000000000000000111010101101101;
assign LUT_3[63943] = 32'b00000000000000001110000001001010;
assign LUT_3[63944] = 32'b00000000000000001101011001011001;
assign LUT_3[63945] = 32'b00000000000000010100000100110110;
assign LUT_3[63946] = 32'b00000000000000001111100000111101;
assign LUT_3[63947] = 32'b00000000000000010110001100011010;
assign LUT_3[63948] = 32'b00000000000000001010100111001111;
assign LUT_3[63949] = 32'b00000000000000010001010010101100;
assign LUT_3[63950] = 32'b00000000000000001100101110110011;
assign LUT_3[63951] = 32'b00000000000000010011011010010000;
assign LUT_3[63952] = 32'b00000000000000001011010011010110;
assign LUT_3[63953] = 32'b00000000000000010001111110110011;
assign LUT_3[63954] = 32'b00000000000000001101011010111010;
assign LUT_3[63955] = 32'b00000000000000010100000110010111;
assign LUT_3[63956] = 32'b00000000000000001000100001001100;
assign LUT_3[63957] = 32'b00000000000000001111001100101001;
assign LUT_3[63958] = 32'b00000000000000001010101000110000;
assign LUT_3[63959] = 32'b00000000000000010001010100001101;
assign LUT_3[63960] = 32'b00000000000000010000101100011100;
assign LUT_3[63961] = 32'b00000000000000010111010111111001;
assign LUT_3[63962] = 32'b00000000000000010010110100000000;
assign LUT_3[63963] = 32'b00000000000000011001011111011101;
assign LUT_3[63964] = 32'b00000000000000001101111010010010;
assign LUT_3[63965] = 32'b00000000000000010100100101101111;
assign LUT_3[63966] = 32'b00000000000000010000000001110110;
assign LUT_3[63967] = 32'b00000000000000010110101101010011;
assign LUT_3[63968] = 32'b00000000000000001001001110110011;
assign LUT_3[63969] = 32'b00000000000000001111111010010000;
assign LUT_3[63970] = 32'b00000000000000001011010110010111;
assign LUT_3[63971] = 32'b00000000000000010010000001110100;
assign LUT_3[63972] = 32'b00000000000000000110011100101001;
assign LUT_3[63973] = 32'b00000000000000001101001000000110;
assign LUT_3[63974] = 32'b00000000000000001000100100001101;
assign LUT_3[63975] = 32'b00000000000000001111001111101010;
assign LUT_3[63976] = 32'b00000000000000001110100111111001;
assign LUT_3[63977] = 32'b00000000000000010101010011010110;
assign LUT_3[63978] = 32'b00000000000000010000101111011101;
assign LUT_3[63979] = 32'b00000000000000010111011010111010;
assign LUT_3[63980] = 32'b00000000000000001011110101101111;
assign LUT_3[63981] = 32'b00000000000000010010100001001100;
assign LUT_3[63982] = 32'b00000000000000001101111101010011;
assign LUT_3[63983] = 32'b00000000000000010100101000110000;
assign LUT_3[63984] = 32'b00000000000000001100100001110110;
assign LUT_3[63985] = 32'b00000000000000010011001101010011;
assign LUT_3[63986] = 32'b00000000000000001110101001011010;
assign LUT_3[63987] = 32'b00000000000000010101010100110111;
assign LUT_3[63988] = 32'b00000000000000001001101111101100;
assign LUT_3[63989] = 32'b00000000000000010000011011001001;
assign LUT_3[63990] = 32'b00000000000000001011110111010000;
assign LUT_3[63991] = 32'b00000000000000010010100010101101;
assign LUT_3[63992] = 32'b00000000000000010001111010111100;
assign LUT_3[63993] = 32'b00000000000000011000100110011001;
assign LUT_3[63994] = 32'b00000000000000010100000010100000;
assign LUT_3[63995] = 32'b00000000000000011010101101111101;
assign LUT_3[63996] = 32'b00000000000000001111001000110010;
assign LUT_3[63997] = 32'b00000000000000010101110100001111;
assign LUT_3[63998] = 32'b00000000000000010001010000010110;
assign LUT_3[63999] = 32'b00000000000000010111111011110011;
assign LUT_3[64000] = 32'b00000000000000001101000010010101;
assign LUT_3[64001] = 32'b00000000000000010011101101110010;
assign LUT_3[64002] = 32'b00000000000000001111001001111001;
assign LUT_3[64003] = 32'b00000000000000010101110101010110;
assign LUT_3[64004] = 32'b00000000000000001010010000001011;
assign LUT_3[64005] = 32'b00000000000000010000111011101000;
assign LUT_3[64006] = 32'b00000000000000001100010111101111;
assign LUT_3[64007] = 32'b00000000000000010011000011001100;
assign LUT_3[64008] = 32'b00000000000000010010011011011011;
assign LUT_3[64009] = 32'b00000000000000011001000110111000;
assign LUT_3[64010] = 32'b00000000000000010100100010111111;
assign LUT_3[64011] = 32'b00000000000000011011001110011100;
assign LUT_3[64012] = 32'b00000000000000001111101001010001;
assign LUT_3[64013] = 32'b00000000000000010110010100101110;
assign LUT_3[64014] = 32'b00000000000000010001110000110101;
assign LUT_3[64015] = 32'b00000000000000011000011100010010;
assign LUT_3[64016] = 32'b00000000000000010000010101011000;
assign LUT_3[64017] = 32'b00000000000000010111000000110101;
assign LUT_3[64018] = 32'b00000000000000010010011100111100;
assign LUT_3[64019] = 32'b00000000000000011001001000011001;
assign LUT_3[64020] = 32'b00000000000000001101100011001110;
assign LUT_3[64021] = 32'b00000000000000010100001110101011;
assign LUT_3[64022] = 32'b00000000000000001111101010110010;
assign LUT_3[64023] = 32'b00000000000000010110010110001111;
assign LUT_3[64024] = 32'b00000000000000010101101110011110;
assign LUT_3[64025] = 32'b00000000000000011100011001111011;
assign LUT_3[64026] = 32'b00000000000000010111110110000010;
assign LUT_3[64027] = 32'b00000000000000011110100001011111;
assign LUT_3[64028] = 32'b00000000000000010010111100010100;
assign LUT_3[64029] = 32'b00000000000000011001100111110001;
assign LUT_3[64030] = 32'b00000000000000010101000011111000;
assign LUT_3[64031] = 32'b00000000000000011011101111010101;
assign LUT_3[64032] = 32'b00000000000000001110010000110101;
assign LUT_3[64033] = 32'b00000000000000010100111100010010;
assign LUT_3[64034] = 32'b00000000000000010000011000011001;
assign LUT_3[64035] = 32'b00000000000000010111000011110110;
assign LUT_3[64036] = 32'b00000000000000001011011110101011;
assign LUT_3[64037] = 32'b00000000000000010010001010001000;
assign LUT_3[64038] = 32'b00000000000000001101100110001111;
assign LUT_3[64039] = 32'b00000000000000010100010001101100;
assign LUT_3[64040] = 32'b00000000000000010011101001111011;
assign LUT_3[64041] = 32'b00000000000000011010010101011000;
assign LUT_3[64042] = 32'b00000000000000010101110001011111;
assign LUT_3[64043] = 32'b00000000000000011100011100111100;
assign LUT_3[64044] = 32'b00000000000000010000110111110001;
assign LUT_3[64045] = 32'b00000000000000010111100011001110;
assign LUT_3[64046] = 32'b00000000000000010010111111010101;
assign LUT_3[64047] = 32'b00000000000000011001101010110010;
assign LUT_3[64048] = 32'b00000000000000010001100011111000;
assign LUT_3[64049] = 32'b00000000000000011000001111010101;
assign LUT_3[64050] = 32'b00000000000000010011101011011100;
assign LUT_3[64051] = 32'b00000000000000011010010110111001;
assign LUT_3[64052] = 32'b00000000000000001110110001101110;
assign LUT_3[64053] = 32'b00000000000000010101011101001011;
assign LUT_3[64054] = 32'b00000000000000010000111001010010;
assign LUT_3[64055] = 32'b00000000000000010111100100101111;
assign LUT_3[64056] = 32'b00000000000000010110111100111110;
assign LUT_3[64057] = 32'b00000000000000011101101000011011;
assign LUT_3[64058] = 32'b00000000000000011001000100100010;
assign LUT_3[64059] = 32'b00000000000000011111101111111111;
assign LUT_3[64060] = 32'b00000000000000010100001010110100;
assign LUT_3[64061] = 32'b00000000000000011010110110010001;
assign LUT_3[64062] = 32'b00000000000000010110010010011000;
assign LUT_3[64063] = 32'b00000000000000011100111101110101;
assign LUT_3[64064] = 32'b00000000000000001100111011000000;
assign LUT_3[64065] = 32'b00000000000000010011100110011101;
assign LUT_3[64066] = 32'b00000000000000001111000010100100;
assign LUT_3[64067] = 32'b00000000000000010101101110000001;
assign LUT_3[64068] = 32'b00000000000000001010001000110110;
assign LUT_3[64069] = 32'b00000000000000010000110100010011;
assign LUT_3[64070] = 32'b00000000000000001100010000011010;
assign LUT_3[64071] = 32'b00000000000000010010111011110111;
assign LUT_3[64072] = 32'b00000000000000010010010100000110;
assign LUT_3[64073] = 32'b00000000000000011000111111100011;
assign LUT_3[64074] = 32'b00000000000000010100011011101010;
assign LUT_3[64075] = 32'b00000000000000011011000111000111;
assign LUT_3[64076] = 32'b00000000000000001111100001111100;
assign LUT_3[64077] = 32'b00000000000000010110001101011001;
assign LUT_3[64078] = 32'b00000000000000010001101001100000;
assign LUT_3[64079] = 32'b00000000000000011000010100111101;
assign LUT_3[64080] = 32'b00000000000000010000001110000011;
assign LUT_3[64081] = 32'b00000000000000010110111001100000;
assign LUT_3[64082] = 32'b00000000000000010010010101100111;
assign LUT_3[64083] = 32'b00000000000000011001000001000100;
assign LUT_3[64084] = 32'b00000000000000001101011011111001;
assign LUT_3[64085] = 32'b00000000000000010100000111010110;
assign LUT_3[64086] = 32'b00000000000000001111100011011101;
assign LUT_3[64087] = 32'b00000000000000010110001110111010;
assign LUT_3[64088] = 32'b00000000000000010101100111001001;
assign LUT_3[64089] = 32'b00000000000000011100010010100110;
assign LUT_3[64090] = 32'b00000000000000010111101110101101;
assign LUT_3[64091] = 32'b00000000000000011110011010001010;
assign LUT_3[64092] = 32'b00000000000000010010110100111111;
assign LUT_3[64093] = 32'b00000000000000011001100000011100;
assign LUT_3[64094] = 32'b00000000000000010100111100100011;
assign LUT_3[64095] = 32'b00000000000000011011101000000000;
assign LUT_3[64096] = 32'b00000000000000001110001001100000;
assign LUT_3[64097] = 32'b00000000000000010100110100111101;
assign LUT_3[64098] = 32'b00000000000000010000010001000100;
assign LUT_3[64099] = 32'b00000000000000010110111100100001;
assign LUT_3[64100] = 32'b00000000000000001011010111010110;
assign LUT_3[64101] = 32'b00000000000000010010000010110011;
assign LUT_3[64102] = 32'b00000000000000001101011110111010;
assign LUT_3[64103] = 32'b00000000000000010100001010010111;
assign LUT_3[64104] = 32'b00000000000000010011100010100110;
assign LUT_3[64105] = 32'b00000000000000011010001110000011;
assign LUT_3[64106] = 32'b00000000000000010101101010001010;
assign LUT_3[64107] = 32'b00000000000000011100010101100111;
assign LUT_3[64108] = 32'b00000000000000010000110000011100;
assign LUT_3[64109] = 32'b00000000000000010111011011111001;
assign LUT_3[64110] = 32'b00000000000000010010111000000000;
assign LUT_3[64111] = 32'b00000000000000011001100011011101;
assign LUT_3[64112] = 32'b00000000000000010001011100100011;
assign LUT_3[64113] = 32'b00000000000000011000001000000000;
assign LUT_3[64114] = 32'b00000000000000010011100100000111;
assign LUT_3[64115] = 32'b00000000000000011010001111100100;
assign LUT_3[64116] = 32'b00000000000000001110101010011001;
assign LUT_3[64117] = 32'b00000000000000010101010101110110;
assign LUT_3[64118] = 32'b00000000000000010000110001111101;
assign LUT_3[64119] = 32'b00000000000000010111011101011010;
assign LUT_3[64120] = 32'b00000000000000010110110101101001;
assign LUT_3[64121] = 32'b00000000000000011101100001000110;
assign LUT_3[64122] = 32'b00000000000000011000111101001101;
assign LUT_3[64123] = 32'b00000000000000011111101000101010;
assign LUT_3[64124] = 32'b00000000000000010100000011011111;
assign LUT_3[64125] = 32'b00000000000000011010101110111100;
assign LUT_3[64126] = 32'b00000000000000010110001011000011;
assign LUT_3[64127] = 32'b00000000000000011100110110100000;
assign LUT_3[64128] = 32'b00000000000000001111001101010011;
assign LUT_3[64129] = 32'b00000000000000010101111000110000;
assign LUT_3[64130] = 32'b00000000000000010001010100110111;
assign LUT_3[64131] = 32'b00000000000000011000000000010100;
assign LUT_3[64132] = 32'b00000000000000001100011011001001;
assign LUT_3[64133] = 32'b00000000000000010011000110100110;
assign LUT_3[64134] = 32'b00000000000000001110100010101101;
assign LUT_3[64135] = 32'b00000000000000010101001110001010;
assign LUT_3[64136] = 32'b00000000000000010100100110011001;
assign LUT_3[64137] = 32'b00000000000000011011010001110110;
assign LUT_3[64138] = 32'b00000000000000010110101101111101;
assign LUT_3[64139] = 32'b00000000000000011101011001011010;
assign LUT_3[64140] = 32'b00000000000000010001110100001111;
assign LUT_3[64141] = 32'b00000000000000011000011111101100;
assign LUT_3[64142] = 32'b00000000000000010011111011110011;
assign LUT_3[64143] = 32'b00000000000000011010100111010000;
assign LUT_3[64144] = 32'b00000000000000010010100000010110;
assign LUT_3[64145] = 32'b00000000000000011001001011110011;
assign LUT_3[64146] = 32'b00000000000000010100100111111010;
assign LUT_3[64147] = 32'b00000000000000011011010011010111;
assign LUT_3[64148] = 32'b00000000000000001111101110001100;
assign LUT_3[64149] = 32'b00000000000000010110011001101001;
assign LUT_3[64150] = 32'b00000000000000010001110101110000;
assign LUT_3[64151] = 32'b00000000000000011000100001001101;
assign LUT_3[64152] = 32'b00000000000000010111111001011100;
assign LUT_3[64153] = 32'b00000000000000011110100100111001;
assign LUT_3[64154] = 32'b00000000000000011010000001000000;
assign LUT_3[64155] = 32'b00000000000000100000101100011101;
assign LUT_3[64156] = 32'b00000000000000010101000111010010;
assign LUT_3[64157] = 32'b00000000000000011011110010101111;
assign LUT_3[64158] = 32'b00000000000000010111001110110110;
assign LUT_3[64159] = 32'b00000000000000011101111010010011;
assign LUT_3[64160] = 32'b00000000000000010000011011110011;
assign LUT_3[64161] = 32'b00000000000000010111000111010000;
assign LUT_3[64162] = 32'b00000000000000010010100011010111;
assign LUT_3[64163] = 32'b00000000000000011001001110110100;
assign LUT_3[64164] = 32'b00000000000000001101101001101001;
assign LUT_3[64165] = 32'b00000000000000010100010101000110;
assign LUT_3[64166] = 32'b00000000000000001111110001001101;
assign LUT_3[64167] = 32'b00000000000000010110011100101010;
assign LUT_3[64168] = 32'b00000000000000010101110100111001;
assign LUT_3[64169] = 32'b00000000000000011100100000010110;
assign LUT_3[64170] = 32'b00000000000000010111111100011101;
assign LUT_3[64171] = 32'b00000000000000011110100111111010;
assign LUT_3[64172] = 32'b00000000000000010011000010101111;
assign LUT_3[64173] = 32'b00000000000000011001101110001100;
assign LUT_3[64174] = 32'b00000000000000010101001010010011;
assign LUT_3[64175] = 32'b00000000000000011011110101110000;
assign LUT_3[64176] = 32'b00000000000000010011101110110110;
assign LUT_3[64177] = 32'b00000000000000011010011010010011;
assign LUT_3[64178] = 32'b00000000000000010101110110011010;
assign LUT_3[64179] = 32'b00000000000000011100100001110111;
assign LUT_3[64180] = 32'b00000000000000010000111100101100;
assign LUT_3[64181] = 32'b00000000000000010111101000001001;
assign LUT_3[64182] = 32'b00000000000000010011000100010000;
assign LUT_3[64183] = 32'b00000000000000011001101111101101;
assign LUT_3[64184] = 32'b00000000000000011001000111111100;
assign LUT_3[64185] = 32'b00000000000000011111110011011001;
assign LUT_3[64186] = 32'b00000000000000011011001111100000;
assign LUT_3[64187] = 32'b00000000000000100001111010111101;
assign LUT_3[64188] = 32'b00000000000000010110010101110010;
assign LUT_3[64189] = 32'b00000000000000011101000001001111;
assign LUT_3[64190] = 32'b00000000000000011000011101010110;
assign LUT_3[64191] = 32'b00000000000000011111001000110011;
assign LUT_3[64192] = 32'b00000000000000001111000101111110;
assign LUT_3[64193] = 32'b00000000000000010101110001011011;
assign LUT_3[64194] = 32'b00000000000000010001001101100010;
assign LUT_3[64195] = 32'b00000000000000010111111000111111;
assign LUT_3[64196] = 32'b00000000000000001100010011110100;
assign LUT_3[64197] = 32'b00000000000000010010111111010001;
assign LUT_3[64198] = 32'b00000000000000001110011011011000;
assign LUT_3[64199] = 32'b00000000000000010101000110110101;
assign LUT_3[64200] = 32'b00000000000000010100011111000100;
assign LUT_3[64201] = 32'b00000000000000011011001010100001;
assign LUT_3[64202] = 32'b00000000000000010110100110101000;
assign LUT_3[64203] = 32'b00000000000000011101010010000101;
assign LUT_3[64204] = 32'b00000000000000010001101100111010;
assign LUT_3[64205] = 32'b00000000000000011000011000010111;
assign LUT_3[64206] = 32'b00000000000000010011110100011110;
assign LUT_3[64207] = 32'b00000000000000011010011111111011;
assign LUT_3[64208] = 32'b00000000000000010010011001000001;
assign LUT_3[64209] = 32'b00000000000000011001000100011110;
assign LUT_3[64210] = 32'b00000000000000010100100000100101;
assign LUT_3[64211] = 32'b00000000000000011011001100000010;
assign LUT_3[64212] = 32'b00000000000000001111100110110111;
assign LUT_3[64213] = 32'b00000000000000010110010010010100;
assign LUT_3[64214] = 32'b00000000000000010001101110011011;
assign LUT_3[64215] = 32'b00000000000000011000011001111000;
assign LUT_3[64216] = 32'b00000000000000010111110010000111;
assign LUT_3[64217] = 32'b00000000000000011110011101100100;
assign LUT_3[64218] = 32'b00000000000000011001111001101011;
assign LUT_3[64219] = 32'b00000000000000100000100101001000;
assign LUT_3[64220] = 32'b00000000000000010100111111111101;
assign LUT_3[64221] = 32'b00000000000000011011101011011010;
assign LUT_3[64222] = 32'b00000000000000010111000111100001;
assign LUT_3[64223] = 32'b00000000000000011101110010111110;
assign LUT_3[64224] = 32'b00000000000000010000010100011110;
assign LUT_3[64225] = 32'b00000000000000010110111111111011;
assign LUT_3[64226] = 32'b00000000000000010010011100000010;
assign LUT_3[64227] = 32'b00000000000000011001000111011111;
assign LUT_3[64228] = 32'b00000000000000001101100010010100;
assign LUT_3[64229] = 32'b00000000000000010100001101110001;
assign LUT_3[64230] = 32'b00000000000000001111101001111000;
assign LUT_3[64231] = 32'b00000000000000010110010101010101;
assign LUT_3[64232] = 32'b00000000000000010101101101100100;
assign LUT_3[64233] = 32'b00000000000000011100011001000001;
assign LUT_3[64234] = 32'b00000000000000010111110101001000;
assign LUT_3[64235] = 32'b00000000000000011110100000100101;
assign LUT_3[64236] = 32'b00000000000000010010111011011010;
assign LUT_3[64237] = 32'b00000000000000011001100110110111;
assign LUT_3[64238] = 32'b00000000000000010101000010111110;
assign LUT_3[64239] = 32'b00000000000000011011101110011011;
assign LUT_3[64240] = 32'b00000000000000010011100111100001;
assign LUT_3[64241] = 32'b00000000000000011010010010111110;
assign LUT_3[64242] = 32'b00000000000000010101101111000101;
assign LUT_3[64243] = 32'b00000000000000011100011010100010;
assign LUT_3[64244] = 32'b00000000000000010000110101010111;
assign LUT_3[64245] = 32'b00000000000000010111100000110100;
assign LUT_3[64246] = 32'b00000000000000010010111100111011;
assign LUT_3[64247] = 32'b00000000000000011001101000011000;
assign LUT_3[64248] = 32'b00000000000000011001000000100111;
assign LUT_3[64249] = 32'b00000000000000011111101100000100;
assign LUT_3[64250] = 32'b00000000000000011011001000001011;
assign LUT_3[64251] = 32'b00000000000000100001110011101000;
assign LUT_3[64252] = 32'b00000000000000010110001110011101;
assign LUT_3[64253] = 32'b00000000000000011100111001111010;
assign LUT_3[64254] = 32'b00000000000000011000010110000001;
assign LUT_3[64255] = 32'b00000000000000011111000001011110;
assign LUT_3[64256] = 32'b00000000000000001001010001110110;
assign LUT_3[64257] = 32'b00000000000000001111111101010011;
assign LUT_3[64258] = 32'b00000000000000001011011001011010;
assign LUT_3[64259] = 32'b00000000000000010010000100110111;
assign LUT_3[64260] = 32'b00000000000000000110011111101100;
assign LUT_3[64261] = 32'b00000000000000001101001011001001;
assign LUT_3[64262] = 32'b00000000000000001000100111010000;
assign LUT_3[64263] = 32'b00000000000000001111010010101101;
assign LUT_3[64264] = 32'b00000000000000001110101010111100;
assign LUT_3[64265] = 32'b00000000000000010101010110011001;
assign LUT_3[64266] = 32'b00000000000000010000110010100000;
assign LUT_3[64267] = 32'b00000000000000010111011101111101;
assign LUT_3[64268] = 32'b00000000000000001011111000110010;
assign LUT_3[64269] = 32'b00000000000000010010100100001111;
assign LUT_3[64270] = 32'b00000000000000001110000000010110;
assign LUT_3[64271] = 32'b00000000000000010100101011110011;
assign LUT_3[64272] = 32'b00000000000000001100100100111001;
assign LUT_3[64273] = 32'b00000000000000010011010000010110;
assign LUT_3[64274] = 32'b00000000000000001110101100011101;
assign LUT_3[64275] = 32'b00000000000000010101010111111010;
assign LUT_3[64276] = 32'b00000000000000001001110010101111;
assign LUT_3[64277] = 32'b00000000000000010000011110001100;
assign LUT_3[64278] = 32'b00000000000000001011111010010011;
assign LUT_3[64279] = 32'b00000000000000010010100101110000;
assign LUT_3[64280] = 32'b00000000000000010001111101111111;
assign LUT_3[64281] = 32'b00000000000000011000101001011100;
assign LUT_3[64282] = 32'b00000000000000010100000101100011;
assign LUT_3[64283] = 32'b00000000000000011010110001000000;
assign LUT_3[64284] = 32'b00000000000000001111001011110101;
assign LUT_3[64285] = 32'b00000000000000010101110111010010;
assign LUT_3[64286] = 32'b00000000000000010001010011011001;
assign LUT_3[64287] = 32'b00000000000000010111111110110110;
assign LUT_3[64288] = 32'b00000000000000001010100000010110;
assign LUT_3[64289] = 32'b00000000000000010001001011110011;
assign LUT_3[64290] = 32'b00000000000000001100100111111010;
assign LUT_3[64291] = 32'b00000000000000010011010011010111;
assign LUT_3[64292] = 32'b00000000000000000111101110001100;
assign LUT_3[64293] = 32'b00000000000000001110011001101001;
assign LUT_3[64294] = 32'b00000000000000001001110101110000;
assign LUT_3[64295] = 32'b00000000000000010000100001001101;
assign LUT_3[64296] = 32'b00000000000000001111111001011100;
assign LUT_3[64297] = 32'b00000000000000010110100100111001;
assign LUT_3[64298] = 32'b00000000000000010010000001000000;
assign LUT_3[64299] = 32'b00000000000000011000101100011101;
assign LUT_3[64300] = 32'b00000000000000001101000111010010;
assign LUT_3[64301] = 32'b00000000000000010011110010101111;
assign LUT_3[64302] = 32'b00000000000000001111001110110110;
assign LUT_3[64303] = 32'b00000000000000010101111010010011;
assign LUT_3[64304] = 32'b00000000000000001101110011011001;
assign LUT_3[64305] = 32'b00000000000000010100011110110110;
assign LUT_3[64306] = 32'b00000000000000001111111010111101;
assign LUT_3[64307] = 32'b00000000000000010110100110011010;
assign LUT_3[64308] = 32'b00000000000000001011000001001111;
assign LUT_3[64309] = 32'b00000000000000010001101100101100;
assign LUT_3[64310] = 32'b00000000000000001101001000110011;
assign LUT_3[64311] = 32'b00000000000000010011110100010000;
assign LUT_3[64312] = 32'b00000000000000010011001100011111;
assign LUT_3[64313] = 32'b00000000000000011001110111111100;
assign LUT_3[64314] = 32'b00000000000000010101010100000011;
assign LUT_3[64315] = 32'b00000000000000011011111111100000;
assign LUT_3[64316] = 32'b00000000000000010000011010010101;
assign LUT_3[64317] = 32'b00000000000000010111000101110010;
assign LUT_3[64318] = 32'b00000000000000010010100001111001;
assign LUT_3[64319] = 32'b00000000000000011001001101010110;
assign LUT_3[64320] = 32'b00000000000000001001001010100001;
assign LUT_3[64321] = 32'b00000000000000001111110101111110;
assign LUT_3[64322] = 32'b00000000000000001011010010000101;
assign LUT_3[64323] = 32'b00000000000000010001111101100010;
assign LUT_3[64324] = 32'b00000000000000000110011000010111;
assign LUT_3[64325] = 32'b00000000000000001101000011110100;
assign LUT_3[64326] = 32'b00000000000000001000011111111011;
assign LUT_3[64327] = 32'b00000000000000001111001011011000;
assign LUT_3[64328] = 32'b00000000000000001110100011100111;
assign LUT_3[64329] = 32'b00000000000000010101001111000100;
assign LUT_3[64330] = 32'b00000000000000010000101011001011;
assign LUT_3[64331] = 32'b00000000000000010111010110101000;
assign LUT_3[64332] = 32'b00000000000000001011110001011101;
assign LUT_3[64333] = 32'b00000000000000010010011100111010;
assign LUT_3[64334] = 32'b00000000000000001101111001000001;
assign LUT_3[64335] = 32'b00000000000000010100100100011110;
assign LUT_3[64336] = 32'b00000000000000001100011101100100;
assign LUT_3[64337] = 32'b00000000000000010011001001000001;
assign LUT_3[64338] = 32'b00000000000000001110100101001000;
assign LUT_3[64339] = 32'b00000000000000010101010000100101;
assign LUT_3[64340] = 32'b00000000000000001001101011011010;
assign LUT_3[64341] = 32'b00000000000000010000010110110111;
assign LUT_3[64342] = 32'b00000000000000001011110010111110;
assign LUT_3[64343] = 32'b00000000000000010010011110011011;
assign LUT_3[64344] = 32'b00000000000000010001110110101010;
assign LUT_3[64345] = 32'b00000000000000011000100010000111;
assign LUT_3[64346] = 32'b00000000000000010011111110001110;
assign LUT_3[64347] = 32'b00000000000000011010101001101011;
assign LUT_3[64348] = 32'b00000000000000001111000100100000;
assign LUT_3[64349] = 32'b00000000000000010101101111111101;
assign LUT_3[64350] = 32'b00000000000000010001001100000100;
assign LUT_3[64351] = 32'b00000000000000010111110111100001;
assign LUT_3[64352] = 32'b00000000000000001010011001000001;
assign LUT_3[64353] = 32'b00000000000000010001000100011110;
assign LUT_3[64354] = 32'b00000000000000001100100000100101;
assign LUT_3[64355] = 32'b00000000000000010011001100000010;
assign LUT_3[64356] = 32'b00000000000000000111100110110111;
assign LUT_3[64357] = 32'b00000000000000001110010010010100;
assign LUT_3[64358] = 32'b00000000000000001001101110011011;
assign LUT_3[64359] = 32'b00000000000000010000011001111000;
assign LUT_3[64360] = 32'b00000000000000001111110010000111;
assign LUT_3[64361] = 32'b00000000000000010110011101100100;
assign LUT_3[64362] = 32'b00000000000000010001111001101011;
assign LUT_3[64363] = 32'b00000000000000011000100101001000;
assign LUT_3[64364] = 32'b00000000000000001100111111111101;
assign LUT_3[64365] = 32'b00000000000000010011101011011010;
assign LUT_3[64366] = 32'b00000000000000001111000111100001;
assign LUT_3[64367] = 32'b00000000000000010101110010111110;
assign LUT_3[64368] = 32'b00000000000000001101101100000100;
assign LUT_3[64369] = 32'b00000000000000010100010111100001;
assign LUT_3[64370] = 32'b00000000000000001111110011101000;
assign LUT_3[64371] = 32'b00000000000000010110011111000101;
assign LUT_3[64372] = 32'b00000000000000001010111001111010;
assign LUT_3[64373] = 32'b00000000000000010001100101010111;
assign LUT_3[64374] = 32'b00000000000000001101000001011110;
assign LUT_3[64375] = 32'b00000000000000010011101100111011;
assign LUT_3[64376] = 32'b00000000000000010011000101001010;
assign LUT_3[64377] = 32'b00000000000000011001110000100111;
assign LUT_3[64378] = 32'b00000000000000010101001100101110;
assign LUT_3[64379] = 32'b00000000000000011011111000001011;
assign LUT_3[64380] = 32'b00000000000000010000010011000000;
assign LUT_3[64381] = 32'b00000000000000010110111110011101;
assign LUT_3[64382] = 32'b00000000000000010010011010100100;
assign LUT_3[64383] = 32'b00000000000000011001000110000001;
assign LUT_3[64384] = 32'b00000000000000001011011100110100;
assign LUT_3[64385] = 32'b00000000000000010010001000010001;
assign LUT_3[64386] = 32'b00000000000000001101100100011000;
assign LUT_3[64387] = 32'b00000000000000010100001111110101;
assign LUT_3[64388] = 32'b00000000000000001000101010101010;
assign LUT_3[64389] = 32'b00000000000000001111010110000111;
assign LUT_3[64390] = 32'b00000000000000001010110010001110;
assign LUT_3[64391] = 32'b00000000000000010001011101101011;
assign LUT_3[64392] = 32'b00000000000000010000110101111010;
assign LUT_3[64393] = 32'b00000000000000010111100001010111;
assign LUT_3[64394] = 32'b00000000000000010010111101011110;
assign LUT_3[64395] = 32'b00000000000000011001101000111011;
assign LUT_3[64396] = 32'b00000000000000001110000011110000;
assign LUT_3[64397] = 32'b00000000000000010100101111001101;
assign LUT_3[64398] = 32'b00000000000000010000001011010100;
assign LUT_3[64399] = 32'b00000000000000010110110110110001;
assign LUT_3[64400] = 32'b00000000000000001110101111110111;
assign LUT_3[64401] = 32'b00000000000000010101011011010100;
assign LUT_3[64402] = 32'b00000000000000010000110111011011;
assign LUT_3[64403] = 32'b00000000000000010111100010111000;
assign LUT_3[64404] = 32'b00000000000000001011111101101101;
assign LUT_3[64405] = 32'b00000000000000010010101001001010;
assign LUT_3[64406] = 32'b00000000000000001110000101010001;
assign LUT_3[64407] = 32'b00000000000000010100110000101110;
assign LUT_3[64408] = 32'b00000000000000010100001000111101;
assign LUT_3[64409] = 32'b00000000000000011010110100011010;
assign LUT_3[64410] = 32'b00000000000000010110010000100001;
assign LUT_3[64411] = 32'b00000000000000011100111011111110;
assign LUT_3[64412] = 32'b00000000000000010001010110110011;
assign LUT_3[64413] = 32'b00000000000000011000000010010000;
assign LUT_3[64414] = 32'b00000000000000010011011110010111;
assign LUT_3[64415] = 32'b00000000000000011010001001110100;
assign LUT_3[64416] = 32'b00000000000000001100101011010100;
assign LUT_3[64417] = 32'b00000000000000010011010110110001;
assign LUT_3[64418] = 32'b00000000000000001110110010111000;
assign LUT_3[64419] = 32'b00000000000000010101011110010101;
assign LUT_3[64420] = 32'b00000000000000001001111001001010;
assign LUT_3[64421] = 32'b00000000000000010000100100100111;
assign LUT_3[64422] = 32'b00000000000000001100000000101110;
assign LUT_3[64423] = 32'b00000000000000010010101100001011;
assign LUT_3[64424] = 32'b00000000000000010010000100011010;
assign LUT_3[64425] = 32'b00000000000000011000101111110111;
assign LUT_3[64426] = 32'b00000000000000010100001011111110;
assign LUT_3[64427] = 32'b00000000000000011010110111011011;
assign LUT_3[64428] = 32'b00000000000000001111010010010000;
assign LUT_3[64429] = 32'b00000000000000010101111101101101;
assign LUT_3[64430] = 32'b00000000000000010001011001110100;
assign LUT_3[64431] = 32'b00000000000000011000000101010001;
assign LUT_3[64432] = 32'b00000000000000001111111110010111;
assign LUT_3[64433] = 32'b00000000000000010110101001110100;
assign LUT_3[64434] = 32'b00000000000000010010000101111011;
assign LUT_3[64435] = 32'b00000000000000011000110001011000;
assign LUT_3[64436] = 32'b00000000000000001101001100001101;
assign LUT_3[64437] = 32'b00000000000000010011110111101010;
assign LUT_3[64438] = 32'b00000000000000001111010011110001;
assign LUT_3[64439] = 32'b00000000000000010101111111001110;
assign LUT_3[64440] = 32'b00000000000000010101010111011101;
assign LUT_3[64441] = 32'b00000000000000011100000010111010;
assign LUT_3[64442] = 32'b00000000000000010111011111000001;
assign LUT_3[64443] = 32'b00000000000000011110001010011110;
assign LUT_3[64444] = 32'b00000000000000010010100101010011;
assign LUT_3[64445] = 32'b00000000000000011001010000110000;
assign LUT_3[64446] = 32'b00000000000000010100101100110111;
assign LUT_3[64447] = 32'b00000000000000011011011000010100;
assign LUT_3[64448] = 32'b00000000000000001011010101011111;
assign LUT_3[64449] = 32'b00000000000000010010000000111100;
assign LUT_3[64450] = 32'b00000000000000001101011101000011;
assign LUT_3[64451] = 32'b00000000000000010100001000100000;
assign LUT_3[64452] = 32'b00000000000000001000100011010101;
assign LUT_3[64453] = 32'b00000000000000001111001110110010;
assign LUT_3[64454] = 32'b00000000000000001010101010111001;
assign LUT_3[64455] = 32'b00000000000000010001010110010110;
assign LUT_3[64456] = 32'b00000000000000010000101110100101;
assign LUT_3[64457] = 32'b00000000000000010111011010000010;
assign LUT_3[64458] = 32'b00000000000000010010110110001001;
assign LUT_3[64459] = 32'b00000000000000011001100001100110;
assign LUT_3[64460] = 32'b00000000000000001101111100011011;
assign LUT_3[64461] = 32'b00000000000000010100100111111000;
assign LUT_3[64462] = 32'b00000000000000010000000011111111;
assign LUT_3[64463] = 32'b00000000000000010110101111011100;
assign LUT_3[64464] = 32'b00000000000000001110101000100010;
assign LUT_3[64465] = 32'b00000000000000010101010011111111;
assign LUT_3[64466] = 32'b00000000000000010000110000000110;
assign LUT_3[64467] = 32'b00000000000000010111011011100011;
assign LUT_3[64468] = 32'b00000000000000001011110110011000;
assign LUT_3[64469] = 32'b00000000000000010010100001110101;
assign LUT_3[64470] = 32'b00000000000000001101111101111100;
assign LUT_3[64471] = 32'b00000000000000010100101001011001;
assign LUT_3[64472] = 32'b00000000000000010100000001101000;
assign LUT_3[64473] = 32'b00000000000000011010101101000101;
assign LUT_3[64474] = 32'b00000000000000010110001001001100;
assign LUT_3[64475] = 32'b00000000000000011100110100101001;
assign LUT_3[64476] = 32'b00000000000000010001001111011110;
assign LUT_3[64477] = 32'b00000000000000010111111010111011;
assign LUT_3[64478] = 32'b00000000000000010011010111000010;
assign LUT_3[64479] = 32'b00000000000000011010000010011111;
assign LUT_3[64480] = 32'b00000000000000001100100011111111;
assign LUT_3[64481] = 32'b00000000000000010011001111011100;
assign LUT_3[64482] = 32'b00000000000000001110101011100011;
assign LUT_3[64483] = 32'b00000000000000010101010111000000;
assign LUT_3[64484] = 32'b00000000000000001001110001110101;
assign LUT_3[64485] = 32'b00000000000000010000011101010010;
assign LUT_3[64486] = 32'b00000000000000001011111001011001;
assign LUT_3[64487] = 32'b00000000000000010010100100110110;
assign LUT_3[64488] = 32'b00000000000000010001111101000101;
assign LUT_3[64489] = 32'b00000000000000011000101000100010;
assign LUT_3[64490] = 32'b00000000000000010100000100101001;
assign LUT_3[64491] = 32'b00000000000000011010110000000110;
assign LUT_3[64492] = 32'b00000000000000001111001010111011;
assign LUT_3[64493] = 32'b00000000000000010101110110011000;
assign LUT_3[64494] = 32'b00000000000000010001010010011111;
assign LUT_3[64495] = 32'b00000000000000010111111101111100;
assign LUT_3[64496] = 32'b00000000000000001111110111000010;
assign LUT_3[64497] = 32'b00000000000000010110100010011111;
assign LUT_3[64498] = 32'b00000000000000010001111110100110;
assign LUT_3[64499] = 32'b00000000000000011000101010000011;
assign LUT_3[64500] = 32'b00000000000000001101000100111000;
assign LUT_3[64501] = 32'b00000000000000010011110000010101;
assign LUT_3[64502] = 32'b00000000000000001111001100011100;
assign LUT_3[64503] = 32'b00000000000000010101110111111001;
assign LUT_3[64504] = 32'b00000000000000010101010000001000;
assign LUT_3[64505] = 32'b00000000000000011011111011100101;
assign LUT_3[64506] = 32'b00000000000000010111010111101100;
assign LUT_3[64507] = 32'b00000000000000011110000011001001;
assign LUT_3[64508] = 32'b00000000000000010010011101111110;
assign LUT_3[64509] = 32'b00000000000000011001001001011011;
assign LUT_3[64510] = 32'b00000000000000010100100101100010;
assign LUT_3[64511] = 32'b00000000000000011011010000111111;
assign LUT_3[64512] = 32'b00000000000000010000010010000110;
assign LUT_3[64513] = 32'b00000000000000010110111101100011;
assign LUT_3[64514] = 32'b00000000000000010010011001101010;
assign LUT_3[64515] = 32'b00000000000000011001000101000111;
assign LUT_3[64516] = 32'b00000000000000001101011111111100;
assign LUT_3[64517] = 32'b00000000000000010100001011011001;
assign LUT_3[64518] = 32'b00000000000000001111100111100000;
assign LUT_3[64519] = 32'b00000000000000010110010010111101;
assign LUT_3[64520] = 32'b00000000000000010101101011001100;
assign LUT_3[64521] = 32'b00000000000000011100010110101001;
assign LUT_3[64522] = 32'b00000000000000010111110010110000;
assign LUT_3[64523] = 32'b00000000000000011110011110001101;
assign LUT_3[64524] = 32'b00000000000000010010111001000010;
assign LUT_3[64525] = 32'b00000000000000011001100100011111;
assign LUT_3[64526] = 32'b00000000000000010101000000100110;
assign LUT_3[64527] = 32'b00000000000000011011101100000011;
assign LUT_3[64528] = 32'b00000000000000010011100101001001;
assign LUT_3[64529] = 32'b00000000000000011010010000100110;
assign LUT_3[64530] = 32'b00000000000000010101101100101101;
assign LUT_3[64531] = 32'b00000000000000011100011000001010;
assign LUT_3[64532] = 32'b00000000000000010000110010111111;
assign LUT_3[64533] = 32'b00000000000000010111011110011100;
assign LUT_3[64534] = 32'b00000000000000010010111010100011;
assign LUT_3[64535] = 32'b00000000000000011001100110000000;
assign LUT_3[64536] = 32'b00000000000000011000111110001111;
assign LUT_3[64537] = 32'b00000000000000011111101001101100;
assign LUT_3[64538] = 32'b00000000000000011011000101110011;
assign LUT_3[64539] = 32'b00000000000000100001110001010000;
assign LUT_3[64540] = 32'b00000000000000010110001100000101;
assign LUT_3[64541] = 32'b00000000000000011100110111100010;
assign LUT_3[64542] = 32'b00000000000000011000010011101001;
assign LUT_3[64543] = 32'b00000000000000011110111111000110;
assign LUT_3[64544] = 32'b00000000000000010001100000100110;
assign LUT_3[64545] = 32'b00000000000000011000001100000011;
assign LUT_3[64546] = 32'b00000000000000010011101000001010;
assign LUT_3[64547] = 32'b00000000000000011010010011100111;
assign LUT_3[64548] = 32'b00000000000000001110101110011100;
assign LUT_3[64549] = 32'b00000000000000010101011001111001;
assign LUT_3[64550] = 32'b00000000000000010000110110000000;
assign LUT_3[64551] = 32'b00000000000000010111100001011101;
assign LUT_3[64552] = 32'b00000000000000010110111001101100;
assign LUT_3[64553] = 32'b00000000000000011101100101001001;
assign LUT_3[64554] = 32'b00000000000000011001000001010000;
assign LUT_3[64555] = 32'b00000000000000011111101100101101;
assign LUT_3[64556] = 32'b00000000000000010100000111100010;
assign LUT_3[64557] = 32'b00000000000000011010110010111111;
assign LUT_3[64558] = 32'b00000000000000010110001111000110;
assign LUT_3[64559] = 32'b00000000000000011100111010100011;
assign LUT_3[64560] = 32'b00000000000000010100110011101001;
assign LUT_3[64561] = 32'b00000000000000011011011111000110;
assign LUT_3[64562] = 32'b00000000000000010110111011001101;
assign LUT_3[64563] = 32'b00000000000000011101100110101010;
assign LUT_3[64564] = 32'b00000000000000010010000001011111;
assign LUT_3[64565] = 32'b00000000000000011000101100111100;
assign LUT_3[64566] = 32'b00000000000000010100001001000011;
assign LUT_3[64567] = 32'b00000000000000011010110100100000;
assign LUT_3[64568] = 32'b00000000000000011010001100101111;
assign LUT_3[64569] = 32'b00000000000000100000111000001100;
assign LUT_3[64570] = 32'b00000000000000011100010100010011;
assign LUT_3[64571] = 32'b00000000000000100010111111110000;
assign LUT_3[64572] = 32'b00000000000000010111011010100101;
assign LUT_3[64573] = 32'b00000000000000011110000110000010;
assign LUT_3[64574] = 32'b00000000000000011001100010001001;
assign LUT_3[64575] = 32'b00000000000000100000001101100110;
assign LUT_3[64576] = 32'b00000000000000010000001010110001;
assign LUT_3[64577] = 32'b00000000000000010110110110001110;
assign LUT_3[64578] = 32'b00000000000000010010010010010101;
assign LUT_3[64579] = 32'b00000000000000011000111101110010;
assign LUT_3[64580] = 32'b00000000000000001101011000100111;
assign LUT_3[64581] = 32'b00000000000000010100000100000100;
assign LUT_3[64582] = 32'b00000000000000001111100000001011;
assign LUT_3[64583] = 32'b00000000000000010110001011101000;
assign LUT_3[64584] = 32'b00000000000000010101100011110111;
assign LUT_3[64585] = 32'b00000000000000011100001111010100;
assign LUT_3[64586] = 32'b00000000000000010111101011011011;
assign LUT_3[64587] = 32'b00000000000000011110010110111000;
assign LUT_3[64588] = 32'b00000000000000010010110001101101;
assign LUT_3[64589] = 32'b00000000000000011001011101001010;
assign LUT_3[64590] = 32'b00000000000000010100111001010001;
assign LUT_3[64591] = 32'b00000000000000011011100100101110;
assign LUT_3[64592] = 32'b00000000000000010011011101110100;
assign LUT_3[64593] = 32'b00000000000000011010001001010001;
assign LUT_3[64594] = 32'b00000000000000010101100101011000;
assign LUT_3[64595] = 32'b00000000000000011100010000110101;
assign LUT_3[64596] = 32'b00000000000000010000101011101010;
assign LUT_3[64597] = 32'b00000000000000010111010111000111;
assign LUT_3[64598] = 32'b00000000000000010010110011001110;
assign LUT_3[64599] = 32'b00000000000000011001011110101011;
assign LUT_3[64600] = 32'b00000000000000011000110110111010;
assign LUT_3[64601] = 32'b00000000000000011111100010010111;
assign LUT_3[64602] = 32'b00000000000000011010111110011110;
assign LUT_3[64603] = 32'b00000000000000100001101001111011;
assign LUT_3[64604] = 32'b00000000000000010110000100110000;
assign LUT_3[64605] = 32'b00000000000000011100110000001101;
assign LUT_3[64606] = 32'b00000000000000011000001100010100;
assign LUT_3[64607] = 32'b00000000000000011110110111110001;
assign LUT_3[64608] = 32'b00000000000000010001011001010001;
assign LUT_3[64609] = 32'b00000000000000011000000100101110;
assign LUT_3[64610] = 32'b00000000000000010011100000110101;
assign LUT_3[64611] = 32'b00000000000000011010001100010010;
assign LUT_3[64612] = 32'b00000000000000001110100111000111;
assign LUT_3[64613] = 32'b00000000000000010101010010100100;
assign LUT_3[64614] = 32'b00000000000000010000101110101011;
assign LUT_3[64615] = 32'b00000000000000010111011010001000;
assign LUT_3[64616] = 32'b00000000000000010110110010010111;
assign LUT_3[64617] = 32'b00000000000000011101011101110100;
assign LUT_3[64618] = 32'b00000000000000011000111001111011;
assign LUT_3[64619] = 32'b00000000000000011111100101011000;
assign LUT_3[64620] = 32'b00000000000000010100000000001101;
assign LUT_3[64621] = 32'b00000000000000011010101011101010;
assign LUT_3[64622] = 32'b00000000000000010110000111110001;
assign LUT_3[64623] = 32'b00000000000000011100110011001110;
assign LUT_3[64624] = 32'b00000000000000010100101100010100;
assign LUT_3[64625] = 32'b00000000000000011011010111110001;
assign LUT_3[64626] = 32'b00000000000000010110110011111000;
assign LUT_3[64627] = 32'b00000000000000011101011111010101;
assign LUT_3[64628] = 32'b00000000000000010001111010001010;
assign LUT_3[64629] = 32'b00000000000000011000100101100111;
assign LUT_3[64630] = 32'b00000000000000010100000001101110;
assign LUT_3[64631] = 32'b00000000000000011010101101001011;
assign LUT_3[64632] = 32'b00000000000000011010000101011010;
assign LUT_3[64633] = 32'b00000000000000100000110000110111;
assign LUT_3[64634] = 32'b00000000000000011100001100111110;
assign LUT_3[64635] = 32'b00000000000000100010111000011011;
assign LUT_3[64636] = 32'b00000000000000010111010011010000;
assign LUT_3[64637] = 32'b00000000000000011101111110101101;
assign LUT_3[64638] = 32'b00000000000000011001011010110100;
assign LUT_3[64639] = 32'b00000000000000100000000110010001;
assign LUT_3[64640] = 32'b00000000000000010010011101000100;
assign LUT_3[64641] = 32'b00000000000000011001001000100001;
assign LUT_3[64642] = 32'b00000000000000010100100100101000;
assign LUT_3[64643] = 32'b00000000000000011011010000000101;
assign LUT_3[64644] = 32'b00000000000000001111101010111010;
assign LUT_3[64645] = 32'b00000000000000010110010110010111;
assign LUT_3[64646] = 32'b00000000000000010001110010011110;
assign LUT_3[64647] = 32'b00000000000000011000011101111011;
assign LUT_3[64648] = 32'b00000000000000010111110110001010;
assign LUT_3[64649] = 32'b00000000000000011110100001100111;
assign LUT_3[64650] = 32'b00000000000000011001111101101110;
assign LUT_3[64651] = 32'b00000000000000100000101001001011;
assign LUT_3[64652] = 32'b00000000000000010101000100000000;
assign LUT_3[64653] = 32'b00000000000000011011101111011101;
assign LUT_3[64654] = 32'b00000000000000010111001011100100;
assign LUT_3[64655] = 32'b00000000000000011101110111000001;
assign LUT_3[64656] = 32'b00000000000000010101110000000111;
assign LUT_3[64657] = 32'b00000000000000011100011011100100;
assign LUT_3[64658] = 32'b00000000000000010111110111101011;
assign LUT_3[64659] = 32'b00000000000000011110100011001000;
assign LUT_3[64660] = 32'b00000000000000010010111101111101;
assign LUT_3[64661] = 32'b00000000000000011001101001011010;
assign LUT_3[64662] = 32'b00000000000000010101000101100001;
assign LUT_3[64663] = 32'b00000000000000011011110000111110;
assign LUT_3[64664] = 32'b00000000000000011011001001001101;
assign LUT_3[64665] = 32'b00000000000000100001110100101010;
assign LUT_3[64666] = 32'b00000000000000011101010000110001;
assign LUT_3[64667] = 32'b00000000000000100011111100001110;
assign LUT_3[64668] = 32'b00000000000000011000010111000011;
assign LUT_3[64669] = 32'b00000000000000011111000010100000;
assign LUT_3[64670] = 32'b00000000000000011010011110100111;
assign LUT_3[64671] = 32'b00000000000000100001001010000100;
assign LUT_3[64672] = 32'b00000000000000010011101011100100;
assign LUT_3[64673] = 32'b00000000000000011010010111000001;
assign LUT_3[64674] = 32'b00000000000000010101110011001000;
assign LUT_3[64675] = 32'b00000000000000011100011110100101;
assign LUT_3[64676] = 32'b00000000000000010000111001011010;
assign LUT_3[64677] = 32'b00000000000000010111100100110111;
assign LUT_3[64678] = 32'b00000000000000010011000000111110;
assign LUT_3[64679] = 32'b00000000000000011001101100011011;
assign LUT_3[64680] = 32'b00000000000000011001000100101010;
assign LUT_3[64681] = 32'b00000000000000011111110000000111;
assign LUT_3[64682] = 32'b00000000000000011011001100001110;
assign LUT_3[64683] = 32'b00000000000000100001110111101011;
assign LUT_3[64684] = 32'b00000000000000010110010010100000;
assign LUT_3[64685] = 32'b00000000000000011100111101111101;
assign LUT_3[64686] = 32'b00000000000000011000011010000100;
assign LUT_3[64687] = 32'b00000000000000011111000101100001;
assign LUT_3[64688] = 32'b00000000000000010110111110100111;
assign LUT_3[64689] = 32'b00000000000000011101101010000100;
assign LUT_3[64690] = 32'b00000000000000011001000110001011;
assign LUT_3[64691] = 32'b00000000000000011111110001101000;
assign LUT_3[64692] = 32'b00000000000000010100001100011101;
assign LUT_3[64693] = 32'b00000000000000011010110111111010;
assign LUT_3[64694] = 32'b00000000000000010110010100000001;
assign LUT_3[64695] = 32'b00000000000000011100111111011110;
assign LUT_3[64696] = 32'b00000000000000011100010111101101;
assign LUT_3[64697] = 32'b00000000000000100011000011001010;
assign LUT_3[64698] = 32'b00000000000000011110011111010001;
assign LUT_3[64699] = 32'b00000000000000100101001010101110;
assign LUT_3[64700] = 32'b00000000000000011001100101100011;
assign LUT_3[64701] = 32'b00000000000000100000010001000000;
assign LUT_3[64702] = 32'b00000000000000011011101101000111;
assign LUT_3[64703] = 32'b00000000000000100010011000100100;
assign LUT_3[64704] = 32'b00000000000000010010010101101111;
assign LUT_3[64705] = 32'b00000000000000011001000001001100;
assign LUT_3[64706] = 32'b00000000000000010100011101010011;
assign LUT_3[64707] = 32'b00000000000000011011001000110000;
assign LUT_3[64708] = 32'b00000000000000001111100011100101;
assign LUT_3[64709] = 32'b00000000000000010110001111000010;
assign LUT_3[64710] = 32'b00000000000000010001101011001001;
assign LUT_3[64711] = 32'b00000000000000011000010110100110;
assign LUT_3[64712] = 32'b00000000000000010111101110110101;
assign LUT_3[64713] = 32'b00000000000000011110011010010010;
assign LUT_3[64714] = 32'b00000000000000011001110110011001;
assign LUT_3[64715] = 32'b00000000000000100000100001110110;
assign LUT_3[64716] = 32'b00000000000000010100111100101011;
assign LUT_3[64717] = 32'b00000000000000011011101000001000;
assign LUT_3[64718] = 32'b00000000000000010111000100001111;
assign LUT_3[64719] = 32'b00000000000000011101101111101100;
assign LUT_3[64720] = 32'b00000000000000010101101000110010;
assign LUT_3[64721] = 32'b00000000000000011100010100001111;
assign LUT_3[64722] = 32'b00000000000000010111110000010110;
assign LUT_3[64723] = 32'b00000000000000011110011011110011;
assign LUT_3[64724] = 32'b00000000000000010010110110101000;
assign LUT_3[64725] = 32'b00000000000000011001100010000101;
assign LUT_3[64726] = 32'b00000000000000010100111110001100;
assign LUT_3[64727] = 32'b00000000000000011011101001101001;
assign LUT_3[64728] = 32'b00000000000000011011000001111000;
assign LUT_3[64729] = 32'b00000000000000100001101101010101;
assign LUT_3[64730] = 32'b00000000000000011101001001011100;
assign LUT_3[64731] = 32'b00000000000000100011110100111001;
assign LUT_3[64732] = 32'b00000000000000011000001111101110;
assign LUT_3[64733] = 32'b00000000000000011110111011001011;
assign LUT_3[64734] = 32'b00000000000000011010010111010010;
assign LUT_3[64735] = 32'b00000000000000100001000010101111;
assign LUT_3[64736] = 32'b00000000000000010011100100001111;
assign LUT_3[64737] = 32'b00000000000000011010001111101100;
assign LUT_3[64738] = 32'b00000000000000010101101011110011;
assign LUT_3[64739] = 32'b00000000000000011100010111010000;
assign LUT_3[64740] = 32'b00000000000000010000110010000101;
assign LUT_3[64741] = 32'b00000000000000010111011101100010;
assign LUT_3[64742] = 32'b00000000000000010010111001101001;
assign LUT_3[64743] = 32'b00000000000000011001100101000110;
assign LUT_3[64744] = 32'b00000000000000011000111101010101;
assign LUT_3[64745] = 32'b00000000000000011111101000110010;
assign LUT_3[64746] = 32'b00000000000000011011000100111001;
assign LUT_3[64747] = 32'b00000000000000100001110000010110;
assign LUT_3[64748] = 32'b00000000000000010110001011001011;
assign LUT_3[64749] = 32'b00000000000000011100110110101000;
assign LUT_3[64750] = 32'b00000000000000011000010010101111;
assign LUT_3[64751] = 32'b00000000000000011110111110001100;
assign LUT_3[64752] = 32'b00000000000000010110110111010010;
assign LUT_3[64753] = 32'b00000000000000011101100010101111;
assign LUT_3[64754] = 32'b00000000000000011000111110110110;
assign LUT_3[64755] = 32'b00000000000000011111101010010011;
assign LUT_3[64756] = 32'b00000000000000010100000101001000;
assign LUT_3[64757] = 32'b00000000000000011010110000100101;
assign LUT_3[64758] = 32'b00000000000000010110001100101100;
assign LUT_3[64759] = 32'b00000000000000011100111000001001;
assign LUT_3[64760] = 32'b00000000000000011100010000011000;
assign LUT_3[64761] = 32'b00000000000000100010111011110101;
assign LUT_3[64762] = 32'b00000000000000011110010111111100;
assign LUT_3[64763] = 32'b00000000000000100101000011011001;
assign LUT_3[64764] = 32'b00000000000000011001011110001110;
assign LUT_3[64765] = 32'b00000000000000100000001001101011;
assign LUT_3[64766] = 32'b00000000000000011011100101110010;
assign LUT_3[64767] = 32'b00000000000000100010010001001111;
assign LUT_3[64768] = 32'b00000000000000001100100001100111;
assign LUT_3[64769] = 32'b00000000000000010011001101000100;
assign LUT_3[64770] = 32'b00000000000000001110101001001011;
assign LUT_3[64771] = 32'b00000000000000010101010100101000;
assign LUT_3[64772] = 32'b00000000000000001001101111011101;
assign LUT_3[64773] = 32'b00000000000000010000011010111010;
assign LUT_3[64774] = 32'b00000000000000001011110111000001;
assign LUT_3[64775] = 32'b00000000000000010010100010011110;
assign LUT_3[64776] = 32'b00000000000000010001111010101101;
assign LUT_3[64777] = 32'b00000000000000011000100110001010;
assign LUT_3[64778] = 32'b00000000000000010100000010010001;
assign LUT_3[64779] = 32'b00000000000000011010101101101110;
assign LUT_3[64780] = 32'b00000000000000001111001000100011;
assign LUT_3[64781] = 32'b00000000000000010101110100000000;
assign LUT_3[64782] = 32'b00000000000000010001010000000111;
assign LUT_3[64783] = 32'b00000000000000010111111011100100;
assign LUT_3[64784] = 32'b00000000000000001111110100101010;
assign LUT_3[64785] = 32'b00000000000000010110100000000111;
assign LUT_3[64786] = 32'b00000000000000010001111100001110;
assign LUT_3[64787] = 32'b00000000000000011000100111101011;
assign LUT_3[64788] = 32'b00000000000000001101000010100000;
assign LUT_3[64789] = 32'b00000000000000010011101101111101;
assign LUT_3[64790] = 32'b00000000000000001111001010000100;
assign LUT_3[64791] = 32'b00000000000000010101110101100001;
assign LUT_3[64792] = 32'b00000000000000010101001101110000;
assign LUT_3[64793] = 32'b00000000000000011011111001001101;
assign LUT_3[64794] = 32'b00000000000000010111010101010100;
assign LUT_3[64795] = 32'b00000000000000011110000000110001;
assign LUT_3[64796] = 32'b00000000000000010010011011100110;
assign LUT_3[64797] = 32'b00000000000000011001000111000011;
assign LUT_3[64798] = 32'b00000000000000010100100011001010;
assign LUT_3[64799] = 32'b00000000000000011011001110100111;
assign LUT_3[64800] = 32'b00000000000000001101110000000111;
assign LUT_3[64801] = 32'b00000000000000010100011011100100;
assign LUT_3[64802] = 32'b00000000000000001111110111101011;
assign LUT_3[64803] = 32'b00000000000000010110100011001000;
assign LUT_3[64804] = 32'b00000000000000001010111101111101;
assign LUT_3[64805] = 32'b00000000000000010001101001011010;
assign LUT_3[64806] = 32'b00000000000000001101000101100001;
assign LUT_3[64807] = 32'b00000000000000010011110000111110;
assign LUT_3[64808] = 32'b00000000000000010011001001001101;
assign LUT_3[64809] = 32'b00000000000000011001110100101010;
assign LUT_3[64810] = 32'b00000000000000010101010000110001;
assign LUT_3[64811] = 32'b00000000000000011011111100001110;
assign LUT_3[64812] = 32'b00000000000000010000010111000011;
assign LUT_3[64813] = 32'b00000000000000010111000010100000;
assign LUT_3[64814] = 32'b00000000000000010010011110100111;
assign LUT_3[64815] = 32'b00000000000000011001001010000100;
assign LUT_3[64816] = 32'b00000000000000010001000011001010;
assign LUT_3[64817] = 32'b00000000000000010111101110100111;
assign LUT_3[64818] = 32'b00000000000000010011001010101110;
assign LUT_3[64819] = 32'b00000000000000011001110110001011;
assign LUT_3[64820] = 32'b00000000000000001110010001000000;
assign LUT_3[64821] = 32'b00000000000000010100111100011101;
assign LUT_3[64822] = 32'b00000000000000010000011000100100;
assign LUT_3[64823] = 32'b00000000000000010111000100000001;
assign LUT_3[64824] = 32'b00000000000000010110011100010000;
assign LUT_3[64825] = 32'b00000000000000011101000111101101;
assign LUT_3[64826] = 32'b00000000000000011000100011110100;
assign LUT_3[64827] = 32'b00000000000000011111001111010001;
assign LUT_3[64828] = 32'b00000000000000010011101010000110;
assign LUT_3[64829] = 32'b00000000000000011010010101100011;
assign LUT_3[64830] = 32'b00000000000000010101110001101010;
assign LUT_3[64831] = 32'b00000000000000011100011101000111;
assign LUT_3[64832] = 32'b00000000000000001100011010010010;
assign LUT_3[64833] = 32'b00000000000000010011000101101111;
assign LUT_3[64834] = 32'b00000000000000001110100001110110;
assign LUT_3[64835] = 32'b00000000000000010101001101010011;
assign LUT_3[64836] = 32'b00000000000000001001101000001000;
assign LUT_3[64837] = 32'b00000000000000010000010011100101;
assign LUT_3[64838] = 32'b00000000000000001011101111101100;
assign LUT_3[64839] = 32'b00000000000000010010011011001001;
assign LUT_3[64840] = 32'b00000000000000010001110011011000;
assign LUT_3[64841] = 32'b00000000000000011000011110110101;
assign LUT_3[64842] = 32'b00000000000000010011111010111100;
assign LUT_3[64843] = 32'b00000000000000011010100110011001;
assign LUT_3[64844] = 32'b00000000000000001111000001001110;
assign LUT_3[64845] = 32'b00000000000000010101101100101011;
assign LUT_3[64846] = 32'b00000000000000010001001000110010;
assign LUT_3[64847] = 32'b00000000000000010111110100001111;
assign LUT_3[64848] = 32'b00000000000000001111101101010101;
assign LUT_3[64849] = 32'b00000000000000010110011000110010;
assign LUT_3[64850] = 32'b00000000000000010001110100111001;
assign LUT_3[64851] = 32'b00000000000000011000100000010110;
assign LUT_3[64852] = 32'b00000000000000001100111011001011;
assign LUT_3[64853] = 32'b00000000000000010011100110101000;
assign LUT_3[64854] = 32'b00000000000000001111000010101111;
assign LUT_3[64855] = 32'b00000000000000010101101110001100;
assign LUT_3[64856] = 32'b00000000000000010101000110011011;
assign LUT_3[64857] = 32'b00000000000000011011110001111000;
assign LUT_3[64858] = 32'b00000000000000010111001101111111;
assign LUT_3[64859] = 32'b00000000000000011101111001011100;
assign LUT_3[64860] = 32'b00000000000000010010010100010001;
assign LUT_3[64861] = 32'b00000000000000011000111111101110;
assign LUT_3[64862] = 32'b00000000000000010100011011110101;
assign LUT_3[64863] = 32'b00000000000000011011000111010010;
assign LUT_3[64864] = 32'b00000000000000001101101000110010;
assign LUT_3[64865] = 32'b00000000000000010100010100001111;
assign LUT_3[64866] = 32'b00000000000000001111110000010110;
assign LUT_3[64867] = 32'b00000000000000010110011011110011;
assign LUT_3[64868] = 32'b00000000000000001010110110101000;
assign LUT_3[64869] = 32'b00000000000000010001100010000101;
assign LUT_3[64870] = 32'b00000000000000001100111110001100;
assign LUT_3[64871] = 32'b00000000000000010011101001101001;
assign LUT_3[64872] = 32'b00000000000000010011000001111000;
assign LUT_3[64873] = 32'b00000000000000011001101101010101;
assign LUT_3[64874] = 32'b00000000000000010101001001011100;
assign LUT_3[64875] = 32'b00000000000000011011110100111001;
assign LUT_3[64876] = 32'b00000000000000010000001111101110;
assign LUT_3[64877] = 32'b00000000000000010110111011001011;
assign LUT_3[64878] = 32'b00000000000000010010010111010010;
assign LUT_3[64879] = 32'b00000000000000011001000010101111;
assign LUT_3[64880] = 32'b00000000000000010000111011110101;
assign LUT_3[64881] = 32'b00000000000000010111100111010010;
assign LUT_3[64882] = 32'b00000000000000010011000011011001;
assign LUT_3[64883] = 32'b00000000000000011001101110110110;
assign LUT_3[64884] = 32'b00000000000000001110001001101011;
assign LUT_3[64885] = 32'b00000000000000010100110101001000;
assign LUT_3[64886] = 32'b00000000000000010000010001001111;
assign LUT_3[64887] = 32'b00000000000000010110111100101100;
assign LUT_3[64888] = 32'b00000000000000010110010100111011;
assign LUT_3[64889] = 32'b00000000000000011101000000011000;
assign LUT_3[64890] = 32'b00000000000000011000011100011111;
assign LUT_3[64891] = 32'b00000000000000011111000111111100;
assign LUT_3[64892] = 32'b00000000000000010011100010110001;
assign LUT_3[64893] = 32'b00000000000000011010001110001110;
assign LUT_3[64894] = 32'b00000000000000010101101010010101;
assign LUT_3[64895] = 32'b00000000000000011100010101110010;
assign LUT_3[64896] = 32'b00000000000000001110101100100101;
assign LUT_3[64897] = 32'b00000000000000010101011000000010;
assign LUT_3[64898] = 32'b00000000000000010000110100001001;
assign LUT_3[64899] = 32'b00000000000000010111011111100110;
assign LUT_3[64900] = 32'b00000000000000001011111010011011;
assign LUT_3[64901] = 32'b00000000000000010010100101111000;
assign LUT_3[64902] = 32'b00000000000000001110000001111111;
assign LUT_3[64903] = 32'b00000000000000010100101101011100;
assign LUT_3[64904] = 32'b00000000000000010100000101101011;
assign LUT_3[64905] = 32'b00000000000000011010110001001000;
assign LUT_3[64906] = 32'b00000000000000010110001101001111;
assign LUT_3[64907] = 32'b00000000000000011100111000101100;
assign LUT_3[64908] = 32'b00000000000000010001010011100001;
assign LUT_3[64909] = 32'b00000000000000010111111110111110;
assign LUT_3[64910] = 32'b00000000000000010011011011000101;
assign LUT_3[64911] = 32'b00000000000000011010000110100010;
assign LUT_3[64912] = 32'b00000000000000010001111111101000;
assign LUT_3[64913] = 32'b00000000000000011000101011000101;
assign LUT_3[64914] = 32'b00000000000000010100000111001100;
assign LUT_3[64915] = 32'b00000000000000011010110010101001;
assign LUT_3[64916] = 32'b00000000000000001111001101011110;
assign LUT_3[64917] = 32'b00000000000000010101111000111011;
assign LUT_3[64918] = 32'b00000000000000010001010101000010;
assign LUT_3[64919] = 32'b00000000000000011000000000011111;
assign LUT_3[64920] = 32'b00000000000000010111011000101110;
assign LUT_3[64921] = 32'b00000000000000011110000100001011;
assign LUT_3[64922] = 32'b00000000000000011001100000010010;
assign LUT_3[64923] = 32'b00000000000000100000001011101111;
assign LUT_3[64924] = 32'b00000000000000010100100110100100;
assign LUT_3[64925] = 32'b00000000000000011011010010000001;
assign LUT_3[64926] = 32'b00000000000000010110101110001000;
assign LUT_3[64927] = 32'b00000000000000011101011001100101;
assign LUT_3[64928] = 32'b00000000000000001111111011000101;
assign LUT_3[64929] = 32'b00000000000000010110100110100010;
assign LUT_3[64930] = 32'b00000000000000010010000010101001;
assign LUT_3[64931] = 32'b00000000000000011000101110000110;
assign LUT_3[64932] = 32'b00000000000000001101001000111011;
assign LUT_3[64933] = 32'b00000000000000010011110100011000;
assign LUT_3[64934] = 32'b00000000000000001111010000011111;
assign LUT_3[64935] = 32'b00000000000000010101111011111100;
assign LUT_3[64936] = 32'b00000000000000010101010100001011;
assign LUT_3[64937] = 32'b00000000000000011011111111101000;
assign LUT_3[64938] = 32'b00000000000000010111011011101111;
assign LUT_3[64939] = 32'b00000000000000011110000111001100;
assign LUT_3[64940] = 32'b00000000000000010010100010000001;
assign LUT_3[64941] = 32'b00000000000000011001001101011110;
assign LUT_3[64942] = 32'b00000000000000010100101001100101;
assign LUT_3[64943] = 32'b00000000000000011011010101000010;
assign LUT_3[64944] = 32'b00000000000000010011001110001000;
assign LUT_3[64945] = 32'b00000000000000011001111001100101;
assign LUT_3[64946] = 32'b00000000000000010101010101101100;
assign LUT_3[64947] = 32'b00000000000000011100000001001001;
assign LUT_3[64948] = 32'b00000000000000010000011011111110;
assign LUT_3[64949] = 32'b00000000000000010111000111011011;
assign LUT_3[64950] = 32'b00000000000000010010100011100010;
assign LUT_3[64951] = 32'b00000000000000011001001110111111;
assign LUT_3[64952] = 32'b00000000000000011000100111001110;
assign LUT_3[64953] = 32'b00000000000000011111010010101011;
assign LUT_3[64954] = 32'b00000000000000011010101110110010;
assign LUT_3[64955] = 32'b00000000000000100001011010001111;
assign LUT_3[64956] = 32'b00000000000000010101110101000100;
assign LUT_3[64957] = 32'b00000000000000011100100000100001;
assign LUT_3[64958] = 32'b00000000000000010111111100101000;
assign LUT_3[64959] = 32'b00000000000000011110101000000101;
assign LUT_3[64960] = 32'b00000000000000001110100101010000;
assign LUT_3[64961] = 32'b00000000000000010101010000101101;
assign LUT_3[64962] = 32'b00000000000000010000101100110100;
assign LUT_3[64963] = 32'b00000000000000010111011000010001;
assign LUT_3[64964] = 32'b00000000000000001011110011000110;
assign LUT_3[64965] = 32'b00000000000000010010011110100011;
assign LUT_3[64966] = 32'b00000000000000001101111010101010;
assign LUT_3[64967] = 32'b00000000000000010100100110000111;
assign LUT_3[64968] = 32'b00000000000000010011111110010110;
assign LUT_3[64969] = 32'b00000000000000011010101001110011;
assign LUT_3[64970] = 32'b00000000000000010110000101111010;
assign LUT_3[64971] = 32'b00000000000000011100110001010111;
assign LUT_3[64972] = 32'b00000000000000010001001100001100;
assign LUT_3[64973] = 32'b00000000000000010111110111101001;
assign LUT_3[64974] = 32'b00000000000000010011010011110000;
assign LUT_3[64975] = 32'b00000000000000011001111111001101;
assign LUT_3[64976] = 32'b00000000000000010001111000010011;
assign LUT_3[64977] = 32'b00000000000000011000100011110000;
assign LUT_3[64978] = 32'b00000000000000010011111111110111;
assign LUT_3[64979] = 32'b00000000000000011010101011010100;
assign LUT_3[64980] = 32'b00000000000000001111000110001001;
assign LUT_3[64981] = 32'b00000000000000010101110001100110;
assign LUT_3[64982] = 32'b00000000000000010001001101101101;
assign LUT_3[64983] = 32'b00000000000000010111111001001010;
assign LUT_3[64984] = 32'b00000000000000010111010001011001;
assign LUT_3[64985] = 32'b00000000000000011101111100110110;
assign LUT_3[64986] = 32'b00000000000000011001011000111101;
assign LUT_3[64987] = 32'b00000000000000100000000100011010;
assign LUT_3[64988] = 32'b00000000000000010100011111001111;
assign LUT_3[64989] = 32'b00000000000000011011001010101100;
assign LUT_3[64990] = 32'b00000000000000010110100110110011;
assign LUT_3[64991] = 32'b00000000000000011101010010010000;
assign LUT_3[64992] = 32'b00000000000000001111110011110000;
assign LUT_3[64993] = 32'b00000000000000010110011111001101;
assign LUT_3[64994] = 32'b00000000000000010001111011010100;
assign LUT_3[64995] = 32'b00000000000000011000100110110001;
assign LUT_3[64996] = 32'b00000000000000001101000001100110;
assign LUT_3[64997] = 32'b00000000000000010011101101000011;
assign LUT_3[64998] = 32'b00000000000000001111001001001010;
assign LUT_3[64999] = 32'b00000000000000010101110100100111;
assign LUT_3[65000] = 32'b00000000000000010101001100110110;
assign LUT_3[65001] = 32'b00000000000000011011111000010011;
assign LUT_3[65002] = 32'b00000000000000010111010100011010;
assign LUT_3[65003] = 32'b00000000000000011101111111110111;
assign LUT_3[65004] = 32'b00000000000000010010011010101100;
assign LUT_3[65005] = 32'b00000000000000011001000110001001;
assign LUT_3[65006] = 32'b00000000000000010100100010010000;
assign LUT_3[65007] = 32'b00000000000000011011001101101101;
assign LUT_3[65008] = 32'b00000000000000010011000110110011;
assign LUT_3[65009] = 32'b00000000000000011001110010010000;
assign LUT_3[65010] = 32'b00000000000000010101001110010111;
assign LUT_3[65011] = 32'b00000000000000011011111001110100;
assign LUT_3[65012] = 32'b00000000000000010000010100101001;
assign LUT_3[65013] = 32'b00000000000000010111000000000110;
assign LUT_3[65014] = 32'b00000000000000010010011100001101;
assign LUT_3[65015] = 32'b00000000000000011001000111101010;
assign LUT_3[65016] = 32'b00000000000000011000011111111001;
assign LUT_3[65017] = 32'b00000000000000011111001011010110;
assign LUT_3[65018] = 32'b00000000000000011010100111011101;
assign LUT_3[65019] = 32'b00000000000000100001010010111010;
assign LUT_3[65020] = 32'b00000000000000010101101101101111;
assign LUT_3[65021] = 32'b00000000000000011100011001001100;
assign LUT_3[65022] = 32'b00000000000000010111110101010011;
assign LUT_3[65023] = 32'b00000000000000011110100000110000;
assign LUT_3[65024] = 32'b00000000000000010011100111010010;
assign LUT_3[65025] = 32'b00000000000000011010010010101111;
assign LUT_3[65026] = 32'b00000000000000010101101110110110;
assign LUT_3[65027] = 32'b00000000000000011100011010010011;
assign LUT_3[65028] = 32'b00000000000000010000110101001000;
assign LUT_3[65029] = 32'b00000000000000010111100000100101;
assign LUT_3[65030] = 32'b00000000000000010010111100101100;
assign LUT_3[65031] = 32'b00000000000000011001101000001001;
assign LUT_3[65032] = 32'b00000000000000011001000000011000;
assign LUT_3[65033] = 32'b00000000000000011111101011110101;
assign LUT_3[65034] = 32'b00000000000000011011000111111100;
assign LUT_3[65035] = 32'b00000000000000100001110011011001;
assign LUT_3[65036] = 32'b00000000000000010110001110001110;
assign LUT_3[65037] = 32'b00000000000000011100111001101011;
assign LUT_3[65038] = 32'b00000000000000011000010101110010;
assign LUT_3[65039] = 32'b00000000000000011111000001001111;
assign LUT_3[65040] = 32'b00000000000000010110111010010101;
assign LUT_3[65041] = 32'b00000000000000011101100101110010;
assign LUT_3[65042] = 32'b00000000000000011001000001111001;
assign LUT_3[65043] = 32'b00000000000000011111101101010110;
assign LUT_3[65044] = 32'b00000000000000010100001000001011;
assign LUT_3[65045] = 32'b00000000000000011010110011101000;
assign LUT_3[65046] = 32'b00000000000000010110001111101111;
assign LUT_3[65047] = 32'b00000000000000011100111011001100;
assign LUT_3[65048] = 32'b00000000000000011100010011011011;
assign LUT_3[65049] = 32'b00000000000000100010111110111000;
assign LUT_3[65050] = 32'b00000000000000011110011010111111;
assign LUT_3[65051] = 32'b00000000000000100101000110011100;
assign LUT_3[65052] = 32'b00000000000000011001100001010001;
assign LUT_3[65053] = 32'b00000000000000100000001100101110;
assign LUT_3[65054] = 32'b00000000000000011011101000110101;
assign LUT_3[65055] = 32'b00000000000000100010010100010010;
assign LUT_3[65056] = 32'b00000000000000010100110101110010;
assign LUT_3[65057] = 32'b00000000000000011011100001001111;
assign LUT_3[65058] = 32'b00000000000000010110111101010110;
assign LUT_3[65059] = 32'b00000000000000011101101000110011;
assign LUT_3[65060] = 32'b00000000000000010010000011101000;
assign LUT_3[65061] = 32'b00000000000000011000101111000101;
assign LUT_3[65062] = 32'b00000000000000010100001011001100;
assign LUT_3[65063] = 32'b00000000000000011010110110101001;
assign LUT_3[65064] = 32'b00000000000000011010001110111000;
assign LUT_3[65065] = 32'b00000000000000100000111010010101;
assign LUT_3[65066] = 32'b00000000000000011100010110011100;
assign LUT_3[65067] = 32'b00000000000000100011000001111001;
assign LUT_3[65068] = 32'b00000000000000010111011100101110;
assign LUT_3[65069] = 32'b00000000000000011110001000001011;
assign LUT_3[65070] = 32'b00000000000000011001100100010010;
assign LUT_3[65071] = 32'b00000000000000100000001111101111;
assign LUT_3[65072] = 32'b00000000000000011000001000110101;
assign LUT_3[65073] = 32'b00000000000000011110110100010010;
assign LUT_3[65074] = 32'b00000000000000011010010000011001;
assign LUT_3[65075] = 32'b00000000000000100000111011110110;
assign LUT_3[65076] = 32'b00000000000000010101010110101011;
assign LUT_3[65077] = 32'b00000000000000011100000010001000;
assign LUT_3[65078] = 32'b00000000000000010111011110001111;
assign LUT_3[65079] = 32'b00000000000000011110001001101100;
assign LUT_3[65080] = 32'b00000000000000011101100001111011;
assign LUT_3[65081] = 32'b00000000000000100100001101011000;
assign LUT_3[65082] = 32'b00000000000000011111101001011111;
assign LUT_3[65083] = 32'b00000000000000100110010100111100;
assign LUT_3[65084] = 32'b00000000000000011010101111110001;
assign LUT_3[65085] = 32'b00000000000000100001011011001110;
assign LUT_3[65086] = 32'b00000000000000011100110111010101;
assign LUT_3[65087] = 32'b00000000000000100011100010110010;
assign LUT_3[65088] = 32'b00000000000000010011011111111101;
assign LUT_3[65089] = 32'b00000000000000011010001011011010;
assign LUT_3[65090] = 32'b00000000000000010101100111100001;
assign LUT_3[65091] = 32'b00000000000000011100010010111110;
assign LUT_3[65092] = 32'b00000000000000010000101101110011;
assign LUT_3[65093] = 32'b00000000000000010111011001010000;
assign LUT_3[65094] = 32'b00000000000000010010110101010111;
assign LUT_3[65095] = 32'b00000000000000011001100000110100;
assign LUT_3[65096] = 32'b00000000000000011000111001000011;
assign LUT_3[65097] = 32'b00000000000000011111100100100000;
assign LUT_3[65098] = 32'b00000000000000011011000000100111;
assign LUT_3[65099] = 32'b00000000000000100001101100000100;
assign LUT_3[65100] = 32'b00000000000000010110000110111001;
assign LUT_3[65101] = 32'b00000000000000011100110010010110;
assign LUT_3[65102] = 32'b00000000000000011000001110011101;
assign LUT_3[65103] = 32'b00000000000000011110111001111010;
assign LUT_3[65104] = 32'b00000000000000010110110011000000;
assign LUT_3[65105] = 32'b00000000000000011101011110011101;
assign LUT_3[65106] = 32'b00000000000000011000111010100100;
assign LUT_3[65107] = 32'b00000000000000011111100110000001;
assign LUT_3[65108] = 32'b00000000000000010100000000110110;
assign LUT_3[65109] = 32'b00000000000000011010101100010011;
assign LUT_3[65110] = 32'b00000000000000010110001000011010;
assign LUT_3[65111] = 32'b00000000000000011100110011110111;
assign LUT_3[65112] = 32'b00000000000000011100001100000110;
assign LUT_3[65113] = 32'b00000000000000100010110111100011;
assign LUT_3[65114] = 32'b00000000000000011110010011101010;
assign LUT_3[65115] = 32'b00000000000000100100111111000111;
assign LUT_3[65116] = 32'b00000000000000011001011001111100;
assign LUT_3[65117] = 32'b00000000000000100000000101011001;
assign LUT_3[65118] = 32'b00000000000000011011100001100000;
assign LUT_3[65119] = 32'b00000000000000100010001100111101;
assign LUT_3[65120] = 32'b00000000000000010100101110011101;
assign LUT_3[65121] = 32'b00000000000000011011011001111010;
assign LUT_3[65122] = 32'b00000000000000010110110110000001;
assign LUT_3[65123] = 32'b00000000000000011101100001011110;
assign LUT_3[65124] = 32'b00000000000000010001111100010011;
assign LUT_3[65125] = 32'b00000000000000011000100111110000;
assign LUT_3[65126] = 32'b00000000000000010100000011110111;
assign LUT_3[65127] = 32'b00000000000000011010101111010100;
assign LUT_3[65128] = 32'b00000000000000011010000111100011;
assign LUT_3[65129] = 32'b00000000000000100000110011000000;
assign LUT_3[65130] = 32'b00000000000000011100001111000111;
assign LUT_3[65131] = 32'b00000000000000100010111010100100;
assign LUT_3[65132] = 32'b00000000000000010111010101011001;
assign LUT_3[65133] = 32'b00000000000000011110000000110110;
assign LUT_3[65134] = 32'b00000000000000011001011100111101;
assign LUT_3[65135] = 32'b00000000000000100000001000011010;
assign LUT_3[65136] = 32'b00000000000000011000000001100000;
assign LUT_3[65137] = 32'b00000000000000011110101100111101;
assign LUT_3[65138] = 32'b00000000000000011010001001000100;
assign LUT_3[65139] = 32'b00000000000000100000110100100001;
assign LUT_3[65140] = 32'b00000000000000010101001111010110;
assign LUT_3[65141] = 32'b00000000000000011011111010110011;
assign LUT_3[65142] = 32'b00000000000000010111010110111010;
assign LUT_3[65143] = 32'b00000000000000011110000010010111;
assign LUT_3[65144] = 32'b00000000000000011101011010100110;
assign LUT_3[65145] = 32'b00000000000000100100000110000011;
assign LUT_3[65146] = 32'b00000000000000011111100010001010;
assign LUT_3[65147] = 32'b00000000000000100110001101100111;
assign LUT_3[65148] = 32'b00000000000000011010101000011100;
assign LUT_3[65149] = 32'b00000000000000100001010011111001;
assign LUT_3[65150] = 32'b00000000000000011100110000000000;
assign LUT_3[65151] = 32'b00000000000000100011011011011101;
assign LUT_3[65152] = 32'b00000000000000010101110010010000;
assign LUT_3[65153] = 32'b00000000000000011100011101101101;
assign LUT_3[65154] = 32'b00000000000000010111111001110100;
assign LUT_3[65155] = 32'b00000000000000011110100101010001;
assign LUT_3[65156] = 32'b00000000000000010011000000000110;
assign LUT_3[65157] = 32'b00000000000000011001101011100011;
assign LUT_3[65158] = 32'b00000000000000010101000111101010;
assign LUT_3[65159] = 32'b00000000000000011011110011000111;
assign LUT_3[65160] = 32'b00000000000000011011001011010110;
assign LUT_3[65161] = 32'b00000000000000100001110110110011;
assign LUT_3[65162] = 32'b00000000000000011101010010111010;
assign LUT_3[65163] = 32'b00000000000000100011111110010111;
assign LUT_3[65164] = 32'b00000000000000011000011001001100;
assign LUT_3[65165] = 32'b00000000000000011111000100101001;
assign LUT_3[65166] = 32'b00000000000000011010100000110000;
assign LUT_3[65167] = 32'b00000000000000100001001100001101;
assign LUT_3[65168] = 32'b00000000000000011001000101010011;
assign LUT_3[65169] = 32'b00000000000000011111110000110000;
assign LUT_3[65170] = 32'b00000000000000011011001100110111;
assign LUT_3[65171] = 32'b00000000000000100001111000010100;
assign LUT_3[65172] = 32'b00000000000000010110010011001001;
assign LUT_3[65173] = 32'b00000000000000011100111110100110;
assign LUT_3[65174] = 32'b00000000000000011000011010101101;
assign LUT_3[65175] = 32'b00000000000000011111000110001010;
assign LUT_3[65176] = 32'b00000000000000011110011110011001;
assign LUT_3[65177] = 32'b00000000000000100101001001110110;
assign LUT_3[65178] = 32'b00000000000000100000100101111101;
assign LUT_3[65179] = 32'b00000000000000100111010001011010;
assign LUT_3[65180] = 32'b00000000000000011011101100001111;
assign LUT_3[65181] = 32'b00000000000000100010010111101100;
assign LUT_3[65182] = 32'b00000000000000011101110011110011;
assign LUT_3[65183] = 32'b00000000000000100100011111010000;
assign LUT_3[65184] = 32'b00000000000000010111000000110000;
assign LUT_3[65185] = 32'b00000000000000011101101100001101;
assign LUT_3[65186] = 32'b00000000000000011001001000010100;
assign LUT_3[65187] = 32'b00000000000000011111110011110001;
assign LUT_3[65188] = 32'b00000000000000010100001110100110;
assign LUT_3[65189] = 32'b00000000000000011010111010000011;
assign LUT_3[65190] = 32'b00000000000000010110010110001010;
assign LUT_3[65191] = 32'b00000000000000011101000001100111;
assign LUT_3[65192] = 32'b00000000000000011100011001110110;
assign LUT_3[65193] = 32'b00000000000000100011000101010011;
assign LUT_3[65194] = 32'b00000000000000011110100001011010;
assign LUT_3[65195] = 32'b00000000000000100101001100110111;
assign LUT_3[65196] = 32'b00000000000000011001100111101100;
assign LUT_3[65197] = 32'b00000000000000100000010011001001;
assign LUT_3[65198] = 32'b00000000000000011011101111010000;
assign LUT_3[65199] = 32'b00000000000000100010011010101101;
assign LUT_3[65200] = 32'b00000000000000011010010011110011;
assign LUT_3[65201] = 32'b00000000000000100000111111010000;
assign LUT_3[65202] = 32'b00000000000000011100011011010111;
assign LUT_3[65203] = 32'b00000000000000100011000110110100;
assign LUT_3[65204] = 32'b00000000000000010111100001101001;
assign LUT_3[65205] = 32'b00000000000000011110001101000110;
assign LUT_3[65206] = 32'b00000000000000011001101001001101;
assign LUT_3[65207] = 32'b00000000000000100000010100101010;
assign LUT_3[65208] = 32'b00000000000000011111101100111001;
assign LUT_3[65209] = 32'b00000000000000100110011000010110;
assign LUT_3[65210] = 32'b00000000000000100001110100011101;
assign LUT_3[65211] = 32'b00000000000000101000011111111010;
assign LUT_3[65212] = 32'b00000000000000011100111010101111;
assign LUT_3[65213] = 32'b00000000000000100011100110001100;
assign LUT_3[65214] = 32'b00000000000000011111000010010011;
assign LUT_3[65215] = 32'b00000000000000100101101101110000;
assign LUT_3[65216] = 32'b00000000000000010101101010111011;
assign LUT_3[65217] = 32'b00000000000000011100010110011000;
assign LUT_3[65218] = 32'b00000000000000010111110010011111;
assign LUT_3[65219] = 32'b00000000000000011110011101111100;
assign LUT_3[65220] = 32'b00000000000000010010111000110001;
assign LUT_3[65221] = 32'b00000000000000011001100100001110;
assign LUT_3[65222] = 32'b00000000000000010101000000010101;
assign LUT_3[65223] = 32'b00000000000000011011101011110010;
assign LUT_3[65224] = 32'b00000000000000011011000100000001;
assign LUT_3[65225] = 32'b00000000000000100001101111011110;
assign LUT_3[65226] = 32'b00000000000000011101001011100101;
assign LUT_3[65227] = 32'b00000000000000100011110111000010;
assign LUT_3[65228] = 32'b00000000000000011000010001110111;
assign LUT_3[65229] = 32'b00000000000000011110111101010100;
assign LUT_3[65230] = 32'b00000000000000011010011001011011;
assign LUT_3[65231] = 32'b00000000000000100001000100111000;
assign LUT_3[65232] = 32'b00000000000000011000111101111110;
assign LUT_3[65233] = 32'b00000000000000011111101001011011;
assign LUT_3[65234] = 32'b00000000000000011011000101100010;
assign LUT_3[65235] = 32'b00000000000000100001110000111111;
assign LUT_3[65236] = 32'b00000000000000010110001011110100;
assign LUT_3[65237] = 32'b00000000000000011100110111010001;
assign LUT_3[65238] = 32'b00000000000000011000010011011000;
assign LUT_3[65239] = 32'b00000000000000011110111110110101;
assign LUT_3[65240] = 32'b00000000000000011110010111000100;
assign LUT_3[65241] = 32'b00000000000000100101000010100001;
assign LUT_3[65242] = 32'b00000000000000100000011110101000;
assign LUT_3[65243] = 32'b00000000000000100111001010000101;
assign LUT_3[65244] = 32'b00000000000000011011100100111010;
assign LUT_3[65245] = 32'b00000000000000100010010000010111;
assign LUT_3[65246] = 32'b00000000000000011101101100011110;
assign LUT_3[65247] = 32'b00000000000000100100010111111011;
assign LUT_3[65248] = 32'b00000000000000010110111001011011;
assign LUT_3[65249] = 32'b00000000000000011101100100111000;
assign LUT_3[65250] = 32'b00000000000000011001000000111111;
assign LUT_3[65251] = 32'b00000000000000011111101100011100;
assign LUT_3[65252] = 32'b00000000000000010100000111010001;
assign LUT_3[65253] = 32'b00000000000000011010110010101110;
assign LUT_3[65254] = 32'b00000000000000010110001110110101;
assign LUT_3[65255] = 32'b00000000000000011100111010010010;
assign LUT_3[65256] = 32'b00000000000000011100010010100001;
assign LUT_3[65257] = 32'b00000000000000100010111101111110;
assign LUT_3[65258] = 32'b00000000000000011110011010000101;
assign LUT_3[65259] = 32'b00000000000000100101000101100010;
assign LUT_3[65260] = 32'b00000000000000011001100000010111;
assign LUT_3[65261] = 32'b00000000000000100000001011110100;
assign LUT_3[65262] = 32'b00000000000000011011100111111011;
assign LUT_3[65263] = 32'b00000000000000100010010011011000;
assign LUT_3[65264] = 32'b00000000000000011010001100011110;
assign LUT_3[65265] = 32'b00000000000000100000110111111011;
assign LUT_3[65266] = 32'b00000000000000011100010100000010;
assign LUT_3[65267] = 32'b00000000000000100010111111011111;
assign LUT_3[65268] = 32'b00000000000000010111011010010100;
assign LUT_3[65269] = 32'b00000000000000011110000101110001;
assign LUT_3[65270] = 32'b00000000000000011001100001111000;
assign LUT_3[65271] = 32'b00000000000000100000001101010101;
assign LUT_3[65272] = 32'b00000000000000011111100101100100;
assign LUT_3[65273] = 32'b00000000000000100110010001000001;
assign LUT_3[65274] = 32'b00000000000000100001101101001000;
assign LUT_3[65275] = 32'b00000000000000101000011000100101;
assign LUT_3[65276] = 32'b00000000000000011100110011011010;
assign LUT_3[65277] = 32'b00000000000000100011011110110111;
assign LUT_3[65278] = 32'b00000000000000011110111010111110;
assign LUT_3[65279] = 32'b00000000000000100101100110011011;
assign LUT_3[65280] = 32'b00000000000000001111110110110011;
assign LUT_3[65281] = 32'b00000000000000010110100010010000;
assign LUT_3[65282] = 32'b00000000000000010001111110010111;
assign LUT_3[65283] = 32'b00000000000000011000101001110100;
assign LUT_3[65284] = 32'b00000000000000001101000100101001;
assign LUT_3[65285] = 32'b00000000000000010011110000000110;
assign LUT_3[65286] = 32'b00000000000000001111001100001101;
assign LUT_3[65287] = 32'b00000000000000010101110111101010;
assign LUT_3[65288] = 32'b00000000000000010101001111111001;
assign LUT_3[65289] = 32'b00000000000000011011111011010110;
assign LUT_3[65290] = 32'b00000000000000010111010111011101;
assign LUT_3[65291] = 32'b00000000000000011110000010111010;
assign LUT_3[65292] = 32'b00000000000000010010011101101111;
assign LUT_3[65293] = 32'b00000000000000011001001001001100;
assign LUT_3[65294] = 32'b00000000000000010100100101010011;
assign LUT_3[65295] = 32'b00000000000000011011010000110000;
assign LUT_3[65296] = 32'b00000000000000010011001001110110;
assign LUT_3[65297] = 32'b00000000000000011001110101010011;
assign LUT_3[65298] = 32'b00000000000000010101010001011010;
assign LUT_3[65299] = 32'b00000000000000011011111100110111;
assign LUT_3[65300] = 32'b00000000000000010000010111101100;
assign LUT_3[65301] = 32'b00000000000000010111000011001001;
assign LUT_3[65302] = 32'b00000000000000010010011111010000;
assign LUT_3[65303] = 32'b00000000000000011001001010101101;
assign LUT_3[65304] = 32'b00000000000000011000100010111100;
assign LUT_3[65305] = 32'b00000000000000011111001110011001;
assign LUT_3[65306] = 32'b00000000000000011010101010100000;
assign LUT_3[65307] = 32'b00000000000000100001010101111101;
assign LUT_3[65308] = 32'b00000000000000010101110000110010;
assign LUT_3[65309] = 32'b00000000000000011100011100001111;
assign LUT_3[65310] = 32'b00000000000000010111111000010110;
assign LUT_3[65311] = 32'b00000000000000011110100011110011;
assign LUT_3[65312] = 32'b00000000000000010001000101010011;
assign LUT_3[65313] = 32'b00000000000000010111110000110000;
assign LUT_3[65314] = 32'b00000000000000010011001100110111;
assign LUT_3[65315] = 32'b00000000000000011001111000010100;
assign LUT_3[65316] = 32'b00000000000000001110010011001001;
assign LUT_3[65317] = 32'b00000000000000010100111110100110;
assign LUT_3[65318] = 32'b00000000000000010000011010101101;
assign LUT_3[65319] = 32'b00000000000000010111000110001010;
assign LUT_3[65320] = 32'b00000000000000010110011110011001;
assign LUT_3[65321] = 32'b00000000000000011101001001110110;
assign LUT_3[65322] = 32'b00000000000000011000100101111101;
assign LUT_3[65323] = 32'b00000000000000011111010001011010;
assign LUT_3[65324] = 32'b00000000000000010011101100001111;
assign LUT_3[65325] = 32'b00000000000000011010010111101100;
assign LUT_3[65326] = 32'b00000000000000010101110011110011;
assign LUT_3[65327] = 32'b00000000000000011100011111010000;
assign LUT_3[65328] = 32'b00000000000000010100011000010110;
assign LUT_3[65329] = 32'b00000000000000011011000011110011;
assign LUT_3[65330] = 32'b00000000000000010110011111111010;
assign LUT_3[65331] = 32'b00000000000000011101001011010111;
assign LUT_3[65332] = 32'b00000000000000010001100110001100;
assign LUT_3[65333] = 32'b00000000000000011000010001101001;
assign LUT_3[65334] = 32'b00000000000000010011101101110000;
assign LUT_3[65335] = 32'b00000000000000011010011001001101;
assign LUT_3[65336] = 32'b00000000000000011001110001011100;
assign LUT_3[65337] = 32'b00000000000000100000011100111001;
assign LUT_3[65338] = 32'b00000000000000011011111001000000;
assign LUT_3[65339] = 32'b00000000000000100010100100011101;
assign LUT_3[65340] = 32'b00000000000000010110111111010010;
assign LUT_3[65341] = 32'b00000000000000011101101010101111;
assign LUT_3[65342] = 32'b00000000000000011001000110110110;
assign LUT_3[65343] = 32'b00000000000000011111110010010011;
assign LUT_3[65344] = 32'b00000000000000001111101111011110;
assign LUT_3[65345] = 32'b00000000000000010110011010111011;
assign LUT_3[65346] = 32'b00000000000000010001110111000010;
assign LUT_3[65347] = 32'b00000000000000011000100010011111;
assign LUT_3[65348] = 32'b00000000000000001100111101010100;
assign LUT_3[65349] = 32'b00000000000000010011101000110001;
assign LUT_3[65350] = 32'b00000000000000001111000100111000;
assign LUT_3[65351] = 32'b00000000000000010101110000010101;
assign LUT_3[65352] = 32'b00000000000000010101001000100100;
assign LUT_3[65353] = 32'b00000000000000011011110100000001;
assign LUT_3[65354] = 32'b00000000000000010111010000001000;
assign LUT_3[65355] = 32'b00000000000000011101111011100101;
assign LUT_3[65356] = 32'b00000000000000010010010110011010;
assign LUT_3[65357] = 32'b00000000000000011001000001110111;
assign LUT_3[65358] = 32'b00000000000000010100011101111110;
assign LUT_3[65359] = 32'b00000000000000011011001001011011;
assign LUT_3[65360] = 32'b00000000000000010011000010100001;
assign LUT_3[65361] = 32'b00000000000000011001101101111110;
assign LUT_3[65362] = 32'b00000000000000010101001010000101;
assign LUT_3[65363] = 32'b00000000000000011011110101100010;
assign LUT_3[65364] = 32'b00000000000000010000010000010111;
assign LUT_3[65365] = 32'b00000000000000010110111011110100;
assign LUT_3[65366] = 32'b00000000000000010010010111111011;
assign LUT_3[65367] = 32'b00000000000000011001000011011000;
assign LUT_3[65368] = 32'b00000000000000011000011011100111;
assign LUT_3[65369] = 32'b00000000000000011111000111000100;
assign LUT_3[65370] = 32'b00000000000000011010100011001011;
assign LUT_3[65371] = 32'b00000000000000100001001110101000;
assign LUT_3[65372] = 32'b00000000000000010101101001011101;
assign LUT_3[65373] = 32'b00000000000000011100010100111010;
assign LUT_3[65374] = 32'b00000000000000010111110001000001;
assign LUT_3[65375] = 32'b00000000000000011110011100011110;
assign LUT_3[65376] = 32'b00000000000000010000111101111110;
assign LUT_3[65377] = 32'b00000000000000010111101001011011;
assign LUT_3[65378] = 32'b00000000000000010011000101100010;
assign LUT_3[65379] = 32'b00000000000000011001110000111111;
assign LUT_3[65380] = 32'b00000000000000001110001011110100;
assign LUT_3[65381] = 32'b00000000000000010100110111010001;
assign LUT_3[65382] = 32'b00000000000000010000010011011000;
assign LUT_3[65383] = 32'b00000000000000010110111110110101;
assign LUT_3[65384] = 32'b00000000000000010110010111000100;
assign LUT_3[65385] = 32'b00000000000000011101000010100001;
assign LUT_3[65386] = 32'b00000000000000011000011110101000;
assign LUT_3[65387] = 32'b00000000000000011111001010000101;
assign LUT_3[65388] = 32'b00000000000000010011100100111010;
assign LUT_3[65389] = 32'b00000000000000011010010000010111;
assign LUT_3[65390] = 32'b00000000000000010101101100011110;
assign LUT_3[65391] = 32'b00000000000000011100010111111011;
assign LUT_3[65392] = 32'b00000000000000010100010001000001;
assign LUT_3[65393] = 32'b00000000000000011010111100011110;
assign LUT_3[65394] = 32'b00000000000000010110011000100101;
assign LUT_3[65395] = 32'b00000000000000011101000100000010;
assign LUT_3[65396] = 32'b00000000000000010001011110110111;
assign LUT_3[65397] = 32'b00000000000000011000001010010100;
assign LUT_3[65398] = 32'b00000000000000010011100110011011;
assign LUT_3[65399] = 32'b00000000000000011010010001111000;
assign LUT_3[65400] = 32'b00000000000000011001101010000111;
assign LUT_3[65401] = 32'b00000000000000100000010101100100;
assign LUT_3[65402] = 32'b00000000000000011011110001101011;
assign LUT_3[65403] = 32'b00000000000000100010011101001000;
assign LUT_3[65404] = 32'b00000000000000010110110111111101;
assign LUT_3[65405] = 32'b00000000000000011101100011011010;
assign LUT_3[65406] = 32'b00000000000000011000111111100001;
assign LUT_3[65407] = 32'b00000000000000011111101010111110;
assign LUT_3[65408] = 32'b00000000000000010010000001110001;
assign LUT_3[65409] = 32'b00000000000000011000101101001110;
assign LUT_3[65410] = 32'b00000000000000010100001001010101;
assign LUT_3[65411] = 32'b00000000000000011010110100110010;
assign LUT_3[65412] = 32'b00000000000000001111001111100111;
assign LUT_3[65413] = 32'b00000000000000010101111011000100;
assign LUT_3[65414] = 32'b00000000000000010001010111001011;
assign LUT_3[65415] = 32'b00000000000000011000000010101000;
assign LUT_3[65416] = 32'b00000000000000010111011010110111;
assign LUT_3[65417] = 32'b00000000000000011110000110010100;
assign LUT_3[65418] = 32'b00000000000000011001100010011011;
assign LUT_3[65419] = 32'b00000000000000100000001101111000;
assign LUT_3[65420] = 32'b00000000000000010100101000101101;
assign LUT_3[65421] = 32'b00000000000000011011010100001010;
assign LUT_3[65422] = 32'b00000000000000010110110000010001;
assign LUT_3[65423] = 32'b00000000000000011101011011101110;
assign LUT_3[65424] = 32'b00000000000000010101010100110100;
assign LUT_3[65425] = 32'b00000000000000011100000000010001;
assign LUT_3[65426] = 32'b00000000000000010111011100011000;
assign LUT_3[65427] = 32'b00000000000000011110000111110101;
assign LUT_3[65428] = 32'b00000000000000010010100010101010;
assign LUT_3[65429] = 32'b00000000000000011001001110000111;
assign LUT_3[65430] = 32'b00000000000000010100101010001110;
assign LUT_3[65431] = 32'b00000000000000011011010101101011;
assign LUT_3[65432] = 32'b00000000000000011010101101111010;
assign LUT_3[65433] = 32'b00000000000000100001011001010111;
assign LUT_3[65434] = 32'b00000000000000011100110101011110;
assign LUT_3[65435] = 32'b00000000000000100011100000111011;
assign LUT_3[65436] = 32'b00000000000000010111111011110000;
assign LUT_3[65437] = 32'b00000000000000011110100111001101;
assign LUT_3[65438] = 32'b00000000000000011010000011010100;
assign LUT_3[65439] = 32'b00000000000000100000101110110001;
assign LUT_3[65440] = 32'b00000000000000010011010000010001;
assign LUT_3[65441] = 32'b00000000000000011001111011101110;
assign LUT_3[65442] = 32'b00000000000000010101010111110101;
assign LUT_3[65443] = 32'b00000000000000011100000011010010;
assign LUT_3[65444] = 32'b00000000000000010000011110000111;
assign LUT_3[65445] = 32'b00000000000000010111001001100100;
assign LUT_3[65446] = 32'b00000000000000010010100101101011;
assign LUT_3[65447] = 32'b00000000000000011001010001001000;
assign LUT_3[65448] = 32'b00000000000000011000101001010111;
assign LUT_3[65449] = 32'b00000000000000011111010100110100;
assign LUT_3[65450] = 32'b00000000000000011010110000111011;
assign LUT_3[65451] = 32'b00000000000000100001011100011000;
assign LUT_3[65452] = 32'b00000000000000010101110111001101;
assign LUT_3[65453] = 32'b00000000000000011100100010101010;
assign LUT_3[65454] = 32'b00000000000000010111111110110001;
assign LUT_3[65455] = 32'b00000000000000011110101010001110;
assign LUT_3[65456] = 32'b00000000000000010110100011010100;
assign LUT_3[65457] = 32'b00000000000000011101001110110001;
assign LUT_3[65458] = 32'b00000000000000011000101010111000;
assign LUT_3[65459] = 32'b00000000000000011111010110010101;
assign LUT_3[65460] = 32'b00000000000000010011110001001010;
assign LUT_3[65461] = 32'b00000000000000011010011100100111;
assign LUT_3[65462] = 32'b00000000000000010101111000101110;
assign LUT_3[65463] = 32'b00000000000000011100100100001011;
assign LUT_3[65464] = 32'b00000000000000011011111100011010;
assign LUT_3[65465] = 32'b00000000000000100010100111110111;
assign LUT_3[65466] = 32'b00000000000000011110000011111110;
assign LUT_3[65467] = 32'b00000000000000100100101111011011;
assign LUT_3[65468] = 32'b00000000000000011001001010010000;
assign LUT_3[65469] = 32'b00000000000000011111110101101101;
assign LUT_3[65470] = 32'b00000000000000011011010001110100;
assign LUT_3[65471] = 32'b00000000000000100001111101010001;
assign LUT_3[65472] = 32'b00000000000000010001111010011100;
assign LUT_3[65473] = 32'b00000000000000011000100101111001;
assign LUT_3[65474] = 32'b00000000000000010100000010000000;
assign LUT_3[65475] = 32'b00000000000000011010101101011101;
assign LUT_3[65476] = 32'b00000000000000001111001000010010;
assign LUT_3[65477] = 32'b00000000000000010101110011101111;
assign LUT_3[65478] = 32'b00000000000000010001001111110110;
assign LUT_3[65479] = 32'b00000000000000010111111011010011;
assign LUT_3[65480] = 32'b00000000000000010111010011100010;
assign LUT_3[65481] = 32'b00000000000000011101111110111111;
assign LUT_3[65482] = 32'b00000000000000011001011011000110;
assign LUT_3[65483] = 32'b00000000000000100000000110100011;
assign LUT_3[65484] = 32'b00000000000000010100100001011000;
assign LUT_3[65485] = 32'b00000000000000011011001100110101;
assign LUT_3[65486] = 32'b00000000000000010110101000111100;
assign LUT_3[65487] = 32'b00000000000000011101010100011001;
assign LUT_3[65488] = 32'b00000000000000010101001101011111;
assign LUT_3[65489] = 32'b00000000000000011011111000111100;
assign LUT_3[65490] = 32'b00000000000000010111010101000011;
assign LUT_3[65491] = 32'b00000000000000011110000000100000;
assign LUT_3[65492] = 32'b00000000000000010010011011010101;
assign LUT_3[65493] = 32'b00000000000000011001000110110010;
assign LUT_3[65494] = 32'b00000000000000010100100010111001;
assign LUT_3[65495] = 32'b00000000000000011011001110010110;
assign LUT_3[65496] = 32'b00000000000000011010100110100101;
assign LUT_3[65497] = 32'b00000000000000100001010010000010;
assign LUT_3[65498] = 32'b00000000000000011100101110001001;
assign LUT_3[65499] = 32'b00000000000000100011011001100110;
assign LUT_3[65500] = 32'b00000000000000010111110100011011;
assign LUT_3[65501] = 32'b00000000000000011110011111111000;
assign LUT_3[65502] = 32'b00000000000000011001111011111111;
assign LUT_3[65503] = 32'b00000000000000100000100111011100;
assign LUT_3[65504] = 32'b00000000000000010011001000111100;
assign LUT_3[65505] = 32'b00000000000000011001110100011001;
assign LUT_3[65506] = 32'b00000000000000010101010000100000;
assign LUT_3[65507] = 32'b00000000000000011011111011111101;
assign LUT_3[65508] = 32'b00000000000000010000010110110010;
assign LUT_3[65509] = 32'b00000000000000010111000010001111;
assign LUT_3[65510] = 32'b00000000000000010010011110010110;
assign LUT_3[65511] = 32'b00000000000000011001001001110011;
assign LUT_3[65512] = 32'b00000000000000011000100010000010;
assign LUT_3[65513] = 32'b00000000000000011111001101011111;
assign LUT_3[65514] = 32'b00000000000000011010101001100110;
assign LUT_3[65515] = 32'b00000000000000100001010101000011;
assign LUT_3[65516] = 32'b00000000000000010101101111111000;
assign LUT_3[65517] = 32'b00000000000000011100011011010101;
assign LUT_3[65518] = 32'b00000000000000010111110111011100;
assign LUT_3[65519] = 32'b00000000000000011110100010111001;
assign LUT_3[65520] = 32'b00000000000000010110011011111111;
assign LUT_3[65521] = 32'b00000000000000011101000111011100;
assign LUT_3[65522] = 32'b00000000000000011000100011100011;
assign LUT_3[65523] = 32'b00000000000000011111001111000000;
assign LUT_3[65524] = 32'b00000000000000010011101001110101;
assign LUT_3[65525] = 32'b00000000000000011010010101010010;
assign LUT_3[65526] = 32'b00000000000000010101110001011001;
assign LUT_3[65527] = 32'b00000000000000011100011100110110;
assign LUT_3[65528] = 32'b00000000000000011011110101000101;
assign LUT_3[65529] = 32'b00000000000000100010100000100010;
assign LUT_3[65530] = 32'b00000000000000011101111100101001;
assign LUT_3[65531] = 32'b00000000000000100100101000000110;
assign LUT_3[65532] = 32'b00000000000000011001000010111011;
assign LUT_3[65533] = 32'b00000000000000011111101110011000;
assign LUT_3[65534] = 32'b00000000000000011011001010011111;
assign LUT_3[65535] = 32'b00000000000000100001110101111100;
endmodule
