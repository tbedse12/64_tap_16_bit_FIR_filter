module DA_table_1(table_in_1 , table_out_1);
input  unsigned [15:0]table_in_1;
output [31:0]table_out_1;
wire   [31:0]LUT_1[65535:0]; 
wire   [31:0]table_out_1; 
assign table_out_1 = LUT_1[table_in_1];
assign LUT_1[0] = 32'b00000000000000000000000000000000;
assign LUT_1[1] = 32'b11111111111111111001010001111100;
assign LUT_1[2] = 32'b11111111111111111011101110010001;
assign LUT_1[3] = 32'b11111111111111110101000000001101;
assign LUT_1[4] = 32'b00000000000000000111111001010111;
assign LUT_1[5] = 32'b00000000000000000001001011010011;
assign LUT_1[6] = 32'b00000000000000000011100111101000;
assign LUT_1[7] = 32'b11111111111111111100111001100100;
assign LUT_1[8] = 32'b11111111111111111111001101110101;
assign LUT_1[9] = 32'b11111111111111111000011111110001;
assign LUT_1[10] = 32'b11111111111111111010111100000110;
assign LUT_1[11] = 32'b11111111111111110100001110000010;
assign LUT_1[12] = 32'b00000000000000000111000111001100;
assign LUT_1[13] = 32'b00000000000000000000011001001000;
assign LUT_1[14] = 32'b00000000000000000010110101011101;
assign LUT_1[15] = 32'b11111111111111111100000111011001;
assign LUT_1[16] = 32'b00000000000000000001111011100010;
assign LUT_1[17] = 32'b11111111111111111011001101011110;
assign LUT_1[18] = 32'b11111111111111111101101001110011;
assign LUT_1[19] = 32'b11111111111111110110111011101111;
assign LUT_1[20] = 32'b00000000000000001001110100111001;
assign LUT_1[21] = 32'b00000000000000000011000110110101;
assign LUT_1[22] = 32'b00000000000000000101100011001010;
assign LUT_1[23] = 32'b11111111111111111110110101000110;
assign LUT_1[24] = 32'b00000000000000000001001001010111;
assign LUT_1[25] = 32'b11111111111111111010011011010011;
assign LUT_1[26] = 32'b11111111111111111100110111101000;
assign LUT_1[27] = 32'b11111111111111110110001001100100;
assign LUT_1[28] = 32'b00000000000000001001000010101110;
assign LUT_1[29] = 32'b00000000000000000010010100101010;
assign LUT_1[30] = 32'b00000000000000000100110000111111;
assign LUT_1[31] = 32'b11111111111111111110000010111011;
assign LUT_1[32] = 32'b00000000000000000000111010111111;
assign LUT_1[33] = 32'b11111111111111111010001100111011;
assign LUT_1[34] = 32'b11111111111111111100101001010000;
assign LUT_1[35] = 32'b11111111111111110101111011001100;
assign LUT_1[36] = 32'b00000000000000001000110100010110;
assign LUT_1[37] = 32'b00000000000000000010000110010010;
assign LUT_1[38] = 32'b00000000000000000100100010100111;
assign LUT_1[39] = 32'b11111111111111111101110100100011;
assign LUT_1[40] = 32'b00000000000000000000001000110100;
assign LUT_1[41] = 32'b11111111111111111001011010110000;
assign LUT_1[42] = 32'b11111111111111111011110111000101;
assign LUT_1[43] = 32'b11111111111111110101001001000001;
assign LUT_1[44] = 32'b00000000000000001000000010001011;
assign LUT_1[45] = 32'b00000000000000000001010100000111;
assign LUT_1[46] = 32'b00000000000000000011110000011100;
assign LUT_1[47] = 32'b11111111111111111101000010011000;
assign LUT_1[48] = 32'b00000000000000000010110110100001;
assign LUT_1[49] = 32'b11111111111111111100001000011101;
assign LUT_1[50] = 32'b11111111111111111110100100110010;
assign LUT_1[51] = 32'b11111111111111110111110110101110;
assign LUT_1[52] = 32'b00000000000000001010101111111000;
assign LUT_1[53] = 32'b00000000000000000100000001110100;
assign LUT_1[54] = 32'b00000000000000000110011110001001;
assign LUT_1[55] = 32'b11111111111111111111110000000101;
assign LUT_1[56] = 32'b00000000000000000010000100010110;
assign LUT_1[57] = 32'b11111111111111111011010110010010;
assign LUT_1[58] = 32'b11111111111111111101110010100111;
assign LUT_1[59] = 32'b11111111111111110111000100100011;
assign LUT_1[60] = 32'b00000000000000001001111101101101;
assign LUT_1[61] = 32'b00000000000000000011001111101001;
assign LUT_1[62] = 32'b00000000000000000101101011111110;
assign LUT_1[63] = 32'b11111111111111111110111101111010;
assign LUT_1[64] = 32'b00000000000000000001111101101000;
assign LUT_1[65] = 32'b11111111111111111011001111100100;
assign LUT_1[66] = 32'b11111111111111111101101011111001;
assign LUT_1[67] = 32'b11111111111111110110111101110101;
assign LUT_1[68] = 32'b00000000000000001001110110111111;
assign LUT_1[69] = 32'b00000000000000000011001000111011;
assign LUT_1[70] = 32'b00000000000000000101100101010000;
assign LUT_1[71] = 32'b11111111111111111110110111001100;
assign LUT_1[72] = 32'b00000000000000000001001011011101;
assign LUT_1[73] = 32'b11111111111111111010011101011001;
assign LUT_1[74] = 32'b11111111111111111100111001101110;
assign LUT_1[75] = 32'b11111111111111110110001011101010;
assign LUT_1[76] = 32'b00000000000000001001000100110100;
assign LUT_1[77] = 32'b00000000000000000010010110110000;
assign LUT_1[78] = 32'b00000000000000000100110011000101;
assign LUT_1[79] = 32'b11111111111111111110000101000001;
assign LUT_1[80] = 32'b00000000000000000011111001001010;
assign LUT_1[81] = 32'b11111111111111111101001011000110;
assign LUT_1[82] = 32'b11111111111111111111100111011011;
assign LUT_1[83] = 32'b11111111111111111000111001010111;
assign LUT_1[84] = 32'b00000000000000001011110010100001;
assign LUT_1[85] = 32'b00000000000000000101000100011101;
assign LUT_1[86] = 32'b00000000000000000111100000110010;
assign LUT_1[87] = 32'b00000000000000000000110010101110;
assign LUT_1[88] = 32'b00000000000000000011000110111111;
assign LUT_1[89] = 32'b11111111111111111100011000111011;
assign LUT_1[90] = 32'b11111111111111111110110101010000;
assign LUT_1[91] = 32'b11111111111111111000000111001100;
assign LUT_1[92] = 32'b00000000000000001011000000010110;
assign LUT_1[93] = 32'b00000000000000000100010010010010;
assign LUT_1[94] = 32'b00000000000000000110101110100111;
assign LUT_1[95] = 32'b00000000000000000000000000100011;
assign LUT_1[96] = 32'b00000000000000000010111000100111;
assign LUT_1[97] = 32'b11111111111111111100001010100011;
assign LUT_1[98] = 32'b11111111111111111110100110111000;
assign LUT_1[99] = 32'b11111111111111110111111000110100;
assign LUT_1[100] = 32'b00000000000000001010110001111110;
assign LUT_1[101] = 32'b00000000000000000100000011111010;
assign LUT_1[102] = 32'b00000000000000000110100000001111;
assign LUT_1[103] = 32'b11111111111111111111110010001011;
assign LUT_1[104] = 32'b00000000000000000010000110011100;
assign LUT_1[105] = 32'b11111111111111111011011000011000;
assign LUT_1[106] = 32'b11111111111111111101110100101101;
assign LUT_1[107] = 32'b11111111111111110111000110101001;
assign LUT_1[108] = 32'b00000000000000001001111111110011;
assign LUT_1[109] = 32'b00000000000000000011010001101111;
assign LUT_1[110] = 32'b00000000000000000101101110000100;
assign LUT_1[111] = 32'b11111111111111111111000000000000;
assign LUT_1[112] = 32'b00000000000000000100110100001001;
assign LUT_1[113] = 32'b11111111111111111110000110000101;
assign LUT_1[114] = 32'b00000000000000000000100010011010;
assign LUT_1[115] = 32'b11111111111111111001110100010110;
assign LUT_1[116] = 32'b00000000000000001100101101100000;
assign LUT_1[117] = 32'b00000000000000000101111111011100;
assign LUT_1[118] = 32'b00000000000000001000011011110001;
assign LUT_1[119] = 32'b00000000000000000001101101101101;
assign LUT_1[120] = 32'b00000000000000000100000001111110;
assign LUT_1[121] = 32'b11111111111111111101010011111010;
assign LUT_1[122] = 32'b11111111111111111111110000001111;
assign LUT_1[123] = 32'b11111111111111111001000010001011;
assign LUT_1[124] = 32'b00000000000000001011111011010101;
assign LUT_1[125] = 32'b00000000000000000101001101010001;
assign LUT_1[126] = 32'b00000000000000000111101001100110;
assign LUT_1[127] = 32'b00000000000000000000111011100010;
assign LUT_1[128] = 32'b00000000000000000011000000000011;
assign LUT_1[129] = 32'b11111111111111111100010001111111;
assign LUT_1[130] = 32'b11111111111111111110101110010100;
assign LUT_1[131] = 32'b11111111111111111000000000010000;
assign LUT_1[132] = 32'b00000000000000001010111001011010;
assign LUT_1[133] = 32'b00000000000000000100001011010110;
assign LUT_1[134] = 32'b00000000000000000110100111101011;
assign LUT_1[135] = 32'b11111111111111111111111001100111;
assign LUT_1[136] = 32'b00000000000000000010001101111000;
assign LUT_1[137] = 32'b11111111111111111011011111110100;
assign LUT_1[138] = 32'b11111111111111111101111100001001;
assign LUT_1[139] = 32'b11111111111111110111001110000101;
assign LUT_1[140] = 32'b00000000000000001010000111001111;
assign LUT_1[141] = 32'b00000000000000000011011001001011;
assign LUT_1[142] = 32'b00000000000000000101110101100000;
assign LUT_1[143] = 32'b11111111111111111111000111011100;
assign LUT_1[144] = 32'b00000000000000000100111011100101;
assign LUT_1[145] = 32'b11111111111111111110001101100001;
assign LUT_1[146] = 32'b00000000000000000000101001110110;
assign LUT_1[147] = 32'b11111111111111111001111011110010;
assign LUT_1[148] = 32'b00000000000000001100110100111100;
assign LUT_1[149] = 32'b00000000000000000110000110111000;
assign LUT_1[150] = 32'b00000000000000001000100011001101;
assign LUT_1[151] = 32'b00000000000000000001110101001001;
assign LUT_1[152] = 32'b00000000000000000100001001011010;
assign LUT_1[153] = 32'b11111111111111111101011011010110;
assign LUT_1[154] = 32'b11111111111111111111110111101011;
assign LUT_1[155] = 32'b11111111111111111001001001100111;
assign LUT_1[156] = 32'b00000000000000001100000010110001;
assign LUT_1[157] = 32'b00000000000000000101010100101101;
assign LUT_1[158] = 32'b00000000000000000111110001000010;
assign LUT_1[159] = 32'b00000000000000000001000010111110;
assign LUT_1[160] = 32'b00000000000000000011111011000010;
assign LUT_1[161] = 32'b11111111111111111101001100111110;
assign LUT_1[162] = 32'b11111111111111111111101001010011;
assign LUT_1[163] = 32'b11111111111111111000111011001111;
assign LUT_1[164] = 32'b00000000000000001011110100011001;
assign LUT_1[165] = 32'b00000000000000000101000110010101;
assign LUT_1[166] = 32'b00000000000000000111100010101010;
assign LUT_1[167] = 32'b00000000000000000000110100100110;
assign LUT_1[168] = 32'b00000000000000000011001000110111;
assign LUT_1[169] = 32'b11111111111111111100011010110011;
assign LUT_1[170] = 32'b11111111111111111110110111001000;
assign LUT_1[171] = 32'b11111111111111111000001001000100;
assign LUT_1[172] = 32'b00000000000000001011000010001110;
assign LUT_1[173] = 32'b00000000000000000100010100001010;
assign LUT_1[174] = 32'b00000000000000000110110000011111;
assign LUT_1[175] = 32'b00000000000000000000000010011011;
assign LUT_1[176] = 32'b00000000000000000101110110100100;
assign LUT_1[177] = 32'b11111111111111111111001000100000;
assign LUT_1[178] = 32'b00000000000000000001100100110101;
assign LUT_1[179] = 32'b11111111111111111010110110110001;
assign LUT_1[180] = 32'b00000000000000001101101111111011;
assign LUT_1[181] = 32'b00000000000000000111000001110111;
assign LUT_1[182] = 32'b00000000000000001001011110001100;
assign LUT_1[183] = 32'b00000000000000000010110000001000;
assign LUT_1[184] = 32'b00000000000000000101000100011001;
assign LUT_1[185] = 32'b11111111111111111110010110010101;
assign LUT_1[186] = 32'b00000000000000000000110010101010;
assign LUT_1[187] = 32'b11111111111111111010000100100110;
assign LUT_1[188] = 32'b00000000000000001100111101110000;
assign LUT_1[189] = 32'b00000000000000000110001111101100;
assign LUT_1[190] = 32'b00000000000000001000101100000001;
assign LUT_1[191] = 32'b00000000000000000001111101111101;
assign LUT_1[192] = 32'b00000000000000000100111101101011;
assign LUT_1[193] = 32'b11111111111111111110001111100111;
assign LUT_1[194] = 32'b00000000000000000000101011111100;
assign LUT_1[195] = 32'b11111111111111111001111101111000;
assign LUT_1[196] = 32'b00000000000000001100110111000010;
assign LUT_1[197] = 32'b00000000000000000110001000111110;
assign LUT_1[198] = 32'b00000000000000001000100101010011;
assign LUT_1[199] = 32'b00000000000000000001110111001111;
assign LUT_1[200] = 32'b00000000000000000100001011100000;
assign LUT_1[201] = 32'b11111111111111111101011101011100;
assign LUT_1[202] = 32'b11111111111111111111111001110001;
assign LUT_1[203] = 32'b11111111111111111001001011101101;
assign LUT_1[204] = 32'b00000000000000001100000100110111;
assign LUT_1[205] = 32'b00000000000000000101010110110011;
assign LUT_1[206] = 32'b00000000000000000111110011001000;
assign LUT_1[207] = 32'b00000000000000000001000101000100;
assign LUT_1[208] = 32'b00000000000000000110111001001101;
assign LUT_1[209] = 32'b00000000000000000000001011001001;
assign LUT_1[210] = 32'b00000000000000000010100111011110;
assign LUT_1[211] = 32'b11111111111111111011111001011010;
assign LUT_1[212] = 32'b00000000000000001110110010100100;
assign LUT_1[213] = 32'b00000000000000001000000100100000;
assign LUT_1[214] = 32'b00000000000000001010100000110101;
assign LUT_1[215] = 32'b00000000000000000011110010110001;
assign LUT_1[216] = 32'b00000000000000000110000111000010;
assign LUT_1[217] = 32'b11111111111111111111011000111110;
assign LUT_1[218] = 32'b00000000000000000001110101010011;
assign LUT_1[219] = 32'b11111111111111111011000111001111;
assign LUT_1[220] = 32'b00000000000000001110000000011001;
assign LUT_1[221] = 32'b00000000000000000111010010010101;
assign LUT_1[222] = 32'b00000000000000001001101110101010;
assign LUT_1[223] = 32'b00000000000000000011000000100110;
assign LUT_1[224] = 32'b00000000000000000101111000101010;
assign LUT_1[225] = 32'b11111111111111111111001010100110;
assign LUT_1[226] = 32'b00000000000000000001100110111011;
assign LUT_1[227] = 32'b11111111111111111010111000110111;
assign LUT_1[228] = 32'b00000000000000001101110010000001;
assign LUT_1[229] = 32'b00000000000000000111000011111101;
assign LUT_1[230] = 32'b00000000000000001001100000010010;
assign LUT_1[231] = 32'b00000000000000000010110010001110;
assign LUT_1[232] = 32'b00000000000000000101000110011111;
assign LUT_1[233] = 32'b11111111111111111110011000011011;
assign LUT_1[234] = 32'b00000000000000000000110100110000;
assign LUT_1[235] = 32'b11111111111111111010000110101100;
assign LUT_1[236] = 32'b00000000000000001100111111110110;
assign LUT_1[237] = 32'b00000000000000000110010001110010;
assign LUT_1[238] = 32'b00000000000000001000101110000111;
assign LUT_1[239] = 32'b00000000000000000010000000000011;
assign LUT_1[240] = 32'b00000000000000000111110100001100;
assign LUT_1[241] = 32'b00000000000000000001000110001000;
assign LUT_1[242] = 32'b00000000000000000011100010011101;
assign LUT_1[243] = 32'b11111111111111111100110100011001;
assign LUT_1[244] = 32'b00000000000000001111101101100011;
assign LUT_1[245] = 32'b00000000000000001000111111011111;
assign LUT_1[246] = 32'b00000000000000001011011011110100;
assign LUT_1[247] = 32'b00000000000000000100101101110000;
assign LUT_1[248] = 32'b00000000000000000111000010000001;
assign LUT_1[249] = 32'b00000000000000000000010011111101;
assign LUT_1[250] = 32'b00000000000000000010110000010010;
assign LUT_1[251] = 32'b11111111111111111100000010001110;
assign LUT_1[252] = 32'b00000000000000001110111011011000;
assign LUT_1[253] = 32'b00000000000000001000001101010100;
assign LUT_1[254] = 32'b00000000000000001010101001101001;
assign LUT_1[255] = 32'b00000000000000000011111011100101;
assign LUT_1[256] = 32'b11111111111111111101110100001100;
assign LUT_1[257] = 32'b11111111111111110111000110001000;
assign LUT_1[258] = 32'b11111111111111111001100010011101;
assign LUT_1[259] = 32'b11111111111111110010110100011001;
assign LUT_1[260] = 32'b00000000000000000101101101100011;
assign LUT_1[261] = 32'b11111111111111111110111111011111;
assign LUT_1[262] = 32'b00000000000000000001011011110100;
assign LUT_1[263] = 32'b11111111111111111010101101110000;
assign LUT_1[264] = 32'b11111111111111111101000010000001;
assign LUT_1[265] = 32'b11111111111111110110010011111101;
assign LUT_1[266] = 32'b11111111111111111000110000010010;
assign LUT_1[267] = 32'b11111111111111110010000010001110;
assign LUT_1[268] = 32'b00000000000000000100111011011000;
assign LUT_1[269] = 32'b11111111111111111110001101010100;
assign LUT_1[270] = 32'b00000000000000000000101001101001;
assign LUT_1[271] = 32'b11111111111111111001111011100101;
assign LUT_1[272] = 32'b11111111111111111111101111101110;
assign LUT_1[273] = 32'b11111111111111111001000001101010;
assign LUT_1[274] = 32'b11111111111111111011011101111111;
assign LUT_1[275] = 32'b11111111111111110100101111111011;
assign LUT_1[276] = 32'b00000000000000000111101001000101;
assign LUT_1[277] = 32'b00000000000000000000111011000001;
assign LUT_1[278] = 32'b00000000000000000011010111010110;
assign LUT_1[279] = 32'b11111111111111111100101001010010;
assign LUT_1[280] = 32'b11111111111111111110111101100011;
assign LUT_1[281] = 32'b11111111111111111000001111011111;
assign LUT_1[282] = 32'b11111111111111111010101011110100;
assign LUT_1[283] = 32'b11111111111111110011111101110000;
assign LUT_1[284] = 32'b00000000000000000110110110111010;
assign LUT_1[285] = 32'b00000000000000000000001000110110;
assign LUT_1[286] = 32'b00000000000000000010100101001011;
assign LUT_1[287] = 32'b11111111111111111011110111000111;
assign LUT_1[288] = 32'b11111111111111111110101111001011;
assign LUT_1[289] = 32'b11111111111111111000000001000111;
assign LUT_1[290] = 32'b11111111111111111010011101011100;
assign LUT_1[291] = 32'b11111111111111110011101111011000;
assign LUT_1[292] = 32'b00000000000000000110101000100010;
assign LUT_1[293] = 32'b11111111111111111111111010011110;
assign LUT_1[294] = 32'b00000000000000000010010110110011;
assign LUT_1[295] = 32'b11111111111111111011101000101111;
assign LUT_1[296] = 32'b11111111111111111101111101000000;
assign LUT_1[297] = 32'b11111111111111110111001110111100;
assign LUT_1[298] = 32'b11111111111111111001101011010001;
assign LUT_1[299] = 32'b11111111111111110010111101001101;
assign LUT_1[300] = 32'b00000000000000000101110110010111;
assign LUT_1[301] = 32'b11111111111111111111001000010011;
assign LUT_1[302] = 32'b00000000000000000001100100101000;
assign LUT_1[303] = 32'b11111111111111111010110110100100;
assign LUT_1[304] = 32'b00000000000000000000101010101101;
assign LUT_1[305] = 32'b11111111111111111001111100101001;
assign LUT_1[306] = 32'b11111111111111111100011000111110;
assign LUT_1[307] = 32'b11111111111111110101101010111010;
assign LUT_1[308] = 32'b00000000000000001000100100000100;
assign LUT_1[309] = 32'b00000000000000000001110110000000;
assign LUT_1[310] = 32'b00000000000000000100010010010101;
assign LUT_1[311] = 32'b11111111111111111101100100010001;
assign LUT_1[312] = 32'b11111111111111111111111000100010;
assign LUT_1[313] = 32'b11111111111111111001001010011110;
assign LUT_1[314] = 32'b11111111111111111011100110110011;
assign LUT_1[315] = 32'b11111111111111110100111000101111;
assign LUT_1[316] = 32'b00000000000000000111110001111001;
assign LUT_1[317] = 32'b00000000000000000001000011110101;
assign LUT_1[318] = 32'b00000000000000000011100000001010;
assign LUT_1[319] = 32'b11111111111111111100110010000110;
assign LUT_1[320] = 32'b11111111111111111111110001110100;
assign LUT_1[321] = 32'b11111111111111111001000011110000;
assign LUT_1[322] = 32'b11111111111111111011100000000101;
assign LUT_1[323] = 32'b11111111111111110100110010000001;
assign LUT_1[324] = 32'b00000000000000000111101011001011;
assign LUT_1[325] = 32'b00000000000000000000111101000111;
assign LUT_1[326] = 32'b00000000000000000011011001011100;
assign LUT_1[327] = 32'b11111111111111111100101011011000;
assign LUT_1[328] = 32'b11111111111111111110111111101001;
assign LUT_1[329] = 32'b11111111111111111000010001100101;
assign LUT_1[330] = 32'b11111111111111111010101101111010;
assign LUT_1[331] = 32'b11111111111111110011111111110110;
assign LUT_1[332] = 32'b00000000000000000110111001000000;
assign LUT_1[333] = 32'b00000000000000000000001010111100;
assign LUT_1[334] = 32'b00000000000000000010100111010001;
assign LUT_1[335] = 32'b11111111111111111011111001001101;
assign LUT_1[336] = 32'b00000000000000000001101101010110;
assign LUT_1[337] = 32'b11111111111111111010111111010010;
assign LUT_1[338] = 32'b11111111111111111101011011100111;
assign LUT_1[339] = 32'b11111111111111110110101101100011;
assign LUT_1[340] = 32'b00000000000000001001100110101101;
assign LUT_1[341] = 32'b00000000000000000010111000101001;
assign LUT_1[342] = 32'b00000000000000000101010100111110;
assign LUT_1[343] = 32'b11111111111111111110100110111010;
assign LUT_1[344] = 32'b00000000000000000000111011001011;
assign LUT_1[345] = 32'b11111111111111111010001101000111;
assign LUT_1[346] = 32'b11111111111111111100101001011100;
assign LUT_1[347] = 32'b11111111111111110101111011011000;
assign LUT_1[348] = 32'b00000000000000001000110100100010;
assign LUT_1[349] = 32'b00000000000000000010000110011110;
assign LUT_1[350] = 32'b00000000000000000100100010110011;
assign LUT_1[351] = 32'b11111111111111111101110100101111;
assign LUT_1[352] = 32'b00000000000000000000101100110011;
assign LUT_1[353] = 32'b11111111111111111001111110101111;
assign LUT_1[354] = 32'b11111111111111111100011011000100;
assign LUT_1[355] = 32'b11111111111111110101101101000000;
assign LUT_1[356] = 32'b00000000000000001000100110001010;
assign LUT_1[357] = 32'b00000000000000000001111000000110;
assign LUT_1[358] = 32'b00000000000000000100010100011011;
assign LUT_1[359] = 32'b11111111111111111101100110010111;
assign LUT_1[360] = 32'b11111111111111111111111010101000;
assign LUT_1[361] = 32'b11111111111111111001001100100100;
assign LUT_1[362] = 32'b11111111111111111011101000111001;
assign LUT_1[363] = 32'b11111111111111110100111010110101;
assign LUT_1[364] = 32'b00000000000000000111110011111111;
assign LUT_1[365] = 32'b00000000000000000001000101111011;
assign LUT_1[366] = 32'b00000000000000000011100010010000;
assign LUT_1[367] = 32'b11111111111111111100110100001100;
assign LUT_1[368] = 32'b00000000000000000010101000010101;
assign LUT_1[369] = 32'b11111111111111111011111010010001;
assign LUT_1[370] = 32'b11111111111111111110010110100110;
assign LUT_1[371] = 32'b11111111111111110111101000100010;
assign LUT_1[372] = 32'b00000000000000001010100001101100;
assign LUT_1[373] = 32'b00000000000000000011110011101000;
assign LUT_1[374] = 32'b00000000000000000110001111111101;
assign LUT_1[375] = 32'b11111111111111111111100001111001;
assign LUT_1[376] = 32'b00000000000000000001110110001010;
assign LUT_1[377] = 32'b11111111111111111011001000000110;
assign LUT_1[378] = 32'b11111111111111111101100100011011;
assign LUT_1[379] = 32'b11111111111111110110110110010111;
assign LUT_1[380] = 32'b00000000000000001001101111100001;
assign LUT_1[381] = 32'b00000000000000000011000001011101;
assign LUT_1[382] = 32'b00000000000000000101011101110010;
assign LUT_1[383] = 32'b11111111111111111110101111101110;
assign LUT_1[384] = 32'b00000000000000000000110100001111;
assign LUT_1[385] = 32'b11111111111111111010000110001011;
assign LUT_1[386] = 32'b11111111111111111100100010100000;
assign LUT_1[387] = 32'b11111111111111110101110100011100;
assign LUT_1[388] = 32'b00000000000000001000101101100110;
assign LUT_1[389] = 32'b00000000000000000001111111100010;
assign LUT_1[390] = 32'b00000000000000000100011011110111;
assign LUT_1[391] = 32'b11111111111111111101101101110011;
assign LUT_1[392] = 32'b00000000000000000000000010000100;
assign LUT_1[393] = 32'b11111111111111111001010100000000;
assign LUT_1[394] = 32'b11111111111111111011110000010101;
assign LUT_1[395] = 32'b11111111111111110101000010010001;
assign LUT_1[396] = 32'b00000000000000000111111011011011;
assign LUT_1[397] = 32'b00000000000000000001001101010111;
assign LUT_1[398] = 32'b00000000000000000011101001101100;
assign LUT_1[399] = 32'b11111111111111111100111011101000;
assign LUT_1[400] = 32'b00000000000000000010101111110001;
assign LUT_1[401] = 32'b11111111111111111100000001101101;
assign LUT_1[402] = 32'b11111111111111111110011110000010;
assign LUT_1[403] = 32'b11111111111111110111101111111110;
assign LUT_1[404] = 32'b00000000000000001010101001001000;
assign LUT_1[405] = 32'b00000000000000000011111011000100;
assign LUT_1[406] = 32'b00000000000000000110010111011001;
assign LUT_1[407] = 32'b11111111111111111111101001010101;
assign LUT_1[408] = 32'b00000000000000000001111101100110;
assign LUT_1[409] = 32'b11111111111111111011001111100010;
assign LUT_1[410] = 32'b11111111111111111101101011110111;
assign LUT_1[411] = 32'b11111111111111110110111101110011;
assign LUT_1[412] = 32'b00000000000000001001110110111101;
assign LUT_1[413] = 32'b00000000000000000011001000111001;
assign LUT_1[414] = 32'b00000000000000000101100101001110;
assign LUT_1[415] = 32'b11111111111111111110110111001010;
assign LUT_1[416] = 32'b00000000000000000001101111001110;
assign LUT_1[417] = 32'b11111111111111111011000001001010;
assign LUT_1[418] = 32'b11111111111111111101011101011111;
assign LUT_1[419] = 32'b11111111111111110110101111011011;
assign LUT_1[420] = 32'b00000000000000001001101000100101;
assign LUT_1[421] = 32'b00000000000000000010111010100001;
assign LUT_1[422] = 32'b00000000000000000101010110110110;
assign LUT_1[423] = 32'b11111111111111111110101000110010;
assign LUT_1[424] = 32'b00000000000000000000111101000011;
assign LUT_1[425] = 32'b11111111111111111010001110111111;
assign LUT_1[426] = 32'b11111111111111111100101011010100;
assign LUT_1[427] = 32'b11111111111111110101111101010000;
assign LUT_1[428] = 32'b00000000000000001000110110011010;
assign LUT_1[429] = 32'b00000000000000000010001000010110;
assign LUT_1[430] = 32'b00000000000000000100100100101011;
assign LUT_1[431] = 32'b11111111111111111101110110100111;
assign LUT_1[432] = 32'b00000000000000000011101010110000;
assign LUT_1[433] = 32'b11111111111111111100111100101100;
assign LUT_1[434] = 32'b11111111111111111111011001000001;
assign LUT_1[435] = 32'b11111111111111111000101010111101;
assign LUT_1[436] = 32'b00000000000000001011100100000111;
assign LUT_1[437] = 32'b00000000000000000100110110000011;
assign LUT_1[438] = 32'b00000000000000000111010010011000;
assign LUT_1[439] = 32'b00000000000000000000100100010100;
assign LUT_1[440] = 32'b00000000000000000010111000100101;
assign LUT_1[441] = 32'b11111111111111111100001010100001;
assign LUT_1[442] = 32'b11111111111111111110100110110110;
assign LUT_1[443] = 32'b11111111111111110111111000110010;
assign LUT_1[444] = 32'b00000000000000001010110001111100;
assign LUT_1[445] = 32'b00000000000000000100000011111000;
assign LUT_1[446] = 32'b00000000000000000110100000001101;
assign LUT_1[447] = 32'b11111111111111111111110010001001;
assign LUT_1[448] = 32'b00000000000000000010110001110111;
assign LUT_1[449] = 32'b11111111111111111100000011110011;
assign LUT_1[450] = 32'b11111111111111111110100000001000;
assign LUT_1[451] = 32'b11111111111111110111110010000100;
assign LUT_1[452] = 32'b00000000000000001010101011001110;
assign LUT_1[453] = 32'b00000000000000000011111101001010;
assign LUT_1[454] = 32'b00000000000000000110011001011111;
assign LUT_1[455] = 32'b11111111111111111111101011011011;
assign LUT_1[456] = 32'b00000000000000000001111111101100;
assign LUT_1[457] = 32'b11111111111111111011010001101000;
assign LUT_1[458] = 32'b11111111111111111101101101111101;
assign LUT_1[459] = 32'b11111111111111110110111111111001;
assign LUT_1[460] = 32'b00000000000000001001111001000011;
assign LUT_1[461] = 32'b00000000000000000011001010111111;
assign LUT_1[462] = 32'b00000000000000000101100111010100;
assign LUT_1[463] = 32'b11111111111111111110111001010000;
assign LUT_1[464] = 32'b00000000000000000100101101011001;
assign LUT_1[465] = 32'b11111111111111111101111111010101;
assign LUT_1[466] = 32'b00000000000000000000011011101010;
assign LUT_1[467] = 32'b11111111111111111001101101100110;
assign LUT_1[468] = 32'b00000000000000001100100110110000;
assign LUT_1[469] = 32'b00000000000000000101111000101100;
assign LUT_1[470] = 32'b00000000000000001000010101000001;
assign LUT_1[471] = 32'b00000000000000000001100110111101;
assign LUT_1[472] = 32'b00000000000000000011111011001110;
assign LUT_1[473] = 32'b11111111111111111101001101001010;
assign LUT_1[474] = 32'b11111111111111111111101001011111;
assign LUT_1[475] = 32'b11111111111111111000111011011011;
assign LUT_1[476] = 32'b00000000000000001011110100100101;
assign LUT_1[477] = 32'b00000000000000000101000110100001;
assign LUT_1[478] = 32'b00000000000000000111100010110110;
assign LUT_1[479] = 32'b00000000000000000000110100110010;
assign LUT_1[480] = 32'b00000000000000000011101100110110;
assign LUT_1[481] = 32'b11111111111111111100111110110010;
assign LUT_1[482] = 32'b11111111111111111111011011000111;
assign LUT_1[483] = 32'b11111111111111111000101101000011;
assign LUT_1[484] = 32'b00000000000000001011100110001101;
assign LUT_1[485] = 32'b00000000000000000100111000001001;
assign LUT_1[486] = 32'b00000000000000000111010100011110;
assign LUT_1[487] = 32'b00000000000000000000100110011010;
assign LUT_1[488] = 32'b00000000000000000010111010101011;
assign LUT_1[489] = 32'b11111111111111111100001100100111;
assign LUT_1[490] = 32'b11111111111111111110101000111100;
assign LUT_1[491] = 32'b11111111111111110111111010111000;
assign LUT_1[492] = 32'b00000000000000001010110100000010;
assign LUT_1[493] = 32'b00000000000000000100000101111110;
assign LUT_1[494] = 32'b00000000000000000110100010010011;
assign LUT_1[495] = 32'b11111111111111111111110100001111;
assign LUT_1[496] = 32'b00000000000000000101101000011000;
assign LUT_1[497] = 32'b11111111111111111110111010010100;
assign LUT_1[498] = 32'b00000000000000000001010110101001;
assign LUT_1[499] = 32'b11111111111111111010101000100101;
assign LUT_1[500] = 32'b00000000000000001101100001101111;
assign LUT_1[501] = 32'b00000000000000000110110011101011;
assign LUT_1[502] = 32'b00000000000000001001010000000000;
assign LUT_1[503] = 32'b00000000000000000010100001111100;
assign LUT_1[504] = 32'b00000000000000000100110110001101;
assign LUT_1[505] = 32'b11111111111111111110001000001001;
assign LUT_1[506] = 32'b00000000000000000000100100011110;
assign LUT_1[507] = 32'b11111111111111111001110110011010;
assign LUT_1[508] = 32'b00000000000000001100101111100100;
assign LUT_1[509] = 32'b00000000000000000110000001100000;
assign LUT_1[510] = 32'b00000000000000001000011101110101;
assign LUT_1[511] = 32'b00000000000000000001101111110001;
assign LUT_1[512] = 32'b11111111111111111001101110011101;
assign LUT_1[513] = 32'b11111111111111110011000000011001;
assign LUT_1[514] = 32'b11111111111111110101011100101110;
assign LUT_1[515] = 32'b11111111111111101110101110101010;
assign LUT_1[516] = 32'b00000000000000000001100111110100;
assign LUT_1[517] = 32'b11111111111111111010111001110000;
assign LUT_1[518] = 32'b11111111111111111101010110000101;
assign LUT_1[519] = 32'b11111111111111110110101000000001;
assign LUT_1[520] = 32'b11111111111111111000111100010010;
assign LUT_1[521] = 32'b11111111111111110010001110001110;
assign LUT_1[522] = 32'b11111111111111110100101010100011;
assign LUT_1[523] = 32'b11111111111111101101111100011111;
assign LUT_1[524] = 32'b00000000000000000000110101101001;
assign LUT_1[525] = 32'b11111111111111111010000111100101;
assign LUT_1[526] = 32'b11111111111111111100100011111010;
assign LUT_1[527] = 32'b11111111111111110101110101110110;
assign LUT_1[528] = 32'b11111111111111111011101001111111;
assign LUT_1[529] = 32'b11111111111111110100111011111011;
assign LUT_1[530] = 32'b11111111111111110111011000010000;
assign LUT_1[531] = 32'b11111111111111110000101010001100;
assign LUT_1[532] = 32'b00000000000000000011100011010110;
assign LUT_1[533] = 32'b11111111111111111100110101010010;
assign LUT_1[534] = 32'b11111111111111111111010001100111;
assign LUT_1[535] = 32'b11111111111111111000100011100011;
assign LUT_1[536] = 32'b11111111111111111010110111110100;
assign LUT_1[537] = 32'b11111111111111110100001001110000;
assign LUT_1[538] = 32'b11111111111111110110100110000101;
assign LUT_1[539] = 32'b11111111111111101111111000000001;
assign LUT_1[540] = 32'b00000000000000000010110001001011;
assign LUT_1[541] = 32'b11111111111111111100000011000111;
assign LUT_1[542] = 32'b11111111111111111110011111011100;
assign LUT_1[543] = 32'b11111111111111110111110001011000;
assign LUT_1[544] = 32'b11111111111111111010101001011100;
assign LUT_1[545] = 32'b11111111111111110011111011011000;
assign LUT_1[546] = 32'b11111111111111110110010111101101;
assign LUT_1[547] = 32'b11111111111111101111101001101001;
assign LUT_1[548] = 32'b00000000000000000010100010110011;
assign LUT_1[549] = 32'b11111111111111111011110100101111;
assign LUT_1[550] = 32'b11111111111111111110010001000100;
assign LUT_1[551] = 32'b11111111111111110111100011000000;
assign LUT_1[552] = 32'b11111111111111111001110111010001;
assign LUT_1[553] = 32'b11111111111111110011001001001101;
assign LUT_1[554] = 32'b11111111111111110101100101100010;
assign LUT_1[555] = 32'b11111111111111101110110111011110;
assign LUT_1[556] = 32'b00000000000000000001110000101000;
assign LUT_1[557] = 32'b11111111111111111011000010100100;
assign LUT_1[558] = 32'b11111111111111111101011110111001;
assign LUT_1[559] = 32'b11111111111111110110110000110101;
assign LUT_1[560] = 32'b11111111111111111100100100111110;
assign LUT_1[561] = 32'b11111111111111110101110110111010;
assign LUT_1[562] = 32'b11111111111111111000010011001111;
assign LUT_1[563] = 32'b11111111111111110001100101001011;
assign LUT_1[564] = 32'b00000000000000000100011110010101;
assign LUT_1[565] = 32'b11111111111111111101110000010001;
assign LUT_1[566] = 32'b00000000000000000000001100100110;
assign LUT_1[567] = 32'b11111111111111111001011110100010;
assign LUT_1[568] = 32'b11111111111111111011110010110011;
assign LUT_1[569] = 32'b11111111111111110101000100101111;
assign LUT_1[570] = 32'b11111111111111110111100001000100;
assign LUT_1[571] = 32'b11111111111111110000110011000000;
assign LUT_1[572] = 32'b00000000000000000011101100001010;
assign LUT_1[573] = 32'b11111111111111111100111110000110;
assign LUT_1[574] = 32'b11111111111111111111011010011011;
assign LUT_1[575] = 32'b11111111111111111000101100010111;
assign LUT_1[576] = 32'b11111111111111111011101100000101;
assign LUT_1[577] = 32'b11111111111111110100111110000001;
assign LUT_1[578] = 32'b11111111111111110111011010010110;
assign LUT_1[579] = 32'b11111111111111110000101100010010;
assign LUT_1[580] = 32'b00000000000000000011100101011100;
assign LUT_1[581] = 32'b11111111111111111100110111011000;
assign LUT_1[582] = 32'b11111111111111111111010011101101;
assign LUT_1[583] = 32'b11111111111111111000100101101001;
assign LUT_1[584] = 32'b11111111111111111010111001111010;
assign LUT_1[585] = 32'b11111111111111110100001011110110;
assign LUT_1[586] = 32'b11111111111111110110101000001011;
assign LUT_1[587] = 32'b11111111111111101111111010000111;
assign LUT_1[588] = 32'b00000000000000000010110011010001;
assign LUT_1[589] = 32'b11111111111111111100000101001101;
assign LUT_1[590] = 32'b11111111111111111110100001100010;
assign LUT_1[591] = 32'b11111111111111110111110011011110;
assign LUT_1[592] = 32'b11111111111111111101100111100111;
assign LUT_1[593] = 32'b11111111111111110110111001100011;
assign LUT_1[594] = 32'b11111111111111111001010101111000;
assign LUT_1[595] = 32'b11111111111111110010100111110100;
assign LUT_1[596] = 32'b00000000000000000101100000111110;
assign LUT_1[597] = 32'b11111111111111111110110010111010;
assign LUT_1[598] = 32'b00000000000000000001001111001111;
assign LUT_1[599] = 32'b11111111111111111010100001001011;
assign LUT_1[600] = 32'b11111111111111111100110101011100;
assign LUT_1[601] = 32'b11111111111111110110000111011000;
assign LUT_1[602] = 32'b11111111111111111000100011101101;
assign LUT_1[603] = 32'b11111111111111110001110101101001;
assign LUT_1[604] = 32'b00000000000000000100101110110011;
assign LUT_1[605] = 32'b11111111111111111110000000101111;
assign LUT_1[606] = 32'b00000000000000000000011101000100;
assign LUT_1[607] = 32'b11111111111111111001101111000000;
assign LUT_1[608] = 32'b11111111111111111100100111000100;
assign LUT_1[609] = 32'b11111111111111110101111001000000;
assign LUT_1[610] = 32'b11111111111111111000010101010101;
assign LUT_1[611] = 32'b11111111111111110001100111010001;
assign LUT_1[612] = 32'b00000000000000000100100000011011;
assign LUT_1[613] = 32'b11111111111111111101110010010111;
assign LUT_1[614] = 32'b00000000000000000000001110101100;
assign LUT_1[615] = 32'b11111111111111111001100000101000;
assign LUT_1[616] = 32'b11111111111111111011110100111001;
assign LUT_1[617] = 32'b11111111111111110101000110110101;
assign LUT_1[618] = 32'b11111111111111110111100011001010;
assign LUT_1[619] = 32'b11111111111111110000110101000110;
assign LUT_1[620] = 32'b00000000000000000011101110010000;
assign LUT_1[621] = 32'b11111111111111111101000000001100;
assign LUT_1[622] = 32'b11111111111111111111011100100001;
assign LUT_1[623] = 32'b11111111111111111000101110011101;
assign LUT_1[624] = 32'b11111111111111111110100010100110;
assign LUT_1[625] = 32'b11111111111111110111110100100010;
assign LUT_1[626] = 32'b11111111111111111010010000110111;
assign LUT_1[627] = 32'b11111111111111110011100010110011;
assign LUT_1[628] = 32'b00000000000000000110011011111101;
assign LUT_1[629] = 32'b11111111111111111111101101111001;
assign LUT_1[630] = 32'b00000000000000000010001010001110;
assign LUT_1[631] = 32'b11111111111111111011011100001010;
assign LUT_1[632] = 32'b11111111111111111101110000011011;
assign LUT_1[633] = 32'b11111111111111110111000010010111;
assign LUT_1[634] = 32'b11111111111111111001011110101100;
assign LUT_1[635] = 32'b11111111111111110010110000101000;
assign LUT_1[636] = 32'b00000000000000000101101001110010;
assign LUT_1[637] = 32'b11111111111111111110111011101110;
assign LUT_1[638] = 32'b00000000000000000001011000000011;
assign LUT_1[639] = 32'b11111111111111111010101001111111;
assign LUT_1[640] = 32'b11111111111111111100101110100000;
assign LUT_1[641] = 32'b11111111111111110110000000011100;
assign LUT_1[642] = 32'b11111111111111111000011100110001;
assign LUT_1[643] = 32'b11111111111111110001101110101101;
assign LUT_1[644] = 32'b00000000000000000100100111110111;
assign LUT_1[645] = 32'b11111111111111111101111001110011;
assign LUT_1[646] = 32'b00000000000000000000010110001000;
assign LUT_1[647] = 32'b11111111111111111001101000000100;
assign LUT_1[648] = 32'b11111111111111111011111100010101;
assign LUT_1[649] = 32'b11111111111111110101001110010001;
assign LUT_1[650] = 32'b11111111111111110111101010100110;
assign LUT_1[651] = 32'b11111111111111110000111100100010;
assign LUT_1[652] = 32'b00000000000000000011110101101100;
assign LUT_1[653] = 32'b11111111111111111101000111101000;
assign LUT_1[654] = 32'b11111111111111111111100011111101;
assign LUT_1[655] = 32'b11111111111111111000110101111001;
assign LUT_1[656] = 32'b11111111111111111110101010000010;
assign LUT_1[657] = 32'b11111111111111110111111011111110;
assign LUT_1[658] = 32'b11111111111111111010011000010011;
assign LUT_1[659] = 32'b11111111111111110011101010001111;
assign LUT_1[660] = 32'b00000000000000000110100011011001;
assign LUT_1[661] = 32'b11111111111111111111110101010101;
assign LUT_1[662] = 32'b00000000000000000010010001101010;
assign LUT_1[663] = 32'b11111111111111111011100011100110;
assign LUT_1[664] = 32'b11111111111111111101110111110111;
assign LUT_1[665] = 32'b11111111111111110111001001110011;
assign LUT_1[666] = 32'b11111111111111111001100110001000;
assign LUT_1[667] = 32'b11111111111111110010111000000100;
assign LUT_1[668] = 32'b00000000000000000101110001001110;
assign LUT_1[669] = 32'b11111111111111111111000011001010;
assign LUT_1[670] = 32'b00000000000000000001011111011111;
assign LUT_1[671] = 32'b11111111111111111010110001011011;
assign LUT_1[672] = 32'b11111111111111111101101001011111;
assign LUT_1[673] = 32'b11111111111111110110111011011011;
assign LUT_1[674] = 32'b11111111111111111001010111110000;
assign LUT_1[675] = 32'b11111111111111110010101001101100;
assign LUT_1[676] = 32'b00000000000000000101100010110110;
assign LUT_1[677] = 32'b11111111111111111110110100110010;
assign LUT_1[678] = 32'b00000000000000000001010001000111;
assign LUT_1[679] = 32'b11111111111111111010100011000011;
assign LUT_1[680] = 32'b11111111111111111100110111010100;
assign LUT_1[681] = 32'b11111111111111110110001001010000;
assign LUT_1[682] = 32'b11111111111111111000100101100101;
assign LUT_1[683] = 32'b11111111111111110001110111100001;
assign LUT_1[684] = 32'b00000000000000000100110000101011;
assign LUT_1[685] = 32'b11111111111111111110000010100111;
assign LUT_1[686] = 32'b00000000000000000000011110111100;
assign LUT_1[687] = 32'b11111111111111111001110000111000;
assign LUT_1[688] = 32'b11111111111111111111100101000001;
assign LUT_1[689] = 32'b11111111111111111000110110111101;
assign LUT_1[690] = 32'b11111111111111111011010011010010;
assign LUT_1[691] = 32'b11111111111111110100100101001110;
assign LUT_1[692] = 32'b00000000000000000111011110011000;
assign LUT_1[693] = 32'b00000000000000000000110000010100;
assign LUT_1[694] = 32'b00000000000000000011001100101001;
assign LUT_1[695] = 32'b11111111111111111100011110100101;
assign LUT_1[696] = 32'b11111111111111111110110010110110;
assign LUT_1[697] = 32'b11111111111111111000000100110010;
assign LUT_1[698] = 32'b11111111111111111010100001000111;
assign LUT_1[699] = 32'b11111111111111110011110011000011;
assign LUT_1[700] = 32'b00000000000000000110101100001101;
assign LUT_1[701] = 32'b11111111111111111111111110001001;
assign LUT_1[702] = 32'b00000000000000000010011010011110;
assign LUT_1[703] = 32'b11111111111111111011101100011010;
assign LUT_1[704] = 32'b11111111111111111110101100001000;
assign LUT_1[705] = 32'b11111111111111110111111110000100;
assign LUT_1[706] = 32'b11111111111111111010011010011001;
assign LUT_1[707] = 32'b11111111111111110011101100010101;
assign LUT_1[708] = 32'b00000000000000000110100101011111;
assign LUT_1[709] = 32'b11111111111111111111110111011011;
assign LUT_1[710] = 32'b00000000000000000010010011110000;
assign LUT_1[711] = 32'b11111111111111111011100101101100;
assign LUT_1[712] = 32'b11111111111111111101111001111101;
assign LUT_1[713] = 32'b11111111111111110111001011111001;
assign LUT_1[714] = 32'b11111111111111111001101000001110;
assign LUT_1[715] = 32'b11111111111111110010111010001010;
assign LUT_1[716] = 32'b00000000000000000101110011010100;
assign LUT_1[717] = 32'b11111111111111111111000101010000;
assign LUT_1[718] = 32'b00000000000000000001100001100101;
assign LUT_1[719] = 32'b11111111111111111010110011100001;
assign LUT_1[720] = 32'b00000000000000000000100111101010;
assign LUT_1[721] = 32'b11111111111111111001111001100110;
assign LUT_1[722] = 32'b11111111111111111100010101111011;
assign LUT_1[723] = 32'b11111111111111110101100111110111;
assign LUT_1[724] = 32'b00000000000000001000100001000001;
assign LUT_1[725] = 32'b00000000000000000001110010111101;
assign LUT_1[726] = 32'b00000000000000000100001111010010;
assign LUT_1[727] = 32'b11111111111111111101100001001110;
assign LUT_1[728] = 32'b11111111111111111111110101011111;
assign LUT_1[729] = 32'b11111111111111111001000111011011;
assign LUT_1[730] = 32'b11111111111111111011100011110000;
assign LUT_1[731] = 32'b11111111111111110100110101101100;
assign LUT_1[732] = 32'b00000000000000000111101110110110;
assign LUT_1[733] = 32'b00000000000000000001000000110010;
assign LUT_1[734] = 32'b00000000000000000011011101000111;
assign LUT_1[735] = 32'b11111111111111111100101111000011;
assign LUT_1[736] = 32'b11111111111111111111100111000111;
assign LUT_1[737] = 32'b11111111111111111000111001000011;
assign LUT_1[738] = 32'b11111111111111111011010101011000;
assign LUT_1[739] = 32'b11111111111111110100100111010100;
assign LUT_1[740] = 32'b00000000000000000111100000011110;
assign LUT_1[741] = 32'b00000000000000000000110010011010;
assign LUT_1[742] = 32'b00000000000000000011001110101111;
assign LUT_1[743] = 32'b11111111111111111100100000101011;
assign LUT_1[744] = 32'b11111111111111111110110100111100;
assign LUT_1[745] = 32'b11111111111111111000000110111000;
assign LUT_1[746] = 32'b11111111111111111010100011001101;
assign LUT_1[747] = 32'b11111111111111110011110101001001;
assign LUT_1[748] = 32'b00000000000000000110101110010011;
assign LUT_1[749] = 32'b00000000000000000000000000001111;
assign LUT_1[750] = 32'b00000000000000000010011100100100;
assign LUT_1[751] = 32'b11111111111111111011101110100000;
assign LUT_1[752] = 32'b00000000000000000001100010101001;
assign LUT_1[753] = 32'b11111111111111111010110100100101;
assign LUT_1[754] = 32'b11111111111111111101010000111010;
assign LUT_1[755] = 32'b11111111111111110110100010110110;
assign LUT_1[756] = 32'b00000000000000001001011100000000;
assign LUT_1[757] = 32'b00000000000000000010101101111100;
assign LUT_1[758] = 32'b00000000000000000101001010010001;
assign LUT_1[759] = 32'b11111111111111111110011100001101;
assign LUT_1[760] = 32'b00000000000000000000110000011110;
assign LUT_1[761] = 32'b11111111111111111010000010011010;
assign LUT_1[762] = 32'b11111111111111111100011110101111;
assign LUT_1[763] = 32'b11111111111111110101110000101011;
assign LUT_1[764] = 32'b00000000000000001000101001110101;
assign LUT_1[765] = 32'b00000000000000000001111011110001;
assign LUT_1[766] = 32'b00000000000000000100011000000110;
assign LUT_1[767] = 32'b11111111111111111101101010000010;
assign LUT_1[768] = 32'b11111111111111110111100010101001;
assign LUT_1[769] = 32'b11111111111111110000110100100101;
assign LUT_1[770] = 32'b11111111111111110011010000111010;
assign LUT_1[771] = 32'b11111111111111101100100010110110;
assign LUT_1[772] = 32'b11111111111111111111011100000000;
assign LUT_1[773] = 32'b11111111111111111000101101111100;
assign LUT_1[774] = 32'b11111111111111111011001010010001;
assign LUT_1[775] = 32'b11111111111111110100011100001101;
assign LUT_1[776] = 32'b11111111111111110110110000011110;
assign LUT_1[777] = 32'b11111111111111110000000010011010;
assign LUT_1[778] = 32'b11111111111111110010011110101111;
assign LUT_1[779] = 32'b11111111111111101011110000101011;
assign LUT_1[780] = 32'b11111111111111111110101001110101;
assign LUT_1[781] = 32'b11111111111111110111111011110001;
assign LUT_1[782] = 32'b11111111111111111010011000000110;
assign LUT_1[783] = 32'b11111111111111110011101010000010;
assign LUT_1[784] = 32'b11111111111111111001011110001011;
assign LUT_1[785] = 32'b11111111111111110010110000000111;
assign LUT_1[786] = 32'b11111111111111110101001100011100;
assign LUT_1[787] = 32'b11111111111111101110011110011000;
assign LUT_1[788] = 32'b00000000000000000001010111100010;
assign LUT_1[789] = 32'b11111111111111111010101001011110;
assign LUT_1[790] = 32'b11111111111111111101000101110011;
assign LUT_1[791] = 32'b11111111111111110110010111101111;
assign LUT_1[792] = 32'b11111111111111111000101100000000;
assign LUT_1[793] = 32'b11111111111111110001111101111100;
assign LUT_1[794] = 32'b11111111111111110100011010010001;
assign LUT_1[795] = 32'b11111111111111101101101100001101;
assign LUT_1[796] = 32'b00000000000000000000100101010111;
assign LUT_1[797] = 32'b11111111111111111001110111010011;
assign LUT_1[798] = 32'b11111111111111111100010011101000;
assign LUT_1[799] = 32'b11111111111111110101100101100100;
assign LUT_1[800] = 32'b11111111111111111000011101101000;
assign LUT_1[801] = 32'b11111111111111110001101111100100;
assign LUT_1[802] = 32'b11111111111111110100001011111001;
assign LUT_1[803] = 32'b11111111111111101101011101110101;
assign LUT_1[804] = 32'b00000000000000000000010110111111;
assign LUT_1[805] = 32'b11111111111111111001101000111011;
assign LUT_1[806] = 32'b11111111111111111100000101010000;
assign LUT_1[807] = 32'b11111111111111110101010111001100;
assign LUT_1[808] = 32'b11111111111111110111101011011101;
assign LUT_1[809] = 32'b11111111111111110000111101011001;
assign LUT_1[810] = 32'b11111111111111110011011001101110;
assign LUT_1[811] = 32'b11111111111111101100101011101010;
assign LUT_1[812] = 32'b11111111111111111111100100110100;
assign LUT_1[813] = 32'b11111111111111111000110110110000;
assign LUT_1[814] = 32'b11111111111111111011010011000101;
assign LUT_1[815] = 32'b11111111111111110100100101000001;
assign LUT_1[816] = 32'b11111111111111111010011001001010;
assign LUT_1[817] = 32'b11111111111111110011101011000110;
assign LUT_1[818] = 32'b11111111111111110110000111011011;
assign LUT_1[819] = 32'b11111111111111101111011001010111;
assign LUT_1[820] = 32'b00000000000000000010010010100001;
assign LUT_1[821] = 32'b11111111111111111011100100011101;
assign LUT_1[822] = 32'b11111111111111111110000000110010;
assign LUT_1[823] = 32'b11111111111111110111010010101110;
assign LUT_1[824] = 32'b11111111111111111001100110111111;
assign LUT_1[825] = 32'b11111111111111110010111000111011;
assign LUT_1[826] = 32'b11111111111111110101010101010000;
assign LUT_1[827] = 32'b11111111111111101110100111001100;
assign LUT_1[828] = 32'b00000000000000000001100000010110;
assign LUT_1[829] = 32'b11111111111111111010110010010010;
assign LUT_1[830] = 32'b11111111111111111101001110100111;
assign LUT_1[831] = 32'b11111111111111110110100000100011;
assign LUT_1[832] = 32'b11111111111111111001100000010001;
assign LUT_1[833] = 32'b11111111111111110010110010001101;
assign LUT_1[834] = 32'b11111111111111110101001110100010;
assign LUT_1[835] = 32'b11111111111111101110100000011110;
assign LUT_1[836] = 32'b00000000000000000001011001101000;
assign LUT_1[837] = 32'b11111111111111111010101011100100;
assign LUT_1[838] = 32'b11111111111111111101000111111001;
assign LUT_1[839] = 32'b11111111111111110110011001110101;
assign LUT_1[840] = 32'b11111111111111111000101110000110;
assign LUT_1[841] = 32'b11111111111111110010000000000010;
assign LUT_1[842] = 32'b11111111111111110100011100010111;
assign LUT_1[843] = 32'b11111111111111101101101110010011;
assign LUT_1[844] = 32'b00000000000000000000100111011101;
assign LUT_1[845] = 32'b11111111111111111001111001011001;
assign LUT_1[846] = 32'b11111111111111111100010101101110;
assign LUT_1[847] = 32'b11111111111111110101100111101010;
assign LUT_1[848] = 32'b11111111111111111011011011110011;
assign LUT_1[849] = 32'b11111111111111110100101101101111;
assign LUT_1[850] = 32'b11111111111111110111001010000100;
assign LUT_1[851] = 32'b11111111111111110000011100000000;
assign LUT_1[852] = 32'b00000000000000000011010101001010;
assign LUT_1[853] = 32'b11111111111111111100100111000110;
assign LUT_1[854] = 32'b11111111111111111111000011011011;
assign LUT_1[855] = 32'b11111111111111111000010101010111;
assign LUT_1[856] = 32'b11111111111111111010101001101000;
assign LUT_1[857] = 32'b11111111111111110011111011100100;
assign LUT_1[858] = 32'b11111111111111110110010111111001;
assign LUT_1[859] = 32'b11111111111111101111101001110101;
assign LUT_1[860] = 32'b00000000000000000010100010111111;
assign LUT_1[861] = 32'b11111111111111111011110100111011;
assign LUT_1[862] = 32'b11111111111111111110010001010000;
assign LUT_1[863] = 32'b11111111111111110111100011001100;
assign LUT_1[864] = 32'b11111111111111111010011011010000;
assign LUT_1[865] = 32'b11111111111111110011101101001100;
assign LUT_1[866] = 32'b11111111111111110110001001100001;
assign LUT_1[867] = 32'b11111111111111101111011011011101;
assign LUT_1[868] = 32'b00000000000000000010010100100111;
assign LUT_1[869] = 32'b11111111111111111011100110100011;
assign LUT_1[870] = 32'b11111111111111111110000010111000;
assign LUT_1[871] = 32'b11111111111111110111010100110100;
assign LUT_1[872] = 32'b11111111111111111001101001000101;
assign LUT_1[873] = 32'b11111111111111110010111011000001;
assign LUT_1[874] = 32'b11111111111111110101010111010110;
assign LUT_1[875] = 32'b11111111111111101110101001010010;
assign LUT_1[876] = 32'b00000000000000000001100010011100;
assign LUT_1[877] = 32'b11111111111111111010110100011000;
assign LUT_1[878] = 32'b11111111111111111101010000101101;
assign LUT_1[879] = 32'b11111111111111110110100010101001;
assign LUT_1[880] = 32'b11111111111111111100010110110010;
assign LUT_1[881] = 32'b11111111111111110101101000101110;
assign LUT_1[882] = 32'b11111111111111111000000101000011;
assign LUT_1[883] = 32'b11111111111111110001010110111111;
assign LUT_1[884] = 32'b00000000000000000100010000001001;
assign LUT_1[885] = 32'b11111111111111111101100010000101;
assign LUT_1[886] = 32'b11111111111111111111111110011010;
assign LUT_1[887] = 32'b11111111111111111001010000010110;
assign LUT_1[888] = 32'b11111111111111111011100100100111;
assign LUT_1[889] = 32'b11111111111111110100110110100011;
assign LUT_1[890] = 32'b11111111111111110111010010111000;
assign LUT_1[891] = 32'b11111111111111110000100100110100;
assign LUT_1[892] = 32'b00000000000000000011011101111110;
assign LUT_1[893] = 32'b11111111111111111100101111111010;
assign LUT_1[894] = 32'b11111111111111111111001100001111;
assign LUT_1[895] = 32'b11111111111111111000011110001011;
assign LUT_1[896] = 32'b11111111111111111010100010101100;
assign LUT_1[897] = 32'b11111111111111110011110100101000;
assign LUT_1[898] = 32'b11111111111111110110010000111101;
assign LUT_1[899] = 32'b11111111111111101111100010111001;
assign LUT_1[900] = 32'b00000000000000000010011100000011;
assign LUT_1[901] = 32'b11111111111111111011101101111111;
assign LUT_1[902] = 32'b11111111111111111110001010010100;
assign LUT_1[903] = 32'b11111111111111110111011100010000;
assign LUT_1[904] = 32'b11111111111111111001110000100001;
assign LUT_1[905] = 32'b11111111111111110011000010011101;
assign LUT_1[906] = 32'b11111111111111110101011110110010;
assign LUT_1[907] = 32'b11111111111111101110110000101110;
assign LUT_1[908] = 32'b00000000000000000001101001111000;
assign LUT_1[909] = 32'b11111111111111111010111011110100;
assign LUT_1[910] = 32'b11111111111111111101011000001001;
assign LUT_1[911] = 32'b11111111111111110110101010000101;
assign LUT_1[912] = 32'b11111111111111111100011110001110;
assign LUT_1[913] = 32'b11111111111111110101110000001010;
assign LUT_1[914] = 32'b11111111111111111000001100011111;
assign LUT_1[915] = 32'b11111111111111110001011110011011;
assign LUT_1[916] = 32'b00000000000000000100010111100101;
assign LUT_1[917] = 32'b11111111111111111101101001100001;
assign LUT_1[918] = 32'b00000000000000000000000101110110;
assign LUT_1[919] = 32'b11111111111111111001010111110010;
assign LUT_1[920] = 32'b11111111111111111011101100000011;
assign LUT_1[921] = 32'b11111111111111110100111101111111;
assign LUT_1[922] = 32'b11111111111111110111011010010100;
assign LUT_1[923] = 32'b11111111111111110000101100010000;
assign LUT_1[924] = 32'b00000000000000000011100101011010;
assign LUT_1[925] = 32'b11111111111111111100110111010110;
assign LUT_1[926] = 32'b11111111111111111111010011101011;
assign LUT_1[927] = 32'b11111111111111111000100101100111;
assign LUT_1[928] = 32'b11111111111111111011011101101011;
assign LUT_1[929] = 32'b11111111111111110100101111100111;
assign LUT_1[930] = 32'b11111111111111110111001011111100;
assign LUT_1[931] = 32'b11111111111111110000011101111000;
assign LUT_1[932] = 32'b00000000000000000011010111000010;
assign LUT_1[933] = 32'b11111111111111111100101000111110;
assign LUT_1[934] = 32'b11111111111111111111000101010011;
assign LUT_1[935] = 32'b11111111111111111000010111001111;
assign LUT_1[936] = 32'b11111111111111111010101011100000;
assign LUT_1[937] = 32'b11111111111111110011111101011100;
assign LUT_1[938] = 32'b11111111111111110110011001110001;
assign LUT_1[939] = 32'b11111111111111101111101011101101;
assign LUT_1[940] = 32'b00000000000000000010100100110111;
assign LUT_1[941] = 32'b11111111111111111011110110110011;
assign LUT_1[942] = 32'b11111111111111111110010011001000;
assign LUT_1[943] = 32'b11111111111111110111100101000100;
assign LUT_1[944] = 32'b11111111111111111101011001001101;
assign LUT_1[945] = 32'b11111111111111110110101011001001;
assign LUT_1[946] = 32'b11111111111111111001000111011110;
assign LUT_1[947] = 32'b11111111111111110010011001011010;
assign LUT_1[948] = 32'b00000000000000000101010010100100;
assign LUT_1[949] = 32'b11111111111111111110100100100000;
assign LUT_1[950] = 32'b00000000000000000001000000110101;
assign LUT_1[951] = 32'b11111111111111111010010010110001;
assign LUT_1[952] = 32'b11111111111111111100100111000010;
assign LUT_1[953] = 32'b11111111111111110101111000111110;
assign LUT_1[954] = 32'b11111111111111111000010101010011;
assign LUT_1[955] = 32'b11111111111111110001100111001111;
assign LUT_1[956] = 32'b00000000000000000100100000011001;
assign LUT_1[957] = 32'b11111111111111111101110010010101;
assign LUT_1[958] = 32'b00000000000000000000001110101010;
assign LUT_1[959] = 32'b11111111111111111001100000100110;
assign LUT_1[960] = 32'b11111111111111111100100000010100;
assign LUT_1[961] = 32'b11111111111111110101110010010000;
assign LUT_1[962] = 32'b11111111111111111000001110100101;
assign LUT_1[963] = 32'b11111111111111110001100000100001;
assign LUT_1[964] = 32'b00000000000000000100011001101011;
assign LUT_1[965] = 32'b11111111111111111101101011100111;
assign LUT_1[966] = 32'b00000000000000000000000111111100;
assign LUT_1[967] = 32'b11111111111111111001011001111000;
assign LUT_1[968] = 32'b11111111111111111011101110001001;
assign LUT_1[969] = 32'b11111111111111110101000000000101;
assign LUT_1[970] = 32'b11111111111111110111011100011010;
assign LUT_1[971] = 32'b11111111111111110000101110010110;
assign LUT_1[972] = 32'b00000000000000000011100111100000;
assign LUT_1[973] = 32'b11111111111111111100111001011100;
assign LUT_1[974] = 32'b11111111111111111111010101110001;
assign LUT_1[975] = 32'b11111111111111111000100111101101;
assign LUT_1[976] = 32'b11111111111111111110011011110110;
assign LUT_1[977] = 32'b11111111111111110111101101110010;
assign LUT_1[978] = 32'b11111111111111111010001010000111;
assign LUT_1[979] = 32'b11111111111111110011011100000011;
assign LUT_1[980] = 32'b00000000000000000110010101001101;
assign LUT_1[981] = 32'b11111111111111111111100111001001;
assign LUT_1[982] = 32'b00000000000000000010000011011110;
assign LUT_1[983] = 32'b11111111111111111011010101011010;
assign LUT_1[984] = 32'b11111111111111111101101001101011;
assign LUT_1[985] = 32'b11111111111111110110111011100111;
assign LUT_1[986] = 32'b11111111111111111001010111111100;
assign LUT_1[987] = 32'b11111111111111110010101001111000;
assign LUT_1[988] = 32'b00000000000000000101100011000010;
assign LUT_1[989] = 32'b11111111111111111110110100111110;
assign LUT_1[990] = 32'b00000000000000000001010001010011;
assign LUT_1[991] = 32'b11111111111111111010100011001111;
assign LUT_1[992] = 32'b11111111111111111101011011010011;
assign LUT_1[993] = 32'b11111111111111110110101101001111;
assign LUT_1[994] = 32'b11111111111111111001001001100100;
assign LUT_1[995] = 32'b11111111111111110010011011100000;
assign LUT_1[996] = 32'b00000000000000000101010100101010;
assign LUT_1[997] = 32'b11111111111111111110100110100110;
assign LUT_1[998] = 32'b00000000000000000001000010111011;
assign LUT_1[999] = 32'b11111111111111111010010100110111;
assign LUT_1[1000] = 32'b11111111111111111100101001001000;
assign LUT_1[1001] = 32'b11111111111111110101111011000100;
assign LUT_1[1002] = 32'b11111111111111111000010111011001;
assign LUT_1[1003] = 32'b11111111111111110001101001010101;
assign LUT_1[1004] = 32'b00000000000000000100100010011111;
assign LUT_1[1005] = 32'b11111111111111111101110100011011;
assign LUT_1[1006] = 32'b00000000000000000000010000110000;
assign LUT_1[1007] = 32'b11111111111111111001100010101100;
assign LUT_1[1008] = 32'b11111111111111111111010110110101;
assign LUT_1[1009] = 32'b11111111111111111000101000110001;
assign LUT_1[1010] = 32'b11111111111111111011000101000110;
assign LUT_1[1011] = 32'b11111111111111110100010111000010;
assign LUT_1[1012] = 32'b00000000000000000111010000001100;
assign LUT_1[1013] = 32'b00000000000000000000100010001000;
assign LUT_1[1014] = 32'b00000000000000000010111110011101;
assign LUT_1[1015] = 32'b11111111111111111100010000011001;
assign LUT_1[1016] = 32'b11111111111111111110100100101010;
assign LUT_1[1017] = 32'b11111111111111110111110110100110;
assign LUT_1[1018] = 32'b11111111111111111010010010111011;
assign LUT_1[1019] = 32'b11111111111111110011100100110111;
assign LUT_1[1020] = 32'b00000000000000000110011110000001;
assign LUT_1[1021] = 32'b11111111111111111111101111111101;
assign LUT_1[1022] = 32'b00000000000000000010001100010010;
assign LUT_1[1023] = 32'b11111111111111111011011110001110;
assign LUT_1[1024] = 32'b00000000000000000110010110110000;
assign LUT_1[1025] = 32'b11111111111111111111101000101100;
assign LUT_1[1026] = 32'b00000000000000000010000101000001;
assign LUT_1[1027] = 32'b11111111111111111011010110111101;
assign LUT_1[1028] = 32'b00000000000000001110010000000111;
assign LUT_1[1029] = 32'b00000000000000000111100010000011;
assign LUT_1[1030] = 32'b00000000000000001001111110011000;
assign LUT_1[1031] = 32'b00000000000000000011010000010100;
assign LUT_1[1032] = 32'b00000000000000000101100100100101;
assign LUT_1[1033] = 32'b11111111111111111110110110100001;
assign LUT_1[1034] = 32'b00000000000000000001010010110110;
assign LUT_1[1035] = 32'b11111111111111111010100100110010;
assign LUT_1[1036] = 32'b00000000000000001101011101111100;
assign LUT_1[1037] = 32'b00000000000000000110101111111000;
assign LUT_1[1038] = 32'b00000000000000001001001100001101;
assign LUT_1[1039] = 32'b00000000000000000010011110001001;
assign LUT_1[1040] = 32'b00000000000000001000010010010010;
assign LUT_1[1041] = 32'b00000000000000000001100100001110;
assign LUT_1[1042] = 32'b00000000000000000100000000100011;
assign LUT_1[1043] = 32'b11111111111111111101010010011111;
assign LUT_1[1044] = 32'b00000000000000010000001011101001;
assign LUT_1[1045] = 32'b00000000000000001001011101100101;
assign LUT_1[1046] = 32'b00000000000000001011111001111010;
assign LUT_1[1047] = 32'b00000000000000000101001011110110;
assign LUT_1[1048] = 32'b00000000000000000111100000000111;
assign LUT_1[1049] = 32'b00000000000000000000110010000011;
assign LUT_1[1050] = 32'b00000000000000000011001110011000;
assign LUT_1[1051] = 32'b11111111111111111100100000010100;
assign LUT_1[1052] = 32'b00000000000000001111011001011110;
assign LUT_1[1053] = 32'b00000000000000001000101011011010;
assign LUT_1[1054] = 32'b00000000000000001011000111101111;
assign LUT_1[1055] = 32'b00000000000000000100011001101011;
assign LUT_1[1056] = 32'b00000000000000000111010001101111;
assign LUT_1[1057] = 32'b00000000000000000000100011101011;
assign LUT_1[1058] = 32'b00000000000000000011000000000000;
assign LUT_1[1059] = 32'b11111111111111111100010001111100;
assign LUT_1[1060] = 32'b00000000000000001111001011000110;
assign LUT_1[1061] = 32'b00000000000000001000011101000010;
assign LUT_1[1062] = 32'b00000000000000001010111001010111;
assign LUT_1[1063] = 32'b00000000000000000100001011010011;
assign LUT_1[1064] = 32'b00000000000000000110011111100100;
assign LUT_1[1065] = 32'b11111111111111111111110001100000;
assign LUT_1[1066] = 32'b00000000000000000010001101110101;
assign LUT_1[1067] = 32'b11111111111111111011011111110001;
assign LUT_1[1068] = 32'b00000000000000001110011000111011;
assign LUT_1[1069] = 32'b00000000000000000111101010110111;
assign LUT_1[1070] = 32'b00000000000000001010000111001100;
assign LUT_1[1071] = 32'b00000000000000000011011001001000;
assign LUT_1[1072] = 32'b00000000000000001001001101010001;
assign LUT_1[1073] = 32'b00000000000000000010011111001101;
assign LUT_1[1074] = 32'b00000000000000000100111011100010;
assign LUT_1[1075] = 32'b11111111111111111110001101011110;
assign LUT_1[1076] = 32'b00000000000000010001000110101000;
assign LUT_1[1077] = 32'b00000000000000001010011000100100;
assign LUT_1[1078] = 32'b00000000000000001100110100111001;
assign LUT_1[1079] = 32'b00000000000000000110000110110101;
assign LUT_1[1080] = 32'b00000000000000001000011011000110;
assign LUT_1[1081] = 32'b00000000000000000001101101000010;
assign LUT_1[1082] = 32'b00000000000000000100001001010111;
assign LUT_1[1083] = 32'b11111111111111111101011011010011;
assign LUT_1[1084] = 32'b00000000000000010000010100011101;
assign LUT_1[1085] = 32'b00000000000000001001100110011001;
assign LUT_1[1086] = 32'b00000000000000001100000010101110;
assign LUT_1[1087] = 32'b00000000000000000101010100101010;
assign LUT_1[1088] = 32'b00000000000000001000010100011000;
assign LUT_1[1089] = 32'b00000000000000000001100110010100;
assign LUT_1[1090] = 32'b00000000000000000100000010101001;
assign LUT_1[1091] = 32'b11111111111111111101010100100101;
assign LUT_1[1092] = 32'b00000000000000010000001101101111;
assign LUT_1[1093] = 32'b00000000000000001001011111101011;
assign LUT_1[1094] = 32'b00000000000000001011111100000000;
assign LUT_1[1095] = 32'b00000000000000000101001101111100;
assign LUT_1[1096] = 32'b00000000000000000111100010001101;
assign LUT_1[1097] = 32'b00000000000000000000110100001001;
assign LUT_1[1098] = 32'b00000000000000000011010000011110;
assign LUT_1[1099] = 32'b11111111111111111100100010011010;
assign LUT_1[1100] = 32'b00000000000000001111011011100100;
assign LUT_1[1101] = 32'b00000000000000001000101101100000;
assign LUT_1[1102] = 32'b00000000000000001011001001110101;
assign LUT_1[1103] = 32'b00000000000000000100011011110001;
assign LUT_1[1104] = 32'b00000000000000001010001111111010;
assign LUT_1[1105] = 32'b00000000000000000011100001110110;
assign LUT_1[1106] = 32'b00000000000000000101111110001011;
assign LUT_1[1107] = 32'b11111111111111111111010000000111;
assign LUT_1[1108] = 32'b00000000000000010010001001010001;
assign LUT_1[1109] = 32'b00000000000000001011011011001101;
assign LUT_1[1110] = 32'b00000000000000001101110111100010;
assign LUT_1[1111] = 32'b00000000000000000111001001011110;
assign LUT_1[1112] = 32'b00000000000000001001011101101111;
assign LUT_1[1113] = 32'b00000000000000000010101111101011;
assign LUT_1[1114] = 32'b00000000000000000101001100000000;
assign LUT_1[1115] = 32'b11111111111111111110011101111100;
assign LUT_1[1116] = 32'b00000000000000010001010111000110;
assign LUT_1[1117] = 32'b00000000000000001010101001000010;
assign LUT_1[1118] = 32'b00000000000000001101000101010111;
assign LUT_1[1119] = 32'b00000000000000000110010111010011;
assign LUT_1[1120] = 32'b00000000000000001001001111010111;
assign LUT_1[1121] = 32'b00000000000000000010100001010011;
assign LUT_1[1122] = 32'b00000000000000000100111101101000;
assign LUT_1[1123] = 32'b11111111111111111110001111100100;
assign LUT_1[1124] = 32'b00000000000000010001001000101110;
assign LUT_1[1125] = 32'b00000000000000001010011010101010;
assign LUT_1[1126] = 32'b00000000000000001100110110111111;
assign LUT_1[1127] = 32'b00000000000000000110001000111011;
assign LUT_1[1128] = 32'b00000000000000001000011101001100;
assign LUT_1[1129] = 32'b00000000000000000001101111001000;
assign LUT_1[1130] = 32'b00000000000000000100001011011101;
assign LUT_1[1131] = 32'b11111111111111111101011101011001;
assign LUT_1[1132] = 32'b00000000000000010000010110100011;
assign LUT_1[1133] = 32'b00000000000000001001101000011111;
assign LUT_1[1134] = 32'b00000000000000001100000100110100;
assign LUT_1[1135] = 32'b00000000000000000101010110110000;
assign LUT_1[1136] = 32'b00000000000000001011001010111001;
assign LUT_1[1137] = 32'b00000000000000000100011100110101;
assign LUT_1[1138] = 32'b00000000000000000110111001001010;
assign LUT_1[1139] = 32'b00000000000000000000001011000110;
assign LUT_1[1140] = 32'b00000000000000010011000100010000;
assign LUT_1[1141] = 32'b00000000000000001100010110001100;
assign LUT_1[1142] = 32'b00000000000000001110110010100001;
assign LUT_1[1143] = 32'b00000000000000001000000100011101;
assign LUT_1[1144] = 32'b00000000000000001010011000101110;
assign LUT_1[1145] = 32'b00000000000000000011101010101010;
assign LUT_1[1146] = 32'b00000000000000000110000110111111;
assign LUT_1[1147] = 32'b11111111111111111111011000111011;
assign LUT_1[1148] = 32'b00000000000000010010010010000101;
assign LUT_1[1149] = 32'b00000000000000001011100100000001;
assign LUT_1[1150] = 32'b00000000000000001110000000010110;
assign LUT_1[1151] = 32'b00000000000000000111010010010010;
assign LUT_1[1152] = 32'b00000000000000001001010110110011;
assign LUT_1[1153] = 32'b00000000000000000010101000101111;
assign LUT_1[1154] = 32'b00000000000000000101000101000100;
assign LUT_1[1155] = 32'b11111111111111111110010111000000;
assign LUT_1[1156] = 32'b00000000000000010001010000001010;
assign LUT_1[1157] = 32'b00000000000000001010100010000110;
assign LUT_1[1158] = 32'b00000000000000001100111110011011;
assign LUT_1[1159] = 32'b00000000000000000110010000010111;
assign LUT_1[1160] = 32'b00000000000000001000100100101000;
assign LUT_1[1161] = 32'b00000000000000000001110110100100;
assign LUT_1[1162] = 32'b00000000000000000100010010111001;
assign LUT_1[1163] = 32'b11111111111111111101100100110101;
assign LUT_1[1164] = 32'b00000000000000010000011101111111;
assign LUT_1[1165] = 32'b00000000000000001001101111111011;
assign LUT_1[1166] = 32'b00000000000000001100001100010000;
assign LUT_1[1167] = 32'b00000000000000000101011110001100;
assign LUT_1[1168] = 32'b00000000000000001011010010010101;
assign LUT_1[1169] = 32'b00000000000000000100100100010001;
assign LUT_1[1170] = 32'b00000000000000000111000000100110;
assign LUT_1[1171] = 32'b00000000000000000000010010100010;
assign LUT_1[1172] = 32'b00000000000000010011001011101100;
assign LUT_1[1173] = 32'b00000000000000001100011101101000;
assign LUT_1[1174] = 32'b00000000000000001110111001111101;
assign LUT_1[1175] = 32'b00000000000000001000001011111001;
assign LUT_1[1176] = 32'b00000000000000001010100000001010;
assign LUT_1[1177] = 32'b00000000000000000011110010000110;
assign LUT_1[1178] = 32'b00000000000000000110001110011011;
assign LUT_1[1179] = 32'b11111111111111111111100000010111;
assign LUT_1[1180] = 32'b00000000000000010010011001100001;
assign LUT_1[1181] = 32'b00000000000000001011101011011101;
assign LUT_1[1182] = 32'b00000000000000001110000111110010;
assign LUT_1[1183] = 32'b00000000000000000111011001101110;
assign LUT_1[1184] = 32'b00000000000000001010010001110010;
assign LUT_1[1185] = 32'b00000000000000000011100011101110;
assign LUT_1[1186] = 32'b00000000000000000110000000000011;
assign LUT_1[1187] = 32'b11111111111111111111010001111111;
assign LUT_1[1188] = 32'b00000000000000010010001011001001;
assign LUT_1[1189] = 32'b00000000000000001011011101000101;
assign LUT_1[1190] = 32'b00000000000000001101111001011010;
assign LUT_1[1191] = 32'b00000000000000000111001011010110;
assign LUT_1[1192] = 32'b00000000000000001001011111100111;
assign LUT_1[1193] = 32'b00000000000000000010110001100011;
assign LUT_1[1194] = 32'b00000000000000000101001101111000;
assign LUT_1[1195] = 32'b11111111111111111110011111110100;
assign LUT_1[1196] = 32'b00000000000000010001011000111110;
assign LUT_1[1197] = 32'b00000000000000001010101010111010;
assign LUT_1[1198] = 32'b00000000000000001101000111001111;
assign LUT_1[1199] = 32'b00000000000000000110011001001011;
assign LUT_1[1200] = 32'b00000000000000001100001101010100;
assign LUT_1[1201] = 32'b00000000000000000101011111010000;
assign LUT_1[1202] = 32'b00000000000000000111111011100101;
assign LUT_1[1203] = 32'b00000000000000000001001101100001;
assign LUT_1[1204] = 32'b00000000000000010100000110101011;
assign LUT_1[1205] = 32'b00000000000000001101011000100111;
assign LUT_1[1206] = 32'b00000000000000001111110100111100;
assign LUT_1[1207] = 32'b00000000000000001001000110111000;
assign LUT_1[1208] = 32'b00000000000000001011011011001001;
assign LUT_1[1209] = 32'b00000000000000000100101101000101;
assign LUT_1[1210] = 32'b00000000000000000111001001011010;
assign LUT_1[1211] = 32'b00000000000000000000011011010110;
assign LUT_1[1212] = 32'b00000000000000010011010100100000;
assign LUT_1[1213] = 32'b00000000000000001100100110011100;
assign LUT_1[1214] = 32'b00000000000000001111000010110001;
assign LUT_1[1215] = 32'b00000000000000001000010100101101;
assign LUT_1[1216] = 32'b00000000000000001011010100011011;
assign LUT_1[1217] = 32'b00000000000000000100100110010111;
assign LUT_1[1218] = 32'b00000000000000000111000010101100;
assign LUT_1[1219] = 32'b00000000000000000000010100101000;
assign LUT_1[1220] = 32'b00000000000000010011001101110010;
assign LUT_1[1221] = 32'b00000000000000001100011111101110;
assign LUT_1[1222] = 32'b00000000000000001110111100000011;
assign LUT_1[1223] = 32'b00000000000000001000001101111111;
assign LUT_1[1224] = 32'b00000000000000001010100010010000;
assign LUT_1[1225] = 32'b00000000000000000011110100001100;
assign LUT_1[1226] = 32'b00000000000000000110010000100001;
assign LUT_1[1227] = 32'b11111111111111111111100010011101;
assign LUT_1[1228] = 32'b00000000000000010010011011100111;
assign LUT_1[1229] = 32'b00000000000000001011101101100011;
assign LUT_1[1230] = 32'b00000000000000001110001001111000;
assign LUT_1[1231] = 32'b00000000000000000111011011110100;
assign LUT_1[1232] = 32'b00000000000000001101001111111101;
assign LUT_1[1233] = 32'b00000000000000000110100001111001;
assign LUT_1[1234] = 32'b00000000000000001000111110001110;
assign LUT_1[1235] = 32'b00000000000000000010010000001010;
assign LUT_1[1236] = 32'b00000000000000010101001001010100;
assign LUT_1[1237] = 32'b00000000000000001110011011010000;
assign LUT_1[1238] = 32'b00000000000000010000110111100101;
assign LUT_1[1239] = 32'b00000000000000001010001001100001;
assign LUT_1[1240] = 32'b00000000000000001100011101110010;
assign LUT_1[1241] = 32'b00000000000000000101101111101110;
assign LUT_1[1242] = 32'b00000000000000001000001100000011;
assign LUT_1[1243] = 32'b00000000000000000001011101111111;
assign LUT_1[1244] = 32'b00000000000000010100010111001001;
assign LUT_1[1245] = 32'b00000000000000001101101001000101;
assign LUT_1[1246] = 32'b00000000000000010000000101011010;
assign LUT_1[1247] = 32'b00000000000000001001010111010110;
assign LUT_1[1248] = 32'b00000000000000001100001111011010;
assign LUT_1[1249] = 32'b00000000000000000101100001010110;
assign LUT_1[1250] = 32'b00000000000000000111111101101011;
assign LUT_1[1251] = 32'b00000000000000000001001111100111;
assign LUT_1[1252] = 32'b00000000000000010100001000110001;
assign LUT_1[1253] = 32'b00000000000000001101011010101101;
assign LUT_1[1254] = 32'b00000000000000001111110111000010;
assign LUT_1[1255] = 32'b00000000000000001001001000111110;
assign LUT_1[1256] = 32'b00000000000000001011011101001111;
assign LUT_1[1257] = 32'b00000000000000000100101111001011;
assign LUT_1[1258] = 32'b00000000000000000111001011100000;
assign LUT_1[1259] = 32'b00000000000000000000011101011100;
assign LUT_1[1260] = 32'b00000000000000010011010110100110;
assign LUT_1[1261] = 32'b00000000000000001100101000100010;
assign LUT_1[1262] = 32'b00000000000000001111000100110111;
assign LUT_1[1263] = 32'b00000000000000001000010110110011;
assign LUT_1[1264] = 32'b00000000000000001110001010111100;
assign LUT_1[1265] = 32'b00000000000000000111011100111000;
assign LUT_1[1266] = 32'b00000000000000001001111001001101;
assign LUT_1[1267] = 32'b00000000000000000011001011001001;
assign LUT_1[1268] = 32'b00000000000000010110000100010011;
assign LUT_1[1269] = 32'b00000000000000001111010110001111;
assign LUT_1[1270] = 32'b00000000000000010001110010100100;
assign LUT_1[1271] = 32'b00000000000000001011000100100000;
assign LUT_1[1272] = 32'b00000000000000001101011000110001;
assign LUT_1[1273] = 32'b00000000000000000110101010101101;
assign LUT_1[1274] = 32'b00000000000000001001000111000010;
assign LUT_1[1275] = 32'b00000000000000000010011000111110;
assign LUT_1[1276] = 32'b00000000000000010101010010001000;
assign LUT_1[1277] = 32'b00000000000000001110100100000100;
assign LUT_1[1278] = 32'b00000000000000010001000000011001;
assign LUT_1[1279] = 32'b00000000000000001010010010010101;
assign LUT_1[1280] = 32'b00000000000000000100001010111100;
assign LUT_1[1281] = 32'b11111111111111111101011100111000;
assign LUT_1[1282] = 32'b11111111111111111111111001001101;
assign LUT_1[1283] = 32'b11111111111111111001001011001001;
assign LUT_1[1284] = 32'b00000000000000001100000100010011;
assign LUT_1[1285] = 32'b00000000000000000101010110001111;
assign LUT_1[1286] = 32'b00000000000000000111110010100100;
assign LUT_1[1287] = 32'b00000000000000000001000100100000;
assign LUT_1[1288] = 32'b00000000000000000011011000110001;
assign LUT_1[1289] = 32'b11111111111111111100101010101101;
assign LUT_1[1290] = 32'b11111111111111111111000111000010;
assign LUT_1[1291] = 32'b11111111111111111000011000111110;
assign LUT_1[1292] = 32'b00000000000000001011010010001000;
assign LUT_1[1293] = 32'b00000000000000000100100100000100;
assign LUT_1[1294] = 32'b00000000000000000111000000011001;
assign LUT_1[1295] = 32'b00000000000000000000010010010101;
assign LUT_1[1296] = 32'b00000000000000000110000110011110;
assign LUT_1[1297] = 32'b11111111111111111111011000011010;
assign LUT_1[1298] = 32'b00000000000000000001110100101111;
assign LUT_1[1299] = 32'b11111111111111111011000110101011;
assign LUT_1[1300] = 32'b00000000000000001101111111110101;
assign LUT_1[1301] = 32'b00000000000000000111010001110001;
assign LUT_1[1302] = 32'b00000000000000001001101110000110;
assign LUT_1[1303] = 32'b00000000000000000011000000000010;
assign LUT_1[1304] = 32'b00000000000000000101010100010011;
assign LUT_1[1305] = 32'b11111111111111111110100110001111;
assign LUT_1[1306] = 32'b00000000000000000001000010100100;
assign LUT_1[1307] = 32'b11111111111111111010010100100000;
assign LUT_1[1308] = 32'b00000000000000001101001101101010;
assign LUT_1[1309] = 32'b00000000000000000110011111100110;
assign LUT_1[1310] = 32'b00000000000000001000111011111011;
assign LUT_1[1311] = 32'b00000000000000000010001101110111;
assign LUT_1[1312] = 32'b00000000000000000101000101111011;
assign LUT_1[1313] = 32'b11111111111111111110010111110111;
assign LUT_1[1314] = 32'b00000000000000000000110100001100;
assign LUT_1[1315] = 32'b11111111111111111010000110001000;
assign LUT_1[1316] = 32'b00000000000000001100111111010010;
assign LUT_1[1317] = 32'b00000000000000000110010001001110;
assign LUT_1[1318] = 32'b00000000000000001000101101100011;
assign LUT_1[1319] = 32'b00000000000000000001111111011111;
assign LUT_1[1320] = 32'b00000000000000000100010011110000;
assign LUT_1[1321] = 32'b11111111111111111101100101101100;
assign LUT_1[1322] = 32'b00000000000000000000000010000001;
assign LUT_1[1323] = 32'b11111111111111111001010011111101;
assign LUT_1[1324] = 32'b00000000000000001100001101000111;
assign LUT_1[1325] = 32'b00000000000000000101011111000011;
assign LUT_1[1326] = 32'b00000000000000000111111011011000;
assign LUT_1[1327] = 32'b00000000000000000001001101010100;
assign LUT_1[1328] = 32'b00000000000000000111000001011101;
assign LUT_1[1329] = 32'b00000000000000000000010011011001;
assign LUT_1[1330] = 32'b00000000000000000010101111101110;
assign LUT_1[1331] = 32'b11111111111111111100000001101010;
assign LUT_1[1332] = 32'b00000000000000001110111010110100;
assign LUT_1[1333] = 32'b00000000000000001000001100110000;
assign LUT_1[1334] = 32'b00000000000000001010101001000101;
assign LUT_1[1335] = 32'b00000000000000000011111011000001;
assign LUT_1[1336] = 32'b00000000000000000110001111010010;
assign LUT_1[1337] = 32'b11111111111111111111100001001110;
assign LUT_1[1338] = 32'b00000000000000000001111101100011;
assign LUT_1[1339] = 32'b11111111111111111011001111011111;
assign LUT_1[1340] = 32'b00000000000000001110001000101001;
assign LUT_1[1341] = 32'b00000000000000000111011010100101;
assign LUT_1[1342] = 32'b00000000000000001001110110111010;
assign LUT_1[1343] = 32'b00000000000000000011001000110110;
assign LUT_1[1344] = 32'b00000000000000000110001000100100;
assign LUT_1[1345] = 32'b11111111111111111111011010100000;
assign LUT_1[1346] = 32'b00000000000000000001110110110101;
assign LUT_1[1347] = 32'b11111111111111111011001000110001;
assign LUT_1[1348] = 32'b00000000000000001110000001111011;
assign LUT_1[1349] = 32'b00000000000000000111010011110111;
assign LUT_1[1350] = 32'b00000000000000001001110000001100;
assign LUT_1[1351] = 32'b00000000000000000011000010001000;
assign LUT_1[1352] = 32'b00000000000000000101010110011001;
assign LUT_1[1353] = 32'b11111111111111111110101000010101;
assign LUT_1[1354] = 32'b00000000000000000001000100101010;
assign LUT_1[1355] = 32'b11111111111111111010010110100110;
assign LUT_1[1356] = 32'b00000000000000001101001111110000;
assign LUT_1[1357] = 32'b00000000000000000110100001101100;
assign LUT_1[1358] = 32'b00000000000000001000111110000001;
assign LUT_1[1359] = 32'b00000000000000000010001111111101;
assign LUT_1[1360] = 32'b00000000000000001000000100000110;
assign LUT_1[1361] = 32'b00000000000000000001010110000010;
assign LUT_1[1362] = 32'b00000000000000000011110010010111;
assign LUT_1[1363] = 32'b11111111111111111101000100010011;
assign LUT_1[1364] = 32'b00000000000000001111111101011101;
assign LUT_1[1365] = 32'b00000000000000001001001111011001;
assign LUT_1[1366] = 32'b00000000000000001011101011101110;
assign LUT_1[1367] = 32'b00000000000000000100111101101010;
assign LUT_1[1368] = 32'b00000000000000000111010001111011;
assign LUT_1[1369] = 32'b00000000000000000000100011110111;
assign LUT_1[1370] = 32'b00000000000000000011000000001100;
assign LUT_1[1371] = 32'b11111111111111111100010010001000;
assign LUT_1[1372] = 32'b00000000000000001111001011010010;
assign LUT_1[1373] = 32'b00000000000000001000011101001110;
assign LUT_1[1374] = 32'b00000000000000001010111001100011;
assign LUT_1[1375] = 32'b00000000000000000100001011011111;
assign LUT_1[1376] = 32'b00000000000000000111000011100011;
assign LUT_1[1377] = 32'b00000000000000000000010101011111;
assign LUT_1[1378] = 32'b00000000000000000010110001110100;
assign LUT_1[1379] = 32'b11111111111111111100000011110000;
assign LUT_1[1380] = 32'b00000000000000001110111100111010;
assign LUT_1[1381] = 32'b00000000000000001000001110110110;
assign LUT_1[1382] = 32'b00000000000000001010101011001011;
assign LUT_1[1383] = 32'b00000000000000000011111101000111;
assign LUT_1[1384] = 32'b00000000000000000110010001011000;
assign LUT_1[1385] = 32'b11111111111111111111100011010100;
assign LUT_1[1386] = 32'b00000000000000000001111111101001;
assign LUT_1[1387] = 32'b11111111111111111011010001100101;
assign LUT_1[1388] = 32'b00000000000000001110001010101111;
assign LUT_1[1389] = 32'b00000000000000000111011100101011;
assign LUT_1[1390] = 32'b00000000000000001001111001000000;
assign LUT_1[1391] = 32'b00000000000000000011001010111100;
assign LUT_1[1392] = 32'b00000000000000001000111111000101;
assign LUT_1[1393] = 32'b00000000000000000010010001000001;
assign LUT_1[1394] = 32'b00000000000000000100101101010110;
assign LUT_1[1395] = 32'b11111111111111111101111111010010;
assign LUT_1[1396] = 32'b00000000000000010000111000011100;
assign LUT_1[1397] = 32'b00000000000000001010001010011000;
assign LUT_1[1398] = 32'b00000000000000001100100110101101;
assign LUT_1[1399] = 32'b00000000000000000101111000101001;
assign LUT_1[1400] = 32'b00000000000000001000001100111010;
assign LUT_1[1401] = 32'b00000000000000000001011110110110;
assign LUT_1[1402] = 32'b00000000000000000011111011001011;
assign LUT_1[1403] = 32'b11111111111111111101001101000111;
assign LUT_1[1404] = 32'b00000000000000010000000110010001;
assign LUT_1[1405] = 32'b00000000000000001001011000001101;
assign LUT_1[1406] = 32'b00000000000000001011110100100010;
assign LUT_1[1407] = 32'b00000000000000000101000110011110;
assign LUT_1[1408] = 32'b00000000000000000111001010111111;
assign LUT_1[1409] = 32'b00000000000000000000011100111011;
assign LUT_1[1410] = 32'b00000000000000000010111001010000;
assign LUT_1[1411] = 32'b11111111111111111100001011001100;
assign LUT_1[1412] = 32'b00000000000000001111000100010110;
assign LUT_1[1413] = 32'b00000000000000001000010110010010;
assign LUT_1[1414] = 32'b00000000000000001010110010100111;
assign LUT_1[1415] = 32'b00000000000000000100000100100011;
assign LUT_1[1416] = 32'b00000000000000000110011000110100;
assign LUT_1[1417] = 32'b11111111111111111111101010110000;
assign LUT_1[1418] = 32'b00000000000000000010000111000101;
assign LUT_1[1419] = 32'b11111111111111111011011001000001;
assign LUT_1[1420] = 32'b00000000000000001110010010001011;
assign LUT_1[1421] = 32'b00000000000000000111100100000111;
assign LUT_1[1422] = 32'b00000000000000001010000000011100;
assign LUT_1[1423] = 32'b00000000000000000011010010011000;
assign LUT_1[1424] = 32'b00000000000000001001000110100001;
assign LUT_1[1425] = 32'b00000000000000000010011000011101;
assign LUT_1[1426] = 32'b00000000000000000100110100110010;
assign LUT_1[1427] = 32'b11111111111111111110000110101110;
assign LUT_1[1428] = 32'b00000000000000010000111111111000;
assign LUT_1[1429] = 32'b00000000000000001010010001110100;
assign LUT_1[1430] = 32'b00000000000000001100101110001001;
assign LUT_1[1431] = 32'b00000000000000000110000000000101;
assign LUT_1[1432] = 32'b00000000000000001000010100010110;
assign LUT_1[1433] = 32'b00000000000000000001100110010010;
assign LUT_1[1434] = 32'b00000000000000000100000010100111;
assign LUT_1[1435] = 32'b11111111111111111101010100100011;
assign LUT_1[1436] = 32'b00000000000000010000001101101101;
assign LUT_1[1437] = 32'b00000000000000001001011111101001;
assign LUT_1[1438] = 32'b00000000000000001011111011111110;
assign LUT_1[1439] = 32'b00000000000000000101001101111010;
assign LUT_1[1440] = 32'b00000000000000001000000101111110;
assign LUT_1[1441] = 32'b00000000000000000001010111111010;
assign LUT_1[1442] = 32'b00000000000000000011110100001111;
assign LUT_1[1443] = 32'b11111111111111111101000110001011;
assign LUT_1[1444] = 32'b00000000000000001111111111010101;
assign LUT_1[1445] = 32'b00000000000000001001010001010001;
assign LUT_1[1446] = 32'b00000000000000001011101101100110;
assign LUT_1[1447] = 32'b00000000000000000100111111100010;
assign LUT_1[1448] = 32'b00000000000000000111010011110011;
assign LUT_1[1449] = 32'b00000000000000000000100101101111;
assign LUT_1[1450] = 32'b00000000000000000011000010000100;
assign LUT_1[1451] = 32'b11111111111111111100010100000000;
assign LUT_1[1452] = 32'b00000000000000001111001101001010;
assign LUT_1[1453] = 32'b00000000000000001000011111000110;
assign LUT_1[1454] = 32'b00000000000000001010111011011011;
assign LUT_1[1455] = 32'b00000000000000000100001101010111;
assign LUT_1[1456] = 32'b00000000000000001010000001100000;
assign LUT_1[1457] = 32'b00000000000000000011010011011100;
assign LUT_1[1458] = 32'b00000000000000000101101111110001;
assign LUT_1[1459] = 32'b11111111111111111111000001101101;
assign LUT_1[1460] = 32'b00000000000000010001111010110111;
assign LUT_1[1461] = 32'b00000000000000001011001100110011;
assign LUT_1[1462] = 32'b00000000000000001101101001001000;
assign LUT_1[1463] = 32'b00000000000000000110111011000100;
assign LUT_1[1464] = 32'b00000000000000001001001111010101;
assign LUT_1[1465] = 32'b00000000000000000010100001010001;
assign LUT_1[1466] = 32'b00000000000000000100111101100110;
assign LUT_1[1467] = 32'b11111111111111111110001111100010;
assign LUT_1[1468] = 32'b00000000000000010001001000101100;
assign LUT_1[1469] = 32'b00000000000000001010011010101000;
assign LUT_1[1470] = 32'b00000000000000001100110110111101;
assign LUT_1[1471] = 32'b00000000000000000110001000111001;
assign LUT_1[1472] = 32'b00000000000000001001001000100111;
assign LUT_1[1473] = 32'b00000000000000000010011010100011;
assign LUT_1[1474] = 32'b00000000000000000100110110111000;
assign LUT_1[1475] = 32'b11111111111111111110001000110100;
assign LUT_1[1476] = 32'b00000000000000010001000001111110;
assign LUT_1[1477] = 32'b00000000000000001010010011111010;
assign LUT_1[1478] = 32'b00000000000000001100110000001111;
assign LUT_1[1479] = 32'b00000000000000000110000010001011;
assign LUT_1[1480] = 32'b00000000000000001000010110011100;
assign LUT_1[1481] = 32'b00000000000000000001101000011000;
assign LUT_1[1482] = 32'b00000000000000000100000100101101;
assign LUT_1[1483] = 32'b11111111111111111101010110101001;
assign LUT_1[1484] = 32'b00000000000000010000001111110011;
assign LUT_1[1485] = 32'b00000000000000001001100001101111;
assign LUT_1[1486] = 32'b00000000000000001011111110000100;
assign LUT_1[1487] = 32'b00000000000000000101010000000000;
assign LUT_1[1488] = 32'b00000000000000001011000100001001;
assign LUT_1[1489] = 32'b00000000000000000100010110000101;
assign LUT_1[1490] = 32'b00000000000000000110110010011010;
assign LUT_1[1491] = 32'b00000000000000000000000100010110;
assign LUT_1[1492] = 32'b00000000000000010010111101100000;
assign LUT_1[1493] = 32'b00000000000000001100001111011100;
assign LUT_1[1494] = 32'b00000000000000001110101011110001;
assign LUT_1[1495] = 32'b00000000000000000111111101101101;
assign LUT_1[1496] = 32'b00000000000000001010010001111110;
assign LUT_1[1497] = 32'b00000000000000000011100011111010;
assign LUT_1[1498] = 32'b00000000000000000110000000001111;
assign LUT_1[1499] = 32'b11111111111111111111010010001011;
assign LUT_1[1500] = 32'b00000000000000010010001011010101;
assign LUT_1[1501] = 32'b00000000000000001011011101010001;
assign LUT_1[1502] = 32'b00000000000000001101111001100110;
assign LUT_1[1503] = 32'b00000000000000000111001011100010;
assign LUT_1[1504] = 32'b00000000000000001010000011100110;
assign LUT_1[1505] = 32'b00000000000000000011010101100010;
assign LUT_1[1506] = 32'b00000000000000000101110001110111;
assign LUT_1[1507] = 32'b11111111111111111111000011110011;
assign LUT_1[1508] = 32'b00000000000000010001111100111101;
assign LUT_1[1509] = 32'b00000000000000001011001110111001;
assign LUT_1[1510] = 32'b00000000000000001101101011001110;
assign LUT_1[1511] = 32'b00000000000000000110111101001010;
assign LUT_1[1512] = 32'b00000000000000001001010001011011;
assign LUT_1[1513] = 32'b00000000000000000010100011010111;
assign LUT_1[1514] = 32'b00000000000000000100111111101100;
assign LUT_1[1515] = 32'b11111111111111111110010001101000;
assign LUT_1[1516] = 32'b00000000000000010001001010110010;
assign LUT_1[1517] = 32'b00000000000000001010011100101110;
assign LUT_1[1518] = 32'b00000000000000001100111001000011;
assign LUT_1[1519] = 32'b00000000000000000110001010111111;
assign LUT_1[1520] = 32'b00000000000000001011111111001000;
assign LUT_1[1521] = 32'b00000000000000000101010001000100;
assign LUT_1[1522] = 32'b00000000000000000111101101011001;
assign LUT_1[1523] = 32'b00000000000000000000111111010101;
assign LUT_1[1524] = 32'b00000000000000010011111000011111;
assign LUT_1[1525] = 32'b00000000000000001101001010011011;
assign LUT_1[1526] = 32'b00000000000000001111100110110000;
assign LUT_1[1527] = 32'b00000000000000001000111000101100;
assign LUT_1[1528] = 32'b00000000000000001011001100111101;
assign LUT_1[1529] = 32'b00000000000000000100011110111001;
assign LUT_1[1530] = 32'b00000000000000000110111011001110;
assign LUT_1[1531] = 32'b00000000000000000000001101001010;
assign LUT_1[1532] = 32'b00000000000000010011000110010100;
assign LUT_1[1533] = 32'b00000000000000001100011000010000;
assign LUT_1[1534] = 32'b00000000000000001110110100100101;
assign LUT_1[1535] = 32'b00000000000000001000000110100001;
assign LUT_1[1536] = 32'b00000000000000000000000101001101;
assign LUT_1[1537] = 32'b11111111111111111001010111001001;
assign LUT_1[1538] = 32'b11111111111111111011110011011110;
assign LUT_1[1539] = 32'b11111111111111110101000101011010;
assign LUT_1[1540] = 32'b00000000000000000111111110100100;
assign LUT_1[1541] = 32'b00000000000000000001010000100000;
assign LUT_1[1542] = 32'b00000000000000000011101100110101;
assign LUT_1[1543] = 32'b11111111111111111100111110110001;
assign LUT_1[1544] = 32'b11111111111111111111010011000010;
assign LUT_1[1545] = 32'b11111111111111111000100100111110;
assign LUT_1[1546] = 32'b11111111111111111011000001010011;
assign LUT_1[1547] = 32'b11111111111111110100010011001111;
assign LUT_1[1548] = 32'b00000000000000000111001100011001;
assign LUT_1[1549] = 32'b00000000000000000000011110010101;
assign LUT_1[1550] = 32'b00000000000000000010111010101010;
assign LUT_1[1551] = 32'b11111111111111111100001100100110;
assign LUT_1[1552] = 32'b00000000000000000010000000101111;
assign LUT_1[1553] = 32'b11111111111111111011010010101011;
assign LUT_1[1554] = 32'b11111111111111111101101111000000;
assign LUT_1[1555] = 32'b11111111111111110111000000111100;
assign LUT_1[1556] = 32'b00000000000000001001111010000110;
assign LUT_1[1557] = 32'b00000000000000000011001100000010;
assign LUT_1[1558] = 32'b00000000000000000101101000010111;
assign LUT_1[1559] = 32'b11111111111111111110111010010011;
assign LUT_1[1560] = 32'b00000000000000000001001110100100;
assign LUT_1[1561] = 32'b11111111111111111010100000100000;
assign LUT_1[1562] = 32'b11111111111111111100111100110101;
assign LUT_1[1563] = 32'b11111111111111110110001110110001;
assign LUT_1[1564] = 32'b00000000000000001001000111111011;
assign LUT_1[1565] = 32'b00000000000000000010011001110111;
assign LUT_1[1566] = 32'b00000000000000000100110110001100;
assign LUT_1[1567] = 32'b11111111111111111110001000001000;
assign LUT_1[1568] = 32'b00000000000000000001000000001100;
assign LUT_1[1569] = 32'b11111111111111111010010010001000;
assign LUT_1[1570] = 32'b11111111111111111100101110011101;
assign LUT_1[1571] = 32'b11111111111111110110000000011001;
assign LUT_1[1572] = 32'b00000000000000001000111001100011;
assign LUT_1[1573] = 32'b00000000000000000010001011011111;
assign LUT_1[1574] = 32'b00000000000000000100100111110100;
assign LUT_1[1575] = 32'b11111111111111111101111001110000;
assign LUT_1[1576] = 32'b00000000000000000000001110000001;
assign LUT_1[1577] = 32'b11111111111111111001011111111101;
assign LUT_1[1578] = 32'b11111111111111111011111100010010;
assign LUT_1[1579] = 32'b11111111111111110101001110001110;
assign LUT_1[1580] = 32'b00000000000000001000000111011000;
assign LUT_1[1581] = 32'b00000000000000000001011001010100;
assign LUT_1[1582] = 32'b00000000000000000011110101101001;
assign LUT_1[1583] = 32'b11111111111111111101000111100101;
assign LUT_1[1584] = 32'b00000000000000000010111011101110;
assign LUT_1[1585] = 32'b11111111111111111100001101101010;
assign LUT_1[1586] = 32'b11111111111111111110101001111111;
assign LUT_1[1587] = 32'b11111111111111110111111011111011;
assign LUT_1[1588] = 32'b00000000000000001010110101000101;
assign LUT_1[1589] = 32'b00000000000000000100000111000001;
assign LUT_1[1590] = 32'b00000000000000000110100011010110;
assign LUT_1[1591] = 32'b11111111111111111111110101010010;
assign LUT_1[1592] = 32'b00000000000000000010001001100011;
assign LUT_1[1593] = 32'b11111111111111111011011011011111;
assign LUT_1[1594] = 32'b11111111111111111101110111110100;
assign LUT_1[1595] = 32'b11111111111111110111001001110000;
assign LUT_1[1596] = 32'b00000000000000001010000010111010;
assign LUT_1[1597] = 32'b00000000000000000011010100110110;
assign LUT_1[1598] = 32'b00000000000000000101110001001011;
assign LUT_1[1599] = 32'b11111111111111111111000011000111;
assign LUT_1[1600] = 32'b00000000000000000010000010110101;
assign LUT_1[1601] = 32'b11111111111111111011010100110001;
assign LUT_1[1602] = 32'b11111111111111111101110001000110;
assign LUT_1[1603] = 32'b11111111111111110111000011000010;
assign LUT_1[1604] = 32'b00000000000000001001111100001100;
assign LUT_1[1605] = 32'b00000000000000000011001110001000;
assign LUT_1[1606] = 32'b00000000000000000101101010011101;
assign LUT_1[1607] = 32'b11111111111111111110111100011001;
assign LUT_1[1608] = 32'b00000000000000000001010000101010;
assign LUT_1[1609] = 32'b11111111111111111010100010100110;
assign LUT_1[1610] = 32'b11111111111111111100111110111011;
assign LUT_1[1611] = 32'b11111111111111110110010000110111;
assign LUT_1[1612] = 32'b00000000000000001001001010000001;
assign LUT_1[1613] = 32'b00000000000000000010011011111101;
assign LUT_1[1614] = 32'b00000000000000000100111000010010;
assign LUT_1[1615] = 32'b11111111111111111110001010001110;
assign LUT_1[1616] = 32'b00000000000000000011111110010111;
assign LUT_1[1617] = 32'b11111111111111111101010000010011;
assign LUT_1[1618] = 32'b11111111111111111111101100101000;
assign LUT_1[1619] = 32'b11111111111111111000111110100100;
assign LUT_1[1620] = 32'b00000000000000001011110111101110;
assign LUT_1[1621] = 32'b00000000000000000101001001101010;
assign LUT_1[1622] = 32'b00000000000000000111100101111111;
assign LUT_1[1623] = 32'b00000000000000000000110111111011;
assign LUT_1[1624] = 32'b00000000000000000011001100001100;
assign LUT_1[1625] = 32'b11111111111111111100011110001000;
assign LUT_1[1626] = 32'b11111111111111111110111010011101;
assign LUT_1[1627] = 32'b11111111111111111000001100011001;
assign LUT_1[1628] = 32'b00000000000000001011000101100011;
assign LUT_1[1629] = 32'b00000000000000000100010111011111;
assign LUT_1[1630] = 32'b00000000000000000110110011110100;
assign LUT_1[1631] = 32'b00000000000000000000000101110000;
assign LUT_1[1632] = 32'b00000000000000000010111101110100;
assign LUT_1[1633] = 32'b11111111111111111100001111110000;
assign LUT_1[1634] = 32'b11111111111111111110101100000101;
assign LUT_1[1635] = 32'b11111111111111110111111110000001;
assign LUT_1[1636] = 32'b00000000000000001010110111001011;
assign LUT_1[1637] = 32'b00000000000000000100001001000111;
assign LUT_1[1638] = 32'b00000000000000000110100101011100;
assign LUT_1[1639] = 32'b11111111111111111111110111011000;
assign LUT_1[1640] = 32'b00000000000000000010001011101001;
assign LUT_1[1641] = 32'b11111111111111111011011101100101;
assign LUT_1[1642] = 32'b11111111111111111101111001111010;
assign LUT_1[1643] = 32'b11111111111111110111001011110110;
assign LUT_1[1644] = 32'b00000000000000001010000101000000;
assign LUT_1[1645] = 32'b00000000000000000011010110111100;
assign LUT_1[1646] = 32'b00000000000000000101110011010001;
assign LUT_1[1647] = 32'b11111111111111111111000101001101;
assign LUT_1[1648] = 32'b00000000000000000100111001010110;
assign LUT_1[1649] = 32'b11111111111111111110001011010010;
assign LUT_1[1650] = 32'b00000000000000000000100111100111;
assign LUT_1[1651] = 32'b11111111111111111001111001100011;
assign LUT_1[1652] = 32'b00000000000000001100110010101101;
assign LUT_1[1653] = 32'b00000000000000000110000100101001;
assign LUT_1[1654] = 32'b00000000000000001000100000111110;
assign LUT_1[1655] = 32'b00000000000000000001110010111010;
assign LUT_1[1656] = 32'b00000000000000000100000111001011;
assign LUT_1[1657] = 32'b11111111111111111101011001000111;
assign LUT_1[1658] = 32'b11111111111111111111110101011100;
assign LUT_1[1659] = 32'b11111111111111111001000111011000;
assign LUT_1[1660] = 32'b00000000000000001100000000100010;
assign LUT_1[1661] = 32'b00000000000000000101010010011110;
assign LUT_1[1662] = 32'b00000000000000000111101110110011;
assign LUT_1[1663] = 32'b00000000000000000001000000101111;
assign LUT_1[1664] = 32'b00000000000000000011000101010000;
assign LUT_1[1665] = 32'b11111111111111111100010111001100;
assign LUT_1[1666] = 32'b11111111111111111110110011100001;
assign LUT_1[1667] = 32'b11111111111111111000000101011101;
assign LUT_1[1668] = 32'b00000000000000001010111110100111;
assign LUT_1[1669] = 32'b00000000000000000100010000100011;
assign LUT_1[1670] = 32'b00000000000000000110101100111000;
assign LUT_1[1671] = 32'b11111111111111111111111110110100;
assign LUT_1[1672] = 32'b00000000000000000010010011000101;
assign LUT_1[1673] = 32'b11111111111111111011100101000001;
assign LUT_1[1674] = 32'b11111111111111111110000001010110;
assign LUT_1[1675] = 32'b11111111111111110111010011010010;
assign LUT_1[1676] = 32'b00000000000000001010001100011100;
assign LUT_1[1677] = 32'b00000000000000000011011110011000;
assign LUT_1[1678] = 32'b00000000000000000101111010101101;
assign LUT_1[1679] = 32'b11111111111111111111001100101001;
assign LUT_1[1680] = 32'b00000000000000000101000000110010;
assign LUT_1[1681] = 32'b11111111111111111110010010101110;
assign LUT_1[1682] = 32'b00000000000000000000101111000011;
assign LUT_1[1683] = 32'b11111111111111111010000000111111;
assign LUT_1[1684] = 32'b00000000000000001100111010001001;
assign LUT_1[1685] = 32'b00000000000000000110001100000101;
assign LUT_1[1686] = 32'b00000000000000001000101000011010;
assign LUT_1[1687] = 32'b00000000000000000001111010010110;
assign LUT_1[1688] = 32'b00000000000000000100001110100111;
assign LUT_1[1689] = 32'b11111111111111111101100000100011;
assign LUT_1[1690] = 32'b11111111111111111111111100111000;
assign LUT_1[1691] = 32'b11111111111111111001001110110100;
assign LUT_1[1692] = 32'b00000000000000001100000111111110;
assign LUT_1[1693] = 32'b00000000000000000101011001111010;
assign LUT_1[1694] = 32'b00000000000000000111110110001111;
assign LUT_1[1695] = 32'b00000000000000000001001000001011;
assign LUT_1[1696] = 32'b00000000000000000100000000001111;
assign LUT_1[1697] = 32'b11111111111111111101010010001011;
assign LUT_1[1698] = 32'b11111111111111111111101110100000;
assign LUT_1[1699] = 32'b11111111111111111001000000011100;
assign LUT_1[1700] = 32'b00000000000000001011111001100110;
assign LUT_1[1701] = 32'b00000000000000000101001011100010;
assign LUT_1[1702] = 32'b00000000000000000111100111110111;
assign LUT_1[1703] = 32'b00000000000000000000111001110011;
assign LUT_1[1704] = 32'b00000000000000000011001110000100;
assign LUT_1[1705] = 32'b11111111111111111100100000000000;
assign LUT_1[1706] = 32'b11111111111111111110111100010101;
assign LUT_1[1707] = 32'b11111111111111111000001110010001;
assign LUT_1[1708] = 32'b00000000000000001011000111011011;
assign LUT_1[1709] = 32'b00000000000000000100011001010111;
assign LUT_1[1710] = 32'b00000000000000000110110101101100;
assign LUT_1[1711] = 32'b00000000000000000000000111101000;
assign LUT_1[1712] = 32'b00000000000000000101111011110001;
assign LUT_1[1713] = 32'b11111111111111111111001101101101;
assign LUT_1[1714] = 32'b00000000000000000001101010000010;
assign LUT_1[1715] = 32'b11111111111111111010111011111110;
assign LUT_1[1716] = 32'b00000000000000001101110101001000;
assign LUT_1[1717] = 32'b00000000000000000111000111000100;
assign LUT_1[1718] = 32'b00000000000000001001100011011001;
assign LUT_1[1719] = 32'b00000000000000000010110101010101;
assign LUT_1[1720] = 32'b00000000000000000101001001100110;
assign LUT_1[1721] = 32'b11111111111111111110011011100010;
assign LUT_1[1722] = 32'b00000000000000000000110111110111;
assign LUT_1[1723] = 32'b11111111111111111010001001110011;
assign LUT_1[1724] = 32'b00000000000000001101000010111101;
assign LUT_1[1725] = 32'b00000000000000000110010100111001;
assign LUT_1[1726] = 32'b00000000000000001000110001001110;
assign LUT_1[1727] = 32'b00000000000000000010000011001010;
assign LUT_1[1728] = 32'b00000000000000000101000010111000;
assign LUT_1[1729] = 32'b11111111111111111110010100110100;
assign LUT_1[1730] = 32'b00000000000000000000110001001001;
assign LUT_1[1731] = 32'b11111111111111111010000011000101;
assign LUT_1[1732] = 32'b00000000000000001100111100001111;
assign LUT_1[1733] = 32'b00000000000000000110001110001011;
assign LUT_1[1734] = 32'b00000000000000001000101010100000;
assign LUT_1[1735] = 32'b00000000000000000001111100011100;
assign LUT_1[1736] = 32'b00000000000000000100010000101101;
assign LUT_1[1737] = 32'b11111111111111111101100010101001;
assign LUT_1[1738] = 32'b11111111111111111111111110111110;
assign LUT_1[1739] = 32'b11111111111111111001010000111010;
assign LUT_1[1740] = 32'b00000000000000001100001010000100;
assign LUT_1[1741] = 32'b00000000000000000101011100000000;
assign LUT_1[1742] = 32'b00000000000000000111111000010101;
assign LUT_1[1743] = 32'b00000000000000000001001010010001;
assign LUT_1[1744] = 32'b00000000000000000110111110011010;
assign LUT_1[1745] = 32'b00000000000000000000010000010110;
assign LUT_1[1746] = 32'b00000000000000000010101100101011;
assign LUT_1[1747] = 32'b11111111111111111011111110100111;
assign LUT_1[1748] = 32'b00000000000000001110110111110001;
assign LUT_1[1749] = 32'b00000000000000001000001001101101;
assign LUT_1[1750] = 32'b00000000000000001010100110000010;
assign LUT_1[1751] = 32'b00000000000000000011110111111110;
assign LUT_1[1752] = 32'b00000000000000000110001100001111;
assign LUT_1[1753] = 32'b11111111111111111111011110001011;
assign LUT_1[1754] = 32'b00000000000000000001111010100000;
assign LUT_1[1755] = 32'b11111111111111111011001100011100;
assign LUT_1[1756] = 32'b00000000000000001110000101100110;
assign LUT_1[1757] = 32'b00000000000000000111010111100010;
assign LUT_1[1758] = 32'b00000000000000001001110011110111;
assign LUT_1[1759] = 32'b00000000000000000011000101110011;
assign LUT_1[1760] = 32'b00000000000000000101111101110111;
assign LUT_1[1761] = 32'b11111111111111111111001111110011;
assign LUT_1[1762] = 32'b00000000000000000001101100001000;
assign LUT_1[1763] = 32'b11111111111111111010111110000100;
assign LUT_1[1764] = 32'b00000000000000001101110111001110;
assign LUT_1[1765] = 32'b00000000000000000111001001001010;
assign LUT_1[1766] = 32'b00000000000000001001100101011111;
assign LUT_1[1767] = 32'b00000000000000000010110111011011;
assign LUT_1[1768] = 32'b00000000000000000101001011101100;
assign LUT_1[1769] = 32'b11111111111111111110011101101000;
assign LUT_1[1770] = 32'b00000000000000000000111001111101;
assign LUT_1[1771] = 32'b11111111111111111010001011111001;
assign LUT_1[1772] = 32'b00000000000000001101000101000011;
assign LUT_1[1773] = 32'b00000000000000000110010110111111;
assign LUT_1[1774] = 32'b00000000000000001000110011010100;
assign LUT_1[1775] = 32'b00000000000000000010000101010000;
assign LUT_1[1776] = 32'b00000000000000000111111001011001;
assign LUT_1[1777] = 32'b00000000000000000001001011010101;
assign LUT_1[1778] = 32'b00000000000000000011100111101010;
assign LUT_1[1779] = 32'b11111111111111111100111001100110;
assign LUT_1[1780] = 32'b00000000000000001111110010110000;
assign LUT_1[1781] = 32'b00000000000000001001000100101100;
assign LUT_1[1782] = 32'b00000000000000001011100001000001;
assign LUT_1[1783] = 32'b00000000000000000100110010111101;
assign LUT_1[1784] = 32'b00000000000000000111000111001110;
assign LUT_1[1785] = 32'b00000000000000000000011001001010;
assign LUT_1[1786] = 32'b00000000000000000010110101011111;
assign LUT_1[1787] = 32'b11111111111111111100000111011011;
assign LUT_1[1788] = 32'b00000000000000001111000000100101;
assign LUT_1[1789] = 32'b00000000000000001000010010100001;
assign LUT_1[1790] = 32'b00000000000000001010101110110110;
assign LUT_1[1791] = 32'b00000000000000000100000000110010;
assign LUT_1[1792] = 32'b11111111111111111101111001011001;
assign LUT_1[1793] = 32'b11111111111111110111001011010101;
assign LUT_1[1794] = 32'b11111111111111111001100111101010;
assign LUT_1[1795] = 32'b11111111111111110010111001100110;
assign LUT_1[1796] = 32'b00000000000000000101110010110000;
assign LUT_1[1797] = 32'b11111111111111111111000100101100;
assign LUT_1[1798] = 32'b00000000000000000001100001000001;
assign LUT_1[1799] = 32'b11111111111111111010110010111101;
assign LUT_1[1800] = 32'b11111111111111111101000111001110;
assign LUT_1[1801] = 32'b11111111111111110110011001001010;
assign LUT_1[1802] = 32'b11111111111111111000110101011111;
assign LUT_1[1803] = 32'b11111111111111110010000111011011;
assign LUT_1[1804] = 32'b00000000000000000101000000100101;
assign LUT_1[1805] = 32'b11111111111111111110010010100001;
assign LUT_1[1806] = 32'b00000000000000000000101110110110;
assign LUT_1[1807] = 32'b11111111111111111010000000110010;
assign LUT_1[1808] = 32'b11111111111111111111110100111011;
assign LUT_1[1809] = 32'b11111111111111111001000110110111;
assign LUT_1[1810] = 32'b11111111111111111011100011001100;
assign LUT_1[1811] = 32'b11111111111111110100110101001000;
assign LUT_1[1812] = 32'b00000000000000000111101110010010;
assign LUT_1[1813] = 32'b00000000000000000001000000001110;
assign LUT_1[1814] = 32'b00000000000000000011011100100011;
assign LUT_1[1815] = 32'b11111111111111111100101110011111;
assign LUT_1[1816] = 32'b11111111111111111111000010110000;
assign LUT_1[1817] = 32'b11111111111111111000010100101100;
assign LUT_1[1818] = 32'b11111111111111111010110001000001;
assign LUT_1[1819] = 32'b11111111111111110100000010111101;
assign LUT_1[1820] = 32'b00000000000000000110111100000111;
assign LUT_1[1821] = 32'b00000000000000000000001110000011;
assign LUT_1[1822] = 32'b00000000000000000010101010011000;
assign LUT_1[1823] = 32'b11111111111111111011111100010100;
assign LUT_1[1824] = 32'b11111111111111111110110100011000;
assign LUT_1[1825] = 32'b11111111111111111000000110010100;
assign LUT_1[1826] = 32'b11111111111111111010100010101001;
assign LUT_1[1827] = 32'b11111111111111110011110100100101;
assign LUT_1[1828] = 32'b00000000000000000110101101101111;
assign LUT_1[1829] = 32'b11111111111111111111111111101011;
assign LUT_1[1830] = 32'b00000000000000000010011100000000;
assign LUT_1[1831] = 32'b11111111111111111011101101111100;
assign LUT_1[1832] = 32'b11111111111111111110000010001101;
assign LUT_1[1833] = 32'b11111111111111110111010100001001;
assign LUT_1[1834] = 32'b11111111111111111001110000011110;
assign LUT_1[1835] = 32'b11111111111111110011000010011010;
assign LUT_1[1836] = 32'b00000000000000000101111011100100;
assign LUT_1[1837] = 32'b11111111111111111111001101100000;
assign LUT_1[1838] = 32'b00000000000000000001101001110101;
assign LUT_1[1839] = 32'b11111111111111111010111011110001;
assign LUT_1[1840] = 32'b00000000000000000000101111111010;
assign LUT_1[1841] = 32'b11111111111111111010000001110110;
assign LUT_1[1842] = 32'b11111111111111111100011110001011;
assign LUT_1[1843] = 32'b11111111111111110101110000000111;
assign LUT_1[1844] = 32'b00000000000000001000101001010001;
assign LUT_1[1845] = 32'b00000000000000000001111011001101;
assign LUT_1[1846] = 32'b00000000000000000100010111100010;
assign LUT_1[1847] = 32'b11111111111111111101101001011110;
assign LUT_1[1848] = 32'b11111111111111111111111101101111;
assign LUT_1[1849] = 32'b11111111111111111001001111101011;
assign LUT_1[1850] = 32'b11111111111111111011101100000000;
assign LUT_1[1851] = 32'b11111111111111110100111101111100;
assign LUT_1[1852] = 32'b00000000000000000111110111000110;
assign LUT_1[1853] = 32'b00000000000000000001001001000010;
assign LUT_1[1854] = 32'b00000000000000000011100101010111;
assign LUT_1[1855] = 32'b11111111111111111100110111010011;
assign LUT_1[1856] = 32'b11111111111111111111110111000001;
assign LUT_1[1857] = 32'b11111111111111111001001000111101;
assign LUT_1[1858] = 32'b11111111111111111011100101010010;
assign LUT_1[1859] = 32'b11111111111111110100110111001110;
assign LUT_1[1860] = 32'b00000000000000000111110000011000;
assign LUT_1[1861] = 32'b00000000000000000001000010010100;
assign LUT_1[1862] = 32'b00000000000000000011011110101001;
assign LUT_1[1863] = 32'b11111111111111111100110000100101;
assign LUT_1[1864] = 32'b11111111111111111111000100110110;
assign LUT_1[1865] = 32'b11111111111111111000010110110010;
assign LUT_1[1866] = 32'b11111111111111111010110011000111;
assign LUT_1[1867] = 32'b11111111111111110100000101000011;
assign LUT_1[1868] = 32'b00000000000000000110111110001101;
assign LUT_1[1869] = 32'b00000000000000000000010000001001;
assign LUT_1[1870] = 32'b00000000000000000010101100011110;
assign LUT_1[1871] = 32'b11111111111111111011111110011010;
assign LUT_1[1872] = 32'b00000000000000000001110010100011;
assign LUT_1[1873] = 32'b11111111111111111011000100011111;
assign LUT_1[1874] = 32'b11111111111111111101100000110100;
assign LUT_1[1875] = 32'b11111111111111110110110010110000;
assign LUT_1[1876] = 32'b00000000000000001001101011111010;
assign LUT_1[1877] = 32'b00000000000000000010111101110110;
assign LUT_1[1878] = 32'b00000000000000000101011010001011;
assign LUT_1[1879] = 32'b11111111111111111110101100000111;
assign LUT_1[1880] = 32'b00000000000000000001000000011000;
assign LUT_1[1881] = 32'b11111111111111111010010010010100;
assign LUT_1[1882] = 32'b11111111111111111100101110101001;
assign LUT_1[1883] = 32'b11111111111111110110000000100101;
assign LUT_1[1884] = 32'b00000000000000001000111001101111;
assign LUT_1[1885] = 32'b00000000000000000010001011101011;
assign LUT_1[1886] = 32'b00000000000000000100101000000000;
assign LUT_1[1887] = 32'b11111111111111111101111001111100;
assign LUT_1[1888] = 32'b00000000000000000000110010000000;
assign LUT_1[1889] = 32'b11111111111111111010000011111100;
assign LUT_1[1890] = 32'b11111111111111111100100000010001;
assign LUT_1[1891] = 32'b11111111111111110101110010001101;
assign LUT_1[1892] = 32'b00000000000000001000101011010111;
assign LUT_1[1893] = 32'b00000000000000000001111101010011;
assign LUT_1[1894] = 32'b00000000000000000100011001101000;
assign LUT_1[1895] = 32'b11111111111111111101101011100100;
assign LUT_1[1896] = 32'b11111111111111111111111111110101;
assign LUT_1[1897] = 32'b11111111111111111001010001110001;
assign LUT_1[1898] = 32'b11111111111111111011101110000110;
assign LUT_1[1899] = 32'b11111111111111110101000000000010;
assign LUT_1[1900] = 32'b00000000000000000111111001001100;
assign LUT_1[1901] = 32'b00000000000000000001001011001000;
assign LUT_1[1902] = 32'b00000000000000000011100111011101;
assign LUT_1[1903] = 32'b11111111111111111100111001011001;
assign LUT_1[1904] = 32'b00000000000000000010101101100010;
assign LUT_1[1905] = 32'b11111111111111111011111111011110;
assign LUT_1[1906] = 32'b11111111111111111110011011110011;
assign LUT_1[1907] = 32'b11111111111111110111101101101111;
assign LUT_1[1908] = 32'b00000000000000001010100110111001;
assign LUT_1[1909] = 32'b00000000000000000011111000110101;
assign LUT_1[1910] = 32'b00000000000000000110010101001010;
assign LUT_1[1911] = 32'b11111111111111111111100111000110;
assign LUT_1[1912] = 32'b00000000000000000001111011010111;
assign LUT_1[1913] = 32'b11111111111111111011001101010011;
assign LUT_1[1914] = 32'b11111111111111111101101001101000;
assign LUT_1[1915] = 32'b11111111111111110110111011100100;
assign LUT_1[1916] = 32'b00000000000000001001110100101110;
assign LUT_1[1917] = 32'b00000000000000000011000110101010;
assign LUT_1[1918] = 32'b00000000000000000101100010111111;
assign LUT_1[1919] = 32'b11111111111111111110110100111011;
assign LUT_1[1920] = 32'b00000000000000000000111001011100;
assign LUT_1[1921] = 32'b11111111111111111010001011011000;
assign LUT_1[1922] = 32'b11111111111111111100100111101101;
assign LUT_1[1923] = 32'b11111111111111110101111001101001;
assign LUT_1[1924] = 32'b00000000000000001000110010110011;
assign LUT_1[1925] = 32'b00000000000000000010000100101111;
assign LUT_1[1926] = 32'b00000000000000000100100001000100;
assign LUT_1[1927] = 32'b11111111111111111101110011000000;
assign LUT_1[1928] = 32'b00000000000000000000000111010001;
assign LUT_1[1929] = 32'b11111111111111111001011001001101;
assign LUT_1[1930] = 32'b11111111111111111011110101100010;
assign LUT_1[1931] = 32'b11111111111111110101000111011110;
assign LUT_1[1932] = 32'b00000000000000001000000000101000;
assign LUT_1[1933] = 32'b00000000000000000001010010100100;
assign LUT_1[1934] = 32'b00000000000000000011101110111001;
assign LUT_1[1935] = 32'b11111111111111111101000000110101;
assign LUT_1[1936] = 32'b00000000000000000010110100111110;
assign LUT_1[1937] = 32'b11111111111111111100000110111010;
assign LUT_1[1938] = 32'b11111111111111111110100011001111;
assign LUT_1[1939] = 32'b11111111111111110111110101001011;
assign LUT_1[1940] = 32'b00000000000000001010101110010101;
assign LUT_1[1941] = 32'b00000000000000000100000000010001;
assign LUT_1[1942] = 32'b00000000000000000110011100100110;
assign LUT_1[1943] = 32'b11111111111111111111101110100010;
assign LUT_1[1944] = 32'b00000000000000000010000010110011;
assign LUT_1[1945] = 32'b11111111111111111011010100101111;
assign LUT_1[1946] = 32'b11111111111111111101110001000100;
assign LUT_1[1947] = 32'b11111111111111110111000011000000;
assign LUT_1[1948] = 32'b00000000000000001001111100001010;
assign LUT_1[1949] = 32'b00000000000000000011001110000110;
assign LUT_1[1950] = 32'b00000000000000000101101010011011;
assign LUT_1[1951] = 32'b11111111111111111110111100010111;
assign LUT_1[1952] = 32'b00000000000000000001110100011011;
assign LUT_1[1953] = 32'b11111111111111111011000110010111;
assign LUT_1[1954] = 32'b11111111111111111101100010101100;
assign LUT_1[1955] = 32'b11111111111111110110110100101000;
assign LUT_1[1956] = 32'b00000000000000001001101101110010;
assign LUT_1[1957] = 32'b00000000000000000010111111101110;
assign LUT_1[1958] = 32'b00000000000000000101011100000011;
assign LUT_1[1959] = 32'b11111111111111111110101101111111;
assign LUT_1[1960] = 32'b00000000000000000001000010010000;
assign LUT_1[1961] = 32'b11111111111111111010010100001100;
assign LUT_1[1962] = 32'b11111111111111111100110000100001;
assign LUT_1[1963] = 32'b11111111111111110110000010011101;
assign LUT_1[1964] = 32'b00000000000000001000111011100111;
assign LUT_1[1965] = 32'b00000000000000000010001101100011;
assign LUT_1[1966] = 32'b00000000000000000100101001111000;
assign LUT_1[1967] = 32'b11111111111111111101111011110100;
assign LUT_1[1968] = 32'b00000000000000000011101111111101;
assign LUT_1[1969] = 32'b11111111111111111101000001111001;
assign LUT_1[1970] = 32'b11111111111111111111011110001110;
assign LUT_1[1971] = 32'b11111111111111111000110000001010;
assign LUT_1[1972] = 32'b00000000000000001011101001010100;
assign LUT_1[1973] = 32'b00000000000000000100111011010000;
assign LUT_1[1974] = 32'b00000000000000000111010111100101;
assign LUT_1[1975] = 32'b00000000000000000000101001100001;
assign LUT_1[1976] = 32'b00000000000000000010111101110010;
assign LUT_1[1977] = 32'b11111111111111111100001111101110;
assign LUT_1[1978] = 32'b11111111111111111110101100000011;
assign LUT_1[1979] = 32'b11111111111111110111111101111111;
assign LUT_1[1980] = 32'b00000000000000001010110111001001;
assign LUT_1[1981] = 32'b00000000000000000100001001000101;
assign LUT_1[1982] = 32'b00000000000000000110100101011010;
assign LUT_1[1983] = 32'b11111111111111111111110111010110;
assign LUT_1[1984] = 32'b00000000000000000010110111000100;
assign LUT_1[1985] = 32'b11111111111111111100001001000000;
assign LUT_1[1986] = 32'b11111111111111111110100101010101;
assign LUT_1[1987] = 32'b11111111111111110111110111010001;
assign LUT_1[1988] = 32'b00000000000000001010110000011011;
assign LUT_1[1989] = 32'b00000000000000000100000010010111;
assign LUT_1[1990] = 32'b00000000000000000110011110101100;
assign LUT_1[1991] = 32'b11111111111111111111110000101000;
assign LUT_1[1992] = 32'b00000000000000000010000100111001;
assign LUT_1[1993] = 32'b11111111111111111011010110110101;
assign LUT_1[1994] = 32'b11111111111111111101110011001010;
assign LUT_1[1995] = 32'b11111111111111110111000101000110;
assign LUT_1[1996] = 32'b00000000000000001001111110010000;
assign LUT_1[1997] = 32'b00000000000000000011010000001100;
assign LUT_1[1998] = 32'b00000000000000000101101100100001;
assign LUT_1[1999] = 32'b11111111111111111110111110011101;
assign LUT_1[2000] = 32'b00000000000000000100110010100110;
assign LUT_1[2001] = 32'b11111111111111111110000100100010;
assign LUT_1[2002] = 32'b00000000000000000000100000110111;
assign LUT_1[2003] = 32'b11111111111111111001110010110011;
assign LUT_1[2004] = 32'b00000000000000001100101011111101;
assign LUT_1[2005] = 32'b00000000000000000101111101111001;
assign LUT_1[2006] = 32'b00000000000000001000011010001110;
assign LUT_1[2007] = 32'b00000000000000000001101100001010;
assign LUT_1[2008] = 32'b00000000000000000100000000011011;
assign LUT_1[2009] = 32'b11111111111111111101010010010111;
assign LUT_1[2010] = 32'b11111111111111111111101110101100;
assign LUT_1[2011] = 32'b11111111111111111001000000101000;
assign LUT_1[2012] = 32'b00000000000000001011111001110010;
assign LUT_1[2013] = 32'b00000000000000000101001011101110;
assign LUT_1[2014] = 32'b00000000000000000111101000000011;
assign LUT_1[2015] = 32'b00000000000000000000111001111111;
assign LUT_1[2016] = 32'b00000000000000000011110010000011;
assign LUT_1[2017] = 32'b11111111111111111101000011111111;
assign LUT_1[2018] = 32'b11111111111111111111100000010100;
assign LUT_1[2019] = 32'b11111111111111111000110010010000;
assign LUT_1[2020] = 32'b00000000000000001011101011011010;
assign LUT_1[2021] = 32'b00000000000000000100111101010110;
assign LUT_1[2022] = 32'b00000000000000000111011001101011;
assign LUT_1[2023] = 32'b00000000000000000000101011100111;
assign LUT_1[2024] = 32'b00000000000000000010111111111000;
assign LUT_1[2025] = 32'b11111111111111111100010001110100;
assign LUT_1[2026] = 32'b11111111111111111110101110001001;
assign LUT_1[2027] = 32'b11111111111111111000000000000101;
assign LUT_1[2028] = 32'b00000000000000001010111001001111;
assign LUT_1[2029] = 32'b00000000000000000100001011001011;
assign LUT_1[2030] = 32'b00000000000000000110100111100000;
assign LUT_1[2031] = 32'b11111111111111111111111001011100;
assign LUT_1[2032] = 32'b00000000000000000101101101100101;
assign LUT_1[2033] = 32'b11111111111111111110111111100001;
assign LUT_1[2034] = 32'b00000000000000000001011011110110;
assign LUT_1[2035] = 32'b11111111111111111010101101110010;
assign LUT_1[2036] = 32'b00000000000000001101100110111100;
assign LUT_1[2037] = 32'b00000000000000000110111000111000;
assign LUT_1[2038] = 32'b00000000000000001001010101001101;
assign LUT_1[2039] = 32'b00000000000000000010100111001001;
assign LUT_1[2040] = 32'b00000000000000000100111011011010;
assign LUT_1[2041] = 32'b11111111111111111110001101010110;
assign LUT_1[2042] = 32'b00000000000000000000101001101011;
assign LUT_1[2043] = 32'b11111111111111111001111011100111;
assign LUT_1[2044] = 32'b00000000000000001100110100110001;
assign LUT_1[2045] = 32'b00000000000000000110000110101101;
assign LUT_1[2046] = 32'b00000000000000001000100011000010;
assign LUT_1[2047] = 32'b00000000000000000001110100111110;
assign LUT_1[2048] = 32'b00000000000000000001000001111011;
assign LUT_1[2049] = 32'b11111111111111111010010011110111;
assign LUT_1[2050] = 32'b11111111111111111100110000001100;
assign LUT_1[2051] = 32'b11111111111111110110000010001000;
assign LUT_1[2052] = 32'b00000000000000001000111011010010;
assign LUT_1[2053] = 32'b00000000000000000010001101001110;
assign LUT_1[2054] = 32'b00000000000000000100101001100011;
assign LUT_1[2055] = 32'b11111111111111111101111011011111;
assign LUT_1[2056] = 32'b00000000000000000000001111110000;
assign LUT_1[2057] = 32'b11111111111111111001100001101100;
assign LUT_1[2058] = 32'b11111111111111111011111110000001;
assign LUT_1[2059] = 32'b11111111111111110101001111111101;
assign LUT_1[2060] = 32'b00000000000000001000001001000111;
assign LUT_1[2061] = 32'b00000000000000000001011011000011;
assign LUT_1[2062] = 32'b00000000000000000011110111011000;
assign LUT_1[2063] = 32'b11111111111111111101001001010100;
assign LUT_1[2064] = 32'b00000000000000000010111101011101;
assign LUT_1[2065] = 32'b11111111111111111100001111011001;
assign LUT_1[2066] = 32'b11111111111111111110101011101110;
assign LUT_1[2067] = 32'b11111111111111110111111101101010;
assign LUT_1[2068] = 32'b00000000000000001010110110110100;
assign LUT_1[2069] = 32'b00000000000000000100001000110000;
assign LUT_1[2070] = 32'b00000000000000000110100101000101;
assign LUT_1[2071] = 32'b11111111111111111111110111000001;
assign LUT_1[2072] = 32'b00000000000000000010001011010010;
assign LUT_1[2073] = 32'b11111111111111111011011101001110;
assign LUT_1[2074] = 32'b11111111111111111101111001100011;
assign LUT_1[2075] = 32'b11111111111111110111001011011111;
assign LUT_1[2076] = 32'b00000000000000001010000100101001;
assign LUT_1[2077] = 32'b00000000000000000011010110100101;
assign LUT_1[2078] = 32'b00000000000000000101110010111010;
assign LUT_1[2079] = 32'b11111111111111111111000100110110;
assign LUT_1[2080] = 32'b00000000000000000001111100111010;
assign LUT_1[2081] = 32'b11111111111111111011001110110110;
assign LUT_1[2082] = 32'b11111111111111111101101011001011;
assign LUT_1[2083] = 32'b11111111111111110110111101000111;
assign LUT_1[2084] = 32'b00000000000000001001110110010001;
assign LUT_1[2085] = 32'b00000000000000000011001000001101;
assign LUT_1[2086] = 32'b00000000000000000101100100100010;
assign LUT_1[2087] = 32'b11111111111111111110110110011110;
assign LUT_1[2088] = 32'b00000000000000000001001010101111;
assign LUT_1[2089] = 32'b11111111111111111010011100101011;
assign LUT_1[2090] = 32'b11111111111111111100111001000000;
assign LUT_1[2091] = 32'b11111111111111110110001010111100;
assign LUT_1[2092] = 32'b00000000000000001001000100000110;
assign LUT_1[2093] = 32'b00000000000000000010010110000010;
assign LUT_1[2094] = 32'b00000000000000000100110010010111;
assign LUT_1[2095] = 32'b11111111111111111110000100010011;
assign LUT_1[2096] = 32'b00000000000000000011111000011100;
assign LUT_1[2097] = 32'b11111111111111111101001010011000;
assign LUT_1[2098] = 32'b11111111111111111111100110101101;
assign LUT_1[2099] = 32'b11111111111111111000111000101001;
assign LUT_1[2100] = 32'b00000000000000001011110001110011;
assign LUT_1[2101] = 32'b00000000000000000101000011101111;
assign LUT_1[2102] = 32'b00000000000000000111100000000100;
assign LUT_1[2103] = 32'b00000000000000000000110010000000;
assign LUT_1[2104] = 32'b00000000000000000011000110010001;
assign LUT_1[2105] = 32'b11111111111111111100011000001101;
assign LUT_1[2106] = 32'b11111111111111111110110100100010;
assign LUT_1[2107] = 32'b11111111111111111000000110011110;
assign LUT_1[2108] = 32'b00000000000000001010111111101000;
assign LUT_1[2109] = 32'b00000000000000000100010001100100;
assign LUT_1[2110] = 32'b00000000000000000110101101111001;
assign LUT_1[2111] = 32'b11111111111111111111111111110101;
assign LUT_1[2112] = 32'b00000000000000000010111111100011;
assign LUT_1[2113] = 32'b11111111111111111100010001011111;
assign LUT_1[2114] = 32'b11111111111111111110101101110100;
assign LUT_1[2115] = 32'b11111111111111110111111111110000;
assign LUT_1[2116] = 32'b00000000000000001010111000111010;
assign LUT_1[2117] = 32'b00000000000000000100001010110110;
assign LUT_1[2118] = 32'b00000000000000000110100111001011;
assign LUT_1[2119] = 32'b11111111111111111111111001000111;
assign LUT_1[2120] = 32'b00000000000000000010001101011000;
assign LUT_1[2121] = 32'b11111111111111111011011111010100;
assign LUT_1[2122] = 32'b11111111111111111101111011101001;
assign LUT_1[2123] = 32'b11111111111111110111001101100101;
assign LUT_1[2124] = 32'b00000000000000001010000110101111;
assign LUT_1[2125] = 32'b00000000000000000011011000101011;
assign LUT_1[2126] = 32'b00000000000000000101110101000000;
assign LUT_1[2127] = 32'b11111111111111111111000110111100;
assign LUT_1[2128] = 32'b00000000000000000100111011000101;
assign LUT_1[2129] = 32'b11111111111111111110001101000001;
assign LUT_1[2130] = 32'b00000000000000000000101001010110;
assign LUT_1[2131] = 32'b11111111111111111001111011010010;
assign LUT_1[2132] = 32'b00000000000000001100110100011100;
assign LUT_1[2133] = 32'b00000000000000000110000110011000;
assign LUT_1[2134] = 32'b00000000000000001000100010101101;
assign LUT_1[2135] = 32'b00000000000000000001110100101001;
assign LUT_1[2136] = 32'b00000000000000000100001000111010;
assign LUT_1[2137] = 32'b11111111111111111101011010110110;
assign LUT_1[2138] = 32'b11111111111111111111110111001011;
assign LUT_1[2139] = 32'b11111111111111111001001001000111;
assign LUT_1[2140] = 32'b00000000000000001100000010010001;
assign LUT_1[2141] = 32'b00000000000000000101010100001101;
assign LUT_1[2142] = 32'b00000000000000000111110000100010;
assign LUT_1[2143] = 32'b00000000000000000001000010011110;
assign LUT_1[2144] = 32'b00000000000000000011111010100010;
assign LUT_1[2145] = 32'b11111111111111111101001100011110;
assign LUT_1[2146] = 32'b11111111111111111111101000110011;
assign LUT_1[2147] = 32'b11111111111111111000111010101111;
assign LUT_1[2148] = 32'b00000000000000001011110011111001;
assign LUT_1[2149] = 32'b00000000000000000101000101110101;
assign LUT_1[2150] = 32'b00000000000000000111100010001010;
assign LUT_1[2151] = 32'b00000000000000000000110100000110;
assign LUT_1[2152] = 32'b00000000000000000011001000010111;
assign LUT_1[2153] = 32'b11111111111111111100011010010011;
assign LUT_1[2154] = 32'b11111111111111111110110110101000;
assign LUT_1[2155] = 32'b11111111111111111000001000100100;
assign LUT_1[2156] = 32'b00000000000000001011000001101110;
assign LUT_1[2157] = 32'b00000000000000000100010011101010;
assign LUT_1[2158] = 32'b00000000000000000110101111111111;
assign LUT_1[2159] = 32'b00000000000000000000000001111011;
assign LUT_1[2160] = 32'b00000000000000000101110110000100;
assign LUT_1[2161] = 32'b11111111111111111111001000000000;
assign LUT_1[2162] = 32'b00000000000000000001100100010101;
assign LUT_1[2163] = 32'b11111111111111111010110110010001;
assign LUT_1[2164] = 32'b00000000000000001101101111011011;
assign LUT_1[2165] = 32'b00000000000000000111000001010111;
assign LUT_1[2166] = 32'b00000000000000001001011101101100;
assign LUT_1[2167] = 32'b00000000000000000010101111101000;
assign LUT_1[2168] = 32'b00000000000000000101000011111001;
assign LUT_1[2169] = 32'b11111111111111111110010101110101;
assign LUT_1[2170] = 32'b00000000000000000000110010001010;
assign LUT_1[2171] = 32'b11111111111111111010000100000110;
assign LUT_1[2172] = 32'b00000000000000001100111101010000;
assign LUT_1[2173] = 32'b00000000000000000110001111001100;
assign LUT_1[2174] = 32'b00000000000000001000101011100001;
assign LUT_1[2175] = 32'b00000000000000000001111101011101;
assign LUT_1[2176] = 32'b00000000000000000100000001111110;
assign LUT_1[2177] = 32'b11111111111111111101010011111010;
assign LUT_1[2178] = 32'b11111111111111111111110000001111;
assign LUT_1[2179] = 32'b11111111111111111001000010001011;
assign LUT_1[2180] = 32'b00000000000000001011111011010101;
assign LUT_1[2181] = 32'b00000000000000000101001101010001;
assign LUT_1[2182] = 32'b00000000000000000111101001100110;
assign LUT_1[2183] = 32'b00000000000000000000111011100010;
assign LUT_1[2184] = 32'b00000000000000000011001111110011;
assign LUT_1[2185] = 32'b11111111111111111100100001101111;
assign LUT_1[2186] = 32'b11111111111111111110111110000100;
assign LUT_1[2187] = 32'b11111111111111111000010000000000;
assign LUT_1[2188] = 32'b00000000000000001011001001001010;
assign LUT_1[2189] = 32'b00000000000000000100011011000110;
assign LUT_1[2190] = 32'b00000000000000000110110111011011;
assign LUT_1[2191] = 32'b00000000000000000000001001010111;
assign LUT_1[2192] = 32'b00000000000000000101111101100000;
assign LUT_1[2193] = 32'b11111111111111111111001111011100;
assign LUT_1[2194] = 32'b00000000000000000001101011110001;
assign LUT_1[2195] = 32'b11111111111111111010111101101101;
assign LUT_1[2196] = 32'b00000000000000001101110110110111;
assign LUT_1[2197] = 32'b00000000000000000111001000110011;
assign LUT_1[2198] = 32'b00000000000000001001100101001000;
assign LUT_1[2199] = 32'b00000000000000000010110111000100;
assign LUT_1[2200] = 32'b00000000000000000101001011010101;
assign LUT_1[2201] = 32'b11111111111111111110011101010001;
assign LUT_1[2202] = 32'b00000000000000000000111001100110;
assign LUT_1[2203] = 32'b11111111111111111010001011100010;
assign LUT_1[2204] = 32'b00000000000000001101000100101100;
assign LUT_1[2205] = 32'b00000000000000000110010110101000;
assign LUT_1[2206] = 32'b00000000000000001000110010111101;
assign LUT_1[2207] = 32'b00000000000000000010000100111001;
assign LUT_1[2208] = 32'b00000000000000000100111100111101;
assign LUT_1[2209] = 32'b11111111111111111110001110111001;
assign LUT_1[2210] = 32'b00000000000000000000101011001110;
assign LUT_1[2211] = 32'b11111111111111111001111101001010;
assign LUT_1[2212] = 32'b00000000000000001100110110010100;
assign LUT_1[2213] = 32'b00000000000000000110001000010000;
assign LUT_1[2214] = 32'b00000000000000001000100100100101;
assign LUT_1[2215] = 32'b00000000000000000001110110100001;
assign LUT_1[2216] = 32'b00000000000000000100001010110010;
assign LUT_1[2217] = 32'b11111111111111111101011100101110;
assign LUT_1[2218] = 32'b11111111111111111111111001000011;
assign LUT_1[2219] = 32'b11111111111111111001001010111111;
assign LUT_1[2220] = 32'b00000000000000001100000100001001;
assign LUT_1[2221] = 32'b00000000000000000101010110000101;
assign LUT_1[2222] = 32'b00000000000000000111110010011010;
assign LUT_1[2223] = 32'b00000000000000000001000100010110;
assign LUT_1[2224] = 32'b00000000000000000110111000011111;
assign LUT_1[2225] = 32'b00000000000000000000001010011011;
assign LUT_1[2226] = 32'b00000000000000000010100110110000;
assign LUT_1[2227] = 32'b11111111111111111011111000101100;
assign LUT_1[2228] = 32'b00000000000000001110110001110110;
assign LUT_1[2229] = 32'b00000000000000001000000011110010;
assign LUT_1[2230] = 32'b00000000000000001010100000000111;
assign LUT_1[2231] = 32'b00000000000000000011110010000011;
assign LUT_1[2232] = 32'b00000000000000000110000110010100;
assign LUT_1[2233] = 32'b11111111111111111111011000010000;
assign LUT_1[2234] = 32'b00000000000000000001110100100101;
assign LUT_1[2235] = 32'b11111111111111111011000110100001;
assign LUT_1[2236] = 32'b00000000000000001101111111101011;
assign LUT_1[2237] = 32'b00000000000000000111010001100111;
assign LUT_1[2238] = 32'b00000000000000001001101101111100;
assign LUT_1[2239] = 32'b00000000000000000010111111111000;
assign LUT_1[2240] = 32'b00000000000000000101111111100110;
assign LUT_1[2241] = 32'b11111111111111111111010001100010;
assign LUT_1[2242] = 32'b00000000000000000001101101110111;
assign LUT_1[2243] = 32'b11111111111111111010111111110011;
assign LUT_1[2244] = 32'b00000000000000001101111000111101;
assign LUT_1[2245] = 32'b00000000000000000111001010111001;
assign LUT_1[2246] = 32'b00000000000000001001100111001110;
assign LUT_1[2247] = 32'b00000000000000000010111001001010;
assign LUT_1[2248] = 32'b00000000000000000101001101011011;
assign LUT_1[2249] = 32'b11111111111111111110011111010111;
assign LUT_1[2250] = 32'b00000000000000000000111011101100;
assign LUT_1[2251] = 32'b11111111111111111010001101101000;
assign LUT_1[2252] = 32'b00000000000000001101000110110010;
assign LUT_1[2253] = 32'b00000000000000000110011000101110;
assign LUT_1[2254] = 32'b00000000000000001000110101000011;
assign LUT_1[2255] = 32'b00000000000000000010000110111111;
assign LUT_1[2256] = 32'b00000000000000000111111011001000;
assign LUT_1[2257] = 32'b00000000000000000001001101000100;
assign LUT_1[2258] = 32'b00000000000000000011101001011001;
assign LUT_1[2259] = 32'b11111111111111111100111011010101;
assign LUT_1[2260] = 32'b00000000000000001111110100011111;
assign LUT_1[2261] = 32'b00000000000000001001000110011011;
assign LUT_1[2262] = 32'b00000000000000001011100010110000;
assign LUT_1[2263] = 32'b00000000000000000100110100101100;
assign LUT_1[2264] = 32'b00000000000000000111001000111101;
assign LUT_1[2265] = 32'b00000000000000000000011010111001;
assign LUT_1[2266] = 32'b00000000000000000010110111001110;
assign LUT_1[2267] = 32'b11111111111111111100001001001010;
assign LUT_1[2268] = 32'b00000000000000001111000010010100;
assign LUT_1[2269] = 32'b00000000000000001000010100010000;
assign LUT_1[2270] = 32'b00000000000000001010110000100101;
assign LUT_1[2271] = 32'b00000000000000000100000010100001;
assign LUT_1[2272] = 32'b00000000000000000110111010100101;
assign LUT_1[2273] = 32'b00000000000000000000001100100001;
assign LUT_1[2274] = 32'b00000000000000000010101000110110;
assign LUT_1[2275] = 32'b11111111111111111011111010110010;
assign LUT_1[2276] = 32'b00000000000000001110110011111100;
assign LUT_1[2277] = 32'b00000000000000001000000101111000;
assign LUT_1[2278] = 32'b00000000000000001010100010001101;
assign LUT_1[2279] = 32'b00000000000000000011110100001001;
assign LUT_1[2280] = 32'b00000000000000000110001000011010;
assign LUT_1[2281] = 32'b11111111111111111111011010010110;
assign LUT_1[2282] = 32'b00000000000000000001110110101011;
assign LUT_1[2283] = 32'b11111111111111111011001000100111;
assign LUT_1[2284] = 32'b00000000000000001110000001110001;
assign LUT_1[2285] = 32'b00000000000000000111010011101101;
assign LUT_1[2286] = 32'b00000000000000001001110000000010;
assign LUT_1[2287] = 32'b00000000000000000011000001111110;
assign LUT_1[2288] = 32'b00000000000000001000110110000111;
assign LUT_1[2289] = 32'b00000000000000000010001000000011;
assign LUT_1[2290] = 32'b00000000000000000100100100011000;
assign LUT_1[2291] = 32'b11111111111111111101110110010100;
assign LUT_1[2292] = 32'b00000000000000010000101111011110;
assign LUT_1[2293] = 32'b00000000000000001010000001011010;
assign LUT_1[2294] = 32'b00000000000000001100011101101111;
assign LUT_1[2295] = 32'b00000000000000000101101111101011;
assign LUT_1[2296] = 32'b00000000000000001000000011111100;
assign LUT_1[2297] = 32'b00000000000000000001010101111000;
assign LUT_1[2298] = 32'b00000000000000000011110010001101;
assign LUT_1[2299] = 32'b11111111111111111101000100001001;
assign LUT_1[2300] = 32'b00000000000000001111111101010011;
assign LUT_1[2301] = 32'b00000000000000001001001111001111;
assign LUT_1[2302] = 32'b00000000000000001011101011100100;
assign LUT_1[2303] = 32'b00000000000000000100111101100000;
assign LUT_1[2304] = 32'b11111111111111111110110110000111;
assign LUT_1[2305] = 32'b11111111111111111000001000000011;
assign LUT_1[2306] = 32'b11111111111111111010100100011000;
assign LUT_1[2307] = 32'b11111111111111110011110110010100;
assign LUT_1[2308] = 32'b00000000000000000110101111011110;
assign LUT_1[2309] = 32'b00000000000000000000000001011010;
assign LUT_1[2310] = 32'b00000000000000000010011101101111;
assign LUT_1[2311] = 32'b11111111111111111011101111101011;
assign LUT_1[2312] = 32'b11111111111111111110000011111100;
assign LUT_1[2313] = 32'b11111111111111110111010101111000;
assign LUT_1[2314] = 32'b11111111111111111001110010001101;
assign LUT_1[2315] = 32'b11111111111111110011000100001001;
assign LUT_1[2316] = 32'b00000000000000000101111101010011;
assign LUT_1[2317] = 32'b11111111111111111111001111001111;
assign LUT_1[2318] = 32'b00000000000000000001101011100100;
assign LUT_1[2319] = 32'b11111111111111111010111101100000;
assign LUT_1[2320] = 32'b00000000000000000000110001101001;
assign LUT_1[2321] = 32'b11111111111111111010000011100101;
assign LUT_1[2322] = 32'b11111111111111111100011111111010;
assign LUT_1[2323] = 32'b11111111111111110101110001110110;
assign LUT_1[2324] = 32'b00000000000000001000101011000000;
assign LUT_1[2325] = 32'b00000000000000000001111100111100;
assign LUT_1[2326] = 32'b00000000000000000100011001010001;
assign LUT_1[2327] = 32'b11111111111111111101101011001101;
assign LUT_1[2328] = 32'b11111111111111111111111111011110;
assign LUT_1[2329] = 32'b11111111111111111001010001011010;
assign LUT_1[2330] = 32'b11111111111111111011101101101111;
assign LUT_1[2331] = 32'b11111111111111110100111111101011;
assign LUT_1[2332] = 32'b00000000000000000111111000110101;
assign LUT_1[2333] = 32'b00000000000000000001001010110001;
assign LUT_1[2334] = 32'b00000000000000000011100111000110;
assign LUT_1[2335] = 32'b11111111111111111100111001000010;
assign LUT_1[2336] = 32'b11111111111111111111110001000110;
assign LUT_1[2337] = 32'b11111111111111111001000011000010;
assign LUT_1[2338] = 32'b11111111111111111011011111010111;
assign LUT_1[2339] = 32'b11111111111111110100110001010011;
assign LUT_1[2340] = 32'b00000000000000000111101010011101;
assign LUT_1[2341] = 32'b00000000000000000000111100011001;
assign LUT_1[2342] = 32'b00000000000000000011011000101110;
assign LUT_1[2343] = 32'b11111111111111111100101010101010;
assign LUT_1[2344] = 32'b11111111111111111110111110111011;
assign LUT_1[2345] = 32'b11111111111111111000010000110111;
assign LUT_1[2346] = 32'b11111111111111111010101101001100;
assign LUT_1[2347] = 32'b11111111111111110011111111001000;
assign LUT_1[2348] = 32'b00000000000000000110111000010010;
assign LUT_1[2349] = 32'b00000000000000000000001010001110;
assign LUT_1[2350] = 32'b00000000000000000010100110100011;
assign LUT_1[2351] = 32'b11111111111111111011111000011111;
assign LUT_1[2352] = 32'b00000000000000000001101100101000;
assign LUT_1[2353] = 32'b11111111111111111010111110100100;
assign LUT_1[2354] = 32'b11111111111111111101011010111001;
assign LUT_1[2355] = 32'b11111111111111110110101100110101;
assign LUT_1[2356] = 32'b00000000000000001001100101111111;
assign LUT_1[2357] = 32'b00000000000000000010110111111011;
assign LUT_1[2358] = 32'b00000000000000000101010100010000;
assign LUT_1[2359] = 32'b11111111111111111110100110001100;
assign LUT_1[2360] = 32'b00000000000000000000111010011101;
assign LUT_1[2361] = 32'b11111111111111111010001100011001;
assign LUT_1[2362] = 32'b11111111111111111100101000101110;
assign LUT_1[2363] = 32'b11111111111111110101111010101010;
assign LUT_1[2364] = 32'b00000000000000001000110011110100;
assign LUT_1[2365] = 32'b00000000000000000010000101110000;
assign LUT_1[2366] = 32'b00000000000000000100100010000101;
assign LUT_1[2367] = 32'b11111111111111111101110100000001;
assign LUT_1[2368] = 32'b00000000000000000000110011101111;
assign LUT_1[2369] = 32'b11111111111111111010000101101011;
assign LUT_1[2370] = 32'b11111111111111111100100010000000;
assign LUT_1[2371] = 32'b11111111111111110101110011111100;
assign LUT_1[2372] = 32'b00000000000000001000101101000110;
assign LUT_1[2373] = 32'b00000000000000000001111111000010;
assign LUT_1[2374] = 32'b00000000000000000100011011010111;
assign LUT_1[2375] = 32'b11111111111111111101101101010011;
assign LUT_1[2376] = 32'b00000000000000000000000001100100;
assign LUT_1[2377] = 32'b11111111111111111001010011100000;
assign LUT_1[2378] = 32'b11111111111111111011101111110101;
assign LUT_1[2379] = 32'b11111111111111110101000001110001;
assign LUT_1[2380] = 32'b00000000000000000111111010111011;
assign LUT_1[2381] = 32'b00000000000000000001001100110111;
assign LUT_1[2382] = 32'b00000000000000000011101001001100;
assign LUT_1[2383] = 32'b11111111111111111100111011001000;
assign LUT_1[2384] = 32'b00000000000000000010101111010001;
assign LUT_1[2385] = 32'b11111111111111111100000001001101;
assign LUT_1[2386] = 32'b11111111111111111110011101100010;
assign LUT_1[2387] = 32'b11111111111111110111101111011110;
assign LUT_1[2388] = 32'b00000000000000001010101000101000;
assign LUT_1[2389] = 32'b00000000000000000011111010100100;
assign LUT_1[2390] = 32'b00000000000000000110010110111001;
assign LUT_1[2391] = 32'b11111111111111111111101000110101;
assign LUT_1[2392] = 32'b00000000000000000001111101000110;
assign LUT_1[2393] = 32'b11111111111111111011001111000010;
assign LUT_1[2394] = 32'b11111111111111111101101011010111;
assign LUT_1[2395] = 32'b11111111111111110110111101010011;
assign LUT_1[2396] = 32'b00000000000000001001110110011101;
assign LUT_1[2397] = 32'b00000000000000000011001000011001;
assign LUT_1[2398] = 32'b00000000000000000101100100101110;
assign LUT_1[2399] = 32'b11111111111111111110110110101010;
assign LUT_1[2400] = 32'b00000000000000000001101110101110;
assign LUT_1[2401] = 32'b11111111111111111011000000101010;
assign LUT_1[2402] = 32'b11111111111111111101011100111111;
assign LUT_1[2403] = 32'b11111111111111110110101110111011;
assign LUT_1[2404] = 32'b00000000000000001001101000000101;
assign LUT_1[2405] = 32'b00000000000000000010111010000001;
assign LUT_1[2406] = 32'b00000000000000000101010110010110;
assign LUT_1[2407] = 32'b11111111111111111110101000010010;
assign LUT_1[2408] = 32'b00000000000000000000111100100011;
assign LUT_1[2409] = 32'b11111111111111111010001110011111;
assign LUT_1[2410] = 32'b11111111111111111100101010110100;
assign LUT_1[2411] = 32'b11111111111111110101111100110000;
assign LUT_1[2412] = 32'b00000000000000001000110101111010;
assign LUT_1[2413] = 32'b00000000000000000010000111110110;
assign LUT_1[2414] = 32'b00000000000000000100100100001011;
assign LUT_1[2415] = 32'b11111111111111111101110110000111;
assign LUT_1[2416] = 32'b00000000000000000011101010010000;
assign LUT_1[2417] = 32'b11111111111111111100111100001100;
assign LUT_1[2418] = 32'b11111111111111111111011000100001;
assign LUT_1[2419] = 32'b11111111111111111000101010011101;
assign LUT_1[2420] = 32'b00000000000000001011100011100111;
assign LUT_1[2421] = 32'b00000000000000000100110101100011;
assign LUT_1[2422] = 32'b00000000000000000111010001111000;
assign LUT_1[2423] = 32'b00000000000000000000100011110100;
assign LUT_1[2424] = 32'b00000000000000000010111000000101;
assign LUT_1[2425] = 32'b11111111111111111100001010000001;
assign LUT_1[2426] = 32'b11111111111111111110100110010110;
assign LUT_1[2427] = 32'b11111111111111110111111000010010;
assign LUT_1[2428] = 32'b00000000000000001010110001011100;
assign LUT_1[2429] = 32'b00000000000000000100000011011000;
assign LUT_1[2430] = 32'b00000000000000000110011111101101;
assign LUT_1[2431] = 32'b11111111111111111111110001101001;
assign LUT_1[2432] = 32'b00000000000000000001110110001010;
assign LUT_1[2433] = 32'b11111111111111111011001000000110;
assign LUT_1[2434] = 32'b11111111111111111101100100011011;
assign LUT_1[2435] = 32'b11111111111111110110110110010111;
assign LUT_1[2436] = 32'b00000000000000001001101111100001;
assign LUT_1[2437] = 32'b00000000000000000011000001011101;
assign LUT_1[2438] = 32'b00000000000000000101011101110010;
assign LUT_1[2439] = 32'b11111111111111111110101111101110;
assign LUT_1[2440] = 32'b00000000000000000001000011111111;
assign LUT_1[2441] = 32'b11111111111111111010010101111011;
assign LUT_1[2442] = 32'b11111111111111111100110010010000;
assign LUT_1[2443] = 32'b11111111111111110110000100001100;
assign LUT_1[2444] = 32'b00000000000000001000111101010110;
assign LUT_1[2445] = 32'b00000000000000000010001111010010;
assign LUT_1[2446] = 32'b00000000000000000100101011100111;
assign LUT_1[2447] = 32'b11111111111111111101111101100011;
assign LUT_1[2448] = 32'b00000000000000000011110001101100;
assign LUT_1[2449] = 32'b11111111111111111101000011101000;
assign LUT_1[2450] = 32'b11111111111111111111011111111101;
assign LUT_1[2451] = 32'b11111111111111111000110001111001;
assign LUT_1[2452] = 32'b00000000000000001011101011000011;
assign LUT_1[2453] = 32'b00000000000000000100111100111111;
assign LUT_1[2454] = 32'b00000000000000000111011001010100;
assign LUT_1[2455] = 32'b00000000000000000000101011010000;
assign LUT_1[2456] = 32'b00000000000000000010111111100001;
assign LUT_1[2457] = 32'b11111111111111111100010001011101;
assign LUT_1[2458] = 32'b11111111111111111110101101110010;
assign LUT_1[2459] = 32'b11111111111111110111111111101110;
assign LUT_1[2460] = 32'b00000000000000001010111000111000;
assign LUT_1[2461] = 32'b00000000000000000100001010110100;
assign LUT_1[2462] = 32'b00000000000000000110100111001001;
assign LUT_1[2463] = 32'b11111111111111111111111001000101;
assign LUT_1[2464] = 32'b00000000000000000010110001001001;
assign LUT_1[2465] = 32'b11111111111111111100000011000101;
assign LUT_1[2466] = 32'b11111111111111111110011111011010;
assign LUT_1[2467] = 32'b11111111111111110111110001010110;
assign LUT_1[2468] = 32'b00000000000000001010101010100000;
assign LUT_1[2469] = 32'b00000000000000000011111100011100;
assign LUT_1[2470] = 32'b00000000000000000110011000110001;
assign LUT_1[2471] = 32'b11111111111111111111101010101101;
assign LUT_1[2472] = 32'b00000000000000000001111110111110;
assign LUT_1[2473] = 32'b11111111111111111011010000111010;
assign LUT_1[2474] = 32'b11111111111111111101101101001111;
assign LUT_1[2475] = 32'b11111111111111110110111111001011;
assign LUT_1[2476] = 32'b00000000000000001001111000010101;
assign LUT_1[2477] = 32'b00000000000000000011001010010001;
assign LUT_1[2478] = 32'b00000000000000000101100110100110;
assign LUT_1[2479] = 32'b11111111111111111110111000100010;
assign LUT_1[2480] = 32'b00000000000000000100101100101011;
assign LUT_1[2481] = 32'b11111111111111111101111110100111;
assign LUT_1[2482] = 32'b00000000000000000000011010111100;
assign LUT_1[2483] = 32'b11111111111111111001101100111000;
assign LUT_1[2484] = 32'b00000000000000001100100110000010;
assign LUT_1[2485] = 32'b00000000000000000101110111111110;
assign LUT_1[2486] = 32'b00000000000000001000010100010011;
assign LUT_1[2487] = 32'b00000000000000000001100110001111;
assign LUT_1[2488] = 32'b00000000000000000011111010100000;
assign LUT_1[2489] = 32'b11111111111111111101001100011100;
assign LUT_1[2490] = 32'b11111111111111111111101000110001;
assign LUT_1[2491] = 32'b11111111111111111000111010101101;
assign LUT_1[2492] = 32'b00000000000000001011110011110111;
assign LUT_1[2493] = 32'b00000000000000000101000101110011;
assign LUT_1[2494] = 32'b00000000000000000111100010001000;
assign LUT_1[2495] = 32'b00000000000000000000110100000100;
assign LUT_1[2496] = 32'b00000000000000000011110011110010;
assign LUT_1[2497] = 32'b11111111111111111101000101101110;
assign LUT_1[2498] = 32'b11111111111111111111100010000011;
assign LUT_1[2499] = 32'b11111111111111111000110011111111;
assign LUT_1[2500] = 32'b00000000000000001011101101001001;
assign LUT_1[2501] = 32'b00000000000000000100111111000101;
assign LUT_1[2502] = 32'b00000000000000000111011011011010;
assign LUT_1[2503] = 32'b00000000000000000000101101010110;
assign LUT_1[2504] = 32'b00000000000000000011000001100111;
assign LUT_1[2505] = 32'b11111111111111111100010011100011;
assign LUT_1[2506] = 32'b11111111111111111110101111111000;
assign LUT_1[2507] = 32'b11111111111111111000000001110100;
assign LUT_1[2508] = 32'b00000000000000001010111010111110;
assign LUT_1[2509] = 32'b00000000000000000100001100111010;
assign LUT_1[2510] = 32'b00000000000000000110101001001111;
assign LUT_1[2511] = 32'b11111111111111111111111011001011;
assign LUT_1[2512] = 32'b00000000000000000101101111010100;
assign LUT_1[2513] = 32'b11111111111111111111000001010000;
assign LUT_1[2514] = 32'b00000000000000000001011101100101;
assign LUT_1[2515] = 32'b11111111111111111010101111100001;
assign LUT_1[2516] = 32'b00000000000000001101101000101011;
assign LUT_1[2517] = 32'b00000000000000000110111010100111;
assign LUT_1[2518] = 32'b00000000000000001001010110111100;
assign LUT_1[2519] = 32'b00000000000000000010101000111000;
assign LUT_1[2520] = 32'b00000000000000000100111101001001;
assign LUT_1[2521] = 32'b11111111111111111110001111000101;
assign LUT_1[2522] = 32'b00000000000000000000101011011010;
assign LUT_1[2523] = 32'b11111111111111111001111101010110;
assign LUT_1[2524] = 32'b00000000000000001100110110100000;
assign LUT_1[2525] = 32'b00000000000000000110001000011100;
assign LUT_1[2526] = 32'b00000000000000001000100100110001;
assign LUT_1[2527] = 32'b00000000000000000001110110101101;
assign LUT_1[2528] = 32'b00000000000000000100101110110001;
assign LUT_1[2529] = 32'b11111111111111111110000000101101;
assign LUT_1[2530] = 32'b00000000000000000000011101000010;
assign LUT_1[2531] = 32'b11111111111111111001101110111110;
assign LUT_1[2532] = 32'b00000000000000001100101000001000;
assign LUT_1[2533] = 32'b00000000000000000101111010000100;
assign LUT_1[2534] = 32'b00000000000000001000010110011001;
assign LUT_1[2535] = 32'b00000000000000000001101000010101;
assign LUT_1[2536] = 32'b00000000000000000011111100100110;
assign LUT_1[2537] = 32'b11111111111111111101001110100010;
assign LUT_1[2538] = 32'b11111111111111111111101010110111;
assign LUT_1[2539] = 32'b11111111111111111000111100110011;
assign LUT_1[2540] = 32'b00000000000000001011110101111101;
assign LUT_1[2541] = 32'b00000000000000000101000111111001;
assign LUT_1[2542] = 32'b00000000000000000111100100001110;
assign LUT_1[2543] = 32'b00000000000000000000110110001010;
assign LUT_1[2544] = 32'b00000000000000000110101010010011;
assign LUT_1[2545] = 32'b11111111111111111111111100001111;
assign LUT_1[2546] = 32'b00000000000000000010011000100100;
assign LUT_1[2547] = 32'b11111111111111111011101010100000;
assign LUT_1[2548] = 32'b00000000000000001110100011101010;
assign LUT_1[2549] = 32'b00000000000000000111110101100110;
assign LUT_1[2550] = 32'b00000000000000001010010001111011;
assign LUT_1[2551] = 32'b00000000000000000011100011110111;
assign LUT_1[2552] = 32'b00000000000000000101111000001000;
assign LUT_1[2553] = 32'b11111111111111111111001010000100;
assign LUT_1[2554] = 32'b00000000000000000001100110011001;
assign LUT_1[2555] = 32'b11111111111111111010111000010101;
assign LUT_1[2556] = 32'b00000000000000001101110001011111;
assign LUT_1[2557] = 32'b00000000000000000111000011011011;
assign LUT_1[2558] = 32'b00000000000000001001011111110000;
assign LUT_1[2559] = 32'b00000000000000000010110001101100;
assign LUT_1[2560] = 32'b11111111111111111010110000011000;
assign LUT_1[2561] = 32'b11111111111111110100000010010100;
assign LUT_1[2562] = 32'b11111111111111110110011110101001;
assign LUT_1[2563] = 32'b11111111111111101111110000100101;
assign LUT_1[2564] = 32'b00000000000000000010101001101111;
assign LUT_1[2565] = 32'b11111111111111111011111011101011;
assign LUT_1[2566] = 32'b11111111111111111110011000000000;
assign LUT_1[2567] = 32'b11111111111111110111101001111100;
assign LUT_1[2568] = 32'b11111111111111111001111110001101;
assign LUT_1[2569] = 32'b11111111111111110011010000001001;
assign LUT_1[2570] = 32'b11111111111111110101101100011110;
assign LUT_1[2571] = 32'b11111111111111101110111110011010;
assign LUT_1[2572] = 32'b00000000000000000001110111100100;
assign LUT_1[2573] = 32'b11111111111111111011001001100000;
assign LUT_1[2574] = 32'b11111111111111111101100101110101;
assign LUT_1[2575] = 32'b11111111111111110110110111110001;
assign LUT_1[2576] = 32'b11111111111111111100101011111010;
assign LUT_1[2577] = 32'b11111111111111110101111101110110;
assign LUT_1[2578] = 32'b11111111111111111000011010001011;
assign LUT_1[2579] = 32'b11111111111111110001101100000111;
assign LUT_1[2580] = 32'b00000000000000000100100101010001;
assign LUT_1[2581] = 32'b11111111111111111101110111001101;
assign LUT_1[2582] = 32'b00000000000000000000010011100010;
assign LUT_1[2583] = 32'b11111111111111111001100101011110;
assign LUT_1[2584] = 32'b11111111111111111011111001101111;
assign LUT_1[2585] = 32'b11111111111111110101001011101011;
assign LUT_1[2586] = 32'b11111111111111110111101000000000;
assign LUT_1[2587] = 32'b11111111111111110000111001111100;
assign LUT_1[2588] = 32'b00000000000000000011110011000110;
assign LUT_1[2589] = 32'b11111111111111111101000101000010;
assign LUT_1[2590] = 32'b11111111111111111111100001010111;
assign LUT_1[2591] = 32'b11111111111111111000110011010011;
assign LUT_1[2592] = 32'b11111111111111111011101011010111;
assign LUT_1[2593] = 32'b11111111111111110100111101010011;
assign LUT_1[2594] = 32'b11111111111111110111011001101000;
assign LUT_1[2595] = 32'b11111111111111110000101011100100;
assign LUT_1[2596] = 32'b00000000000000000011100100101110;
assign LUT_1[2597] = 32'b11111111111111111100110110101010;
assign LUT_1[2598] = 32'b11111111111111111111010010111111;
assign LUT_1[2599] = 32'b11111111111111111000100100111011;
assign LUT_1[2600] = 32'b11111111111111111010111001001100;
assign LUT_1[2601] = 32'b11111111111111110100001011001000;
assign LUT_1[2602] = 32'b11111111111111110110100111011101;
assign LUT_1[2603] = 32'b11111111111111101111111001011001;
assign LUT_1[2604] = 32'b00000000000000000010110010100011;
assign LUT_1[2605] = 32'b11111111111111111100000100011111;
assign LUT_1[2606] = 32'b11111111111111111110100000110100;
assign LUT_1[2607] = 32'b11111111111111110111110010110000;
assign LUT_1[2608] = 32'b11111111111111111101100110111001;
assign LUT_1[2609] = 32'b11111111111111110110111000110101;
assign LUT_1[2610] = 32'b11111111111111111001010101001010;
assign LUT_1[2611] = 32'b11111111111111110010100111000110;
assign LUT_1[2612] = 32'b00000000000000000101100000010000;
assign LUT_1[2613] = 32'b11111111111111111110110010001100;
assign LUT_1[2614] = 32'b00000000000000000001001110100001;
assign LUT_1[2615] = 32'b11111111111111111010100000011101;
assign LUT_1[2616] = 32'b11111111111111111100110100101110;
assign LUT_1[2617] = 32'b11111111111111110110000110101010;
assign LUT_1[2618] = 32'b11111111111111111000100010111111;
assign LUT_1[2619] = 32'b11111111111111110001110100111011;
assign LUT_1[2620] = 32'b00000000000000000100101110000101;
assign LUT_1[2621] = 32'b11111111111111111110000000000001;
assign LUT_1[2622] = 32'b00000000000000000000011100010110;
assign LUT_1[2623] = 32'b11111111111111111001101110010010;
assign LUT_1[2624] = 32'b11111111111111111100101110000000;
assign LUT_1[2625] = 32'b11111111111111110101111111111100;
assign LUT_1[2626] = 32'b11111111111111111000011100010001;
assign LUT_1[2627] = 32'b11111111111111110001101110001101;
assign LUT_1[2628] = 32'b00000000000000000100100111010111;
assign LUT_1[2629] = 32'b11111111111111111101111001010011;
assign LUT_1[2630] = 32'b00000000000000000000010101101000;
assign LUT_1[2631] = 32'b11111111111111111001100111100100;
assign LUT_1[2632] = 32'b11111111111111111011111011110101;
assign LUT_1[2633] = 32'b11111111111111110101001101110001;
assign LUT_1[2634] = 32'b11111111111111110111101010000110;
assign LUT_1[2635] = 32'b11111111111111110000111100000010;
assign LUT_1[2636] = 32'b00000000000000000011110101001100;
assign LUT_1[2637] = 32'b11111111111111111101000111001000;
assign LUT_1[2638] = 32'b11111111111111111111100011011101;
assign LUT_1[2639] = 32'b11111111111111111000110101011001;
assign LUT_1[2640] = 32'b11111111111111111110101001100010;
assign LUT_1[2641] = 32'b11111111111111110111111011011110;
assign LUT_1[2642] = 32'b11111111111111111010010111110011;
assign LUT_1[2643] = 32'b11111111111111110011101001101111;
assign LUT_1[2644] = 32'b00000000000000000110100010111001;
assign LUT_1[2645] = 32'b11111111111111111111110100110101;
assign LUT_1[2646] = 32'b00000000000000000010010001001010;
assign LUT_1[2647] = 32'b11111111111111111011100011000110;
assign LUT_1[2648] = 32'b11111111111111111101110111010111;
assign LUT_1[2649] = 32'b11111111111111110111001001010011;
assign LUT_1[2650] = 32'b11111111111111111001100101101000;
assign LUT_1[2651] = 32'b11111111111111110010110111100100;
assign LUT_1[2652] = 32'b00000000000000000101110000101110;
assign LUT_1[2653] = 32'b11111111111111111111000010101010;
assign LUT_1[2654] = 32'b00000000000000000001011110111111;
assign LUT_1[2655] = 32'b11111111111111111010110000111011;
assign LUT_1[2656] = 32'b11111111111111111101101000111111;
assign LUT_1[2657] = 32'b11111111111111110110111010111011;
assign LUT_1[2658] = 32'b11111111111111111001010111010000;
assign LUT_1[2659] = 32'b11111111111111110010101001001100;
assign LUT_1[2660] = 32'b00000000000000000101100010010110;
assign LUT_1[2661] = 32'b11111111111111111110110100010010;
assign LUT_1[2662] = 32'b00000000000000000001010000100111;
assign LUT_1[2663] = 32'b11111111111111111010100010100011;
assign LUT_1[2664] = 32'b11111111111111111100110110110100;
assign LUT_1[2665] = 32'b11111111111111110110001000110000;
assign LUT_1[2666] = 32'b11111111111111111000100101000101;
assign LUT_1[2667] = 32'b11111111111111110001110111000001;
assign LUT_1[2668] = 32'b00000000000000000100110000001011;
assign LUT_1[2669] = 32'b11111111111111111110000010000111;
assign LUT_1[2670] = 32'b00000000000000000000011110011100;
assign LUT_1[2671] = 32'b11111111111111111001110000011000;
assign LUT_1[2672] = 32'b11111111111111111111100100100001;
assign LUT_1[2673] = 32'b11111111111111111000110110011101;
assign LUT_1[2674] = 32'b11111111111111111011010010110010;
assign LUT_1[2675] = 32'b11111111111111110100100100101110;
assign LUT_1[2676] = 32'b00000000000000000111011101111000;
assign LUT_1[2677] = 32'b00000000000000000000101111110100;
assign LUT_1[2678] = 32'b00000000000000000011001100001001;
assign LUT_1[2679] = 32'b11111111111111111100011110000101;
assign LUT_1[2680] = 32'b11111111111111111110110010010110;
assign LUT_1[2681] = 32'b11111111111111111000000100010010;
assign LUT_1[2682] = 32'b11111111111111111010100000100111;
assign LUT_1[2683] = 32'b11111111111111110011110010100011;
assign LUT_1[2684] = 32'b00000000000000000110101011101101;
assign LUT_1[2685] = 32'b11111111111111111111111101101001;
assign LUT_1[2686] = 32'b00000000000000000010011001111110;
assign LUT_1[2687] = 32'b11111111111111111011101011111010;
assign LUT_1[2688] = 32'b11111111111111111101110000011011;
assign LUT_1[2689] = 32'b11111111111111110111000010010111;
assign LUT_1[2690] = 32'b11111111111111111001011110101100;
assign LUT_1[2691] = 32'b11111111111111110010110000101000;
assign LUT_1[2692] = 32'b00000000000000000101101001110010;
assign LUT_1[2693] = 32'b11111111111111111110111011101110;
assign LUT_1[2694] = 32'b00000000000000000001011000000011;
assign LUT_1[2695] = 32'b11111111111111111010101001111111;
assign LUT_1[2696] = 32'b11111111111111111100111110010000;
assign LUT_1[2697] = 32'b11111111111111110110010000001100;
assign LUT_1[2698] = 32'b11111111111111111000101100100001;
assign LUT_1[2699] = 32'b11111111111111110001111110011101;
assign LUT_1[2700] = 32'b00000000000000000100110111100111;
assign LUT_1[2701] = 32'b11111111111111111110001001100011;
assign LUT_1[2702] = 32'b00000000000000000000100101111000;
assign LUT_1[2703] = 32'b11111111111111111001110111110100;
assign LUT_1[2704] = 32'b11111111111111111111101011111101;
assign LUT_1[2705] = 32'b11111111111111111000111101111001;
assign LUT_1[2706] = 32'b11111111111111111011011010001110;
assign LUT_1[2707] = 32'b11111111111111110100101100001010;
assign LUT_1[2708] = 32'b00000000000000000111100101010100;
assign LUT_1[2709] = 32'b00000000000000000000110111010000;
assign LUT_1[2710] = 32'b00000000000000000011010011100101;
assign LUT_1[2711] = 32'b11111111111111111100100101100001;
assign LUT_1[2712] = 32'b11111111111111111110111001110010;
assign LUT_1[2713] = 32'b11111111111111111000001011101110;
assign LUT_1[2714] = 32'b11111111111111111010101000000011;
assign LUT_1[2715] = 32'b11111111111111110011111001111111;
assign LUT_1[2716] = 32'b00000000000000000110110011001001;
assign LUT_1[2717] = 32'b00000000000000000000000101000101;
assign LUT_1[2718] = 32'b00000000000000000010100001011010;
assign LUT_1[2719] = 32'b11111111111111111011110011010110;
assign LUT_1[2720] = 32'b11111111111111111110101011011010;
assign LUT_1[2721] = 32'b11111111111111110111111101010110;
assign LUT_1[2722] = 32'b11111111111111111010011001101011;
assign LUT_1[2723] = 32'b11111111111111110011101011100111;
assign LUT_1[2724] = 32'b00000000000000000110100100110001;
assign LUT_1[2725] = 32'b11111111111111111111110110101101;
assign LUT_1[2726] = 32'b00000000000000000010010011000010;
assign LUT_1[2727] = 32'b11111111111111111011100100111110;
assign LUT_1[2728] = 32'b11111111111111111101111001001111;
assign LUT_1[2729] = 32'b11111111111111110111001011001011;
assign LUT_1[2730] = 32'b11111111111111111001100111100000;
assign LUT_1[2731] = 32'b11111111111111110010111001011100;
assign LUT_1[2732] = 32'b00000000000000000101110010100110;
assign LUT_1[2733] = 32'b11111111111111111111000100100010;
assign LUT_1[2734] = 32'b00000000000000000001100000110111;
assign LUT_1[2735] = 32'b11111111111111111010110010110011;
assign LUT_1[2736] = 32'b00000000000000000000100110111100;
assign LUT_1[2737] = 32'b11111111111111111001111000111000;
assign LUT_1[2738] = 32'b11111111111111111100010101001101;
assign LUT_1[2739] = 32'b11111111111111110101100111001001;
assign LUT_1[2740] = 32'b00000000000000001000100000010011;
assign LUT_1[2741] = 32'b00000000000000000001110010001111;
assign LUT_1[2742] = 32'b00000000000000000100001110100100;
assign LUT_1[2743] = 32'b11111111111111111101100000100000;
assign LUT_1[2744] = 32'b11111111111111111111110100110001;
assign LUT_1[2745] = 32'b11111111111111111001000110101101;
assign LUT_1[2746] = 32'b11111111111111111011100011000010;
assign LUT_1[2747] = 32'b11111111111111110100110100111110;
assign LUT_1[2748] = 32'b00000000000000000111101110001000;
assign LUT_1[2749] = 32'b00000000000000000001000000000100;
assign LUT_1[2750] = 32'b00000000000000000011011100011001;
assign LUT_1[2751] = 32'b11111111111111111100101110010101;
assign LUT_1[2752] = 32'b11111111111111111111101110000011;
assign LUT_1[2753] = 32'b11111111111111111000111111111111;
assign LUT_1[2754] = 32'b11111111111111111011011100010100;
assign LUT_1[2755] = 32'b11111111111111110100101110010000;
assign LUT_1[2756] = 32'b00000000000000000111100111011010;
assign LUT_1[2757] = 32'b00000000000000000000111001010110;
assign LUT_1[2758] = 32'b00000000000000000011010101101011;
assign LUT_1[2759] = 32'b11111111111111111100100111100111;
assign LUT_1[2760] = 32'b11111111111111111110111011111000;
assign LUT_1[2761] = 32'b11111111111111111000001101110100;
assign LUT_1[2762] = 32'b11111111111111111010101010001001;
assign LUT_1[2763] = 32'b11111111111111110011111100000101;
assign LUT_1[2764] = 32'b00000000000000000110110101001111;
assign LUT_1[2765] = 32'b00000000000000000000000111001011;
assign LUT_1[2766] = 32'b00000000000000000010100011100000;
assign LUT_1[2767] = 32'b11111111111111111011110101011100;
assign LUT_1[2768] = 32'b00000000000000000001101001100101;
assign LUT_1[2769] = 32'b11111111111111111010111011100001;
assign LUT_1[2770] = 32'b11111111111111111101010111110110;
assign LUT_1[2771] = 32'b11111111111111110110101001110010;
assign LUT_1[2772] = 32'b00000000000000001001100010111100;
assign LUT_1[2773] = 32'b00000000000000000010110100111000;
assign LUT_1[2774] = 32'b00000000000000000101010001001101;
assign LUT_1[2775] = 32'b11111111111111111110100011001001;
assign LUT_1[2776] = 32'b00000000000000000000110111011010;
assign LUT_1[2777] = 32'b11111111111111111010001001010110;
assign LUT_1[2778] = 32'b11111111111111111100100101101011;
assign LUT_1[2779] = 32'b11111111111111110101110111100111;
assign LUT_1[2780] = 32'b00000000000000001000110000110001;
assign LUT_1[2781] = 32'b00000000000000000010000010101101;
assign LUT_1[2782] = 32'b00000000000000000100011111000010;
assign LUT_1[2783] = 32'b11111111111111111101110000111110;
assign LUT_1[2784] = 32'b00000000000000000000101001000010;
assign LUT_1[2785] = 32'b11111111111111111001111010111110;
assign LUT_1[2786] = 32'b11111111111111111100010111010011;
assign LUT_1[2787] = 32'b11111111111111110101101001001111;
assign LUT_1[2788] = 32'b00000000000000001000100010011001;
assign LUT_1[2789] = 32'b00000000000000000001110100010101;
assign LUT_1[2790] = 32'b00000000000000000100010000101010;
assign LUT_1[2791] = 32'b11111111111111111101100010100110;
assign LUT_1[2792] = 32'b11111111111111111111110110110111;
assign LUT_1[2793] = 32'b11111111111111111001001000110011;
assign LUT_1[2794] = 32'b11111111111111111011100101001000;
assign LUT_1[2795] = 32'b11111111111111110100110111000100;
assign LUT_1[2796] = 32'b00000000000000000111110000001110;
assign LUT_1[2797] = 32'b00000000000000000001000010001010;
assign LUT_1[2798] = 32'b00000000000000000011011110011111;
assign LUT_1[2799] = 32'b11111111111111111100110000011011;
assign LUT_1[2800] = 32'b00000000000000000010100100100100;
assign LUT_1[2801] = 32'b11111111111111111011110110100000;
assign LUT_1[2802] = 32'b11111111111111111110010010110101;
assign LUT_1[2803] = 32'b11111111111111110111100100110001;
assign LUT_1[2804] = 32'b00000000000000001010011101111011;
assign LUT_1[2805] = 32'b00000000000000000011101111110111;
assign LUT_1[2806] = 32'b00000000000000000110001100001100;
assign LUT_1[2807] = 32'b11111111111111111111011110001000;
assign LUT_1[2808] = 32'b00000000000000000001110010011001;
assign LUT_1[2809] = 32'b11111111111111111011000100010101;
assign LUT_1[2810] = 32'b11111111111111111101100000101010;
assign LUT_1[2811] = 32'b11111111111111110110110010100110;
assign LUT_1[2812] = 32'b00000000000000001001101011110000;
assign LUT_1[2813] = 32'b00000000000000000010111101101100;
assign LUT_1[2814] = 32'b00000000000000000101011010000001;
assign LUT_1[2815] = 32'b11111111111111111110101011111101;
assign LUT_1[2816] = 32'b11111111111111111000100100100100;
assign LUT_1[2817] = 32'b11111111111111110001110110100000;
assign LUT_1[2818] = 32'b11111111111111110100010010110101;
assign LUT_1[2819] = 32'b11111111111111101101100100110001;
assign LUT_1[2820] = 32'b00000000000000000000011101111011;
assign LUT_1[2821] = 32'b11111111111111111001101111110111;
assign LUT_1[2822] = 32'b11111111111111111100001100001100;
assign LUT_1[2823] = 32'b11111111111111110101011110001000;
assign LUT_1[2824] = 32'b11111111111111110111110010011001;
assign LUT_1[2825] = 32'b11111111111111110001000100010101;
assign LUT_1[2826] = 32'b11111111111111110011100000101010;
assign LUT_1[2827] = 32'b11111111111111101100110010100110;
assign LUT_1[2828] = 32'b11111111111111111111101011110000;
assign LUT_1[2829] = 32'b11111111111111111000111101101100;
assign LUT_1[2830] = 32'b11111111111111111011011010000001;
assign LUT_1[2831] = 32'b11111111111111110100101011111101;
assign LUT_1[2832] = 32'b11111111111111111010100000000110;
assign LUT_1[2833] = 32'b11111111111111110011110010000010;
assign LUT_1[2834] = 32'b11111111111111110110001110010111;
assign LUT_1[2835] = 32'b11111111111111101111100000010011;
assign LUT_1[2836] = 32'b00000000000000000010011001011101;
assign LUT_1[2837] = 32'b11111111111111111011101011011001;
assign LUT_1[2838] = 32'b11111111111111111110000111101110;
assign LUT_1[2839] = 32'b11111111111111110111011001101010;
assign LUT_1[2840] = 32'b11111111111111111001101101111011;
assign LUT_1[2841] = 32'b11111111111111110010111111110111;
assign LUT_1[2842] = 32'b11111111111111110101011100001100;
assign LUT_1[2843] = 32'b11111111111111101110101110001000;
assign LUT_1[2844] = 32'b00000000000000000001100111010010;
assign LUT_1[2845] = 32'b11111111111111111010111001001110;
assign LUT_1[2846] = 32'b11111111111111111101010101100011;
assign LUT_1[2847] = 32'b11111111111111110110100111011111;
assign LUT_1[2848] = 32'b11111111111111111001011111100011;
assign LUT_1[2849] = 32'b11111111111111110010110001011111;
assign LUT_1[2850] = 32'b11111111111111110101001101110100;
assign LUT_1[2851] = 32'b11111111111111101110011111110000;
assign LUT_1[2852] = 32'b00000000000000000001011000111010;
assign LUT_1[2853] = 32'b11111111111111111010101010110110;
assign LUT_1[2854] = 32'b11111111111111111101000111001011;
assign LUT_1[2855] = 32'b11111111111111110110011001000111;
assign LUT_1[2856] = 32'b11111111111111111000101101011000;
assign LUT_1[2857] = 32'b11111111111111110001111111010100;
assign LUT_1[2858] = 32'b11111111111111110100011011101001;
assign LUT_1[2859] = 32'b11111111111111101101101101100101;
assign LUT_1[2860] = 32'b00000000000000000000100110101111;
assign LUT_1[2861] = 32'b11111111111111111001111000101011;
assign LUT_1[2862] = 32'b11111111111111111100010101000000;
assign LUT_1[2863] = 32'b11111111111111110101100110111100;
assign LUT_1[2864] = 32'b11111111111111111011011011000101;
assign LUT_1[2865] = 32'b11111111111111110100101101000001;
assign LUT_1[2866] = 32'b11111111111111110111001001010110;
assign LUT_1[2867] = 32'b11111111111111110000011011010010;
assign LUT_1[2868] = 32'b00000000000000000011010100011100;
assign LUT_1[2869] = 32'b11111111111111111100100110011000;
assign LUT_1[2870] = 32'b11111111111111111111000010101101;
assign LUT_1[2871] = 32'b11111111111111111000010100101001;
assign LUT_1[2872] = 32'b11111111111111111010101000111010;
assign LUT_1[2873] = 32'b11111111111111110011111010110110;
assign LUT_1[2874] = 32'b11111111111111110110010111001011;
assign LUT_1[2875] = 32'b11111111111111101111101001000111;
assign LUT_1[2876] = 32'b00000000000000000010100010010001;
assign LUT_1[2877] = 32'b11111111111111111011110100001101;
assign LUT_1[2878] = 32'b11111111111111111110010000100010;
assign LUT_1[2879] = 32'b11111111111111110111100010011110;
assign LUT_1[2880] = 32'b11111111111111111010100010001100;
assign LUT_1[2881] = 32'b11111111111111110011110100001000;
assign LUT_1[2882] = 32'b11111111111111110110010000011101;
assign LUT_1[2883] = 32'b11111111111111101111100010011001;
assign LUT_1[2884] = 32'b00000000000000000010011011100011;
assign LUT_1[2885] = 32'b11111111111111111011101101011111;
assign LUT_1[2886] = 32'b11111111111111111110001001110100;
assign LUT_1[2887] = 32'b11111111111111110111011011110000;
assign LUT_1[2888] = 32'b11111111111111111001110000000001;
assign LUT_1[2889] = 32'b11111111111111110011000001111101;
assign LUT_1[2890] = 32'b11111111111111110101011110010010;
assign LUT_1[2891] = 32'b11111111111111101110110000001110;
assign LUT_1[2892] = 32'b00000000000000000001101001011000;
assign LUT_1[2893] = 32'b11111111111111111010111011010100;
assign LUT_1[2894] = 32'b11111111111111111101010111101001;
assign LUT_1[2895] = 32'b11111111111111110110101001100101;
assign LUT_1[2896] = 32'b11111111111111111100011101101110;
assign LUT_1[2897] = 32'b11111111111111110101101111101010;
assign LUT_1[2898] = 32'b11111111111111111000001011111111;
assign LUT_1[2899] = 32'b11111111111111110001011101111011;
assign LUT_1[2900] = 32'b00000000000000000100010111000101;
assign LUT_1[2901] = 32'b11111111111111111101101001000001;
assign LUT_1[2902] = 32'b00000000000000000000000101010110;
assign LUT_1[2903] = 32'b11111111111111111001010111010010;
assign LUT_1[2904] = 32'b11111111111111111011101011100011;
assign LUT_1[2905] = 32'b11111111111111110100111101011111;
assign LUT_1[2906] = 32'b11111111111111110111011001110100;
assign LUT_1[2907] = 32'b11111111111111110000101011110000;
assign LUT_1[2908] = 32'b00000000000000000011100100111010;
assign LUT_1[2909] = 32'b11111111111111111100110110110110;
assign LUT_1[2910] = 32'b11111111111111111111010011001011;
assign LUT_1[2911] = 32'b11111111111111111000100101000111;
assign LUT_1[2912] = 32'b11111111111111111011011101001011;
assign LUT_1[2913] = 32'b11111111111111110100101111000111;
assign LUT_1[2914] = 32'b11111111111111110111001011011100;
assign LUT_1[2915] = 32'b11111111111111110000011101011000;
assign LUT_1[2916] = 32'b00000000000000000011010110100010;
assign LUT_1[2917] = 32'b11111111111111111100101000011110;
assign LUT_1[2918] = 32'b11111111111111111111000100110011;
assign LUT_1[2919] = 32'b11111111111111111000010110101111;
assign LUT_1[2920] = 32'b11111111111111111010101011000000;
assign LUT_1[2921] = 32'b11111111111111110011111100111100;
assign LUT_1[2922] = 32'b11111111111111110110011001010001;
assign LUT_1[2923] = 32'b11111111111111101111101011001101;
assign LUT_1[2924] = 32'b00000000000000000010100100010111;
assign LUT_1[2925] = 32'b11111111111111111011110110010011;
assign LUT_1[2926] = 32'b11111111111111111110010010101000;
assign LUT_1[2927] = 32'b11111111111111110111100100100100;
assign LUT_1[2928] = 32'b11111111111111111101011000101101;
assign LUT_1[2929] = 32'b11111111111111110110101010101001;
assign LUT_1[2930] = 32'b11111111111111111001000110111110;
assign LUT_1[2931] = 32'b11111111111111110010011000111010;
assign LUT_1[2932] = 32'b00000000000000000101010010000100;
assign LUT_1[2933] = 32'b11111111111111111110100100000000;
assign LUT_1[2934] = 32'b00000000000000000001000000010101;
assign LUT_1[2935] = 32'b11111111111111111010010010010001;
assign LUT_1[2936] = 32'b11111111111111111100100110100010;
assign LUT_1[2937] = 32'b11111111111111110101111000011110;
assign LUT_1[2938] = 32'b11111111111111111000010100110011;
assign LUT_1[2939] = 32'b11111111111111110001100110101111;
assign LUT_1[2940] = 32'b00000000000000000100011111111001;
assign LUT_1[2941] = 32'b11111111111111111101110001110101;
assign LUT_1[2942] = 32'b00000000000000000000001110001010;
assign LUT_1[2943] = 32'b11111111111111111001100000000110;
assign LUT_1[2944] = 32'b11111111111111111011100100100111;
assign LUT_1[2945] = 32'b11111111111111110100110110100011;
assign LUT_1[2946] = 32'b11111111111111110111010010111000;
assign LUT_1[2947] = 32'b11111111111111110000100100110100;
assign LUT_1[2948] = 32'b00000000000000000011011101111110;
assign LUT_1[2949] = 32'b11111111111111111100101111111010;
assign LUT_1[2950] = 32'b11111111111111111111001100001111;
assign LUT_1[2951] = 32'b11111111111111111000011110001011;
assign LUT_1[2952] = 32'b11111111111111111010110010011100;
assign LUT_1[2953] = 32'b11111111111111110100000100011000;
assign LUT_1[2954] = 32'b11111111111111110110100000101101;
assign LUT_1[2955] = 32'b11111111111111101111110010101001;
assign LUT_1[2956] = 32'b00000000000000000010101011110011;
assign LUT_1[2957] = 32'b11111111111111111011111101101111;
assign LUT_1[2958] = 32'b11111111111111111110011010000100;
assign LUT_1[2959] = 32'b11111111111111110111101100000000;
assign LUT_1[2960] = 32'b11111111111111111101100000001001;
assign LUT_1[2961] = 32'b11111111111111110110110010000101;
assign LUT_1[2962] = 32'b11111111111111111001001110011010;
assign LUT_1[2963] = 32'b11111111111111110010100000010110;
assign LUT_1[2964] = 32'b00000000000000000101011001100000;
assign LUT_1[2965] = 32'b11111111111111111110101011011100;
assign LUT_1[2966] = 32'b00000000000000000001000111110001;
assign LUT_1[2967] = 32'b11111111111111111010011001101101;
assign LUT_1[2968] = 32'b11111111111111111100101101111110;
assign LUT_1[2969] = 32'b11111111111111110101111111111010;
assign LUT_1[2970] = 32'b11111111111111111000011100001111;
assign LUT_1[2971] = 32'b11111111111111110001101110001011;
assign LUT_1[2972] = 32'b00000000000000000100100111010101;
assign LUT_1[2973] = 32'b11111111111111111101111001010001;
assign LUT_1[2974] = 32'b00000000000000000000010101100110;
assign LUT_1[2975] = 32'b11111111111111111001100111100010;
assign LUT_1[2976] = 32'b11111111111111111100011111100110;
assign LUT_1[2977] = 32'b11111111111111110101110001100010;
assign LUT_1[2978] = 32'b11111111111111111000001101110111;
assign LUT_1[2979] = 32'b11111111111111110001011111110011;
assign LUT_1[2980] = 32'b00000000000000000100011000111101;
assign LUT_1[2981] = 32'b11111111111111111101101010111001;
assign LUT_1[2982] = 32'b00000000000000000000000111001110;
assign LUT_1[2983] = 32'b11111111111111111001011001001010;
assign LUT_1[2984] = 32'b11111111111111111011101101011011;
assign LUT_1[2985] = 32'b11111111111111110100111111010111;
assign LUT_1[2986] = 32'b11111111111111110111011011101100;
assign LUT_1[2987] = 32'b11111111111111110000101101101000;
assign LUT_1[2988] = 32'b00000000000000000011100110110010;
assign LUT_1[2989] = 32'b11111111111111111100111000101110;
assign LUT_1[2990] = 32'b11111111111111111111010101000011;
assign LUT_1[2991] = 32'b11111111111111111000100110111111;
assign LUT_1[2992] = 32'b11111111111111111110011011001000;
assign LUT_1[2993] = 32'b11111111111111110111101101000100;
assign LUT_1[2994] = 32'b11111111111111111010001001011001;
assign LUT_1[2995] = 32'b11111111111111110011011011010101;
assign LUT_1[2996] = 32'b00000000000000000110010100011111;
assign LUT_1[2997] = 32'b11111111111111111111100110011011;
assign LUT_1[2998] = 32'b00000000000000000010000010110000;
assign LUT_1[2999] = 32'b11111111111111111011010100101100;
assign LUT_1[3000] = 32'b11111111111111111101101000111101;
assign LUT_1[3001] = 32'b11111111111111110110111010111001;
assign LUT_1[3002] = 32'b11111111111111111001010111001110;
assign LUT_1[3003] = 32'b11111111111111110010101001001010;
assign LUT_1[3004] = 32'b00000000000000000101100010010100;
assign LUT_1[3005] = 32'b11111111111111111110110100010000;
assign LUT_1[3006] = 32'b00000000000000000001010000100101;
assign LUT_1[3007] = 32'b11111111111111111010100010100001;
assign LUT_1[3008] = 32'b11111111111111111101100010001111;
assign LUT_1[3009] = 32'b11111111111111110110110100001011;
assign LUT_1[3010] = 32'b11111111111111111001010000100000;
assign LUT_1[3011] = 32'b11111111111111110010100010011100;
assign LUT_1[3012] = 32'b00000000000000000101011011100110;
assign LUT_1[3013] = 32'b11111111111111111110101101100010;
assign LUT_1[3014] = 32'b00000000000000000001001001110111;
assign LUT_1[3015] = 32'b11111111111111111010011011110011;
assign LUT_1[3016] = 32'b11111111111111111100110000000100;
assign LUT_1[3017] = 32'b11111111111111110110000010000000;
assign LUT_1[3018] = 32'b11111111111111111000011110010101;
assign LUT_1[3019] = 32'b11111111111111110001110000010001;
assign LUT_1[3020] = 32'b00000000000000000100101001011011;
assign LUT_1[3021] = 32'b11111111111111111101111011010111;
assign LUT_1[3022] = 32'b00000000000000000000010111101100;
assign LUT_1[3023] = 32'b11111111111111111001101001101000;
assign LUT_1[3024] = 32'b11111111111111111111011101110001;
assign LUT_1[3025] = 32'b11111111111111111000101111101101;
assign LUT_1[3026] = 32'b11111111111111111011001100000010;
assign LUT_1[3027] = 32'b11111111111111110100011101111110;
assign LUT_1[3028] = 32'b00000000000000000111010111001000;
assign LUT_1[3029] = 32'b00000000000000000000101001000100;
assign LUT_1[3030] = 32'b00000000000000000011000101011001;
assign LUT_1[3031] = 32'b11111111111111111100010111010101;
assign LUT_1[3032] = 32'b11111111111111111110101011100110;
assign LUT_1[3033] = 32'b11111111111111110111111101100010;
assign LUT_1[3034] = 32'b11111111111111111010011001110111;
assign LUT_1[3035] = 32'b11111111111111110011101011110011;
assign LUT_1[3036] = 32'b00000000000000000110100100111101;
assign LUT_1[3037] = 32'b11111111111111111111110110111001;
assign LUT_1[3038] = 32'b00000000000000000010010011001110;
assign LUT_1[3039] = 32'b11111111111111111011100101001010;
assign LUT_1[3040] = 32'b11111111111111111110011101001110;
assign LUT_1[3041] = 32'b11111111111111110111101111001010;
assign LUT_1[3042] = 32'b11111111111111111010001011011111;
assign LUT_1[3043] = 32'b11111111111111110011011101011011;
assign LUT_1[3044] = 32'b00000000000000000110010110100101;
assign LUT_1[3045] = 32'b11111111111111111111101000100001;
assign LUT_1[3046] = 32'b00000000000000000010000100110110;
assign LUT_1[3047] = 32'b11111111111111111011010110110010;
assign LUT_1[3048] = 32'b11111111111111111101101011000011;
assign LUT_1[3049] = 32'b11111111111111110110111100111111;
assign LUT_1[3050] = 32'b11111111111111111001011001010100;
assign LUT_1[3051] = 32'b11111111111111110010101011010000;
assign LUT_1[3052] = 32'b00000000000000000101100100011010;
assign LUT_1[3053] = 32'b11111111111111111110110110010110;
assign LUT_1[3054] = 32'b00000000000000000001010010101011;
assign LUT_1[3055] = 32'b11111111111111111010100100100111;
assign LUT_1[3056] = 32'b00000000000000000000011000110000;
assign LUT_1[3057] = 32'b11111111111111111001101010101100;
assign LUT_1[3058] = 32'b11111111111111111100000111000001;
assign LUT_1[3059] = 32'b11111111111111110101011000111101;
assign LUT_1[3060] = 32'b00000000000000001000010010000111;
assign LUT_1[3061] = 32'b00000000000000000001100100000011;
assign LUT_1[3062] = 32'b00000000000000000100000000011000;
assign LUT_1[3063] = 32'b11111111111111111101010010010100;
assign LUT_1[3064] = 32'b11111111111111111111100110100101;
assign LUT_1[3065] = 32'b11111111111111111000111000100001;
assign LUT_1[3066] = 32'b11111111111111111011010100110110;
assign LUT_1[3067] = 32'b11111111111111110100100110110010;
assign LUT_1[3068] = 32'b00000000000000000111011111111100;
assign LUT_1[3069] = 32'b00000000000000000000110001111000;
assign LUT_1[3070] = 32'b00000000000000000011001110001101;
assign LUT_1[3071] = 32'b11111111111111111100100000001001;
assign LUT_1[3072] = 32'b00000000000000000111011000101011;
assign LUT_1[3073] = 32'b00000000000000000000101010100111;
assign LUT_1[3074] = 32'b00000000000000000011000110111100;
assign LUT_1[3075] = 32'b11111111111111111100011000111000;
assign LUT_1[3076] = 32'b00000000000000001111010010000010;
assign LUT_1[3077] = 32'b00000000000000001000100011111110;
assign LUT_1[3078] = 32'b00000000000000001011000000010011;
assign LUT_1[3079] = 32'b00000000000000000100010010001111;
assign LUT_1[3080] = 32'b00000000000000000110100110100000;
assign LUT_1[3081] = 32'b11111111111111111111111000011100;
assign LUT_1[3082] = 32'b00000000000000000010010100110001;
assign LUT_1[3083] = 32'b11111111111111111011100110101101;
assign LUT_1[3084] = 32'b00000000000000001110011111110111;
assign LUT_1[3085] = 32'b00000000000000000111110001110011;
assign LUT_1[3086] = 32'b00000000000000001010001110001000;
assign LUT_1[3087] = 32'b00000000000000000011100000000100;
assign LUT_1[3088] = 32'b00000000000000001001010100001101;
assign LUT_1[3089] = 32'b00000000000000000010100110001001;
assign LUT_1[3090] = 32'b00000000000000000101000010011110;
assign LUT_1[3091] = 32'b11111111111111111110010100011010;
assign LUT_1[3092] = 32'b00000000000000010001001101100100;
assign LUT_1[3093] = 32'b00000000000000001010011111100000;
assign LUT_1[3094] = 32'b00000000000000001100111011110101;
assign LUT_1[3095] = 32'b00000000000000000110001101110001;
assign LUT_1[3096] = 32'b00000000000000001000100010000010;
assign LUT_1[3097] = 32'b00000000000000000001110011111110;
assign LUT_1[3098] = 32'b00000000000000000100010000010011;
assign LUT_1[3099] = 32'b11111111111111111101100010001111;
assign LUT_1[3100] = 32'b00000000000000010000011011011001;
assign LUT_1[3101] = 32'b00000000000000001001101101010101;
assign LUT_1[3102] = 32'b00000000000000001100001001101010;
assign LUT_1[3103] = 32'b00000000000000000101011011100110;
assign LUT_1[3104] = 32'b00000000000000001000010011101010;
assign LUT_1[3105] = 32'b00000000000000000001100101100110;
assign LUT_1[3106] = 32'b00000000000000000100000001111011;
assign LUT_1[3107] = 32'b11111111111111111101010011110111;
assign LUT_1[3108] = 32'b00000000000000010000001101000001;
assign LUT_1[3109] = 32'b00000000000000001001011110111101;
assign LUT_1[3110] = 32'b00000000000000001011111011010010;
assign LUT_1[3111] = 32'b00000000000000000101001101001110;
assign LUT_1[3112] = 32'b00000000000000000111100001011111;
assign LUT_1[3113] = 32'b00000000000000000000110011011011;
assign LUT_1[3114] = 32'b00000000000000000011001111110000;
assign LUT_1[3115] = 32'b11111111111111111100100001101100;
assign LUT_1[3116] = 32'b00000000000000001111011010110110;
assign LUT_1[3117] = 32'b00000000000000001000101100110010;
assign LUT_1[3118] = 32'b00000000000000001011001001000111;
assign LUT_1[3119] = 32'b00000000000000000100011011000011;
assign LUT_1[3120] = 32'b00000000000000001010001111001100;
assign LUT_1[3121] = 32'b00000000000000000011100001001000;
assign LUT_1[3122] = 32'b00000000000000000101111101011101;
assign LUT_1[3123] = 32'b11111111111111111111001111011001;
assign LUT_1[3124] = 32'b00000000000000010010001000100011;
assign LUT_1[3125] = 32'b00000000000000001011011010011111;
assign LUT_1[3126] = 32'b00000000000000001101110110110100;
assign LUT_1[3127] = 32'b00000000000000000111001000110000;
assign LUT_1[3128] = 32'b00000000000000001001011101000001;
assign LUT_1[3129] = 32'b00000000000000000010101110111101;
assign LUT_1[3130] = 32'b00000000000000000101001011010010;
assign LUT_1[3131] = 32'b11111111111111111110011101001110;
assign LUT_1[3132] = 32'b00000000000000010001010110011000;
assign LUT_1[3133] = 32'b00000000000000001010101000010100;
assign LUT_1[3134] = 32'b00000000000000001101000100101001;
assign LUT_1[3135] = 32'b00000000000000000110010110100101;
assign LUT_1[3136] = 32'b00000000000000001001010110010011;
assign LUT_1[3137] = 32'b00000000000000000010101000001111;
assign LUT_1[3138] = 32'b00000000000000000101000100100100;
assign LUT_1[3139] = 32'b11111111111111111110010110100000;
assign LUT_1[3140] = 32'b00000000000000010001001111101010;
assign LUT_1[3141] = 32'b00000000000000001010100001100110;
assign LUT_1[3142] = 32'b00000000000000001100111101111011;
assign LUT_1[3143] = 32'b00000000000000000110001111110111;
assign LUT_1[3144] = 32'b00000000000000001000100100001000;
assign LUT_1[3145] = 32'b00000000000000000001110110000100;
assign LUT_1[3146] = 32'b00000000000000000100010010011001;
assign LUT_1[3147] = 32'b11111111111111111101100100010101;
assign LUT_1[3148] = 32'b00000000000000010000011101011111;
assign LUT_1[3149] = 32'b00000000000000001001101111011011;
assign LUT_1[3150] = 32'b00000000000000001100001011110000;
assign LUT_1[3151] = 32'b00000000000000000101011101101100;
assign LUT_1[3152] = 32'b00000000000000001011010001110101;
assign LUT_1[3153] = 32'b00000000000000000100100011110001;
assign LUT_1[3154] = 32'b00000000000000000111000000000110;
assign LUT_1[3155] = 32'b00000000000000000000010010000010;
assign LUT_1[3156] = 32'b00000000000000010011001011001100;
assign LUT_1[3157] = 32'b00000000000000001100011101001000;
assign LUT_1[3158] = 32'b00000000000000001110111001011101;
assign LUT_1[3159] = 32'b00000000000000001000001011011001;
assign LUT_1[3160] = 32'b00000000000000001010011111101010;
assign LUT_1[3161] = 32'b00000000000000000011110001100110;
assign LUT_1[3162] = 32'b00000000000000000110001101111011;
assign LUT_1[3163] = 32'b11111111111111111111011111110111;
assign LUT_1[3164] = 32'b00000000000000010010011001000001;
assign LUT_1[3165] = 32'b00000000000000001011101010111101;
assign LUT_1[3166] = 32'b00000000000000001110000111010010;
assign LUT_1[3167] = 32'b00000000000000000111011001001110;
assign LUT_1[3168] = 32'b00000000000000001010010001010010;
assign LUT_1[3169] = 32'b00000000000000000011100011001110;
assign LUT_1[3170] = 32'b00000000000000000101111111100011;
assign LUT_1[3171] = 32'b11111111111111111111010001011111;
assign LUT_1[3172] = 32'b00000000000000010010001010101001;
assign LUT_1[3173] = 32'b00000000000000001011011100100101;
assign LUT_1[3174] = 32'b00000000000000001101111000111010;
assign LUT_1[3175] = 32'b00000000000000000111001010110110;
assign LUT_1[3176] = 32'b00000000000000001001011111000111;
assign LUT_1[3177] = 32'b00000000000000000010110001000011;
assign LUT_1[3178] = 32'b00000000000000000101001101011000;
assign LUT_1[3179] = 32'b11111111111111111110011111010100;
assign LUT_1[3180] = 32'b00000000000000010001011000011110;
assign LUT_1[3181] = 32'b00000000000000001010101010011010;
assign LUT_1[3182] = 32'b00000000000000001101000110101111;
assign LUT_1[3183] = 32'b00000000000000000110011000101011;
assign LUT_1[3184] = 32'b00000000000000001100001100110100;
assign LUT_1[3185] = 32'b00000000000000000101011110110000;
assign LUT_1[3186] = 32'b00000000000000000111111011000101;
assign LUT_1[3187] = 32'b00000000000000000001001101000001;
assign LUT_1[3188] = 32'b00000000000000010100000110001011;
assign LUT_1[3189] = 32'b00000000000000001101011000000111;
assign LUT_1[3190] = 32'b00000000000000001111110100011100;
assign LUT_1[3191] = 32'b00000000000000001001000110011000;
assign LUT_1[3192] = 32'b00000000000000001011011010101001;
assign LUT_1[3193] = 32'b00000000000000000100101100100101;
assign LUT_1[3194] = 32'b00000000000000000111001000111010;
assign LUT_1[3195] = 32'b00000000000000000000011010110110;
assign LUT_1[3196] = 32'b00000000000000010011010100000000;
assign LUT_1[3197] = 32'b00000000000000001100100101111100;
assign LUT_1[3198] = 32'b00000000000000001111000010010001;
assign LUT_1[3199] = 32'b00000000000000001000010100001101;
assign LUT_1[3200] = 32'b00000000000000001010011000101110;
assign LUT_1[3201] = 32'b00000000000000000011101010101010;
assign LUT_1[3202] = 32'b00000000000000000110000110111111;
assign LUT_1[3203] = 32'b11111111111111111111011000111011;
assign LUT_1[3204] = 32'b00000000000000010010010010000101;
assign LUT_1[3205] = 32'b00000000000000001011100100000001;
assign LUT_1[3206] = 32'b00000000000000001110000000010110;
assign LUT_1[3207] = 32'b00000000000000000111010010010010;
assign LUT_1[3208] = 32'b00000000000000001001100110100011;
assign LUT_1[3209] = 32'b00000000000000000010111000011111;
assign LUT_1[3210] = 32'b00000000000000000101010100110100;
assign LUT_1[3211] = 32'b11111111111111111110100110110000;
assign LUT_1[3212] = 32'b00000000000000010001011111111010;
assign LUT_1[3213] = 32'b00000000000000001010110001110110;
assign LUT_1[3214] = 32'b00000000000000001101001110001011;
assign LUT_1[3215] = 32'b00000000000000000110100000000111;
assign LUT_1[3216] = 32'b00000000000000001100010100010000;
assign LUT_1[3217] = 32'b00000000000000000101100110001100;
assign LUT_1[3218] = 32'b00000000000000001000000010100001;
assign LUT_1[3219] = 32'b00000000000000000001010100011101;
assign LUT_1[3220] = 32'b00000000000000010100001101100111;
assign LUT_1[3221] = 32'b00000000000000001101011111100011;
assign LUT_1[3222] = 32'b00000000000000001111111011111000;
assign LUT_1[3223] = 32'b00000000000000001001001101110100;
assign LUT_1[3224] = 32'b00000000000000001011100010000101;
assign LUT_1[3225] = 32'b00000000000000000100110100000001;
assign LUT_1[3226] = 32'b00000000000000000111010000010110;
assign LUT_1[3227] = 32'b00000000000000000000100010010010;
assign LUT_1[3228] = 32'b00000000000000010011011011011100;
assign LUT_1[3229] = 32'b00000000000000001100101101011000;
assign LUT_1[3230] = 32'b00000000000000001111001001101101;
assign LUT_1[3231] = 32'b00000000000000001000011011101001;
assign LUT_1[3232] = 32'b00000000000000001011010011101101;
assign LUT_1[3233] = 32'b00000000000000000100100101101001;
assign LUT_1[3234] = 32'b00000000000000000111000001111110;
assign LUT_1[3235] = 32'b00000000000000000000010011111010;
assign LUT_1[3236] = 32'b00000000000000010011001101000100;
assign LUT_1[3237] = 32'b00000000000000001100011111000000;
assign LUT_1[3238] = 32'b00000000000000001110111011010101;
assign LUT_1[3239] = 32'b00000000000000001000001101010001;
assign LUT_1[3240] = 32'b00000000000000001010100001100010;
assign LUT_1[3241] = 32'b00000000000000000011110011011110;
assign LUT_1[3242] = 32'b00000000000000000110001111110011;
assign LUT_1[3243] = 32'b11111111111111111111100001101111;
assign LUT_1[3244] = 32'b00000000000000010010011010111001;
assign LUT_1[3245] = 32'b00000000000000001011101100110101;
assign LUT_1[3246] = 32'b00000000000000001110001001001010;
assign LUT_1[3247] = 32'b00000000000000000111011011000110;
assign LUT_1[3248] = 32'b00000000000000001101001111001111;
assign LUT_1[3249] = 32'b00000000000000000110100001001011;
assign LUT_1[3250] = 32'b00000000000000001000111101100000;
assign LUT_1[3251] = 32'b00000000000000000010001111011100;
assign LUT_1[3252] = 32'b00000000000000010101001000100110;
assign LUT_1[3253] = 32'b00000000000000001110011010100010;
assign LUT_1[3254] = 32'b00000000000000010000110110110111;
assign LUT_1[3255] = 32'b00000000000000001010001000110011;
assign LUT_1[3256] = 32'b00000000000000001100011101000100;
assign LUT_1[3257] = 32'b00000000000000000101101111000000;
assign LUT_1[3258] = 32'b00000000000000001000001011010101;
assign LUT_1[3259] = 32'b00000000000000000001011101010001;
assign LUT_1[3260] = 32'b00000000000000010100010110011011;
assign LUT_1[3261] = 32'b00000000000000001101101000010111;
assign LUT_1[3262] = 32'b00000000000000010000000100101100;
assign LUT_1[3263] = 32'b00000000000000001001010110101000;
assign LUT_1[3264] = 32'b00000000000000001100010110010110;
assign LUT_1[3265] = 32'b00000000000000000101101000010010;
assign LUT_1[3266] = 32'b00000000000000001000000100100111;
assign LUT_1[3267] = 32'b00000000000000000001010110100011;
assign LUT_1[3268] = 32'b00000000000000010100001111101101;
assign LUT_1[3269] = 32'b00000000000000001101100001101001;
assign LUT_1[3270] = 32'b00000000000000001111111101111110;
assign LUT_1[3271] = 32'b00000000000000001001001111111010;
assign LUT_1[3272] = 32'b00000000000000001011100100001011;
assign LUT_1[3273] = 32'b00000000000000000100110110000111;
assign LUT_1[3274] = 32'b00000000000000000111010010011100;
assign LUT_1[3275] = 32'b00000000000000000000100100011000;
assign LUT_1[3276] = 32'b00000000000000010011011101100010;
assign LUT_1[3277] = 32'b00000000000000001100101111011110;
assign LUT_1[3278] = 32'b00000000000000001111001011110011;
assign LUT_1[3279] = 32'b00000000000000001000011101101111;
assign LUT_1[3280] = 32'b00000000000000001110010001111000;
assign LUT_1[3281] = 32'b00000000000000000111100011110100;
assign LUT_1[3282] = 32'b00000000000000001010000000001001;
assign LUT_1[3283] = 32'b00000000000000000011010010000101;
assign LUT_1[3284] = 32'b00000000000000010110001011001111;
assign LUT_1[3285] = 32'b00000000000000001111011101001011;
assign LUT_1[3286] = 32'b00000000000000010001111001100000;
assign LUT_1[3287] = 32'b00000000000000001011001011011100;
assign LUT_1[3288] = 32'b00000000000000001101011111101101;
assign LUT_1[3289] = 32'b00000000000000000110110001101001;
assign LUT_1[3290] = 32'b00000000000000001001001101111110;
assign LUT_1[3291] = 32'b00000000000000000010011111111010;
assign LUT_1[3292] = 32'b00000000000000010101011001000100;
assign LUT_1[3293] = 32'b00000000000000001110101011000000;
assign LUT_1[3294] = 32'b00000000000000010001000111010101;
assign LUT_1[3295] = 32'b00000000000000001010011001010001;
assign LUT_1[3296] = 32'b00000000000000001101010001010101;
assign LUT_1[3297] = 32'b00000000000000000110100011010001;
assign LUT_1[3298] = 32'b00000000000000001000111111100110;
assign LUT_1[3299] = 32'b00000000000000000010010001100010;
assign LUT_1[3300] = 32'b00000000000000010101001010101100;
assign LUT_1[3301] = 32'b00000000000000001110011100101000;
assign LUT_1[3302] = 32'b00000000000000010000111000111101;
assign LUT_1[3303] = 32'b00000000000000001010001010111001;
assign LUT_1[3304] = 32'b00000000000000001100011111001010;
assign LUT_1[3305] = 32'b00000000000000000101110001000110;
assign LUT_1[3306] = 32'b00000000000000001000001101011011;
assign LUT_1[3307] = 32'b00000000000000000001011111010111;
assign LUT_1[3308] = 32'b00000000000000010100011000100001;
assign LUT_1[3309] = 32'b00000000000000001101101010011101;
assign LUT_1[3310] = 32'b00000000000000010000000110110010;
assign LUT_1[3311] = 32'b00000000000000001001011000101110;
assign LUT_1[3312] = 32'b00000000000000001111001100110111;
assign LUT_1[3313] = 32'b00000000000000001000011110110011;
assign LUT_1[3314] = 32'b00000000000000001010111011001000;
assign LUT_1[3315] = 32'b00000000000000000100001101000100;
assign LUT_1[3316] = 32'b00000000000000010111000110001110;
assign LUT_1[3317] = 32'b00000000000000010000011000001010;
assign LUT_1[3318] = 32'b00000000000000010010110100011111;
assign LUT_1[3319] = 32'b00000000000000001100000110011011;
assign LUT_1[3320] = 32'b00000000000000001110011010101100;
assign LUT_1[3321] = 32'b00000000000000000111101100101000;
assign LUT_1[3322] = 32'b00000000000000001010001000111101;
assign LUT_1[3323] = 32'b00000000000000000011011010111001;
assign LUT_1[3324] = 32'b00000000000000010110010100000011;
assign LUT_1[3325] = 32'b00000000000000001111100101111111;
assign LUT_1[3326] = 32'b00000000000000010010000010010100;
assign LUT_1[3327] = 32'b00000000000000001011010100010000;
assign LUT_1[3328] = 32'b00000000000000000101001100110111;
assign LUT_1[3329] = 32'b11111111111111111110011110110011;
assign LUT_1[3330] = 32'b00000000000000000000111011001000;
assign LUT_1[3331] = 32'b11111111111111111010001101000100;
assign LUT_1[3332] = 32'b00000000000000001101000110001110;
assign LUT_1[3333] = 32'b00000000000000000110011000001010;
assign LUT_1[3334] = 32'b00000000000000001000110100011111;
assign LUT_1[3335] = 32'b00000000000000000010000110011011;
assign LUT_1[3336] = 32'b00000000000000000100011010101100;
assign LUT_1[3337] = 32'b11111111111111111101101100101000;
assign LUT_1[3338] = 32'b00000000000000000000001000111101;
assign LUT_1[3339] = 32'b11111111111111111001011010111001;
assign LUT_1[3340] = 32'b00000000000000001100010100000011;
assign LUT_1[3341] = 32'b00000000000000000101100101111111;
assign LUT_1[3342] = 32'b00000000000000001000000010010100;
assign LUT_1[3343] = 32'b00000000000000000001010100010000;
assign LUT_1[3344] = 32'b00000000000000000111001000011001;
assign LUT_1[3345] = 32'b00000000000000000000011010010101;
assign LUT_1[3346] = 32'b00000000000000000010110110101010;
assign LUT_1[3347] = 32'b11111111111111111100001000100110;
assign LUT_1[3348] = 32'b00000000000000001111000001110000;
assign LUT_1[3349] = 32'b00000000000000001000010011101100;
assign LUT_1[3350] = 32'b00000000000000001010110000000001;
assign LUT_1[3351] = 32'b00000000000000000100000001111101;
assign LUT_1[3352] = 32'b00000000000000000110010110001110;
assign LUT_1[3353] = 32'b11111111111111111111101000001010;
assign LUT_1[3354] = 32'b00000000000000000010000100011111;
assign LUT_1[3355] = 32'b11111111111111111011010110011011;
assign LUT_1[3356] = 32'b00000000000000001110001111100101;
assign LUT_1[3357] = 32'b00000000000000000111100001100001;
assign LUT_1[3358] = 32'b00000000000000001001111101110110;
assign LUT_1[3359] = 32'b00000000000000000011001111110010;
assign LUT_1[3360] = 32'b00000000000000000110000111110110;
assign LUT_1[3361] = 32'b11111111111111111111011001110010;
assign LUT_1[3362] = 32'b00000000000000000001110110000111;
assign LUT_1[3363] = 32'b11111111111111111011001000000011;
assign LUT_1[3364] = 32'b00000000000000001110000001001101;
assign LUT_1[3365] = 32'b00000000000000000111010011001001;
assign LUT_1[3366] = 32'b00000000000000001001101111011110;
assign LUT_1[3367] = 32'b00000000000000000011000001011010;
assign LUT_1[3368] = 32'b00000000000000000101010101101011;
assign LUT_1[3369] = 32'b11111111111111111110100111100111;
assign LUT_1[3370] = 32'b00000000000000000001000011111100;
assign LUT_1[3371] = 32'b11111111111111111010010101111000;
assign LUT_1[3372] = 32'b00000000000000001101001111000010;
assign LUT_1[3373] = 32'b00000000000000000110100000111110;
assign LUT_1[3374] = 32'b00000000000000001000111101010011;
assign LUT_1[3375] = 32'b00000000000000000010001111001111;
assign LUT_1[3376] = 32'b00000000000000001000000011011000;
assign LUT_1[3377] = 32'b00000000000000000001010101010100;
assign LUT_1[3378] = 32'b00000000000000000011110001101001;
assign LUT_1[3379] = 32'b11111111111111111101000011100101;
assign LUT_1[3380] = 32'b00000000000000001111111100101111;
assign LUT_1[3381] = 32'b00000000000000001001001110101011;
assign LUT_1[3382] = 32'b00000000000000001011101011000000;
assign LUT_1[3383] = 32'b00000000000000000100111100111100;
assign LUT_1[3384] = 32'b00000000000000000111010001001101;
assign LUT_1[3385] = 32'b00000000000000000000100011001001;
assign LUT_1[3386] = 32'b00000000000000000010111111011110;
assign LUT_1[3387] = 32'b11111111111111111100010001011010;
assign LUT_1[3388] = 32'b00000000000000001111001010100100;
assign LUT_1[3389] = 32'b00000000000000001000011100100000;
assign LUT_1[3390] = 32'b00000000000000001010111000110101;
assign LUT_1[3391] = 32'b00000000000000000100001010110001;
assign LUT_1[3392] = 32'b00000000000000000111001010011111;
assign LUT_1[3393] = 32'b00000000000000000000011100011011;
assign LUT_1[3394] = 32'b00000000000000000010111000110000;
assign LUT_1[3395] = 32'b11111111111111111100001010101100;
assign LUT_1[3396] = 32'b00000000000000001111000011110110;
assign LUT_1[3397] = 32'b00000000000000001000010101110010;
assign LUT_1[3398] = 32'b00000000000000001010110010000111;
assign LUT_1[3399] = 32'b00000000000000000100000100000011;
assign LUT_1[3400] = 32'b00000000000000000110011000010100;
assign LUT_1[3401] = 32'b11111111111111111111101010010000;
assign LUT_1[3402] = 32'b00000000000000000010000110100101;
assign LUT_1[3403] = 32'b11111111111111111011011000100001;
assign LUT_1[3404] = 32'b00000000000000001110010001101011;
assign LUT_1[3405] = 32'b00000000000000000111100011100111;
assign LUT_1[3406] = 32'b00000000000000001001111111111100;
assign LUT_1[3407] = 32'b00000000000000000011010001111000;
assign LUT_1[3408] = 32'b00000000000000001001000110000001;
assign LUT_1[3409] = 32'b00000000000000000010010111111101;
assign LUT_1[3410] = 32'b00000000000000000100110100010010;
assign LUT_1[3411] = 32'b11111111111111111110000110001110;
assign LUT_1[3412] = 32'b00000000000000010000111111011000;
assign LUT_1[3413] = 32'b00000000000000001010010001010100;
assign LUT_1[3414] = 32'b00000000000000001100101101101001;
assign LUT_1[3415] = 32'b00000000000000000101111111100101;
assign LUT_1[3416] = 32'b00000000000000001000010011110110;
assign LUT_1[3417] = 32'b00000000000000000001100101110010;
assign LUT_1[3418] = 32'b00000000000000000100000010000111;
assign LUT_1[3419] = 32'b11111111111111111101010100000011;
assign LUT_1[3420] = 32'b00000000000000010000001101001101;
assign LUT_1[3421] = 32'b00000000000000001001011111001001;
assign LUT_1[3422] = 32'b00000000000000001011111011011110;
assign LUT_1[3423] = 32'b00000000000000000101001101011010;
assign LUT_1[3424] = 32'b00000000000000001000000101011110;
assign LUT_1[3425] = 32'b00000000000000000001010111011010;
assign LUT_1[3426] = 32'b00000000000000000011110011101111;
assign LUT_1[3427] = 32'b11111111111111111101000101101011;
assign LUT_1[3428] = 32'b00000000000000001111111110110101;
assign LUT_1[3429] = 32'b00000000000000001001010000110001;
assign LUT_1[3430] = 32'b00000000000000001011101101000110;
assign LUT_1[3431] = 32'b00000000000000000100111111000010;
assign LUT_1[3432] = 32'b00000000000000000111010011010011;
assign LUT_1[3433] = 32'b00000000000000000000100101001111;
assign LUT_1[3434] = 32'b00000000000000000011000001100100;
assign LUT_1[3435] = 32'b11111111111111111100010011100000;
assign LUT_1[3436] = 32'b00000000000000001111001100101010;
assign LUT_1[3437] = 32'b00000000000000001000011110100110;
assign LUT_1[3438] = 32'b00000000000000001010111010111011;
assign LUT_1[3439] = 32'b00000000000000000100001100110111;
assign LUT_1[3440] = 32'b00000000000000001010000001000000;
assign LUT_1[3441] = 32'b00000000000000000011010010111100;
assign LUT_1[3442] = 32'b00000000000000000101101111010001;
assign LUT_1[3443] = 32'b11111111111111111111000001001101;
assign LUT_1[3444] = 32'b00000000000000010001111010010111;
assign LUT_1[3445] = 32'b00000000000000001011001100010011;
assign LUT_1[3446] = 32'b00000000000000001101101000101000;
assign LUT_1[3447] = 32'b00000000000000000110111010100100;
assign LUT_1[3448] = 32'b00000000000000001001001110110101;
assign LUT_1[3449] = 32'b00000000000000000010100000110001;
assign LUT_1[3450] = 32'b00000000000000000100111101000110;
assign LUT_1[3451] = 32'b11111111111111111110001111000010;
assign LUT_1[3452] = 32'b00000000000000010001001000001100;
assign LUT_1[3453] = 32'b00000000000000001010011010001000;
assign LUT_1[3454] = 32'b00000000000000001100110110011101;
assign LUT_1[3455] = 32'b00000000000000000110001000011001;
assign LUT_1[3456] = 32'b00000000000000001000001100111010;
assign LUT_1[3457] = 32'b00000000000000000001011110110110;
assign LUT_1[3458] = 32'b00000000000000000011111011001011;
assign LUT_1[3459] = 32'b11111111111111111101001101000111;
assign LUT_1[3460] = 32'b00000000000000010000000110010001;
assign LUT_1[3461] = 32'b00000000000000001001011000001101;
assign LUT_1[3462] = 32'b00000000000000001011110100100010;
assign LUT_1[3463] = 32'b00000000000000000101000110011110;
assign LUT_1[3464] = 32'b00000000000000000111011010101111;
assign LUT_1[3465] = 32'b00000000000000000000101100101011;
assign LUT_1[3466] = 32'b00000000000000000011001001000000;
assign LUT_1[3467] = 32'b11111111111111111100011010111100;
assign LUT_1[3468] = 32'b00000000000000001111010100000110;
assign LUT_1[3469] = 32'b00000000000000001000100110000010;
assign LUT_1[3470] = 32'b00000000000000001011000010010111;
assign LUT_1[3471] = 32'b00000000000000000100010100010011;
assign LUT_1[3472] = 32'b00000000000000001010001000011100;
assign LUT_1[3473] = 32'b00000000000000000011011010011000;
assign LUT_1[3474] = 32'b00000000000000000101110110101101;
assign LUT_1[3475] = 32'b11111111111111111111001000101001;
assign LUT_1[3476] = 32'b00000000000000010010000001110011;
assign LUT_1[3477] = 32'b00000000000000001011010011101111;
assign LUT_1[3478] = 32'b00000000000000001101110000000100;
assign LUT_1[3479] = 32'b00000000000000000111000010000000;
assign LUT_1[3480] = 32'b00000000000000001001010110010001;
assign LUT_1[3481] = 32'b00000000000000000010101000001101;
assign LUT_1[3482] = 32'b00000000000000000101000100100010;
assign LUT_1[3483] = 32'b11111111111111111110010110011110;
assign LUT_1[3484] = 32'b00000000000000010001001111101000;
assign LUT_1[3485] = 32'b00000000000000001010100001100100;
assign LUT_1[3486] = 32'b00000000000000001100111101111001;
assign LUT_1[3487] = 32'b00000000000000000110001111110101;
assign LUT_1[3488] = 32'b00000000000000001001000111111001;
assign LUT_1[3489] = 32'b00000000000000000010011001110101;
assign LUT_1[3490] = 32'b00000000000000000100110110001010;
assign LUT_1[3491] = 32'b11111111111111111110001000000110;
assign LUT_1[3492] = 32'b00000000000000010001000001010000;
assign LUT_1[3493] = 32'b00000000000000001010010011001100;
assign LUT_1[3494] = 32'b00000000000000001100101111100001;
assign LUT_1[3495] = 32'b00000000000000000110000001011101;
assign LUT_1[3496] = 32'b00000000000000001000010101101110;
assign LUT_1[3497] = 32'b00000000000000000001100111101010;
assign LUT_1[3498] = 32'b00000000000000000100000011111111;
assign LUT_1[3499] = 32'b11111111111111111101010101111011;
assign LUT_1[3500] = 32'b00000000000000010000001111000101;
assign LUT_1[3501] = 32'b00000000000000001001100001000001;
assign LUT_1[3502] = 32'b00000000000000001011111101010110;
assign LUT_1[3503] = 32'b00000000000000000101001111010010;
assign LUT_1[3504] = 32'b00000000000000001011000011011011;
assign LUT_1[3505] = 32'b00000000000000000100010101010111;
assign LUT_1[3506] = 32'b00000000000000000110110001101100;
assign LUT_1[3507] = 32'b00000000000000000000000011101000;
assign LUT_1[3508] = 32'b00000000000000010010111100110010;
assign LUT_1[3509] = 32'b00000000000000001100001110101110;
assign LUT_1[3510] = 32'b00000000000000001110101011000011;
assign LUT_1[3511] = 32'b00000000000000000111111100111111;
assign LUT_1[3512] = 32'b00000000000000001010010001010000;
assign LUT_1[3513] = 32'b00000000000000000011100011001100;
assign LUT_1[3514] = 32'b00000000000000000101111111100001;
assign LUT_1[3515] = 32'b11111111111111111111010001011101;
assign LUT_1[3516] = 32'b00000000000000010010001010100111;
assign LUT_1[3517] = 32'b00000000000000001011011100100011;
assign LUT_1[3518] = 32'b00000000000000001101111000111000;
assign LUT_1[3519] = 32'b00000000000000000111001010110100;
assign LUT_1[3520] = 32'b00000000000000001010001010100010;
assign LUT_1[3521] = 32'b00000000000000000011011100011110;
assign LUT_1[3522] = 32'b00000000000000000101111000110011;
assign LUT_1[3523] = 32'b11111111111111111111001010101111;
assign LUT_1[3524] = 32'b00000000000000010010000011111001;
assign LUT_1[3525] = 32'b00000000000000001011010101110101;
assign LUT_1[3526] = 32'b00000000000000001101110010001010;
assign LUT_1[3527] = 32'b00000000000000000111000100000110;
assign LUT_1[3528] = 32'b00000000000000001001011000010111;
assign LUT_1[3529] = 32'b00000000000000000010101010010011;
assign LUT_1[3530] = 32'b00000000000000000101000110101000;
assign LUT_1[3531] = 32'b11111111111111111110011000100100;
assign LUT_1[3532] = 32'b00000000000000010001010001101110;
assign LUT_1[3533] = 32'b00000000000000001010100011101010;
assign LUT_1[3534] = 32'b00000000000000001100111111111111;
assign LUT_1[3535] = 32'b00000000000000000110010001111011;
assign LUT_1[3536] = 32'b00000000000000001100000110000100;
assign LUT_1[3537] = 32'b00000000000000000101011000000000;
assign LUT_1[3538] = 32'b00000000000000000111110100010101;
assign LUT_1[3539] = 32'b00000000000000000001000110010001;
assign LUT_1[3540] = 32'b00000000000000010011111111011011;
assign LUT_1[3541] = 32'b00000000000000001101010001010111;
assign LUT_1[3542] = 32'b00000000000000001111101101101100;
assign LUT_1[3543] = 32'b00000000000000001000111111101000;
assign LUT_1[3544] = 32'b00000000000000001011010011111001;
assign LUT_1[3545] = 32'b00000000000000000100100101110101;
assign LUT_1[3546] = 32'b00000000000000000111000010001010;
assign LUT_1[3547] = 32'b00000000000000000000010100000110;
assign LUT_1[3548] = 32'b00000000000000010011001101010000;
assign LUT_1[3549] = 32'b00000000000000001100011111001100;
assign LUT_1[3550] = 32'b00000000000000001110111011100001;
assign LUT_1[3551] = 32'b00000000000000001000001101011101;
assign LUT_1[3552] = 32'b00000000000000001011000101100001;
assign LUT_1[3553] = 32'b00000000000000000100010111011101;
assign LUT_1[3554] = 32'b00000000000000000110110011110010;
assign LUT_1[3555] = 32'b00000000000000000000000101101110;
assign LUT_1[3556] = 32'b00000000000000010010111110111000;
assign LUT_1[3557] = 32'b00000000000000001100010000110100;
assign LUT_1[3558] = 32'b00000000000000001110101101001001;
assign LUT_1[3559] = 32'b00000000000000000111111111000101;
assign LUT_1[3560] = 32'b00000000000000001010010011010110;
assign LUT_1[3561] = 32'b00000000000000000011100101010010;
assign LUT_1[3562] = 32'b00000000000000000110000001100111;
assign LUT_1[3563] = 32'b11111111111111111111010011100011;
assign LUT_1[3564] = 32'b00000000000000010010001100101101;
assign LUT_1[3565] = 32'b00000000000000001011011110101001;
assign LUT_1[3566] = 32'b00000000000000001101111010111110;
assign LUT_1[3567] = 32'b00000000000000000111001100111010;
assign LUT_1[3568] = 32'b00000000000000001101000001000011;
assign LUT_1[3569] = 32'b00000000000000000110010010111111;
assign LUT_1[3570] = 32'b00000000000000001000101111010100;
assign LUT_1[3571] = 32'b00000000000000000010000001010000;
assign LUT_1[3572] = 32'b00000000000000010100111010011010;
assign LUT_1[3573] = 32'b00000000000000001110001100010110;
assign LUT_1[3574] = 32'b00000000000000010000101000101011;
assign LUT_1[3575] = 32'b00000000000000001001111010100111;
assign LUT_1[3576] = 32'b00000000000000001100001110111000;
assign LUT_1[3577] = 32'b00000000000000000101100000110100;
assign LUT_1[3578] = 32'b00000000000000000111111101001001;
assign LUT_1[3579] = 32'b00000000000000000001001111000101;
assign LUT_1[3580] = 32'b00000000000000010100001000001111;
assign LUT_1[3581] = 32'b00000000000000001101011010001011;
assign LUT_1[3582] = 32'b00000000000000001111110110100000;
assign LUT_1[3583] = 32'b00000000000000001001001000011100;
assign LUT_1[3584] = 32'b00000000000000000001000111001000;
assign LUT_1[3585] = 32'b11111111111111111010011001000100;
assign LUT_1[3586] = 32'b11111111111111111100110101011001;
assign LUT_1[3587] = 32'b11111111111111110110000111010101;
assign LUT_1[3588] = 32'b00000000000000001001000000011111;
assign LUT_1[3589] = 32'b00000000000000000010010010011011;
assign LUT_1[3590] = 32'b00000000000000000100101110110000;
assign LUT_1[3591] = 32'b11111111111111111110000000101100;
assign LUT_1[3592] = 32'b00000000000000000000010100111101;
assign LUT_1[3593] = 32'b11111111111111111001100110111001;
assign LUT_1[3594] = 32'b11111111111111111100000011001110;
assign LUT_1[3595] = 32'b11111111111111110101010101001010;
assign LUT_1[3596] = 32'b00000000000000001000001110010100;
assign LUT_1[3597] = 32'b00000000000000000001100000010000;
assign LUT_1[3598] = 32'b00000000000000000011111100100101;
assign LUT_1[3599] = 32'b11111111111111111101001110100001;
assign LUT_1[3600] = 32'b00000000000000000011000010101010;
assign LUT_1[3601] = 32'b11111111111111111100010100100110;
assign LUT_1[3602] = 32'b11111111111111111110110000111011;
assign LUT_1[3603] = 32'b11111111111111111000000010110111;
assign LUT_1[3604] = 32'b00000000000000001010111100000001;
assign LUT_1[3605] = 32'b00000000000000000100001101111101;
assign LUT_1[3606] = 32'b00000000000000000110101010010010;
assign LUT_1[3607] = 32'b11111111111111111111111100001110;
assign LUT_1[3608] = 32'b00000000000000000010010000011111;
assign LUT_1[3609] = 32'b11111111111111111011100010011011;
assign LUT_1[3610] = 32'b11111111111111111101111110110000;
assign LUT_1[3611] = 32'b11111111111111110111010000101100;
assign LUT_1[3612] = 32'b00000000000000001010001001110110;
assign LUT_1[3613] = 32'b00000000000000000011011011110010;
assign LUT_1[3614] = 32'b00000000000000000101111000000111;
assign LUT_1[3615] = 32'b11111111111111111111001010000011;
assign LUT_1[3616] = 32'b00000000000000000010000010000111;
assign LUT_1[3617] = 32'b11111111111111111011010100000011;
assign LUT_1[3618] = 32'b11111111111111111101110000011000;
assign LUT_1[3619] = 32'b11111111111111110111000010010100;
assign LUT_1[3620] = 32'b00000000000000001001111011011110;
assign LUT_1[3621] = 32'b00000000000000000011001101011010;
assign LUT_1[3622] = 32'b00000000000000000101101001101111;
assign LUT_1[3623] = 32'b11111111111111111110111011101011;
assign LUT_1[3624] = 32'b00000000000000000001001111111100;
assign LUT_1[3625] = 32'b11111111111111111010100001111000;
assign LUT_1[3626] = 32'b11111111111111111100111110001101;
assign LUT_1[3627] = 32'b11111111111111110110010000001001;
assign LUT_1[3628] = 32'b00000000000000001001001001010011;
assign LUT_1[3629] = 32'b00000000000000000010011011001111;
assign LUT_1[3630] = 32'b00000000000000000100110111100100;
assign LUT_1[3631] = 32'b11111111111111111110001001100000;
assign LUT_1[3632] = 32'b00000000000000000011111101101001;
assign LUT_1[3633] = 32'b11111111111111111101001111100101;
assign LUT_1[3634] = 32'b11111111111111111111101011111010;
assign LUT_1[3635] = 32'b11111111111111111000111101110110;
assign LUT_1[3636] = 32'b00000000000000001011110111000000;
assign LUT_1[3637] = 32'b00000000000000000101001000111100;
assign LUT_1[3638] = 32'b00000000000000000111100101010001;
assign LUT_1[3639] = 32'b00000000000000000000110111001101;
assign LUT_1[3640] = 32'b00000000000000000011001011011110;
assign LUT_1[3641] = 32'b11111111111111111100011101011010;
assign LUT_1[3642] = 32'b11111111111111111110111001101111;
assign LUT_1[3643] = 32'b11111111111111111000001011101011;
assign LUT_1[3644] = 32'b00000000000000001011000100110101;
assign LUT_1[3645] = 32'b00000000000000000100010110110001;
assign LUT_1[3646] = 32'b00000000000000000110110011000110;
assign LUT_1[3647] = 32'b00000000000000000000000101000010;
assign LUT_1[3648] = 32'b00000000000000000011000100110000;
assign LUT_1[3649] = 32'b11111111111111111100010110101100;
assign LUT_1[3650] = 32'b11111111111111111110110011000001;
assign LUT_1[3651] = 32'b11111111111111111000000100111101;
assign LUT_1[3652] = 32'b00000000000000001010111110000111;
assign LUT_1[3653] = 32'b00000000000000000100010000000011;
assign LUT_1[3654] = 32'b00000000000000000110101100011000;
assign LUT_1[3655] = 32'b11111111111111111111111110010100;
assign LUT_1[3656] = 32'b00000000000000000010010010100101;
assign LUT_1[3657] = 32'b11111111111111111011100100100001;
assign LUT_1[3658] = 32'b11111111111111111110000000110110;
assign LUT_1[3659] = 32'b11111111111111110111010010110010;
assign LUT_1[3660] = 32'b00000000000000001010001011111100;
assign LUT_1[3661] = 32'b00000000000000000011011101111000;
assign LUT_1[3662] = 32'b00000000000000000101111010001101;
assign LUT_1[3663] = 32'b11111111111111111111001100001001;
assign LUT_1[3664] = 32'b00000000000000000101000000010010;
assign LUT_1[3665] = 32'b11111111111111111110010010001110;
assign LUT_1[3666] = 32'b00000000000000000000101110100011;
assign LUT_1[3667] = 32'b11111111111111111010000000011111;
assign LUT_1[3668] = 32'b00000000000000001100111001101001;
assign LUT_1[3669] = 32'b00000000000000000110001011100101;
assign LUT_1[3670] = 32'b00000000000000001000100111111010;
assign LUT_1[3671] = 32'b00000000000000000001111001110110;
assign LUT_1[3672] = 32'b00000000000000000100001110000111;
assign LUT_1[3673] = 32'b11111111111111111101100000000011;
assign LUT_1[3674] = 32'b11111111111111111111111100011000;
assign LUT_1[3675] = 32'b11111111111111111001001110010100;
assign LUT_1[3676] = 32'b00000000000000001100000111011110;
assign LUT_1[3677] = 32'b00000000000000000101011001011010;
assign LUT_1[3678] = 32'b00000000000000000111110101101111;
assign LUT_1[3679] = 32'b00000000000000000001000111101011;
assign LUT_1[3680] = 32'b00000000000000000011111111101111;
assign LUT_1[3681] = 32'b11111111111111111101010001101011;
assign LUT_1[3682] = 32'b11111111111111111111101110000000;
assign LUT_1[3683] = 32'b11111111111111111000111111111100;
assign LUT_1[3684] = 32'b00000000000000001011111001000110;
assign LUT_1[3685] = 32'b00000000000000000101001011000010;
assign LUT_1[3686] = 32'b00000000000000000111100111010111;
assign LUT_1[3687] = 32'b00000000000000000000111001010011;
assign LUT_1[3688] = 32'b00000000000000000011001101100100;
assign LUT_1[3689] = 32'b11111111111111111100011111100000;
assign LUT_1[3690] = 32'b11111111111111111110111011110101;
assign LUT_1[3691] = 32'b11111111111111111000001101110001;
assign LUT_1[3692] = 32'b00000000000000001011000110111011;
assign LUT_1[3693] = 32'b00000000000000000100011000110111;
assign LUT_1[3694] = 32'b00000000000000000110110101001100;
assign LUT_1[3695] = 32'b00000000000000000000000111001000;
assign LUT_1[3696] = 32'b00000000000000000101111011010001;
assign LUT_1[3697] = 32'b11111111111111111111001101001101;
assign LUT_1[3698] = 32'b00000000000000000001101001100010;
assign LUT_1[3699] = 32'b11111111111111111010111011011110;
assign LUT_1[3700] = 32'b00000000000000001101110100101000;
assign LUT_1[3701] = 32'b00000000000000000111000110100100;
assign LUT_1[3702] = 32'b00000000000000001001100010111001;
assign LUT_1[3703] = 32'b00000000000000000010110100110101;
assign LUT_1[3704] = 32'b00000000000000000101001001000110;
assign LUT_1[3705] = 32'b11111111111111111110011011000010;
assign LUT_1[3706] = 32'b00000000000000000000110111010111;
assign LUT_1[3707] = 32'b11111111111111111010001001010011;
assign LUT_1[3708] = 32'b00000000000000001101000010011101;
assign LUT_1[3709] = 32'b00000000000000000110010100011001;
assign LUT_1[3710] = 32'b00000000000000001000110000101110;
assign LUT_1[3711] = 32'b00000000000000000010000010101010;
assign LUT_1[3712] = 32'b00000000000000000100000111001011;
assign LUT_1[3713] = 32'b11111111111111111101011001000111;
assign LUT_1[3714] = 32'b11111111111111111111110101011100;
assign LUT_1[3715] = 32'b11111111111111111001000111011000;
assign LUT_1[3716] = 32'b00000000000000001100000000100010;
assign LUT_1[3717] = 32'b00000000000000000101010010011110;
assign LUT_1[3718] = 32'b00000000000000000111101110110011;
assign LUT_1[3719] = 32'b00000000000000000001000000101111;
assign LUT_1[3720] = 32'b00000000000000000011010101000000;
assign LUT_1[3721] = 32'b11111111111111111100100110111100;
assign LUT_1[3722] = 32'b11111111111111111111000011010001;
assign LUT_1[3723] = 32'b11111111111111111000010101001101;
assign LUT_1[3724] = 32'b00000000000000001011001110010111;
assign LUT_1[3725] = 32'b00000000000000000100100000010011;
assign LUT_1[3726] = 32'b00000000000000000110111100101000;
assign LUT_1[3727] = 32'b00000000000000000000001110100100;
assign LUT_1[3728] = 32'b00000000000000000110000010101101;
assign LUT_1[3729] = 32'b11111111111111111111010100101001;
assign LUT_1[3730] = 32'b00000000000000000001110000111110;
assign LUT_1[3731] = 32'b11111111111111111011000010111010;
assign LUT_1[3732] = 32'b00000000000000001101111100000100;
assign LUT_1[3733] = 32'b00000000000000000111001110000000;
assign LUT_1[3734] = 32'b00000000000000001001101010010101;
assign LUT_1[3735] = 32'b00000000000000000010111100010001;
assign LUT_1[3736] = 32'b00000000000000000101010000100010;
assign LUT_1[3737] = 32'b11111111111111111110100010011110;
assign LUT_1[3738] = 32'b00000000000000000000111110110011;
assign LUT_1[3739] = 32'b11111111111111111010010000101111;
assign LUT_1[3740] = 32'b00000000000000001101001001111001;
assign LUT_1[3741] = 32'b00000000000000000110011011110101;
assign LUT_1[3742] = 32'b00000000000000001000111000001010;
assign LUT_1[3743] = 32'b00000000000000000010001010000110;
assign LUT_1[3744] = 32'b00000000000000000101000010001010;
assign LUT_1[3745] = 32'b11111111111111111110010100000110;
assign LUT_1[3746] = 32'b00000000000000000000110000011011;
assign LUT_1[3747] = 32'b11111111111111111010000010010111;
assign LUT_1[3748] = 32'b00000000000000001100111011100001;
assign LUT_1[3749] = 32'b00000000000000000110001101011101;
assign LUT_1[3750] = 32'b00000000000000001000101001110010;
assign LUT_1[3751] = 32'b00000000000000000001111011101110;
assign LUT_1[3752] = 32'b00000000000000000100001111111111;
assign LUT_1[3753] = 32'b11111111111111111101100001111011;
assign LUT_1[3754] = 32'b11111111111111111111111110010000;
assign LUT_1[3755] = 32'b11111111111111111001010000001100;
assign LUT_1[3756] = 32'b00000000000000001100001001010110;
assign LUT_1[3757] = 32'b00000000000000000101011011010010;
assign LUT_1[3758] = 32'b00000000000000000111110111100111;
assign LUT_1[3759] = 32'b00000000000000000001001001100011;
assign LUT_1[3760] = 32'b00000000000000000110111101101100;
assign LUT_1[3761] = 32'b00000000000000000000001111101000;
assign LUT_1[3762] = 32'b00000000000000000010101011111101;
assign LUT_1[3763] = 32'b11111111111111111011111101111001;
assign LUT_1[3764] = 32'b00000000000000001110110111000011;
assign LUT_1[3765] = 32'b00000000000000001000001000111111;
assign LUT_1[3766] = 32'b00000000000000001010100101010100;
assign LUT_1[3767] = 32'b00000000000000000011110111010000;
assign LUT_1[3768] = 32'b00000000000000000110001011100001;
assign LUT_1[3769] = 32'b11111111111111111111011101011101;
assign LUT_1[3770] = 32'b00000000000000000001111001110010;
assign LUT_1[3771] = 32'b11111111111111111011001011101110;
assign LUT_1[3772] = 32'b00000000000000001110000100111000;
assign LUT_1[3773] = 32'b00000000000000000111010110110100;
assign LUT_1[3774] = 32'b00000000000000001001110011001001;
assign LUT_1[3775] = 32'b00000000000000000011000101000101;
assign LUT_1[3776] = 32'b00000000000000000110000100110011;
assign LUT_1[3777] = 32'b11111111111111111111010110101111;
assign LUT_1[3778] = 32'b00000000000000000001110011000100;
assign LUT_1[3779] = 32'b11111111111111111011000101000000;
assign LUT_1[3780] = 32'b00000000000000001101111110001010;
assign LUT_1[3781] = 32'b00000000000000000111010000000110;
assign LUT_1[3782] = 32'b00000000000000001001101100011011;
assign LUT_1[3783] = 32'b00000000000000000010111110010111;
assign LUT_1[3784] = 32'b00000000000000000101010010101000;
assign LUT_1[3785] = 32'b11111111111111111110100100100100;
assign LUT_1[3786] = 32'b00000000000000000001000000111001;
assign LUT_1[3787] = 32'b11111111111111111010010010110101;
assign LUT_1[3788] = 32'b00000000000000001101001011111111;
assign LUT_1[3789] = 32'b00000000000000000110011101111011;
assign LUT_1[3790] = 32'b00000000000000001000111010010000;
assign LUT_1[3791] = 32'b00000000000000000010001100001100;
assign LUT_1[3792] = 32'b00000000000000001000000000010101;
assign LUT_1[3793] = 32'b00000000000000000001010010010001;
assign LUT_1[3794] = 32'b00000000000000000011101110100110;
assign LUT_1[3795] = 32'b11111111111111111101000000100010;
assign LUT_1[3796] = 32'b00000000000000001111111001101100;
assign LUT_1[3797] = 32'b00000000000000001001001011101000;
assign LUT_1[3798] = 32'b00000000000000001011100111111101;
assign LUT_1[3799] = 32'b00000000000000000100111001111001;
assign LUT_1[3800] = 32'b00000000000000000111001110001010;
assign LUT_1[3801] = 32'b00000000000000000000100000000110;
assign LUT_1[3802] = 32'b00000000000000000010111100011011;
assign LUT_1[3803] = 32'b11111111111111111100001110010111;
assign LUT_1[3804] = 32'b00000000000000001111000111100001;
assign LUT_1[3805] = 32'b00000000000000001000011001011101;
assign LUT_1[3806] = 32'b00000000000000001010110101110010;
assign LUT_1[3807] = 32'b00000000000000000100000111101110;
assign LUT_1[3808] = 32'b00000000000000000110111111110010;
assign LUT_1[3809] = 32'b00000000000000000000010001101110;
assign LUT_1[3810] = 32'b00000000000000000010101110000011;
assign LUT_1[3811] = 32'b11111111111111111011111111111111;
assign LUT_1[3812] = 32'b00000000000000001110111001001001;
assign LUT_1[3813] = 32'b00000000000000001000001011000101;
assign LUT_1[3814] = 32'b00000000000000001010100111011010;
assign LUT_1[3815] = 32'b00000000000000000011111001010110;
assign LUT_1[3816] = 32'b00000000000000000110001101100111;
assign LUT_1[3817] = 32'b11111111111111111111011111100011;
assign LUT_1[3818] = 32'b00000000000000000001111011111000;
assign LUT_1[3819] = 32'b11111111111111111011001101110100;
assign LUT_1[3820] = 32'b00000000000000001110000110111110;
assign LUT_1[3821] = 32'b00000000000000000111011000111010;
assign LUT_1[3822] = 32'b00000000000000001001110101001111;
assign LUT_1[3823] = 32'b00000000000000000011000111001011;
assign LUT_1[3824] = 32'b00000000000000001000111011010100;
assign LUT_1[3825] = 32'b00000000000000000010001101010000;
assign LUT_1[3826] = 32'b00000000000000000100101001100101;
assign LUT_1[3827] = 32'b11111111111111111101111011100001;
assign LUT_1[3828] = 32'b00000000000000010000110100101011;
assign LUT_1[3829] = 32'b00000000000000001010000110100111;
assign LUT_1[3830] = 32'b00000000000000001100100010111100;
assign LUT_1[3831] = 32'b00000000000000000101110100111000;
assign LUT_1[3832] = 32'b00000000000000001000001001001001;
assign LUT_1[3833] = 32'b00000000000000000001011011000101;
assign LUT_1[3834] = 32'b00000000000000000011110111011010;
assign LUT_1[3835] = 32'b11111111111111111101001001010110;
assign LUT_1[3836] = 32'b00000000000000010000000010100000;
assign LUT_1[3837] = 32'b00000000000000001001010100011100;
assign LUT_1[3838] = 32'b00000000000000001011110000110001;
assign LUT_1[3839] = 32'b00000000000000000101000010101101;
assign LUT_1[3840] = 32'b11111111111111111110111011010100;
assign LUT_1[3841] = 32'b11111111111111111000001101010000;
assign LUT_1[3842] = 32'b11111111111111111010101001100101;
assign LUT_1[3843] = 32'b11111111111111110011111011100001;
assign LUT_1[3844] = 32'b00000000000000000110110100101011;
assign LUT_1[3845] = 32'b00000000000000000000000110100111;
assign LUT_1[3846] = 32'b00000000000000000010100010111100;
assign LUT_1[3847] = 32'b11111111111111111011110100111000;
assign LUT_1[3848] = 32'b11111111111111111110001001001001;
assign LUT_1[3849] = 32'b11111111111111110111011011000101;
assign LUT_1[3850] = 32'b11111111111111111001110111011010;
assign LUT_1[3851] = 32'b11111111111111110011001001010110;
assign LUT_1[3852] = 32'b00000000000000000110000010100000;
assign LUT_1[3853] = 32'b11111111111111111111010100011100;
assign LUT_1[3854] = 32'b00000000000000000001110000110001;
assign LUT_1[3855] = 32'b11111111111111111011000010101101;
assign LUT_1[3856] = 32'b00000000000000000000110110110110;
assign LUT_1[3857] = 32'b11111111111111111010001000110010;
assign LUT_1[3858] = 32'b11111111111111111100100101000111;
assign LUT_1[3859] = 32'b11111111111111110101110111000011;
assign LUT_1[3860] = 32'b00000000000000001000110000001101;
assign LUT_1[3861] = 32'b00000000000000000010000010001001;
assign LUT_1[3862] = 32'b00000000000000000100011110011110;
assign LUT_1[3863] = 32'b11111111111111111101110000011010;
assign LUT_1[3864] = 32'b00000000000000000000000100101011;
assign LUT_1[3865] = 32'b11111111111111111001010110100111;
assign LUT_1[3866] = 32'b11111111111111111011110010111100;
assign LUT_1[3867] = 32'b11111111111111110101000100111000;
assign LUT_1[3868] = 32'b00000000000000000111111110000010;
assign LUT_1[3869] = 32'b00000000000000000001001111111110;
assign LUT_1[3870] = 32'b00000000000000000011101100010011;
assign LUT_1[3871] = 32'b11111111111111111100111110001111;
assign LUT_1[3872] = 32'b11111111111111111111110110010011;
assign LUT_1[3873] = 32'b11111111111111111001001000001111;
assign LUT_1[3874] = 32'b11111111111111111011100100100100;
assign LUT_1[3875] = 32'b11111111111111110100110110100000;
assign LUT_1[3876] = 32'b00000000000000000111101111101010;
assign LUT_1[3877] = 32'b00000000000000000001000001100110;
assign LUT_1[3878] = 32'b00000000000000000011011101111011;
assign LUT_1[3879] = 32'b11111111111111111100101111110111;
assign LUT_1[3880] = 32'b11111111111111111111000100001000;
assign LUT_1[3881] = 32'b11111111111111111000010110000100;
assign LUT_1[3882] = 32'b11111111111111111010110010011001;
assign LUT_1[3883] = 32'b11111111111111110100000100010101;
assign LUT_1[3884] = 32'b00000000000000000110111101011111;
assign LUT_1[3885] = 32'b00000000000000000000001111011011;
assign LUT_1[3886] = 32'b00000000000000000010101011110000;
assign LUT_1[3887] = 32'b11111111111111111011111101101100;
assign LUT_1[3888] = 32'b00000000000000000001110001110101;
assign LUT_1[3889] = 32'b11111111111111111011000011110001;
assign LUT_1[3890] = 32'b11111111111111111101100000000110;
assign LUT_1[3891] = 32'b11111111111111110110110010000010;
assign LUT_1[3892] = 32'b00000000000000001001101011001100;
assign LUT_1[3893] = 32'b00000000000000000010111101001000;
assign LUT_1[3894] = 32'b00000000000000000101011001011101;
assign LUT_1[3895] = 32'b11111111111111111110101011011001;
assign LUT_1[3896] = 32'b00000000000000000000111111101010;
assign LUT_1[3897] = 32'b11111111111111111010010001100110;
assign LUT_1[3898] = 32'b11111111111111111100101101111011;
assign LUT_1[3899] = 32'b11111111111111110101111111110111;
assign LUT_1[3900] = 32'b00000000000000001000111001000001;
assign LUT_1[3901] = 32'b00000000000000000010001010111101;
assign LUT_1[3902] = 32'b00000000000000000100100111010010;
assign LUT_1[3903] = 32'b11111111111111111101111001001110;
assign LUT_1[3904] = 32'b00000000000000000000111000111100;
assign LUT_1[3905] = 32'b11111111111111111010001010111000;
assign LUT_1[3906] = 32'b11111111111111111100100111001101;
assign LUT_1[3907] = 32'b11111111111111110101111001001001;
assign LUT_1[3908] = 32'b00000000000000001000110010010011;
assign LUT_1[3909] = 32'b00000000000000000010000100001111;
assign LUT_1[3910] = 32'b00000000000000000100100000100100;
assign LUT_1[3911] = 32'b11111111111111111101110010100000;
assign LUT_1[3912] = 32'b00000000000000000000000110110001;
assign LUT_1[3913] = 32'b11111111111111111001011000101101;
assign LUT_1[3914] = 32'b11111111111111111011110101000010;
assign LUT_1[3915] = 32'b11111111111111110101000110111110;
assign LUT_1[3916] = 32'b00000000000000001000000000001000;
assign LUT_1[3917] = 32'b00000000000000000001010010000100;
assign LUT_1[3918] = 32'b00000000000000000011101110011001;
assign LUT_1[3919] = 32'b11111111111111111101000000010101;
assign LUT_1[3920] = 32'b00000000000000000010110100011110;
assign LUT_1[3921] = 32'b11111111111111111100000110011010;
assign LUT_1[3922] = 32'b11111111111111111110100010101111;
assign LUT_1[3923] = 32'b11111111111111110111110100101011;
assign LUT_1[3924] = 32'b00000000000000001010101101110101;
assign LUT_1[3925] = 32'b00000000000000000011111111110001;
assign LUT_1[3926] = 32'b00000000000000000110011100000110;
assign LUT_1[3927] = 32'b11111111111111111111101110000010;
assign LUT_1[3928] = 32'b00000000000000000010000010010011;
assign LUT_1[3929] = 32'b11111111111111111011010100001111;
assign LUT_1[3930] = 32'b11111111111111111101110000100100;
assign LUT_1[3931] = 32'b11111111111111110111000010100000;
assign LUT_1[3932] = 32'b00000000000000001001111011101010;
assign LUT_1[3933] = 32'b00000000000000000011001101100110;
assign LUT_1[3934] = 32'b00000000000000000101101001111011;
assign LUT_1[3935] = 32'b11111111111111111110111011110111;
assign LUT_1[3936] = 32'b00000000000000000001110011111011;
assign LUT_1[3937] = 32'b11111111111111111011000101110111;
assign LUT_1[3938] = 32'b11111111111111111101100010001100;
assign LUT_1[3939] = 32'b11111111111111110110110100001000;
assign LUT_1[3940] = 32'b00000000000000001001101101010010;
assign LUT_1[3941] = 32'b00000000000000000010111111001110;
assign LUT_1[3942] = 32'b00000000000000000101011011100011;
assign LUT_1[3943] = 32'b11111111111111111110101101011111;
assign LUT_1[3944] = 32'b00000000000000000001000001110000;
assign LUT_1[3945] = 32'b11111111111111111010010011101100;
assign LUT_1[3946] = 32'b11111111111111111100110000000001;
assign LUT_1[3947] = 32'b11111111111111110110000001111101;
assign LUT_1[3948] = 32'b00000000000000001000111011000111;
assign LUT_1[3949] = 32'b00000000000000000010001101000011;
assign LUT_1[3950] = 32'b00000000000000000100101001011000;
assign LUT_1[3951] = 32'b11111111111111111101111011010100;
assign LUT_1[3952] = 32'b00000000000000000011101111011101;
assign LUT_1[3953] = 32'b11111111111111111101000001011001;
assign LUT_1[3954] = 32'b11111111111111111111011101101110;
assign LUT_1[3955] = 32'b11111111111111111000101111101010;
assign LUT_1[3956] = 32'b00000000000000001011101000110100;
assign LUT_1[3957] = 32'b00000000000000000100111010110000;
assign LUT_1[3958] = 32'b00000000000000000111010111000101;
assign LUT_1[3959] = 32'b00000000000000000000101001000001;
assign LUT_1[3960] = 32'b00000000000000000010111101010010;
assign LUT_1[3961] = 32'b11111111111111111100001111001110;
assign LUT_1[3962] = 32'b11111111111111111110101011100011;
assign LUT_1[3963] = 32'b11111111111111110111111101011111;
assign LUT_1[3964] = 32'b00000000000000001010110110101001;
assign LUT_1[3965] = 32'b00000000000000000100001000100101;
assign LUT_1[3966] = 32'b00000000000000000110100100111010;
assign LUT_1[3967] = 32'b11111111111111111111110110110110;
assign LUT_1[3968] = 32'b00000000000000000001111011010111;
assign LUT_1[3969] = 32'b11111111111111111011001101010011;
assign LUT_1[3970] = 32'b11111111111111111101101001101000;
assign LUT_1[3971] = 32'b11111111111111110110111011100100;
assign LUT_1[3972] = 32'b00000000000000001001110100101110;
assign LUT_1[3973] = 32'b00000000000000000011000110101010;
assign LUT_1[3974] = 32'b00000000000000000101100010111111;
assign LUT_1[3975] = 32'b11111111111111111110110100111011;
assign LUT_1[3976] = 32'b00000000000000000001001001001100;
assign LUT_1[3977] = 32'b11111111111111111010011011001000;
assign LUT_1[3978] = 32'b11111111111111111100110111011101;
assign LUT_1[3979] = 32'b11111111111111110110001001011001;
assign LUT_1[3980] = 32'b00000000000000001001000010100011;
assign LUT_1[3981] = 32'b00000000000000000010010100011111;
assign LUT_1[3982] = 32'b00000000000000000100110000110100;
assign LUT_1[3983] = 32'b11111111111111111110000010110000;
assign LUT_1[3984] = 32'b00000000000000000011110110111001;
assign LUT_1[3985] = 32'b11111111111111111101001000110101;
assign LUT_1[3986] = 32'b11111111111111111111100101001010;
assign LUT_1[3987] = 32'b11111111111111111000110111000110;
assign LUT_1[3988] = 32'b00000000000000001011110000010000;
assign LUT_1[3989] = 32'b00000000000000000101000010001100;
assign LUT_1[3990] = 32'b00000000000000000111011110100001;
assign LUT_1[3991] = 32'b00000000000000000000110000011101;
assign LUT_1[3992] = 32'b00000000000000000011000100101110;
assign LUT_1[3993] = 32'b11111111111111111100010110101010;
assign LUT_1[3994] = 32'b11111111111111111110110010111111;
assign LUT_1[3995] = 32'b11111111111111111000000100111011;
assign LUT_1[3996] = 32'b00000000000000001010111110000101;
assign LUT_1[3997] = 32'b00000000000000000100010000000001;
assign LUT_1[3998] = 32'b00000000000000000110101100010110;
assign LUT_1[3999] = 32'b11111111111111111111111110010010;
assign LUT_1[4000] = 32'b00000000000000000010110110010110;
assign LUT_1[4001] = 32'b11111111111111111100001000010010;
assign LUT_1[4002] = 32'b11111111111111111110100100100111;
assign LUT_1[4003] = 32'b11111111111111110111110110100011;
assign LUT_1[4004] = 32'b00000000000000001010101111101101;
assign LUT_1[4005] = 32'b00000000000000000100000001101001;
assign LUT_1[4006] = 32'b00000000000000000110011101111110;
assign LUT_1[4007] = 32'b11111111111111111111101111111010;
assign LUT_1[4008] = 32'b00000000000000000010000100001011;
assign LUT_1[4009] = 32'b11111111111111111011010110000111;
assign LUT_1[4010] = 32'b11111111111111111101110010011100;
assign LUT_1[4011] = 32'b11111111111111110111000100011000;
assign LUT_1[4012] = 32'b00000000000000001001111101100010;
assign LUT_1[4013] = 32'b00000000000000000011001111011110;
assign LUT_1[4014] = 32'b00000000000000000101101011110011;
assign LUT_1[4015] = 32'b11111111111111111110111101101111;
assign LUT_1[4016] = 32'b00000000000000000100110001111000;
assign LUT_1[4017] = 32'b11111111111111111110000011110100;
assign LUT_1[4018] = 32'b00000000000000000000100000001001;
assign LUT_1[4019] = 32'b11111111111111111001110010000101;
assign LUT_1[4020] = 32'b00000000000000001100101011001111;
assign LUT_1[4021] = 32'b00000000000000000101111101001011;
assign LUT_1[4022] = 32'b00000000000000001000011001100000;
assign LUT_1[4023] = 32'b00000000000000000001101011011100;
assign LUT_1[4024] = 32'b00000000000000000011111111101101;
assign LUT_1[4025] = 32'b11111111111111111101010001101001;
assign LUT_1[4026] = 32'b11111111111111111111101101111110;
assign LUT_1[4027] = 32'b11111111111111111000111111111010;
assign LUT_1[4028] = 32'b00000000000000001011111001000100;
assign LUT_1[4029] = 32'b00000000000000000101001011000000;
assign LUT_1[4030] = 32'b00000000000000000111100111010101;
assign LUT_1[4031] = 32'b00000000000000000000111001010001;
assign LUT_1[4032] = 32'b00000000000000000011111000111111;
assign LUT_1[4033] = 32'b11111111111111111101001010111011;
assign LUT_1[4034] = 32'b11111111111111111111100111010000;
assign LUT_1[4035] = 32'b11111111111111111000111001001100;
assign LUT_1[4036] = 32'b00000000000000001011110010010110;
assign LUT_1[4037] = 32'b00000000000000000101000100010010;
assign LUT_1[4038] = 32'b00000000000000000111100000100111;
assign LUT_1[4039] = 32'b00000000000000000000110010100011;
assign LUT_1[4040] = 32'b00000000000000000011000110110100;
assign LUT_1[4041] = 32'b11111111111111111100011000110000;
assign LUT_1[4042] = 32'b11111111111111111110110101000101;
assign LUT_1[4043] = 32'b11111111111111111000000111000001;
assign LUT_1[4044] = 32'b00000000000000001011000000001011;
assign LUT_1[4045] = 32'b00000000000000000100010010000111;
assign LUT_1[4046] = 32'b00000000000000000110101110011100;
assign LUT_1[4047] = 32'b00000000000000000000000000011000;
assign LUT_1[4048] = 32'b00000000000000000101110100100001;
assign LUT_1[4049] = 32'b11111111111111111111000110011101;
assign LUT_1[4050] = 32'b00000000000000000001100010110010;
assign LUT_1[4051] = 32'b11111111111111111010110100101110;
assign LUT_1[4052] = 32'b00000000000000001101101101111000;
assign LUT_1[4053] = 32'b00000000000000000110111111110100;
assign LUT_1[4054] = 32'b00000000000000001001011100001001;
assign LUT_1[4055] = 32'b00000000000000000010101110000101;
assign LUT_1[4056] = 32'b00000000000000000101000010010110;
assign LUT_1[4057] = 32'b11111111111111111110010100010010;
assign LUT_1[4058] = 32'b00000000000000000000110000100111;
assign LUT_1[4059] = 32'b11111111111111111010000010100011;
assign LUT_1[4060] = 32'b00000000000000001100111011101101;
assign LUT_1[4061] = 32'b00000000000000000110001101101001;
assign LUT_1[4062] = 32'b00000000000000001000101001111110;
assign LUT_1[4063] = 32'b00000000000000000001111011111010;
assign LUT_1[4064] = 32'b00000000000000000100110011111110;
assign LUT_1[4065] = 32'b11111111111111111110000101111010;
assign LUT_1[4066] = 32'b00000000000000000000100010001111;
assign LUT_1[4067] = 32'b11111111111111111001110100001011;
assign LUT_1[4068] = 32'b00000000000000001100101101010101;
assign LUT_1[4069] = 32'b00000000000000000101111111010001;
assign LUT_1[4070] = 32'b00000000000000001000011011100110;
assign LUT_1[4071] = 32'b00000000000000000001101101100010;
assign LUT_1[4072] = 32'b00000000000000000100000001110011;
assign LUT_1[4073] = 32'b11111111111111111101010011101111;
assign LUT_1[4074] = 32'b11111111111111111111110000000100;
assign LUT_1[4075] = 32'b11111111111111111001000010000000;
assign LUT_1[4076] = 32'b00000000000000001011111011001010;
assign LUT_1[4077] = 32'b00000000000000000101001101000110;
assign LUT_1[4078] = 32'b00000000000000000111101001011011;
assign LUT_1[4079] = 32'b00000000000000000000111011010111;
assign LUT_1[4080] = 32'b00000000000000000110101111100000;
assign LUT_1[4081] = 32'b00000000000000000000000001011100;
assign LUT_1[4082] = 32'b00000000000000000010011101110001;
assign LUT_1[4083] = 32'b11111111111111111011101111101101;
assign LUT_1[4084] = 32'b00000000000000001110101000110111;
assign LUT_1[4085] = 32'b00000000000000000111111010110011;
assign LUT_1[4086] = 32'b00000000000000001010010111001000;
assign LUT_1[4087] = 32'b00000000000000000011101001000100;
assign LUT_1[4088] = 32'b00000000000000000101111101010101;
assign LUT_1[4089] = 32'b11111111111111111111001111010001;
assign LUT_1[4090] = 32'b00000000000000000001101011100110;
assign LUT_1[4091] = 32'b11111111111111111010111101100010;
assign LUT_1[4092] = 32'b00000000000000001101110110101100;
assign LUT_1[4093] = 32'b00000000000000000111001000101000;
assign LUT_1[4094] = 32'b00000000000000001001100100111101;
assign LUT_1[4095] = 32'b00000000000000000010110110111001;
assign LUT_1[4096] = 32'b11111111111111111111110101000110;
assign LUT_1[4097] = 32'b11111111111111111001000111000010;
assign LUT_1[4098] = 32'b11111111111111111011100011010111;
assign LUT_1[4099] = 32'b11111111111111110100110101010011;
assign LUT_1[4100] = 32'b00000000000000000111101110011101;
assign LUT_1[4101] = 32'b00000000000000000001000000011001;
assign LUT_1[4102] = 32'b00000000000000000011011100101110;
assign LUT_1[4103] = 32'b11111111111111111100101110101010;
assign LUT_1[4104] = 32'b11111111111111111111000010111011;
assign LUT_1[4105] = 32'b11111111111111111000010100110111;
assign LUT_1[4106] = 32'b11111111111111111010110001001100;
assign LUT_1[4107] = 32'b11111111111111110100000011001000;
assign LUT_1[4108] = 32'b00000000000000000110111100010010;
assign LUT_1[4109] = 32'b00000000000000000000001110001110;
assign LUT_1[4110] = 32'b00000000000000000010101010100011;
assign LUT_1[4111] = 32'b11111111111111111011111100011111;
assign LUT_1[4112] = 32'b00000000000000000001110000101000;
assign LUT_1[4113] = 32'b11111111111111111011000010100100;
assign LUT_1[4114] = 32'b11111111111111111101011110111001;
assign LUT_1[4115] = 32'b11111111111111110110110000110101;
assign LUT_1[4116] = 32'b00000000000000001001101001111111;
assign LUT_1[4117] = 32'b00000000000000000010111011111011;
assign LUT_1[4118] = 32'b00000000000000000101011000010000;
assign LUT_1[4119] = 32'b11111111111111111110101010001100;
assign LUT_1[4120] = 32'b00000000000000000000111110011101;
assign LUT_1[4121] = 32'b11111111111111111010010000011001;
assign LUT_1[4122] = 32'b11111111111111111100101100101110;
assign LUT_1[4123] = 32'b11111111111111110101111110101010;
assign LUT_1[4124] = 32'b00000000000000001000110111110100;
assign LUT_1[4125] = 32'b00000000000000000010001001110000;
assign LUT_1[4126] = 32'b00000000000000000100100110000101;
assign LUT_1[4127] = 32'b11111111111111111101111000000001;
assign LUT_1[4128] = 32'b00000000000000000000110000000101;
assign LUT_1[4129] = 32'b11111111111111111010000010000001;
assign LUT_1[4130] = 32'b11111111111111111100011110010110;
assign LUT_1[4131] = 32'b11111111111111110101110000010010;
assign LUT_1[4132] = 32'b00000000000000001000101001011100;
assign LUT_1[4133] = 32'b00000000000000000001111011011000;
assign LUT_1[4134] = 32'b00000000000000000100010111101101;
assign LUT_1[4135] = 32'b11111111111111111101101001101001;
assign LUT_1[4136] = 32'b11111111111111111111111101111010;
assign LUT_1[4137] = 32'b11111111111111111001001111110110;
assign LUT_1[4138] = 32'b11111111111111111011101100001011;
assign LUT_1[4139] = 32'b11111111111111110100111110000111;
assign LUT_1[4140] = 32'b00000000000000000111110111010001;
assign LUT_1[4141] = 32'b00000000000000000001001001001101;
assign LUT_1[4142] = 32'b00000000000000000011100101100010;
assign LUT_1[4143] = 32'b11111111111111111100110111011110;
assign LUT_1[4144] = 32'b00000000000000000010101011100111;
assign LUT_1[4145] = 32'b11111111111111111011111101100011;
assign LUT_1[4146] = 32'b11111111111111111110011001111000;
assign LUT_1[4147] = 32'b11111111111111110111101011110100;
assign LUT_1[4148] = 32'b00000000000000001010100100111110;
assign LUT_1[4149] = 32'b00000000000000000011110110111010;
assign LUT_1[4150] = 32'b00000000000000000110010011001111;
assign LUT_1[4151] = 32'b11111111111111111111100101001011;
assign LUT_1[4152] = 32'b00000000000000000001111001011100;
assign LUT_1[4153] = 32'b11111111111111111011001011011000;
assign LUT_1[4154] = 32'b11111111111111111101100111101101;
assign LUT_1[4155] = 32'b11111111111111110110111001101001;
assign LUT_1[4156] = 32'b00000000000000001001110010110011;
assign LUT_1[4157] = 32'b00000000000000000011000100101111;
assign LUT_1[4158] = 32'b00000000000000000101100001000100;
assign LUT_1[4159] = 32'b11111111111111111110110011000000;
assign LUT_1[4160] = 32'b00000000000000000001110010101110;
assign LUT_1[4161] = 32'b11111111111111111011000100101010;
assign LUT_1[4162] = 32'b11111111111111111101100000111111;
assign LUT_1[4163] = 32'b11111111111111110110110010111011;
assign LUT_1[4164] = 32'b00000000000000001001101100000101;
assign LUT_1[4165] = 32'b00000000000000000010111110000001;
assign LUT_1[4166] = 32'b00000000000000000101011010010110;
assign LUT_1[4167] = 32'b11111111111111111110101100010010;
assign LUT_1[4168] = 32'b00000000000000000001000000100011;
assign LUT_1[4169] = 32'b11111111111111111010010010011111;
assign LUT_1[4170] = 32'b11111111111111111100101110110100;
assign LUT_1[4171] = 32'b11111111111111110110000000110000;
assign LUT_1[4172] = 32'b00000000000000001000111001111010;
assign LUT_1[4173] = 32'b00000000000000000010001011110110;
assign LUT_1[4174] = 32'b00000000000000000100101000001011;
assign LUT_1[4175] = 32'b11111111111111111101111010000111;
assign LUT_1[4176] = 32'b00000000000000000011101110010000;
assign LUT_1[4177] = 32'b11111111111111111101000000001100;
assign LUT_1[4178] = 32'b11111111111111111111011100100001;
assign LUT_1[4179] = 32'b11111111111111111000101110011101;
assign LUT_1[4180] = 32'b00000000000000001011100111100111;
assign LUT_1[4181] = 32'b00000000000000000100111001100011;
assign LUT_1[4182] = 32'b00000000000000000111010101111000;
assign LUT_1[4183] = 32'b00000000000000000000100111110100;
assign LUT_1[4184] = 32'b00000000000000000010111100000101;
assign LUT_1[4185] = 32'b11111111111111111100001110000001;
assign LUT_1[4186] = 32'b11111111111111111110101010010110;
assign LUT_1[4187] = 32'b11111111111111110111111100010010;
assign LUT_1[4188] = 32'b00000000000000001010110101011100;
assign LUT_1[4189] = 32'b00000000000000000100000111011000;
assign LUT_1[4190] = 32'b00000000000000000110100011101101;
assign LUT_1[4191] = 32'b11111111111111111111110101101001;
assign LUT_1[4192] = 32'b00000000000000000010101101101101;
assign LUT_1[4193] = 32'b11111111111111111011111111101001;
assign LUT_1[4194] = 32'b11111111111111111110011011111110;
assign LUT_1[4195] = 32'b11111111111111110111101101111010;
assign LUT_1[4196] = 32'b00000000000000001010100111000100;
assign LUT_1[4197] = 32'b00000000000000000011111001000000;
assign LUT_1[4198] = 32'b00000000000000000110010101010101;
assign LUT_1[4199] = 32'b11111111111111111111100111010001;
assign LUT_1[4200] = 32'b00000000000000000001111011100010;
assign LUT_1[4201] = 32'b11111111111111111011001101011110;
assign LUT_1[4202] = 32'b11111111111111111101101001110011;
assign LUT_1[4203] = 32'b11111111111111110110111011101111;
assign LUT_1[4204] = 32'b00000000000000001001110100111001;
assign LUT_1[4205] = 32'b00000000000000000011000110110101;
assign LUT_1[4206] = 32'b00000000000000000101100011001010;
assign LUT_1[4207] = 32'b11111111111111111110110101000110;
assign LUT_1[4208] = 32'b00000000000000000100101001001111;
assign LUT_1[4209] = 32'b11111111111111111101111011001011;
assign LUT_1[4210] = 32'b00000000000000000000010111100000;
assign LUT_1[4211] = 32'b11111111111111111001101001011100;
assign LUT_1[4212] = 32'b00000000000000001100100010100110;
assign LUT_1[4213] = 32'b00000000000000000101110100100010;
assign LUT_1[4214] = 32'b00000000000000001000010000110111;
assign LUT_1[4215] = 32'b00000000000000000001100010110011;
assign LUT_1[4216] = 32'b00000000000000000011110111000100;
assign LUT_1[4217] = 32'b11111111111111111101001001000000;
assign LUT_1[4218] = 32'b11111111111111111111100101010101;
assign LUT_1[4219] = 32'b11111111111111111000110111010001;
assign LUT_1[4220] = 32'b00000000000000001011110000011011;
assign LUT_1[4221] = 32'b00000000000000000101000010010111;
assign LUT_1[4222] = 32'b00000000000000000111011110101100;
assign LUT_1[4223] = 32'b00000000000000000000110000101000;
assign LUT_1[4224] = 32'b00000000000000000010110101001001;
assign LUT_1[4225] = 32'b11111111111111111100000111000101;
assign LUT_1[4226] = 32'b11111111111111111110100011011010;
assign LUT_1[4227] = 32'b11111111111111110111110101010110;
assign LUT_1[4228] = 32'b00000000000000001010101110100000;
assign LUT_1[4229] = 32'b00000000000000000100000000011100;
assign LUT_1[4230] = 32'b00000000000000000110011100110001;
assign LUT_1[4231] = 32'b11111111111111111111101110101101;
assign LUT_1[4232] = 32'b00000000000000000010000010111110;
assign LUT_1[4233] = 32'b11111111111111111011010100111010;
assign LUT_1[4234] = 32'b11111111111111111101110001001111;
assign LUT_1[4235] = 32'b11111111111111110111000011001011;
assign LUT_1[4236] = 32'b00000000000000001001111100010101;
assign LUT_1[4237] = 32'b00000000000000000011001110010001;
assign LUT_1[4238] = 32'b00000000000000000101101010100110;
assign LUT_1[4239] = 32'b11111111111111111110111100100010;
assign LUT_1[4240] = 32'b00000000000000000100110000101011;
assign LUT_1[4241] = 32'b11111111111111111110000010100111;
assign LUT_1[4242] = 32'b00000000000000000000011110111100;
assign LUT_1[4243] = 32'b11111111111111111001110000111000;
assign LUT_1[4244] = 32'b00000000000000001100101010000010;
assign LUT_1[4245] = 32'b00000000000000000101111011111110;
assign LUT_1[4246] = 32'b00000000000000001000011000010011;
assign LUT_1[4247] = 32'b00000000000000000001101010001111;
assign LUT_1[4248] = 32'b00000000000000000011111110100000;
assign LUT_1[4249] = 32'b11111111111111111101010000011100;
assign LUT_1[4250] = 32'b11111111111111111111101100110001;
assign LUT_1[4251] = 32'b11111111111111111000111110101101;
assign LUT_1[4252] = 32'b00000000000000001011110111110111;
assign LUT_1[4253] = 32'b00000000000000000101001001110011;
assign LUT_1[4254] = 32'b00000000000000000111100110001000;
assign LUT_1[4255] = 32'b00000000000000000000111000000100;
assign LUT_1[4256] = 32'b00000000000000000011110000001000;
assign LUT_1[4257] = 32'b11111111111111111101000010000100;
assign LUT_1[4258] = 32'b11111111111111111111011110011001;
assign LUT_1[4259] = 32'b11111111111111111000110000010101;
assign LUT_1[4260] = 32'b00000000000000001011101001011111;
assign LUT_1[4261] = 32'b00000000000000000100111011011011;
assign LUT_1[4262] = 32'b00000000000000000111010111110000;
assign LUT_1[4263] = 32'b00000000000000000000101001101100;
assign LUT_1[4264] = 32'b00000000000000000010111101111101;
assign LUT_1[4265] = 32'b11111111111111111100001111111001;
assign LUT_1[4266] = 32'b11111111111111111110101100001110;
assign LUT_1[4267] = 32'b11111111111111110111111110001010;
assign LUT_1[4268] = 32'b00000000000000001010110111010100;
assign LUT_1[4269] = 32'b00000000000000000100001001010000;
assign LUT_1[4270] = 32'b00000000000000000110100101100101;
assign LUT_1[4271] = 32'b11111111111111111111110111100001;
assign LUT_1[4272] = 32'b00000000000000000101101011101010;
assign LUT_1[4273] = 32'b11111111111111111110111101100110;
assign LUT_1[4274] = 32'b00000000000000000001011001111011;
assign LUT_1[4275] = 32'b11111111111111111010101011110111;
assign LUT_1[4276] = 32'b00000000000000001101100101000001;
assign LUT_1[4277] = 32'b00000000000000000110110110111101;
assign LUT_1[4278] = 32'b00000000000000001001010011010010;
assign LUT_1[4279] = 32'b00000000000000000010100101001110;
assign LUT_1[4280] = 32'b00000000000000000100111001011111;
assign LUT_1[4281] = 32'b11111111111111111110001011011011;
assign LUT_1[4282] = 32'b00000000000000000000100111110000;
assign LUT_1[4283] = 32'b11111111111111111001111001101100;
assign LUT_1[4284] = 32'b00000000000000001100110010110110;
assign LUT_1[4285] = 32'b00000000000000000110000100110010;
assign LUT_1[4286] = 32'b00000000000000001000100001000111;
assign LUT_1[4287] = 32'b00000000000000000001110011000011;
assign LUT_1[4288] = 32'b00000000000000000100110010110001;
assign LUT_1[4289] = 32'b11111111111111111110000100101101;
assign LUT_1[4290] = 32'b00000000000000000000100001000010;
assign LUT_1[4291] = 32'b11111111111111111001110010111110;
assign LUT_1[4292] = 32'b00000000000000001100101100001000;
assign LUT_1[4293] = 32'b00000000000000000101111110000100;
assign LUT_1[4294] = 32'b00000000000000001000011010011001;
assign LUT_1[4295] = 32'b00000000000000000001101100010101;
assign LUT_1[4296] = 32'b00000000000000000100000000100110;
assign LUT_1[4297] = 32'b11111111111111111101010010100010;
assign LUT_1[4298] = 32'b11111111111111111111101110110111;
assign LUT_1[4299] = 32'b11111111111111111001000000110011;
assign LUT_1[4300] = 32'b00000000000000001011111001111101;
assign LUT_1[4301] = 32'b00000000000000000101001011111001;
assign LUT_1[4302] = 32'b00000000000000000111101000001110;
assign LUT_1[4303] = 32'b00000000000000000000111010001010;
assign LUT_1[4304] = 32'b00000000000000000110101110010011;
assign LUT_1[4305] = 32'b00000000000000000000000000001111;
assign LUT_1[4306] = 32'b00000000000000000010011100100100;
assign LUT_1[4307] = 32'b11111111111111111011101110100000;
assign LUT_1[4308] = 32'b00000000000000001110100111101010;
assign LUT_1[4309] = 32'b00000000000000000111111001100110;
assign LUT_1[4310] = 32'b00000000000000001010010101111011;
assign LUT_1[4311] = 32'b00000000000000000011100111110111;
assign LUT_1[4312] = 32'b00000000000000000101111100001000;
assign LUT_1[4313] = 32'b11111111111111111111001110000100;
assign LUT_1[4314] = 32'b00000000000000000001101010011001;
assign LUT_1[4315] = 32'b11111111111111111010111100010101;
assign LUT_1[4316] = 32'b00000000000000001101110101011111;
assign LUT_1[4317] = 32'b00000000000000000111000111011011;
assign LUT_1[4318] = 32'b00000000000000001001100011110000;
assign LUT_1[4319] = 32'b00000000000000000010110101101100;
assign LUT_1[4320] = 32'b00000000000000000101101101110000;
assign LUT_1[4321] = 32'b11111111111111111110111111101100;
assign LUT_1[4322] = 32'b00000000000000000001011100000001;
assign LUT_1[4323] = 32'b11111111111111111010101101111101;
assign LUT_1[4324] = 32'b00000000000000001101100111000111;
assign LUT_1[4325] = 32'b00000000000000000110111001000011;
assign LUT_1[4326] = 32'b00000000000000001001010101011000;
assign LUT_1[4327] = 32'b00000000000000000010100111010100;
assign LUT_1[4328] = 32'b00000000000000000100111011100101;
assign LUT_1[4329] = 32'b11111111111111111110001101100001;
assign LUT_1[4330] = 32'b00000000000000000000101001110110;
assign LUT_1[4331] = 32'b11111111111111111001111011110010;
assign LUT_1[4332] = 32'b00000000000000001100110100111100;
assign LUT_1[4333] = 32'b00000000000000000110000110111000;
assign LUT_1[4334] = 32'b00000000000000001000100011001101;
assign LUT_1[4335] = 32'b00000000000000000001110101001001;
assign LUT_1[4336] = 32'b00000000000000000111101001010010;
assign LUT_1[4337] = 32'b00000000000000000000111011001110;
assign LUT_1[4338] = 32'b00000000000000000011010111100011;
assign LUT_1[4339] = 32'b11111111111111111100101001011111;
assign LUT_1[4340] = 32'b00000000000000001111100010101001;
assign LUT_1[4341] = 32'b00000000000000001000110100100101;
assign LUT_1[4342] = 32'b00000000000000001011010000111010;
assign LUT_1[4343] = 32'b00000000000000000100100010110110;
assign LUT_1[4344] = 32'b00000000000000000110110111000111;
assign LUT_1[4345] = 32'b00000000000000000000001001000011;
assign LUT_1[4346] = 32'b00000000000000000010100101011000;
assign LUT_1[4347] = 32'b11111111111111111011110111010100;
assign LUT_1[4348] = 32'b00000000000000001110110000011110;
assign LUT_1[4349] = 32'b00000000000000001000000010011010;
assign LUT_1[4350] = 32'b00000000000000001010011110101111;
assign LUT_1[4351] = 32'b00000000000000000011110000101011;
assign LUT_1[4352] = 32'b11111111111111111101101001010010;
assign LUT_1[4353] = 32'b11111111111111110110111011001110;
assign LUT_1[4354] = 32'b11111111111111111001010111100011;
assign LUT_1[4355] = 32'b11111111111111110010101001011111;
assign LUT_1[4356] = 32'b00000000000000000101100010101001;
assign LUT_1[4357] = 32'b11111111111111111110110100100101;
assign LUT_1[4358] = 32'b00000000000000000001010000111010;
assign LUT_1[4359] = 32'b11111111111111111010100010110110;
assign LUT_1[4360] = 32'b11111111111111111100110111000111;
assign LUT_1[4361] = 32'b11111111111111110110001001000011;
assign LUT_1[4362] = 32'b11111111111111111000100101011000;
assign LUT_1[4363] = 32'b11111111111111110001110111010100;
assign LUT_1[4364] = 32'b00000000000000000100110000011110;
assign LUT_1[4365] = 32'b11111111111111111110000010011010;
assign LUT_1[4366] = 32'b00000000000000000000011110101111;
assign LUT_1[4367] = 32'b11111111111111111001110000101011;
assign LUT_1[4368] = 32'b11111111111111111111100100110100;
assign LUT_1[4369] = 32'b11111111111111111000110110110000;
assign LUT_1[4370] = 32'b11111111111111111011010011000101;
assign LUT_1[4371] = 32'b11111111111111110100100101000001;
assign LUT_1[4372] = 32'b00000000000000000111011110001011;
assign LUT_1[4373] = 32'b00000000000000000000110000000111;
assign LUT_1[4374] = 32'b00000000000000000011001100011100;
assign LUT_1[4375] = 32'b11111111111111111100011110011000;
assign LUT_1[4376] = 32'b11111111111111111110110010101001;
assign LUT_1[4377] = 32'b11111111111111111000000100100101;
assign LUT_1[4378] = 32'b11111111111111111010100000111010;
assign LUT_1[4379] = 32'b11111111111111110011110010110110;
assign LUT_1[4380] = 32'b00000000000000000110101100000000;
assign LUT_1[4381] = 32'b11111111111111111111111101111100;
assign LUT_1[4382] = 32'b00000000000000000010011010010001;
assign LUT_1[4383] = 32'b11111111111111111011101100001101;
assign LUT_1[4384] = 32'b11111111111111111110100100010001;
assign LUT_1[4385] = 32'b11111111111111110111110110001101;
assign LUT_1[4386] = 32'b11111111111111111010010010100010;
assign LUT_1[4387] = 32'b11111111111111110011100100011110;
assign LUT_1[4388] = 32'b00000000000000000110011101101000;
assign LUT_1[4389] = 32'b11111111111111111111101111100100;
assign LUT_1[4390] = 32'b00000000000000000010001011111001;
assign LUT_1[4391] = 32'b11111111111111111011011101110101;
assign LUT_1[4392] = 32'b11111111111111111101110010000110;
assign LUT_1[4393] = 32'b11111111111111110111000100000010;
assign LUT_1[4394] = 32'b11111111111111111001100000010111;
assign LUT_1[4395] = 32'b11111111111111110010110010010011;
assign LUT_1[4396] = 32'b00000000000000000101101011011101;
assign LUT_1[4397] = 32'b11111111111111111110111101011001;
assign LUT_1[4398] = 32'b00000000000000000001011001101110;
assign LUT_1[4399] = 32'b11111111111111111010101011101010;
assign LUT_1[4400] = 32'b00000000000000000000011111110011;
assign LUT_1[4401] = 32'b11111111111111111001110001101111;
assign LUT_1[4402] = 32'b11111111111111111100001110000100;
assign LUT_1[4403] = 32'b11111111111111110101100000000000;
assign LUT_1[4404] = 32'b00000000000000001000011001001010;
assign LUT_1[4405] = 32'b00000000000000000001101011000110;
assign LUT_1[4406] = 32'b00000000000000000100000111011011;
assign LUT_1[4407] = 32'b11111111111111111101011001010111;
assign LUT_1[4408] = 32'b11111111111111111111101101101000;
assign LUT_1[4409] = 32'b11111111111111111000111111100100;
assign LUT_1[4410] = 32'b11111111111111111011011011111001;
assign LUT_1[4411] = 32'b11111111111111110100101101110101;
assign LUT_1[4412] = 32'b00000000000000000111100110111111;
assign LUT_1[4413] = 32'b00000000000000000000111000111011;
assign LUT_1[4414] = 32'b00000000000000000011010101010000;
assign LUT_1[4415] = 32'b11111111111111111100100111001100;
assign LUT_1[4416] = 32'b11111111111111111111100110111010;
assign LUT_1[4417] = 32'b11111111111111111000111000110110;
assign LUT_1[4418] = 32'b11111111111111111011010101001011;
assign LUT_1[4419] = 32'b11111111111111110100100111000111;
assign LUT_1[4420] = 32'b00000000000000000111100000010001;
assign LUT_1[4421] = 32'b00000000000000000000110010001101;
assign LUT_1[4422] = 32'b00000000000000000011001110100010;
assign LUT_1[4423] = 32'b11111111111111111100100000011110;
assign LUT_1[4424] = 32'b11111111111111111110110100101111;
assign LUT_1[4425] = 32'b11111111111111111000000110101011;
assign LUT_1[4426] = 32'b11111111111111111010100011000000;
assign LUT_1[4427] = 32'b11111111111111110011110100111100;
assign LUT_1[4428] = 32'b00000000000000000110101110000110;
assign LUT_1[4429] = 32'b00000000000000000000000000000010;
assign LUT_1[4430] = 32'b00000000000000000010011100010111;
assign LUT_1[4431] = 32'b11111111111111111011101110010011;
assign LUT_1[4432] = 32'b00000000000000000001100010011100;
assign LUT_1[4433] = 32'b11111111111111111010110100011000;
assign LUT_1[4434] = 32'b11111111111111111101010000101101;
assign LUT_1[4435] = 32'b11111111111111110110100010101001;
assign LUT_1[4436] = 32'b00000000000000001001011011110011;
assign LUT_1[4437] = 32'b00000000000000000010101101101111;
assign LUT_1[4438] = 32'b00000000000000000101001010000100;
assign LUT_1[4439] = 32'b11111111111111111110011100000000;
assign LUT_1[4440] = 32'b00000000000000000000110000010001;
assign LUT_1[4441] = 32'b11111111111111111010000010001101;
assign LUT_1[4442] = 32'b11111111111111111100011110100010;
assign LUT_1[4443] = 32'b11111111111111110101110000011110;
assign LUT_1[4444] = 32'b00000000000000001000101001101000;
assign LUT_1[4445] = 32'b00000000000000000001111011100100;
assign LUT_1[4446] = 32'b00000000000000000100010111111001;
assign LUT_1[4447] = 32'b11111111111111111101101001110101;
assign LUT_1[4448] = 32'b00000000000000000000100001111001;
assign LUT_1[4449] = 32'b11111111111111111001110011110101;
assign LUT_1[4450] = 32'b11111111111111111100010000001010;
assign LUT_1[4451] = 32'b11111111111111110101100010000110;
assign LUT_1[4452] = 32'b00000000000000001000011011010000;
assign LUT_1[4453] = 32'b00000000000000000001101101001100;
assign LUT_1[4454] = 32'b00000000000000000100001001100001;
assign LUT_1[4455] = 32'b11111111111111111101011011011101;
assign LUT_1[4456] = 32'b11111111111111111111101111101110;
assign LUT_1[4457] = 32'b11111111111111111001000001101010;
assign LUT_1[4458] = 32'b11111111111111111011011101111111;
assign LUT_1[4459] = 32'b11111111111111110100101111111011;
assign LUT_1[4460] = 32'b00000000000000000111101001000101;
assign LUT_1[4461] = 32'b00000000000000000000111011000001;
assign LUT_1[4462] = 32'b00000000000000000011010111010110;
assign LUT_1[4463] = 32'b11111111111111111100101001010010;
assign LUT_1[4464] = 32'b00000000000000000010011101011011;
assign LUT_1[4465] = 32'b11111111111111111011101111010111;
assign LUT_1[4466] = 32'b11111111111111111110001011101100;
assign LUT_1[4467] = 32'b11111111111111110111011101101000;
assign LUT_1[4468] = 32'b00000000000000001010010110110010;
assign LUT_1[4469] = 32'b00000000000000000011101000101110;
assign LUT_1[4470] = 32'b00000000000000000110000101000011;
assign LUT_1[4471] = 32'b11111111111111111111010110111111;
assign LUT_1[4472] = 32'b00000000000000000001101011010000;
assign LUT_1[4473] = 32'b11111111111111111010111101001100;
assign LUT_1[4474] = 32'b11111111111111111101011001100001;
assign LUT_1[4475] = 32'b11111111111111110110101011011101;
assign LUT_1[4476] = 32'b00000000000000001001100100100111;
assign LUT_1[4477] = 32'b00000000000000000010110110100011;
assign LUT_1[4478] = 32'b00000000000000000101010010111000;
assign LUT_1[4479] = 32'b11111111111111111110100100110100;
assign LUT_1[4480] = 32'b00000000000000000000101001010101;
assign LUT_1[4481] = 32'b11111111111111111001111011010001;
assign LUT_1[4482] = 32'b11111111111111111100010111100110;
assign LUT_1[4483] = 32'b11111111111111110101101001100010;
assign LUT_1[4484] = 32'b00000000000000001000100010101100;
assign LUT_1[4485] = 32'b00000000000000000001110100101000;
assign LUT_1[4486] = 32'b00000000000000000100010000111101;
assign LUT_1[4487] = 32'b11111111111111111101100010111001;
assign LUT_1[4488] = 32'b11111111111111111111110111001010;
assign LUT_1[4489] = 32'b11111111111111111001001001000110;
assign LUT_1[4490] = 32'b11111111111111111011100101011011;
assign LUT_1[4491] = 32'b11111111111111110100110111010111;
assign LUT_1[4492] = 32'b00000000000000000111110000100001;
assign LUT_1[4493] = 32'b00000000000000000001000010011101;
assign LUT_1[4494] = 32'b00000000000000000011011110110010;
assign LUT_1[4495] = 32'b11111111111111111100110000101110;
assign LUT_1[4496] = 32'b00000000000000000010100100110111;
assign LUT_1[4497] = 32'b11111111111111111011110110110011;
assign LUT_1[4498] = 32'b11111111111111111110010011001000;
assign LUT_1[4499] = 32'b11111111111111110111100101000100;
assign LUT_1[4500] = 32'b00000000000000001010011110001110;
assign LUT_1[4501] = 32'b00000000000000000011110000001010;
assign LUT_1[4502] = 32'b00000000000000000110001100011111;
assign LUT_1[4503] = 32'b11111111111111111111011110011011;
assign LUT_1[4504] = 32'b00000000000000000001110010101100;
assign LUT_1[4505] = 32'b11111111111111111011000100101000;
assign LUT_1[4506] = 32'b11111111111111111101100000111101;
assign LUT_1[4507] = 32'b11111111111111110110110010111001;
assign LUT_1[4508] = 32'b00000000000000001001101100000011;
assign LUT_1[4509] = 32'b00000000000000000010111101111111;
assign LUT_1[4510] = 32'b00000000000000000101011010010100;
assign LUT_1[4511] = 32'b11111111111111111110101100010000;
assign LUT_1[4512] = 32'b00000000000000000001100100010100;
assign LUT_1[4513] = 32'b11111111111111111010110110010000;
assign LUT_1[4514] = 32'b11111111111111111101010010100101;
assign LUT_1[4515] = 32'b11111111111111110110100100100001;
assign LUT_1[4516] = 32'b00000000000000001001011101101011;
assign LUT_1[4517] = 32'b00000000000000000010101111100111;
assign LUT_1[4518] = 32'b00000000000000000101001011111100;
assign LUT_1[4519] = 32'b11111111111111111110011101111000;
assign LUT_1[4520] = 32'b00000000000000000000110010001001;
assign LUT_1[4521] = 32'b11111111111111111010000100000101;
assign LUT_1[4522] = 32'b11111111111111111100100000011010;
assign LUT_1[4523] = 32'b11111111111111110101110010010110;
assign LUT_1[4524] = 32'b00000000000000001000101011100000;
assign LUT_1[4525] = 32'b00000000000000000001111101011100;
assign LUT_1[4526] = 32'b00000000000000000100011001110001;
assign LUT_1[4527] = 32'b11111111111111111101101011101101;
assign LUT_1[4528] = 32'b00000000000000000011011111110110;
assign LUT_1[4529] = 32'b11111111111111111100110001110010;
assign LUT_1[4530] = 32'b11111111111111111111001110000111;
assign LUT_1[4531] = 32'b11111111111111111000100000000011;
assign LUT_1[4532] = 32'b00000000000000001011011001001101;
assign LUT_1[4533] = 32'b00000000000000000100101011001001;
assign LUT_1[4534] = 32'b00000000000000000111000111011110;
assign LUT_1[4535] = 32'b00000000000000000000011001011010;
assign LUT_1[4536] = 32'b00000000000000000010101101101011;
assign LUT_1[4537] = 32'b11111111111111111011111111100111;
assign LUT_1[4538] = 32'b11111111111111111110011011111100;
assign LUT_1[4539] = 32'b11111111111111110111101101111000;
assign LUT_1[4540] = 32'b00000000000000001010100111000010;
assign LUT_1[4541] = 32'b00000000000000000011111000111110;
assign LUT_1[4542] = 32'b00000000000000000110010101010011;
assign LUT_1[4543] = 32'b11111111111111111111100111001111;
assign LUT_1[4544] = 32'b00000000000000000010100110111101;
assign LUT_1[4545] = 32'b11111111111111111011111000111001;
assign LUT_1[4546] = 32'b11111111111111111110010101001110;
assign LUT_1[4547] = 32'b11111111111111110111100111001010;
assign LUT_1[4548] = 32'b00000000000000001010100000010100;
assign LUT_1[4549] = 32'b00000000000000000011110010010000;
assign LUT_1[4550] = 32'b00000000000000000110001110100101;
assign LUT_1[4551] = 32'b11111111111111111111100000100001;
assign LUT_1[4552] = 32'b00000000000000000001110100110010;
assign LUT_1[4553] = 32'b11111111111111111011000110101110;
assign LUT_1[4554] = 32'b11111111111111111101100011000011;
assign LUT_1[4555] = 32'b11111111111111110110110100111111;
assign LUT_1[4556] = 32'b00000000000000001001101110001001;
assign LUT_1[4557] = 32'b00000000000000000011000000000101;
assign LUT_1[4558] = 32'b00000000000000000101011100011010;
assign LUT_1[4559] = 32'b11111111111111111110101110010110;
assign LUT_1[4560] = 32'b00000000000000000100100010011111;
assign LUT_1[4561] = 32'b11111111111111111101110100011011;
assign LUT_1[4562] = 32'b00000000000000000000010000110000;
assign LUT_1[4563] = 32'b11111111111111111001100010101100;
assign LUT_1[4564] = 32'b00000000000000001100011011110110;
assign LUT_1[4565] = 32'b00000000000000000101101101110010;
assign LUT_1[4566] = 32'b00000000000000001000001010000111;
assign LUT_1[4567] = 32'b00000000000000000001011100000011;
assign LUT_1[4568] = 32'b00000000000000000011110000010100;
assign LUT_1[4569] = 32'b11111111111111111101000010010000;
assign LUT_1[4570] = 32'b11111111111111111111011110100101;
assign LUT_1[4571] = 32'b11111111111111111000110000100001;
assign LUT_1[4572] = 32'b00000000000000001011101001101011;
assign LUT_1[4573] = 32'b00000000000000000100111011100111;
assign LUT_1[4574] = 32'b00000000000000000111010111111100;
assign LUT_1[4575] = 32'b00000000000000000000101001111000;
assign LUT_1[4576] = 32'b00000000000000000011100001111100;
assign LUT_1[4577] = 32'b11111111111111111100110011111000;
assign LUT_1[4578] = 32'b11111111111111111111010000001101;
assign LUT_1[4579] = 32'b11111111111111111000100010001001;
assign LUT_1[4580] = 32'b00000000000000001011011011010011;
assign LUT_1[4581] = 32'b00000000000000000100101101001111;
assign LUT_1[4582] = 32'b00000000000000000111001001100100;
assign LUT_1[4583] = 32'b00000000000000000000011011100000;
assign LUT_1[4584] = 32'b00000000000000000010101111110001;
assign LUT_1[4585] = 32'b11111111111111111100000001101101;
assign LUT_1[4586] = 32'b11111111111111111110011110000010;
assign LUT_1[4587] = 32'b11111111111111110111101111111110;
assign LUT_1[4588] = 32'b00000000000000001010101001001000;
assign LUT_1[4589] = 32'b00000000000000000011111011000100;
assign LUT_1[4590] = 32'b00000000000000000110010111011001;
assign LUT_1[4591] = 32'b11111111111111111111101001010101;
assign LUT_1[4592] = 32'b00000000000000000101011101011110;
assign LUT_1[4593] = 32'b11111111111111111110101111011010;
assign LUT_1[4594] = 32'b00000000000000000001001011101111;
assign LUT_1[4595] = 32'b11111111111111111010011101101011;
assign LUT_1[4596] = 32'b00000000000000001101010110110101;
assign LUT_1[4597] = 32'b00000000000000000110101000110001;
assign LUT_1[4598] = 32'b00000000000000001001000101000110;
assign LUT_1[4599] = 32'b00000000000000000010010111000010;
assign LUT_1[4600] = 32'b00000000000000000100101011010011;
assign LUT_1[4601] = 32'b11111111111111111101111101001111;
assign LUT_1[4602] = 32'b00000000000000000000011001100100;
assign LUT_1[4603] = 32'b11111111111111111001101011100000;
assign LUT_1[4604] = 32'b00000000000000001100100100101010;
assign LUT_1[4605] = 32'b00000000000000000101110110100110;
assign LUT_1[4606] = 32'b00000000000000001000010010111011;
assign LUT_1[4607] = 32'b00000000000000000001100100110111;
assign LUT_1[4608] = 32'b11111111111111111001100011100011;
assign LUT_1[4609] = 32'b11111111111111110010110101011111;
assign LUT_1[4610] = 32'b11111111111111110101010001110100;
assign LUT_1[4611] = 32'b11111111111111101110100011110000;
assign LUT_1[4612] = 32'b00000000000000000001011100111010;
assign LUT_1[4613] = 32'b11111111111111111010101110110110;
assign LUT_1[4614] = 32'b11111111111111111101001011001011;
assign LUT_1[4615] = 32'b11111111111111110110011101000111;
assign LUT_1[4616] = 32'b11111111111111111000110001011000;
assign LUT_1[4617] = 32'b11111111111111110010000011010100;
assign LUT_1[4618] = 32'b11111111111111110100011111101001;
assign LUT_1[4619] = 32'b11111111111111101101110001100101;
assign LUT_1[4620] = 32'b00000000000000000000101010101111;
assign LUT_1[4621] = 32'b11111111111111111001111100101011;
assign LUT_1[4622] = 32'b11111111111111111100011001000000;
assign LUT_1[4623] = 32'b11111111111111110101101010111100;
assign LUT_1[4624] = 32'b11111111111111111011011111000101;
assign LUT_1[4625] = 32'b11111111111111110100110001000001;
assign LUT_1[4626] = 32'b11111111111111110111001101010110;
assign LUT_1[4627] = 32'b11111111111111110000011111010010;
assign LUT_1[4628] = 32'b00000000000000000011011000011100;
assign LUT_1[4629] = 32'b11111111111111111100101010011000;
assign LUT_1[4630] = 32'b11111111111111111111000110101101;
assign LUT_1[4631] = 32'b11111111111111111000011000101001;
assign LUT_1[4632] = 32'b11111111111111111010101100111010;
assign LUT_1[4633] = 32'b11111111111111110011111110110110;
assign LUT_1[4634] = 32'b11111111111111110110011011001011;
assign LUT_1[4635] = 32'b11111111111111101111101101000111;
assign LUT_1[4636] = 32'b00000000000000000010100110010001;
assign LUT_1[4637] = 32'b11111111111111111011111000001101;
assign LUT_1[4638] = 32'b11111111111111111110010100100010;
assign LUT_1[4639] = 32'b11111111111111110111100110011110;
assign LUT_1[4640] = 32'b11111111111111111010011110100010;
assign LUT_1[4641] = 32'b11111111111111110011110000011110;
assign LUT_1[4642] = 32'b11111111111111110110001100110011;
assign LUT_1[4643] = 32'b11111111111111101111011110101111;
assign LUT_1[4644] = 32'b00000000000000000010010111111001;
assign LUT_1[4645] = 32'b11111111111111111011101001110101;
assign LUT_1[4646] = 32'b11111111111111111110000110001010;
assign LUT_1[4647] = 32'b11111111111111110111011000000110;
assign LUT_1[4648] = 32'b11111111111111111001101100010111;
assign LUT_1[4649] = 32'b11111111111111110010111110010011;
assign LUT_1[4650] = 32'b11111111111111110101011010101000;
assign LUT_1[4651] = 32'b11111111111111101110101100100100;
assign LUT_1[4652] = 32'b00000000000000000001100101101110;
assign LUT_1[4653] = 32'b11111111111111111010110111101010;
assign LUT_1[4654] = 32'b11111111111111111101010011111111;
assign LUT_1[4655] = 32'b11111111111111110110100101111011;
assign LUT_1[4656] = 32'b11111111111111111100011010000100;
assign LUT_1[4657] = 32'b11111111111111110101101100000000;
assign LUT_1[4658] = 32'b11111111111111111000001000010101;
assign LUT_1[4659] = 32'b11111111111111110001011010010001;
assign LUT_1[4660] = 32'b00000000000000000100010011011011;
assign LUT_1[4661] = 32'b11111111111111111101100101010111;
assign LUT_1[4662] = 32'b00000000000000000000000001101100;
assign LUT_1[4663] = 32'b11111111111111111001010011101000;
assign LUT_1[4664] = 32'b11111111111111111011100111111001;
assign LUT_1[4665] = 32'b11111111111111110100111001110101;
assign LUT_1[4666] = 32'b11111111111111110111010110001010;
assign LUT_1[4667] = 32'b11111111111111110000101000000110;
assign LUT_1[4668] = 32'b00000000000000000011100001010000;
assign LUT_1[4669] = 32'b11111111111111111100110011001100;
assign LUT_1[4670] = 32'b11111111111111111111001111100001;
assign LUT_1[4671] = 32'b11111111111111111000100001011101;
assign LUT_1[4672] = 32'b11111111111111111011100001001011;
assign LUT_1[4673] = 32'b11111111111111110100110011000111;
assign LUT_1[4674] = 32'b11111111111111110111001111011100;
assign LUT_1[4675] = 32'b11111111111111110000100001011000;
assign LUT_1[4676] = 32'b00000000000000000011011010100010;
assign LUT_1[4677] = 32'b11111111111111111100101100011110;
assign LUT_1[4678] = 32'b11111111111111111111001000110011;
assign LUT_1[4679] = 32'b11111111111111111000011010101111;
assign LUT_1[4680] = 32'b11111111111111111010101111000000;
assign LUT_1[4681] = 32'b11111111111111110100000000111100;
assign LUT_1[4682] = 32'b11111111111111110110011101010001;
assign LUT_1[4683] = 32'b11111111111111101111101111001101;
assign LUT_1[4684] = 32'b00000000000000000010101000010111;
assign LUT_1[4685] = 32'b11111111111111111011111010010011;
assign LUT_1[4686] = 32'b11111111111111111110010110101000;
assign LUT_1[4687] = 32'b11111111111111110111101000100100;
assign LUT_1[4688] = 32'b11111111111111111101011100101101;
assign LUT_1[4689] = 32'b11111111111111110110101110101001;
assign LUT_1[4690] = 32'b11111111111111111001001010111110;
assign LUT_1[4691] = 32'b11111111111111110010011100111010;
assign LUT_1[4692] = 32'b00000000000000000101010110000100;
assign LUT_1[4693] = 32'b11111111111111111110101000000000;
assign LUT_1[4694] = 32'b00000000000000000001000100010101;
assign LUT_1[4695] = 32'b11111111111111111010010110010001;
assign LUT_1[4696] = 32'b11111111111111111100101010100010;
assign LUT_1[4697] = 32'b11111111111111110101111100011110;
assign LUT_1[4698] = 32'b11111111111111111000011000110011;
assign LUT_1[4699] = 32'b11111111111111110001101010101111;
assign LUT_1[4700] = 32'b00000000000000000100100011111001;
assign LUT_1[4701] = 32'b11111111111111111101110101110101;
assign LUT_1[4702] = 32'b00000000000000000000010010001010;
assign LUT_1[4703] = 32'b11111111111111111001100100000110;
assign LUT_1[4704] = 32'b11111111111111111100011100001010;
assign LUT_1[4705] = 32'b11111111111111110101101110000110;
assign LUT_1[4706] = 32'b11111111111111111000001010011011;
assign LUT_1[4707] = 32'b11111111111111110001011100010111;
assign LUT_1[4708] = 32'b00000000000000000100010101100001;
assign LUT_1[4709] = 32'b11111111111111111101100111011101;
assign LUT_1[4710] = 32'b00000000000000000000000011110010;
assign LUT_1[4711] = 32'b11111111111111111001010101101110;
assign LUT_1[4712] = 32'b11111111111111111011101001111111;
assign LUT_1[4713] = 32'b11111111111111110100111011111011;
assign LUT_1[4714] = 32'b11111111111111110111011000010000;
assign LUT_1[4715] = 32'b11111111111111110000101010001100;
assign LUT_1[4716] = 32'b00000000000000000011100011010110;
assign LUT_1[4717] = 32'b11111111111111111100110101010010;
assign LUT_1[4718] = 32'b11111111111111111111010001100111;
assign LUT_1[4719] = 32'b11111111111111111000100011100011;
assign LUT_1[4720] = 32'b11111111111111111110010111101100;
assign LUT_1[4721] = 32'b11111111111111110111101001101000;
assign LUT_1[4722] = 32'b11111111111111111010000101111101;
assign LUT_1[4723] = 32'b11111111111111110011010111111001;
assign LUT_1[4724] = 32'b00000000000000000110010001000011;
assign LUT_1[4725] = 32'b11111111111111111111100010111111;
assign LUT_1[4726] = 32'b00000000000000000001111111010100;
assign LUT_1[4727] = 32'b11111111111111111011010001010000;
assign LUT_1[4728] = 32'b11111111111111111101100101100001;
assign LUT_1[4729] = 32'b11111111111111110110110111011101;
assign LUT_1[4730] = 32'b11111111111111111001010011110010;
assign LUT_1[4731] = 32'b11111111111111110010100101101110;
assign LUT_1[4732] = 32'b00000000000000000101011110111000;
assign LUT_1[4733] = 32'b11111111111111111110110000110100;
assign LUT_1[4734] = 32'b00000000000000000001001101001001;
assign LUT_1[4735] = 32'b11111111111111111010011111000101;
assign LUT_1[4736] = 32'b11111111111111111100100011100110;
assign LUT_1[4737] = 32'b11111111111111110101110101100010;
assign LUT_1[4738] = 32'b11111111111111111000010001110111;
assign LUT_1[4739] = 32'b11111111111111110001100011110011;
assign LUT_1[4740] = 32'b00000000000000000100011100111101;
assign LUT_1[4741] = 32'b11111111111111111101101110111001;
assign LUT_1[4742] = 32'b00000000000000000000001011001110;
assign LUT_1[4743] = 32'b11111111111111111001011101001010;
assign LUT_1[4744] = 32'b11111111111111111011110001011011;
assign LUT_1[4745] = 32'b11111111111111110101000011010111;
assign LUT_1[4746] = 32'b11111111111111110111011111101100;
assign LUT_1[4747] = 32'b11111111111111110000110001101000;
assign LUT_1[4748] = 32'b00000000000000000011101010110010;
assign LUT_1[4749] = 32'b11111111111111111100111100101110;
assign LUT_1[4750] = 32'b11111111111111111111011001000011;
assign LUT_1[4751] = 32'b11111111111111111000101010111111;
assign LUT_1[4752] = 32'b11111111111111111110011111001000;
assign LUT_1[4753] = 32'b11111111111111110111110001000100;
assign LUT_1[4754] = 32'b11111111111111111010001101011001;
assign LUT_1[4755] = 32'b11111111111111110011011111010101;
assign LUT_1[4756] = 32'b00000000000000000110011000011111;
assign LUT_1[4757] = 32'b11111111111111111111101010011011;
assign LUT_1[4758] = 32'b00000000000000000010000110110000;
assign LUT_1[4759] = 32'b11111111111111111011011000101100;
assign LUT_1[4760] = 32'b11111111111111111101101100111101;
assign LUT_1[4761] = 32'b11111111111111110110111110111001;
assign LUT_1[4762] = 32'b11111111111111111001011011001110;
assign LUT_1[4763] = 32'b11111111111111110010101101001010;
assign LUT_1[4764] = 32'b00000000000000000101100110010100;
assign LUT_1[4765] = 32'b11111111111111111110111000010000;
assign LUT_1[4766] = 32'b00000000000000000001010100100101;
assign LUT_1[4767] = 32'b11111111111111111010100110100001;
assign LUT_1[4768] = 32'b11111111111111111101011110100101;
assign LUT_1[4769] = 32'b11111111111111110110110000100001;
assign LUT_1[4770] = 32'b11111111111111111001001100110110;
assign LUT_1[4771] = 32'b11111111111111110010011110110010;
assign LUT_1[4772] = 32'b00000000000000000101010111111100;
assign LUT_1[4773] = 32'b11111111111111111110101001111000;
assign LUT_1[4774] = 32'b00000000000000000001000110001101;
assign LUT_1[4775] = 32'b11111111111111111010011000001001;
assign LUT_1[4776] = 32'b11111111111111111100101100011010;
assign LUT_1[4777] = 32'b11111111111111110101111110010110;
assign LUT_1[4778] = 32'b11111111111111111000011010101011;
assign LUT_1[4779] = 32'b11111111111111110001101100100111;
assign LUT_1[4780] = 32'b00000000000000000100100101110001;
assign LUT_1[4781] = 32'b11111111111111111101110111101101;
assign LUT_1[4782] = 32'b00000000000000000000010100000010;
assign LUT_1[4783] = 32'b11111111111111111001100101111110;
assign LUT_1[4784] = 32'b11111111111111111111011010000111;
assign LUT_1[4785] = 32'b11111111111111111000101100000011;
assign LUT_1[4786] = 32'b11111111111111111011001000011000;
assign LUT_1[4787] = 32'b11111111111111110100011010010100;
assign LUT_1[4788] = 32'b00000000000000000111010011011110;
assign LUT_1[4789] = 32'b00000000000000000000100101011010;
assign LUT_1[4790] = 32'b00000000000000000011000001101111;
assign LUT_1[4791] = 32'b11111111111111111100010011101011;
assign LUT_1[4792] = 32'b11111111111111111110100111111100;
assign LUT_1[4793] = 32'b11111111111111110111111001111000;
assign LUT_1[4794] = 32'b11111111111111111010010110001101;
assign LUT_1[4795] = 32'b11111111111111110011101000001001;
assign LUT_1[4796] = 32'b00000000000000000110100001010011;
assign LUT_1[4797] = 32'b11111111111111111111110011001111;
assign LUT_1[4798] = 32'b00000000000000000010001111100100;
assign LUT_1[4799] = 32'b11111111111111111011100001100000;
assign LUT_1[4800] = 32'b11111111111111111110100001001110;
assign LUT_1[4801] = 32'b11111111111111110111110011001010;
assign LUT_1[4802] = 32'b11111111111111111010001111011111;
assign LUT_1[4803] = 32'b11111111111111110011100001011011;
assign LUT_1[4804] = 32'b00000000000000000110011010100101;
assign LUT_1[4805] = 32'b11111111111111111111101100100001;
assign LUT_1[4806] = 32'b00000000000000000010001000110110;
assign LUT_1[4807] = 32'b11111111111111111011011010110010;
assign LUT_1[4808] = 32'b11111111111111111101101111000011;
assign LUT_1[4809] = 32'b11111111111111110111000000111111;
assign LUT_1[4810] = 32'b11111111111111111001011101010100;
assign LUT_1[4811] = 32'b11111111111111110010101111010000;
assign LUT_1[4812] = 32'b00000000000000000101101000011010;
assign LUT_1[4813] = 32'b11111111111111111110111010010110;
assign LUT_1[4814] = 32'b00000000000000000001010110101011;
assign LUT_1[4815] = 32'b11111111111111111010101000100111;
assign LUT_1[4816] = 32'b00000000000000000000011100110000;
assign LUT_1[4817] = 32'b11111111111111111001101110101100;
assign LUT_1[4818] = 32'b11111111111111111100001011000001;
assign LUT_1[4819] = 32'b11111111111111110101011100111101;
assign LUT_1[4820] = 32'b00000000000000001000010110000111;
assign LUT_1[4821] = 32'b00000000000000000001101000000011;
assign LUT_1[4822] = 32'b00000000000000000100000100011000;
assign LUT_1[4823] = 32'b11111111111111111101010110010100;
assign LUT_1[4824] = 32'b11111111111111111111101010100101;
assign LUT_1[4825] = 32'b11111111111111111000111100100001;
assign LUT_1[4826] = 32'b11111111111111111011011000110110;
assign LUT_1[4827] = 32'b11111111111111110100101010110010;
assign LUT_1[4828] = 32'b00000000000000000111100011111100;
assign LUT_1[4829] = 32'b00000000000000000000110101111000;
assign LUT_1[4830] = 32'b00000000000000000011010010001101;
assign LUT_1[4831] = 32'b11111111111111111100100100001001;
assign LUT_1[4832] = 32'b11111111111111111111011100001101;
assign LUT_1[4833] = 32'b11111111111111111000101110001001;
assign LUT_1[4834] = 32'b11111111111111111011001010011110;
assign LUT_1[4835] = 32'b11111111111111110100011100011010;
assign LUT_1[4836] = 32'b00000000000000000111010101100100;
assign LUT_1[4837] = 32'b00000000000000000000100111100000;
assign LUT_1[4838] = 32'b00000000000000000011000011110101;
assign LUT_1[4839] = 32'b11111111111111111100010101110001;
assign LUT_1[4840] = 32'b11111111111111111110101010000010;
assign LUT_1[4841] = 32'b11111111111111110111111011111110;
assign LUT_1[4842] = 32'b11111111111111111010011000010011;
assign LUT_1[4843] = 32'b11111111111111110011101010001111;
assign LUT_1[4844] = 32'b00000000000000000110100011011001;
assign LUT_1[4845] = 32'b11111111111111111111110101010101;
assign LUT_1[4846] = 32'b00000000000000000010010001101010;
assign LUT_1[4847] = 32'b11111111111111111011100011100110;
assign LUT_1[4848] = 32'b00000000000000000001010111101111;
assign LUT_1[4849] = 32'b11111111111111111010101001101011;
assign LUT_1[4850] = 32'b11111111111111111101000110000000;
assign LUT_1[4851] = 32'b11111111111111110110010111111100;
assign LUT_1[4852] = 32'b00000000000000001001010001000110;
assign LUT_1[4853] = 32'b00000000000000000010100011000010;
assign LUT_1[4854] = 32'b00000000000000000100111111010111;
assign LUT_1[4855] = 32'b11111111111111111110010001010011;
assign LUT_1[4856] = 32'b00000000000000000000100101100100;
assign LUT_1[4857] = 32'b11111111111111111001110111100000;
assign LUT_1[4858] = 32'b11111111111111111100010011110101;
assign LUT_1[4859] = 32'b11111111111111110101100101110001;
assign LUT_1[4860] = 32'b00000000000000001000011110111011;
assign LUT_1[4861] = 32'b00000000000000000001110000110111;
assign LUT_1[4862] = 32'b00000000000000000100001101001100;
assign LUT_1[4863] = 32'b11111111111111111101011111001000;
assign LUT_1[4864] = 32'b11111111111111110111010111101111;
assign LUT_1[4865] = 32'b11111111111111110000101001101011;
assign LUT_1[4866] = 32'b11111111111111110011000110000000;
assign LUT_1[4867] = 32'b11111111111111101100010111111100;
assign LUT_1[4868] = 32'b11111111111111111111010001000110;
assign LUT_1[4869] = 32'b11111111111111111000100011000010;
assign LUT_1[4870] = 32'b11111111111111111010111111010111;
assign LUT_1[4871] = 32'b11111111111111110100010001010011;
assign LUT_1[4872] = 32'b11111111111111110110100101100100;
assign LUT_1[4873] = 32'b11111111111111101111110111100000;
assign LUT_1[4874] = 32'b11111111111111110010010011110101;
assign LUT_1[4875] = 32'b11111111111111101011100101110001;
assign LUT_1[4876] = 32'b11111111111111111110011110111011;
assign LUT_1[4877] = 32'b11111111111111110111110000110111;
assign LUT_1[4878] = 32'b11111111111111111010001101001100;
assign LUT_1[4879] = 32'b11111111111111110011011111001000;
assign LUT_1[4880] = 32'b11111111111111111001010011010001;
assign LUT_1[4881] = 32'b11111111111111110010100101001101;
assign LUT_1[4882] = 32'b11111111111111110101000001100010;
assign LUT_1[4883] = 32'b11111111111111101110010011011110;
assign LUT_1[4884] = 32'b00000000000000000001001100101000;
assign LUT_1[4885] = 32'b11111111111111111010011110100100;
assign LUT_1[4886] = 32'b11111111111111111100111010111001;
assign LUT_1[4887] = 32'b11111111111111110110001100110101;
assign LUT_1[4888] = 32'b11111111111111111000100001000110;
assign LUT_1[4889] = 32'b11111111111111110001110011000010;
assign LUT_1[4890] = 32'b11111111111111110100001111010111;
assign LUT_1[4891] = 32'b11111111111111101101100001010011;
assign LUT_1[4892] = 32'b00000000000000000000011010011101;
assign LUT_1[4893] = 32'b11111111111111111001101100011001;
assign LUT_1[4894] = 32'b11111111111111111100001000101110;
assign LUT_1[4895] = 32'b11111111111111110101011010101010;
assign LUT_1[4896] = 32'b11111111111111111000010010101110;
assign LUT_1[4897] = 32'b11111111111111110001100100101010;
assign LUT_1[4898] = 32'b11111111111111110100000000111111;
assign LUT_1[4899] = 32'b11111111111111101101010010111011;
assign LUT_1[4900] = 32'b00000000000000000000001100000101;
assign LUT_1[4901] = 32'b11111111111111111001011110000001;
assign LUT_1[4902] = 32'b11111111111111111011111010010110;
assign LUT_1[4903] = 32'b11111111111111110101001100010010;
assign LUT_1[4904] = 32'b11111111111111110111100000100011;
assign LUT_1[4905] = 32'b11111111111111110000110010011111;
assign LUT_1[4906] = 32'b11111111111111110011001110110100;
assign LUT_1[4907] = 32'b11111111111111101100100000110000;
assign LUT_1[4908] = 32'b11111111111111111111011001111010;
assign LUT_1[4909] = 32'b11111111111111111000101011110110;
assign LUT_1[4910] = 32'b11111111111111111011001000001011;
assign LUT_1[4911] = 32'b11111111111111110100011010000111;
assign LUT_1[4912] = 32'b11111111111111111010001110010000;
assign LUT_1[4913] = 32'b11111111111111110011100000001100;
assign LUT_1[4914] = 32'b11111111111111110101111100100001;
assign LUT_1[4915] = 32'b11111111111111101111001110011101;
assign LUT_1[4916] = 32'b00000000000000000010000111100111;
assign LUT_1[4917] = 32'b11111111111111111011011001100011;
assign LUT_1[4918] = 32'b11111111111111111101110101111000;
assign LUT_1[4919] = 32'b11111111111111110111000111110100;
assign LUT_1[4920] = 32'b11111111111111111001011100000101;
assign LUT_1[4921] = 32'b11111111111111110010101110000001;
assign LUT_1[4922] = 32'b11111111111111110101001010010110;
assign LUT_1[4923] = 32'b11111111111111101110011100010010;
assign LUT_1[4924] = 32'b00000000000000000001010101011100;
assign LUT_1[4925] = 32'b11111111111111111010100111011000;
assign LUT_1[4926] = 32'b11111111111111111101000011101101;
assign LUT_1[4927] = 32'b11111111111111110110010101101001;
assign LUT_1[4928] = 32'b11111111111111111001010101010111;
assign LUT_1[4929] = 32'b11111111111111110010100111010011;
assign LUT_1[4930] = 32'b11111111111111110101000011101000;
assign LUT_1[4931] = 32'b11111111111111101110010101100100;
assign LUT_1[4932] = 32'b00000000000000000001001110101110;
assign LUT_1[4933] = 32'b11111111111111111010100000101010;
assign LUT_1[4934] = 32'b11111111111111111100111100111111;
assign LUT_1[4935] = 32'b11111111111111110110001110111011;
assign LUT_1[4936] = 32'b11111111111111111000100011001100;
assign LUT_1[4937] = 32'b11111111111111110001110101001000;
assign LUT_1[4938] = 32'b11111111111111110100010001011101;
assign LUT_1[4939] = 32'b11111111111111101101100011011001;
assign LUT_1[4940] = 32'b00000000000000000000011100100011;
assign LUT_1[4941] = 32'b11111111111111111001101110011111;
assign LUT_1[4942] = 32'b11111111111111111100001010110100;
assign LUT_1[4943] = 32'b11111111111111110101011100110000;
assign LUT_1[4944] = 32'b11111111111111111011010000111001;
assign LUT_1[4945] = 32'b11111111111111110100100010110101;
assign LUT_1[4946] = 32'b11111111111111110110111111001010;
assign LUT_1[4947] = 32'b11111111111111110000010001000110;
assign LUT_1[4948] = 32'b00000000000000000011001010010000;
assign LUT_1[4949] = 32'b11111111111111111100011100001100;
assign LUT_1[4950] = 32'b11111111111111111110111000100001;
assign LUT_1[4951] = 32'b11111111111111111000001010011101;
assign LUT_1[4952] = 32'b11111111111111111010011110101110;
assign LUT_1[4953] = 32'b11111111111111110011110000101010;
assign LUT_1[4954] = 32'b11111111111111110110001100111111;
assign LUT_1[4955] = 32'b11111111111111101111011110111011;
assign LUT_1[4956] = 32'b00000000000000000010011000000101;
assign LUT_1[4957] = 32'b11111111111111111011101010000001;
assign LUT_1[4958] = 32'b11111111111111111110000110010110;
assign LUT_1[4959] = 32'b11111111111111110111011000010010;
assign LUT_1[4960] = 32'b11111111111111111010010000010110;
assign LUT_1[4961] = 32'b11111111111111110011100010010010;
assign LUT_1[4962] = 32'b11111111111111110101111110100111;
assign LUT_1[4963] = 32'b11111111111111101111010000100011;
assign LUT_1[4964] = 32'b00000000000000000010001001101101;
assign LUT_1[4965] = 32'b11111111111111111011011011101001;
assign LUT_1[4966] = 32'b11111111111111111101110111111110;
assign LUT_1[4967] = 32'b11111111111111110111001001111010;
assign LUT_1[4968] = 32'b11111111111111111001011110001011;
assign LUT_1[4969] = 32'b11111111111111110010110000000111;
assign LUT_1[4970] = 32'b11111111111111110101001100011100;
assign LUT_1[4971] = 32'b11111111111111101110011110011000;
assign LUT_1[4972] = 32'b00000000000000000001010111100010;
assign LUT_1[4973] = 32'b11111111111111111010101001011110;
assign LUT_1[4974] = 32'b11111111111111111101000101110011;
assign LUT_1[4975] = 32'b11111111111111110110010111101111;
assign LUT_1[4976] = 32'b11111111111111111100001011111000;
assign LUT_1[4977] = 32'b11111111111111110101011101110100;
assign LUT_1[4978] = 32'b11111111111111110111111010001001;
assign LUT_1[4979] = 32'b11111111111111110001001100000101;
assign LUT_1[4980] = 32'b00000000000000000100000101001111;
assign LUT_1[4981] = 32'b11111111111111111101010111001011;
assign LUT_1[4982] = 32'b11111111111111111111110011100000;
assign LUT_1[4983] = 32'b11111111111111111001000101011100;
assign LUT_1[4984] = 32'b11111111111111111011011001101101;
assign LUT_1[4985] = 32'b11111111111111110100101011101001;
assign LUT_1[4986] = 32'b11111111111111110111000111111110;
assign LUT_1[4987] = 32'b11111111111111110000011001111010;
assign LUT_1[4988] = 32'b00000000000000000011010011000100;
assign LUT_1[4989] = 32'b11111111111111111100100101000000;
assign LUT_1[4990] = 32'b11111111111111111111000001010101;
assign LUT_1[4991] = 32'b11111111111111111000010011010001;
assign LUT_1[4992] = 32'b11111111111111111010010111110010;
assign LUT_1[4993] = 32'b11111111111111110011101001101110;
assign LUT_1[4994] = 32'b11111111111111110110000110000011;
assign LUT_1[4995] = 32'b11111111111111101111010111111111;
assign LUT_1[4996] = 32'b00000000000000000010010001001001;
assign LUT_1[4997] = 32'b11111111111111111011100011000101;
assign LUT_1[4998] = 32'b11111111111111111101111111011010;
assign LUT_1[4999] = 32'b11111111111111110111010001010110;
assign LUT_1[5000] = 32'b11111111111111111001100101100111;
assign LUT_1[5001] = 32'b11111111111111110010110111100011;
assign LUT_1[5002] = 32'b11111111111111110101010011111000;
assign LUT_1[5003] = 32'b11111111111111101110100101110100;
assign LUT_1[5004] = 32'b00000000000000000001011110111110;
assign LUT_1[5005] = 32'b11111111111111111010110000111010;
assign LUT_1[5006] = 32'b11111111111111111101001101001111;
assign LUT_1[5007] = 32'b11111111111111110110011111001011;
assign LUT_1[5008] = 32'b11111111111111111100010011010100;
assign LUT_1[5009] = 32'b11111111111111110101100101010000;
assign LUT_1[5010] = 32'b11111111111111111000000001100101;
assign LUT_1[5011] = 32'b11111111111111110001010011100001;
assign LUT_1[5012] = 32'b00000000000000000100001100101011;
assign LUT_1[5013] = 32'b11111111111111111101011110100111;
assign LUT_1[5014] = 32'b11111111111111111111111010111100;
assign LUT_1[5015] = 32'b11111111111111111001001100111000;
assign LUT_1[5016] = 32'b11111111111111111011100001001001;
assign LUT_1[5017] = 32'b11111111111111110100110011000101;
assign LUT_1[5018] = 32'b11111111111111110111001111011010;
assign LUT_1[5019] = 32'b11111111111111110000100001010110;
assign LUT_1[5020] = 32'b00000000000000000011011010100000;
assign LUT_1[5021] = 32'b11111111111111111100101100011100;
assign LUT_1[5022] = 32'b11111111111111111111001000110001;
assign LUT_1[5023] = 32'b11111111111111111000011010101101;
assign LUT_1[5024] = 32'b11111111111111111011010010110001;
assign LUT_1[5025] = 32'b11111111111111110100100100101101;
assign LUT_1[5026] = 32'b11111111111111110111000001000010;
assign LUT_1[5027] = 32'b11111111111111110000010010111110;
assign LUT_1[5028] = 32'b00000000000000000011001100001000;
assign LUT_1[5029] = 32'b11111111111111111100011110000100;
assign LUT_1[5030] = 32'b11111111111111111110111010011001;
assign LUT_1[5031] = 32'b11111111111111111000001100010101;
assign LUT_1[5032] = 32'b11111111111111111010100000100110;
assign LUT_1[5033] = 32'b11111111111111110011110010100010;
assign LUT_1[5034] = 32'b11111111111111110110001110110111;
assign LUT_1[5035] = 32'b11111111111111101111100000110011;
assign LUT_1[5036] = 32'b00000000000000000010011001111101;
assign LUT_1[5037] = 32'b11111111111111111011101011111001;
assign LUT_1[5038] = 32'b11111111111111111110001000001110;
assign LUT_1[5039] = 32'b11111111111111110111011010001010;
assign LUT_1[5040] = 32'b11111111111111111101001110010011;
assign LUT_1[5041] = 32'b11111111111111110110100000001111;
assign LUT_1[5042] = 32'b11111111111111111000111100100100;
assign LUT_1[5043] = 32'b11111111111111110010001110100000;
assign LUT_1[5044] = 32'b00000000000000000101000111101010;
assign LUT_1[5045] = 32'b11111111111111111110011001100110;
assign LUT_1[5046] = 32'b00000000000000000000110101111011;
assign LUT_1[5047] = 32'b11111111111111111010000111110111;
assign LUT_1[5048] = 32'b11111111111111111100011100001000;
assign LUT_1[5049] = 32'b11111111111111110101101110000100;
assign LUT_1[5050] = 32'b11111111111111111000001010011001;
assign LUT_1[5051] = 32'b11111111111111110001011100010101;
assign LUT_1[5052] = 32'b00000000000000000100010101011111;
assign LUT_1[5053] = 32'b11111111111111111101100111011011;
assign LUT_1[5054] = 32'b00000000000000000000000011110000;
assign LUT_1[5055] = 32'b11111111111111111001010101101100;
assign LUT_1[5056] = 32'b11111111111111111100010101011010;
assign LUT_1[5057] = 32'b11111111111111110101100111010110;
assign LUT_1[5058] = 32'b11111111111111111000000011101011;
assign LUT_1[5059] = 32'b11111111111111110001010101100111;
assign LUT_1[5060] = 32'b00000000000000000100001110110001;
assign LUT_1[5061] = 32'b11111111111111111101100000101101;
assign LUT_1[5062] = 32'b11111111111111111111111101000010;
assign LUT_1[5063] = 32'b11111111111111111001001110111110;
assign LUT_1[5064] = 32'b11111111111111111011100011001111;
assign LUT_1[5065] = 32'b11111111111111110100110101001011;
assign LUT_1[5066] = 32'b11111111111111110111010001100000;
assign LUT_1[5067] = 32'b11111111111111110000100011011100;
assign LUT_1[5068] = 32'b00000000000000000011011100100110;
assign LUT_1[5069] = 32'b11111111111111111100101110100010;
assign LUT_1[5070] = 32'b11111111111111111111001010110111;
assign LUT_1[5071] = 32'b11111111111111111000011100110011;
assign LUT_1[5072] = 32'b11111111111111111110010000111100;
assign LUT_1[5073] = 32'b11111111111111110111100010111000;
assign LUT_1[5074] = 32'b11111111111111111001111111001101;
assign LUT_1[5075] = 32'b11111111111111110011010001001001;
assign LUT_1[5076] = 32'b00000000000000000110001010010011;
assign LUT_1[5077] = 32'b11111111111111111111011100001111;
assign LUT_1[5078] = 32'b00000000000000000001111000100100;
assign LUT_1[5079] = 32'b11111111111111111011001010100000;
assign LUT_1[5080] = 32'b11111111111111111101011110110001;
assign LUT_1[5081] = 32'b11111111111111110110110000101101;
assign LUT_1[5082] = 32'b11111111111111111001001101000010;
assign LUT_1[5083] = 32'b11111111111111110010011110111110;
assign LUT_1[5084] = 32'b00000000000000000101011000001000;
assign LUT_1[5085] = 32'b11111111111111111110101010000100;
assign LUT_1[5086] = 32'b00000000000000000001000110011001;
assign LUT_1[5087] = 32'b11111111111111111010011000010101;
assign LUT_1[5088] = 32'b11111111111111111101010000011001;
assign LUT_1[5089] = 32'b11111111111111110110100010010101;
assign LUT_1[5090] = 32'b11111111111111111000111110101010;
assign LUT_1[5091] = 32'b11111111111111110010010000100110;
assign LUT_1[5092] = 32'b00000000000000000101001001110000;
assign LUT_1[5093] = 32'b11111111111111111110011011101100;
assign LUT_1[5094] = 32'b00000000000000000000111000000001;
assign LUT_1[5095] = 32'b11111111111111111010001001111101;
assign LUT_1[5096] = 32'b11111111111111111100011110001110;
assign LUT_1[5097] = 32'b11111111111111110101110000001010;
assign LUT_1[5098] = 32'b11111111111111111000001100011111;
assign LUT_1[5099] = 32'b11111111111111110001011110011011;
assign LUT_1[5100] = 32'b00000000000000000100010111100101;
assign LUT_1[5101] = 32'b11111111111111111101101001100001;
assign LUT_1[5102] = 32'b00000000000000000000000101110110;
assign LUT_1[5103] = 32'b11111111111111111001010111110010;
assign LUT_1[5104] = 32'b11111111111111111111001011111011;
assign LUT_1[5105] = 32'b11111111111111111000011101110111;
assign LUT_1[5106] = 32'b11111111111111111010111010001100;
assign LUT_1[5107] = 32'b11111111111111110100001100001000;
assign LUT_1[5108] = 32'b00000000000000000111000101010010;
assign LUT_1[5109] = 32'b00000000000000000000010111001110;
assign LUT_1[5110] = 32'b00000000000000000010110011100011;
assign LUT_1[5111] = 32'b11111111111111111100000101011111;
assign LUT_1[5112] = 32'b11111111111111111110011001110000;
assign LUT_1[5113] = 32'b11111111111111110111101011101100;
assign LUT_1[5114] = 32'b11111111111111111010001000000001;
assign LUT_1[5115] = 32'b11111111111111110011011001111101;
assign LUT_1[5116] = 32'b00000000000000000110010011000111;
assign LUT_1[5117] = 32'b11111111111111111111100101000011;
assign LUT_1[5118] = 32'b00000000000000000010000001011000;
assign LUT_1[5119] = 32'b11111111111111111011010011010100;
assign LUT_1[5120] = 32'b00000000000000000110001011110110;
assign LUT_1[5121] = 32'b11111111111111111111011101110010;
assign LUT_1[5122] = 32'b00000000000000000001111010000111;
assign LUT_1[5123] = 32'b11111111111111111011001100000011;
assign LUT_1[5124] = 32'b00000000000000001110000101001101;
assign LUT_1[5125] = 32'b00000000000000000111010111001001;
assign LUT_1[5126] = 32'b00000000000000001001110011011110;
assign LUT_1[5127] = 32'b00000000000000000011000101011010;
assign LUT_1[5128] = 32'b00000000000000000101011001101011;
assign LUT_1[5129] = 32'b11111111111111111110101011100111;
assign LUT_1[5130] = 32'b00000000000000000001000111111100;
assign LUT_1[5131] = 32'b11111111111111111010011001111000;
assign LUT_1[5132] = 32'b00000000000000001101010011000010;
assign LUT_1[5133] = 32'b00000000000000000110100100111110;
assign LUT_1[5134] = 32'b00000000000000001001000001010011;
assign LUT_1[5135] = 32'b00000000000000000010010011001111;
assign LUT_1[5136] = 32'b00000000000000001000000111011000;
assign LUT_1[5137] = 32'b00000000000000000001011001010100;
assign LUT_1[5138] = 32'b00000000000000000011110101101001;
assign LUT_1[5139] = 32'b11111111111111111101000111100101;
assign LUT_1[5140] = 32'b00000000000000010000000000101111;
assign LUT_1[5141] = 32'b00000000000000001001010010101011;
assign LUT_1[5142] = 32'b00000000000000001011101111000000;
assign LUT_1[5143] = 32'b00000000000000000101000000111100;
assign LUT_1[5144] = 32'b00000000000000000111010101001101;
assign LUT_1[5145] = 32'b00000000000000000000100111001001;
assign LUT_1[5146] = 32'b00000000000000000011000011011110;
assign LUT_1[5147] = 32'b11111111111111111100010101011010;
assign LUT_1[5148] = 32'b00000000000000001111001110100100;
assign LUT_1[5149] = 32'b00000000000000001000100000100000;
assign LUT_1[5150] = 32'b00000000000000001010111100110101;
assign LUT_1[5151] = 32'b00000000000000000100001110110001;
assign LUT_1[5152] = 32'b00000000000000000111000110110101;
assign LUT_1[5153] = 32'b00000000000000000000011000110001;
assign LUT_1[5154] = 32'b00000000000000000010110101000110;
assign LUT_1[5155] = 32'b11111111111111111100000111000010;
assign LUT_1[5156] = 32'b00000000000000001111000000001100;
assign LUT_1[5157] = 32'b00000000000000001000010010001000;
assign LUT_1[5158] = 32'b00000000000000001010101110011101;
assign LUT_1[5159] = 32'b00000000000000000100000000011001;
assign LUT_1[5160] = 32'b00000000000000000110010100101010;
assign LUT_1[5161] = 32'b11111111111111111111100110100110;
assign LUT_1[5162] = 32'b00000000000000000010000010111011;
assign LUT_1[5163] = 32'b11111111111111111011010100110111;
assign LUT_1[5164] = 32'b00000000000000001110001110000001;
assign LUT_1[5165] = 32'b00000000000000000111011111111101;
assign LUT_1[5166] = 32'b00000000000000001001111100010010;
assign LUT_1[5167] = 32'b00000000000000000011001110001110;
assign LUT_1[5168] = 32'b00000000000000001001000010010111;
assign LUT_1[5169] = 32'b00000000000000000010010100010011;
assign LUT_1[5170] = 32'b00000000000000000100110000101000;
assign LUT_1[5171] = 32'b11111111111111111110000010100100;
assign LUT_1[5172] = 32'b00000000000000010000111011101110;
assign LUT_1[5173] = 32'b00000000000000001010001101101010;
assign LUT_1[5174] = 32'b00000000000000001100101001111111;
assign LUT_1[5175] = 32'b00000000000000000101111011111011;
assign LUT_1[5176] = 32'b00000000000000001000010000001100;
assign LUT_1[5177] = 32'b00000000000000000001100010001000;
assign LUT_1[5178] = 32'b00000000000000000011111110011101;
assign LUT_1[5179] = 32'b11111111111111111101010000011001;
assign LUT_1[5180] = 32'b00000000000000010000001001100011;
assign LUT_1[5181] = 32'b00000000000000001001011011011111;
assign LUT_1[5182] = 32'b00000000000000001011110111110100;
assign LUT_1[5183] = 32'b00000000000000000101001001110000;
assign LUT_1[5184] = 32'b00000000000000001000001001011110;
assign LUT_1[5185] = 32'b00000000000000000001011011011010;
assign LUT_1[5186] = 32'b00000000000000000011110111101111;
assign LUT_1[5187] = 32'b11111111111111111101001001101011;
assign LUT_1[5188] = 32'b00000000000000010000000010110101;
assign LUT_1[5189] = 32'b00000000000000001001010100110001;
assign LUT_1[5190] = 32'b00000000000000001011110001000110;
assign LUT_1[5191] = 32'b00000000000000000101000011000010;
assign LUT_1[5192] = 32'b00000000000000000111010111010011;
assign LUT_1[5193] = 32'b00000000000000000000101001001111;
assign LUT_1[5194] = 32'b00000000000000000011000101100100;
assign LUT_1[5195] = 32'b11111111111111111100010111100000;
assign LUT_1[5196] = 32'b00000000000000001111010000101010;
assign LUT_1[5197] = 32'b00000000000000001000100010100110;
assign LUT_1[5198] = 32'b00000000000000001010111110111011;
assign LUT_1[5199] = 32'b00000000000000000100010000110111;
assign LUT_1[5200] = 32'b00000000000000001010000101000000;
assign LUT_1[5201] = 32'b00000000000000000011010110111100;
assign LUT_1[5202] = 32'b00000000000000000101110011010001;
assign LUT_1[5203] = 32'b11111111111111111111000101001101;
assign LUT_1[5204] = 32'b00000000000000010001111110010111;
assign LUT_1[5205] = 32'b00000000000000001011010000010011;
assign LUT_1[5206] = 32'b00000000000000001101101100101000;
assign LUT_1[5207] = 32'b00000000000000000110111110100100;
assign LUT_1[5208] = 32'b00000000000000001001010010110101;
assign LUT_1[5209] = 32'b00000000000000000010100100110001;
assign LUT_1[5210] = 32'b00000000000000000101000001000110;
assign LUT_1[5211] = 32'b11111111111111111110010011000010;
assign LUT_1[5212] = 32'b00000000000000010001001100001100;
assign LUT_1[5213] = 32'b00000000000000001010011110001000;
assign LUT_1[5214] = 32'b00000000000000001100111010011101;
assign LUT_1[5215] = 32'b00000000000000000110001100011001;
assign LUT_1[5216] = 32'b00000000000000001001000100011101;
assign LUT_1[5217] = 32'b00000000000000000010010110011001;
assign LUT_1[5218] = 32'b00000000000000000100110010101110;
assign LUT_1[5219] = 32'b11111111111111111110000100101010;
assign LUT_1[5220] = 32'b00000000000000010000111101110100;
assign LUT_1[5221] = 32'b00000000000000001010001111110000;
assign LUT_1[5222] = 32'b00000000000000001100101100000101;
assign LUT_1[5223] = 32'b00000000000000000101111110000001;
assign LUT_1[5224] = 32'b00000000000000001000010010010010;
assign LUT_1[5225] = 32'b00000000000000000001100100001110;
assign LUT_1[5226] = 32'b00000000000000000100000000100011;
assign LUT_1[5227] = 32'b11111111111111111101010010011111;
assign LUT_1[5228] = 32'b00000000000000010000001011101001;
assign LUT_1[5229] = 32'b00000000000000001001011101100101;
assign LUT_1[5230] = 32'b00000000000000001011111001111010;
assign LUT_1[5231] = 32'b00000000000000000101001011110110;
assign LUT_1[5232] = 32'b00000000000000001010111111111111;
assign LUT_1[5233] = 32'b00000000000000000100010001111011;
assign LUT_1[5234] = 32'b00000000000000000110101110010000;
assign LUT_1[5235] = 32'b00000000000000000000000000001100;
assign LUT_1[5236] = 32'b00000000000000010010111001010110;
assign LUT_1[5237] = 32'b00000000000000001100001011010010;
assign LUT_1[5238] = 32'b00000000000000001110100111100111;
assign LUT_1[5239] = 32'b00000000000000000111111001100011;
assign LUT_1[5240] = 32'b00000000000000001010001101110100;
assign LUT_1[5241] = 32'b00000000000000000011011111110000;
assign LUT_1[5242] = 32'b00000000000000000101111100000101;
assign LUT_1[5243] = 32'b11111111111111111111001110000001;
assign LUT_1[5244] = 32'b00000000000000010010000111001011;
assign LUT_1[5245] = 32'b00000000000000001011011001000111;
assign LUT_1[5246] = 32'b00000000000000001101110101011100;
assign LUT_1[5247] = 32'b00000000000000000111000111011000;
assign LUT_1[5248] = 32'b00000000000000001001001011111001;
assign LUT_1[5249] = 32'b00000000000000000010011101110101;
assign LUT_1[5250] = 32'b00000000000000000100111010001010;
assign LUT_1[5251] = 32'b11111111111111111110001100000110;
assign LUT_1[5252] = 32'b00000000000000010001000101010000;
assign LUT_1[5253] = 32'b00000000000000001010010111001100;
assign LUT_1[5254] = 32'b00000000000000001100110011100001;
assign LUT_1[5255] = 32'b00000000000000000110000101011101;
assign LUT_1[5256] = 32'b00000000000000001000011001101110;
assign LUT_1[5257] = 32'b00000000000000000001101011101010;
assign LUT_1[5258] = 32'b00000000000000000100000111111111;
assign LUT_1[5259] = 32'b11111111111111111101011001111011;
assign LUT_1[5260] = 32'b00000000000000010000010011000101;
assign LUT_1[5261] = 32'b00000000000000001001100101000001;
assign LUT_1[5262] = 32'b00000000000000001100000001010110;
assign LUT_1[5263] = 32'b00000000000000000101010011010010;
assign LUT_1[5264] = 32'b00000000000000001011000111011011;
assign LUT_1[5265] = 32'b00000000000000000100011001010111;
assign LUT_1[5266] = 32'b00000000000000000110110101101100;
assign LUT_1[5267] = 32'b00000000000000000000000111101000;
assign LUT_1[5268] = 32'b00000000000000010011000000110010;
assign LUT_1[5269] = 32'b00000000000000001100010010101110;
assign LUT_1[5270] = 32'b00000000000000001110101111000011;
assign LUT_1[5271] = 32'b00000000000000001000000000111111;
assign LUT_1[5272] = 32'b00000000000000001010010101010000;
assign LUT_1[5273] = 32'b00000000000000000011100111001100;
assign LUT_1[5274] = 32'b00000000000000000110000011100001;
assign LUT_1[5275] = 32'b11111111111111111111010101011101;
assign LUT_1[5276] = 32'b00000000000000010010001110100111;
assign LUT_1[5277] = 32'b00000000000000001011100000100011;
assign LUT_1[5278] = 32'b00000000000000001101111100111000;
assign LUT_1[5279] = 32'b00000000000000000111001110110100;
assign LUT_1[5280] = 32'b00000000000000001010000110111000;
assign LUT_1[5281] = 32'b00000000000000000011011000110100;
assign LUT_1[5282] = 32'b00000000000000000101110101001001;
assign LUT_1[5283] = 32'b11111111111111111111000111000101;
assign LUT_1[5284] = 32'b00000000000000010010000000001111;
assign LUT_1[5285] = 32'b00000000000000001011010010001011;
assign LUT_1[5286] = 32'b00000000000000001101101110100000;
assign LUT_1[5287] = 32'b00000000000000000111000000011100;
assign LUT_1[5288] = 32'b00000000000000001001010100101101;
assign LUT_1[5289] = 32'b00000000000000000010100110101001;
assign LUT_1[5290] = 32'b00000000000000000101000010111110;
assign LUT_1[5291] = 32'b11111111111111111110010100111010;
assign LUT_1[5292] = 32'b00000000000000010001001110000100;
assign LUT_1[5293] = 32'b00000000000000001010100000000000;
assign LUT_1[5294] = 32'b00000000000000001100111100010101;
assign LUT_1[5295] = 32'b00000000000000000110001110010001;
assign LUT_1[5296] = 32'b00000000000000001100000010011010;
assign LUT_1[5297] = 32'b00000000000000000101010100010110;
assign LUT_1[5298] = 32'b00000000000000000111110000101011;
assign LUT_1[5299] = 32'b00000000000000000001000010100111;
assign LUT_1[5300] = 32'b00000000000000010011111011110001;
assign LUT_1[5301] = 32'b00000000000000001101001101101101;
assign LUT_1[5302] = 32'b00000000000000001111101010000010;
assign LUT_1[5303] = 32'b00000000000000001000111011111110;
assign LUT_1[5304] = 32'b00000000000000001011010000001111;
assign LUT_1[5305] = 32'b00000000000000000100100010001011;
assign LUT_1[5306] = 32'b00000000000000000110111110100000;
assign LUT_1[5307] = 32'b00000000000000000000010000011100;
assign LUT_1[5308] = 32'b00000000000000010011001001100110;
assign LUT_1[5309] = 32'b00000000000000001100011011100010;
assign LUT_1[5310] = 32'b00000000000000001110110111110111;
assign LUT_1[5311] = 32'b00000000000000001000001001110011;
assign LUT_1[5312] = 32'b00000000000000001011001001100001;
assign LUT_1[5313] = 32'b00000000000000000100011011011101;
assign LUT_1[5314] = 32'b00000000000000000110110111110010;
assign LUT_1[5315] = 32'b00000000000000000000001001101110;
assign LUT_1[5316] = 32'b00000000000000010011000010111000;
assign LUT_1[5317] = 32'b00000000000000001100010100110100;
assign LUT_1[5318] = 32'b00000000000000001110110001001001;
assign LUT_1[5319] = 32'b00000000000000001000000011000101;
assign LUT_1[5320] = 32'b00000000000000001010010111010110;
assign LUT_1[5321] = 32'b00000000000000000011101001010010;
assign LUT_1[5322] = 32'b00000000000000000110000101100111;
assign LUT_1[5323] = 32'b11111111111111111111010111100011;
assign LUT_1[5324] = 32'b00000000000000010010010000101101;
assign LUT_1[5325] = 32'b00000000000000001011100010101001;
assign LUT_1[5326] = 32'b00000000000000001101111110111110;
assign LUT_1[5327] = 32'b00000000000000000111010000111010;
assign LUT_1[5328] = 32'b00000000000000001101000101000011;
assign LUT_1[5329] = 32'b00000000000000000110010110111111;
assign LUT_1[5330] = 32'b00000000000000001000110011010100;
assign LUT_1[5331] = 32'b00000000000000000010000101010000;
assign LUT_1[5332] = 32'b00000000000000010100111110011010;
assign LUT_1[5333] = 32'b00000000000000001110010000010110;
assign LUT_1[5334] = 32'b00000000000000010000101100101011;
assign LUT_1[5335] = 32'b00000000000000001001111110100111;
assign LUT_1[5336] = 32'b00000000000000001100010010111000;
assign LUT_1[5337] = 32'b00000000000000000101100100110100;
assign LUT_1[5338] = 32'b00000000000000001000000001001001;
assign LUT_1[5339] = 32'b00000000000000000001010011000101;
assign LUT_1[5340] = 32'b00000000000000010100001100001111;
assign LUT_1[5341] = 32'b00000000000000001101011110001011;
assign LUT_1[5342] = 32'b00000000000000001111111010100000;
assign LUT_1[5343] = 32'b00000000000000001001001100011100;
assign LUT_1[5344] = 32'b00000000000000001100000100100000;
assign LUT_1[5345] = 32'b00000000000000000101010110011100;
assign LUT_1[5346] = 32'b00000000000000000111110010110001;
assign LUT_1[5347] = 32'b00000000000000000001000100101101;
assign LUT_1[5348] = 32'b00000000000000010011111101110111;
assign LUT_1[5349] = 32'b00000000000000001101001111110011;
assign LUT_1[5350] = 32'b00000000000000001111101100001000;
assign LUT_1[5351] = 32'b00000000000000001000111110000100;
assign LUT_1[5352] = 32'b00000000000000001011010010010101;
assign LUT_1[5353] = 32'b00000000000000000100100100010001;
assign LUT_1[5354] = 32'b00000000000000000111000000100110;
assign LUT_1[5355] = 32'b00000000000000000000010010100010;
assign LUT_1[5356] = 32'b00000000000000010011001011101100;
assign LUT_1[5357] = 32'b00000000000000001100011101101000;
assign LUT_1[5358] = 32'b00000000000000001110111001111101;
assign LUT_1[5359] = 32'b00000000000000001000001011111001;
assign LUT_1[5360] = 32'b00000000000000001110000000000010;
assign LUT_1[5361] = 32'b00000000000000000111010001111110;
assign LUT_1[5362] = 32'b00000000000000001001101110010011;
assign LUT_1[5363] = 32'b00000000000000000011000000001111;
assign LUT_1[5364] = 32'b00000000000000010101111001011001;
assign LUT_1[5365] = 32'b00000000000000001111001011010101;
assign LUT_1[5366] = 32'b00000000000000010001100111101010;
assign LUT_1[5367] = 32'b00000000000000001010111001100110;
assign LUT_1[5368] = 32'b00000000000000001101001101110111;
assign LUT_1[5369] = 32'b00000000000000000110011111110011;
assign LUT_1[5370] = 32'b00000000000000001000111100001000;
assign LUT_1[5371] = 32'b00000000000000000010001110000100;
assign LUT_1[5372] = 32'b00000000000000010101000111001110;
assign LUT_1[5373] = 32'b00000000000000001110011001001010;
assign LUT_1[5374] = 32'b00000000000000010000110101011111;
assign LUT_1[5375] = 32'b00000000000000001010000111011011;
assign LUT_1[5376] = 32'b00000000000000000100000000000010;
assign LUT_1[5377] = 32'b11111111111111111101010001111110;
assign LUT_1[5378] = 32'b11111111111111111111101110010011;
assign LUT_1[5379] = 32'b11111111111111111001000000001111;
assign LUT_1[5380] = 32'b00000000000000001011111001011001;
assign LUT_1[5381] = 32'b00000000000000000101001011010101;
assign LUT_1[5382] = 32'b00000000000000000111100111101010;
assign LUT_1[5383] = 32'b00000000000000000000111001100110;
assign LUT_1[5384] = 32'b00000000000000000011001101110111;
assign LUT_1[5385] = 32'b11111111111111111100011111110011;
assign LUT_1[5386] = 32'b11111111111111111110111100001000;
assign LUT_1[5387] = 32'b11111111111111111000001110000100;
assign LUT_1[5388] = 32'b00000000000000001011000111001110;
assign LUT_1[5389] = 32'b00000000000000000100011001001010;
assign LUT_1[5390] = 32'b00000000000000000110110101011111;
assign LUT_1[5391] = 32'b00000000000000000000000111011011;
assign LUT_1[5392] = 32'b00000000000000000101111011100100;
assign LUT_1[5393] = 32'b11111111111111111111001101100000;
assign LUT_1[5394] = 32'b00000000000000000001101001110101;
assign LUT_1[5395] = 32'b11111111111111111010111011110001;
assign LUT_1[5396] = 32'b00000000000000001101110100111011;
assign LUT_1[5397] = 32'b00000000000000000111000110110111;
assign LUT_1[5398] = 32'b00000000000000001001100011001100;
assign LUT_1[5399] = 32'b00000000000000000010110101001000;
assign LUT_1[5400] = 32'b00000000000000000101001001011001;
assign LUT_1[5401] = 32'b11111111111111111110011011010101;
assign LUT_1[5402] = 32'b00000000000000000000110111101010;
assign LUT_1[5403] = 32'b11111111111111111010001001100110;
assign LUT_1[5404] = 32'b00000000000000001101000010110000;
assign LUT_1[5405] = 32'b00000000000000000110010100101100;
assign LUT_1[5406] = 32'b00000000000000001000110001000001;
assign LUT_1[5407] = 32'b00000000000000000010000010111101;
assign LUT_1[5408] = 32'b00000000000000000100111011000001;
assign LUT_1[5409] = 32'b11111111111111111110001100111101;
assign LUT_1[5410] = 32'b00000000000000000000101001010010;
assign LUT_1[5411] = 32'b11111111111111111001111011001110;
assign LUT_1[5412] = 32'b00000000000000001100110100011000;
assign LUT_1[5413] = 32'b00000000000000000110000110010100;
assign LUT_1[5414] = 32'b00000000000000001000100010101001;
assign LUT_1[5415] = 32'b00000000000000000001110100100101;
assign LUT_1[5416] = 32'b00000000000000000100001000110110;
assign LUT_1[5417] = 32'b11111111111111111101011010110010;
assign LUT_1[5418] = 32'b11111111111111111111110111000111;
assign LUT_1[5419] = 32'b11111111111111111001001001000011;
assign LUT_1[5420] = 32'b00000000000000001100000010001101;
assign LUT_1[5421] = 32'b00000000000000000101010100001001;
assign LUT_1[5422] = 32'b00000000000000000111110000011110;
assign LUT_1[5423] = 32'b00000000000000000001000010011010;
assign LUT_1[5424] = 32'b00000000000000000110110110100011;
assign LUT_1[5425] = 32'b00000000000000000000001000011111;
assign LUT_1[5426] = 32'b00000000000000000010100100110100;
assign LUT_1[5427] = 32'b11111111111111111011110110110000;
assign LUT_1[5428] = 32'b00000000000000001110101111111010;
assign LUT_1[5429] = 32'b00000000000000001000000001110110;
assign LUT_1[5430] = 32'b00000000000000001010011110001011;
assign LUT_1[5431] = 32'b00000000000000000011110000000111;
assign LUT_1[5432] = 32'b00000000000000000110000100011000;
assign LUT_1[5433] = 32'b11111111111111111111010110010100;
assign LUT_1[5434] = 32'b00000000000000000001110010101001;
assign LUT_1[5435] = 32'b11111111111111111011000100100101;
assign LUT_1[5436] = 32'b00000000000000001101111101101111;
assign LUT_1[5437] = 32'b00000000000000000111001111101011;
assign LUT_1[5438] = 32'b00000000000000001001101100000000;
assign LUT_1[5439] = 32'b00000000000000000010111101111100;
assign LUT_1[5440] = 32'b00000000000000000101111101101010;
assign LUT_1[5441] = 32'b11111111111111111111001111100110;
assign LUT_1[5442] = 32'b00000000000000000001101011111011;
assign LUT_1[5443] = 32'b11111111111111111010111101110111;
assign LUT_1[5444] = 32'b00000000000000001101110111000001;
assign LUT_1[5445] = 32'b00000000000000000111001000111101;
assign LUT_1[5446] = 32'b00000000000000001001100101010010;
assign LUT_1[5447] = 32'b00000000000000000010110111001110;
assign LUT_1[5448] = 32'b00000000000000000101001011011111;
assign LUT_1[5449] = 32'b11111111111111111110011101011011;
assign LUT_1[5450] = 32'b00000000000000000000111001110000;
assign LUT_1[5451] = 32'b11111111111111111010001011101100;
assign LUT_1[5452] = 32'b00000000000000001101000100110110;
assign LUT_1[5453] = 32'b00000000000000000110010110110010;
assign LUT_1[5454] = 32'b00000000000000001000110011000111;
assign LUT_1[5455] = 32'b00000000000000000010000101000011;
assign LUT_1[5456] = 32'b00000000000000000111111001001100;
assign LUT_1[5457] = 32'b00000000000000000001001011001000;
assign LUT_1[5458] = 32'b00000000000000000011100111011101;
assign LUT_1[5459] = 32'b11111111111111111100111001011001;
assign LUT_1[5460] = 32'b00000000000000001111110010100011;
assign LUT_1[5461] = 32'b00000000000000001001000100011111;
assign LUT_1[5462] = 32'b00000000000000001011100000110100;
assign LUT_1[5463] = 32'b00000000000000000100110010110000;
assign LUT_1[5464] = 32'b00000000000000000111000111000001;
assign LUT_1[5465] = 32'b00000000000000000000011000111101;
assign LUT_1[5466] = 32'b00000000000000000010110101010010;
assign LUT_1[5467] = 32'b11111111111111111100000111001110;
assign LUT_1[5468] = 32'b00000000000000001111000000011000;
assign LUT_1[5469] = 32'b00000000000000001000010010010100;
assign LUT_1[5470] = 32'b00000000000000001010101110101001;
assign LUT_1[5471] = 32'b00000000000000000100000000100101;
assign LUT_1[5472] = 32'b00000000000000000110111000101001;
assign LUT_1[5473] = 32'b00000000000000000000001010100101;
assign LUT_1[5474] = 32'b00000000000000000010100110111010;
assign LUT_1[5475] = 32'b11111111111111111011111000110110;
assign LUT_1[5476] = 32'b00000000000000001110110010000000;
assign LUT_1[5477] = 32'b00000000000000001000000011111100;
assign LUT_1[5478] = 32'b00000000000000001010100000010001;
assign LUT_1[5479] = 32'b00000000000000000011110010001101;
assign LUT_1[5480] = 32'b00000000000000000110000110011110;
assign LUT_1[5481] = 32'b11111111111111111111011000011010;
assign LUT_1[5482] = 32'b00000000000000000001110100101111;
assign LUT_1[5483] = 32'b11111111111111111011000110101011;
assign LUT_1[5484] = 32'b00000000000000001101111111110101;
assign LUT_1[5485] = 32'b00000000000000000111010001110001;
assign LUT_1[5486] = 32'b00000000000000001001101110000110;
assign LUT_1[5487] = 32'b00000000000000000011000000000010;
assign LUT_1[5488] = 32'b00000000000000001000110100001011;
assign LUT_1[5489] = 32'b00000000000000000010000110000111;
assign LUT_1[5490] = 32'b00000000000000000100100010011100;
assign LUT_1[5491] = 32'b11111111111111111101110100011000;
assign LUT_1[5492] = 32'b00000000000000010000101101100010;
assign LUT_1[5493] = 32'b00000000000000001001111111011110;
assign LUT_1[5494] = 32'b00000000000000001100011011110011;
assign LUT_1[5495] = 32'b00000000000000000101101101101111;
assign LUT_1[5496] = 32'b00000000000000001000000010000000;
assign LUT_1[5497] = 32'b00000000000000000001010011111100;
assign LUT_1[5498] = 32'b00000000000000000011110000010001;
assign LUT_1[5499] = 32'b11111111111111111101000010001101;
assign LUT_1[5500] = 32'b00000000000000001111111011010111;
assign LUT_1[5501] = 32'b00000000000000001001001101010011;
assign LUT_1[5502] = 32'b00000000000000001011101001101000;
assign LUT_1[5503] = 32'b00000000000000000100111011100100;
assign LUT_1[5504] = 32'b00000000000000000111000000000101;
assign LUT_1[5505] = 32'b00000000000000000000010010000001;
assign LUT_1[5506] = 32'b00000000000000000010101110010110;
assign LUT_1[5507] = 32'b11111111111111111100000000010010;
assign LUT_1[5508] = 32'b00000000000000001110111001011100;
assign LUT_1[5509] = 32'b00000000000000001000001011011000;
assign LUT_1[5510] = 32'b00000000000000001010100111101101;
assign LUT_1[5511] = 32'b00000000000000000011111001101001;
assign LUT_1[5512] = 32'b00000000000000000110001101111010;
assign LUT_1[5513] = 32'b11111111111111111111011111110110;
assign LUT_1[5514] = 32'b00000000000000000001111100001011;
assign LUT_1[5515] = 32'b11111111111111111011001110000111;
assign LUT_1[5516] = 32'b00000000000000001110000111010001;
assign LUT_1[5517] = 32'b00000000000000000111011001001101;
assign LUT_1[5518] = 32'b00000000000000001001110101100010;
assign LUT_1[5519] = 32'b00000000000000000011000111011110;
assign LUT_1[5520] = 32'b00000000000000001000111011100111;
assign LUT_1[5521] = 32'b00000000000000000010001101100011;
assign LUT_1[5522] = 32'b00000000000000000100101001111000;
assign LUT_1[5523] = 32'b11111111111111111101111011110100;
assign LUT_1[5524] = 32'b00000000000000010000110100111110;
assign LUT_1[5525] = 32'b00000000000000001010000110111010;
assign LUT_1[5526] = 32'b00000000000000001100100011001111;
assign LUT_1[5527] = 32'b00000000000000000101110101001011;
assign LUT_1[5528] = 32'b00000000000000001000001001011100;
assign LUT_1[5529] = 32'b00000000000000000001011011011000;
assign LUT_1[5530] = 32'b00000000000000000011110111101101;
assign LUT_1[5531] = 32'b11111111111111111101001001101001;
assign LUT_1[5532] = 32'b00000000000000010000000010110011;
assign LUT_1[5533] = 32'b00000000000000001001010100101111;
assign LUT_1[5534] = 32'b00000000000000001011110001000100;
assign LUT_1[5535] = 32'b00000000000000000101000011000000;
assign LUT_1[5536] = 32'b00000000000000000111111011000100;
assign LUT_1[5537] = 32'b00000000000000000001001101000000;
assign LUT_1[5538] = 32'b00000000000000000011101001010101;
assign LUT_1[5539] = 32'b11111111111111111100111011010001;
assign LUT_1[5540] = 32'b00000000000000001111110100011011;
assign LUT_1[5541] = 32'b00000000000000001001000110010111;
assign LUT_1[5542] = 32'b00000000000000001011100010101100;
assign LUT_1[5543] = 32'b00000000000000000100110100101000;
assign LUT_1[5544] = 32'b00000000000000000111001000111001;
assign LUT_1[5545] = 32'b00000000000000000000011010110101;
assign LUT_1[5546] = 32'b00000000000000000010110111001010;
assign LUT_1[5547] = 32'b11111111111111111100001001000110;
assign LUT_1[5548] = 32'b00000000000000001111000010010000;
assign LUT_1[5549] = 32'b00000000000000001000010100001100;
assign LUT_1[5550] = 32'b00000000000000001010110000100001;
assign LUT_1[5551] = 32'b00000000000000000100000010011101;
assign LUT_1[5552] = 32'b00000000000000001001110110100110;
assign LUT_1[5553] = 32'b00000000000000000011001000100010;
assign LUT_1[5554] = 32'b00000000000000000101100100110111;
assign LUT_1[5555] = 32'b11111111111111111110110110110011;
assign LUT_1[5556] = 32'b00000000000000010001101111111101;
assign LUT_1[5557] = 32'b00000000000000001011000001111001;
assign LUT_1[5558] = 32'b00000000000000001101011110001110;
assign LUT_1[5559] = 32'b00000000000000000110110000001010;
assign LUT_1[5560] = 32'b00000000000000001001000100011011;
assign LUT_1[5561] = 32'b00000000000000000010010110010111;
assign LUT_1[5562] = 32'b00000000000000000100110010101100;
assign LUT_1[5563] = 32'b11111111111111111110000100101000;
assign LUT_1[5564] = 32'b00000000000000010000111101110010;
assign LUT_1[5565] = 32'b00000000000000001010001111101110;
assign LUT_1[5566] = 32'b00000000000000001100101100000011;
assign LUT_1[5567] = 32'b00000000000000000101111101111111;
assign LUT_1[5568] = 32'b00000000000000001000111101101101;
assign LUT_1[5569] = 32'b00000000000000000010001111101001;
assign LUT_1[5570] = 32'b00000000000000000100101011111110;
assign LUT_1[5571] = 32'b11111111111111111101111101111010;
assign LUT_1[5572] = 32'b00000000000000010000110111000100;
assign LUT_1[5573] = 32'b00000000000000001010001001000000;
assign LUT_1[5574] = 32'b00000000000000001100100101010101;
assign LUT_1[5575] = 32'b00000000000000000101110111010001;
assign LUT_1[5576] = 32'b00000000000000001000001011100010;
assign LUT_1[5577] = 32'b00000000000000000001011101011110;
assign LUT_1[5578] = 32'b00000000000000000011111001110011;
assign LUT_1[5579] = 32'b11111111111111111101001011101111;
assign LUT_1[5580] = 32'b00000000000000010000000100111001;
assign LUT_1[5581] = 32'b00000000000000001001010110110101;
assign LUT_1[5582] = 32'b00000000000000001011110011001010;
assign LUT_1[5583] = 32'b00000000000000000101000101000110;
assign LUT_1[5584] = 32'b00000000000000001010111001001111;
assign LUT_1[5585] = 32'b00000000000000000100001011001011;
assign LUT_1[5586] = 32'b00000000000000000110100111100000;
assign LUT_1[5587] = 32'b11111111111111111111111001011100;
assign LUT_1[5588] = 32'b00000000000000010010110010100110;
assign LUT_1[5589] = 32'b00000000000000001100000100100010;
assign LUT_1[5590] = 32'b00000000000000001110100000110111;
assign LUT_1[5591] = 32'b00000000000000000111110010110011;
assign LUT_1[5592] = 32'b00000000000000001010000111000100;
assign LUT_1[5593] = 32'b00000000000000000011011001000000;
assign LUT_1[5594] = 32'b00000000000000000101110101010101;
assign LUT_1[5595] = 32'b11111111111111111111000111010001;
assign LUT_1[5596] = 32'b00000000000000010010000000011011;
assign LUT_1[5597] = 32'b00000000000000001011010010010111;
assign LUT_1[5598] = 32'b00000000000000001101101110101100;
assign LUT_1[5599] = 32'b00000000000000000111000000101000;
assign LUT_1[5600] = 32'b00000000000000001001111000101100;
assign LUT_1[5601] = 32'b00000000000000000011001010101000;
assign LUT_1[5602] = 32'b00000000000000000101100110111101;
assign LUT_1[5603] = 32'b11111111111111111110111000111001;
assign LUT_1[5604] = 32'b00000000000000010001110010000011;
assign LUT_1[5605] = 32'b00000000000000001011000011111111;
assign LUT_1[5606] = 32'b00000000000000001101100000010100;
assign LUT_1[5607] = 32'b00000000000000000110110010010000;
assign LUT_1[5608] = 32'b00000000000000001001000110100001;
assign LUT_1[5609] = 32'b00000000000000000010011000011101;
assign LUT_1[5610] = 32'b00000000000000000100110100110010;
assign LUT_1[5611] = 32'b11111111111111111110000110101110;
assign LUT_1[5612] = 32'b00000000000000010000111111111000;
assign LUT_1[5613] = 32'b00000000000000001010010001110100;
assign LUT_1[5614] = 32'b00000000000000001100101110001001;
assign LUT_1[5615] = 32'b00000000000000000110000000000101;
assign LUT_1[5616] = 32'b00000000000000001011110100001110;
assign LUT_1[5617] = 32'b00000000000000000101000110001010;
assign LUT_1[5618] = 32'b00000000000000000111100010011111;
assign LUT_1[5619] = 32'b00000000000000000000110100011011;
assign LUT_1[5620] = 32'b00000000000000010011101101100101;
assign LUT_1[5621] = 32'b00000000000000001100111111100001;
assign LUT_1[5622] = 32'b00000000000000001111011011110110;
assign LUT_1[5623] = 32'b00000000000000001000101101110010;
assign LUT_1[5624] = 32'b00000000000000001011000010000011;
assign LUT_1[5625] = 32'b00000000000000000100010011111111;
assign LUT_1[5626] = 32'b00000000000000000110110000010100;
assign LUT_1[5627] = 32'b00000000000000000000000010010000;
assign LUT_1[5628] = 32'b00000000000000010010111011011010;
assign LUT_1[5629] = 32'b00000000000000001100001101010110;
assign LUT_1[5630] = 32'b00000000000000001110101001101011;
assign LUT_1[5631] = 32'b00000000000000000111111011100111;
assign LUT_1[5632] = 32'b11111111111111111111111010010011;
assign LUT_1[5633] = 32'b11111111111111111001001100001111;
assign LUT_1[5634] = 32'b11111111111111111011101000100100;
assign LUT_1[5635] = 32'b11111111111111110100111010100000;
assign LUT_1[5636] = 32'b00000000000000000111110011101010;
assign LUT_1[5637] = 32'b00000000000000000001000101100110;
assign LUT_1[5638] = 32'b00000000000000000011100001111011;
assign LUT_1[5639] = 32'b11111111111111111100110011110111;
assign LUT_1[5640] = 32'b11111111111111111111001000001000;
assign LUT_1[5641] = 32'b11111111111111111000011010000100;
assign LUT_1[5642] = 32'b11111111111111111010110110011001;
assign LUT_1[5643] = 32'b11111111111111110100001000010101;
assign LUT_1[5644] = 32'b00000000000000000111000001011111;
assign LUT_1[5645] = 32'b00000000000000000000010011011011;
assign LUT_1[5646] = 32'b00000000000000000010101111110000;
assign LUT_1[5647] = 32'b11111111111111111100000001101100;
assign LUT_1[5648] = 32'b00000000000000000001110101110101;
assign LUT_1[5649] = 32'b11111111111111111011000111110001;
assign LUT_1[5650] = 32'b11111111111111111101100100000110;
assign LUT_1[5651] = 32'b11111111111111110110110110000010;
assign LUT_1[5652] = 32'b00000000000000001001101111001100;
assign LUT_1[5653] = 32'b00000000000000000011000001001000;
assign LUT_1[5654] = 32'b00000000000000000101011101011101;
assign LUT_1[5655] = 32'b11111111111111111110101111011001;
assign LUT_1[5656] = 32'b00000000000000000001000011101010;
assign LUT_1[5657] = 32'b11111111111111111010010101100110;
assign LUT_1[5658] = 32'b11111111111111111100110001111011;
assign LUT_1[5659] = 32'b11111111111111110110000011110111;
assign LUT_1[5660] = 32'b00000000000000001000111101000001;
assign LUT_1[5661] = 32'b00000000000000000010001110111101;
assign LUT_1[5662] = 32'b00000000000000000100101011010010;
assign LUT_1[5663] = 32'b11111111111111111101111101001110;
assign LUT_1[5664] = 32'b00000000000000000000110101010010;
assign LUT_1[5665] = 32'b11111111111111111010000111001110;
assign LUT_1[5666] = 32'b11111111111111111100100011100011;
assign LUT_1[5667] = 32'b11111111111111110101110101011111;
assign LUT_1[5668] = 32'b00000000000000001000101110101001;
assign LUT_1[5669] = 32'b00000000000000000010000000100101;
assign LUT_1[5670] = 32'b00000000000000000100011100111010;
assign LUT_1[5671] = 32'b11111111111111111101101110110110;
assign LUT_1[5672] = 32'b00000000000000000000000011000111;
assign LUT_1[5673] = 32'b11111111111111111001010101000011;
assign LUT_1[5674] = 32'b11111111111111111011110001011000;
assign LUT_1[5675] = 32'b11111111111111110101000011010100;
assign LUT_1[5676] = 32'b00000000000000000111111100011110;
assign LUT_1[5677] = 32'b00000000000000000001001110011010;
assign LUT_1[5678] = 32'b00000000000000000011101010101111;
assign LUT_1[5679] = 32'b11111111111111111100111100101011;
assign LUT_1[5680] = 32'b00000000000000000010110000110100;
assign LUT_1[5681] = 32'b11111111111111111100000010110000;
assign LUT_1[5682] = 32'b11111111111111111110011111000101;
assign LUT_1[5683] = 32'b11111111111111110111110001000001;
assign LUT_1[5684] = 32'b00000000000000001010101010001011;
assign LUT_1[5685] = 32'b00000000000000000011111100000111;
assign LUT_1[5686] = 32'b00000000000000000110011000011100;
assign LUT_1[5687] = 32'b11111111111111111111101010011000;
assign LUT_1[5688] = 32'b00000000000000000001111110101001;
assign LUT_1[5689] = 32'b11111111111111111011010000100101;
assign LUT_1[5690] = 32'b11111111111111111101101100111010;
assign LUT_1[5691] = 32'b11111111111111110110111110110110;
assign LUT_1[5692] = 32'b00000000000000001001111000000000;
assign LUT_1[5693] = 32'b00000000000000000011001001111100;
assign LUT_1[5694] = 32'b00000000000000000101100110010001;
assign LUT_1[5695] = 32'b11111111111111111110111000001101;
assign LUT_1[5696] = 32'b00000000000000000001110111111011;
assign LUT_1[5697] = 32'b11111111111111111011001001110111;
assign LUT_1[5698] = 32'b11111111111111111101100110001100;
assign LUT_1[5699] = 32'b11111111111111110110111000001000;
assign LUT_1[5700] = 32'b00000000000000001001110001010010;
assign LUT_1[5701] = 32'b00000000000000000011000011001110;
assign LUT_1[5702] = 32'b00000000000000000101011111100011;
assign LUT_1[5703] = 32'b11111111111111111110110001011111;
assign LUT_1[5704] = 32'b00000000000000000001000101110000;
assign LUT_1[5705] = 32'b11111111111111111010010111101100;
assign LUT_1[5706] = 32'b11111111111111111100110100000001;
assign LUT_1[5707] = 32'b11111111111111110110000101111101;
assign LUT_1[5708] = 32'b00000000000000001000111111000111;
assign LUT_1[5709] = 32'b00000000000000000010010001000011;
assign LUT_1[5710] = 32'b00000000000000000100101101011000;
assign LUT_1[5711] = 32'b11111111111111111101111111010100;
assign LUT_1[5712] = 32'b00000000000000000011110011011101;
assign LUT_1[5713] = 32'b11111111111111111101000101011001;
assign LUT_1[5714] = 32'b11111111111111111111100001101110;
assign LUT_1[5715] = 32'b11111111111111111000110011101010;
assign LUT_1[5716] = 32'b00000000000000001011101100110100;
assign LUT_1[5717] = 32'b00000000000000000100111110110000;
assign LUT_1[5718] = 32'b00000000000000000111011011000101;
assign LUT_1[5719] = 32'b00000000000000000000101101000001;
assign LUT_1[5720] = 32'b00000000000000000011000001010010;
assign LUT_1[5721] = 32'b11111111111111111100010011001110;
assign LUT_1[5722] = 32'b11111111111111111110101111100011;
assign LUT_1[5723] = 32'b11111111111111111000000001011111;
assign LUT_1[5724] = 32'b00000000000000001010111010101001;
assign LUT_1[5725] = 32'b00000000000000000100001100100101;
assign LUT_1[5726] = 32'b00000000000000000110101000111010;
assign LUT_1[5727] = 32'b11111111111111111111111010110110;
assign LUT_1[5728] = 32'b00000000000000000010110010111010;
assign LUT_1[5729] = 32'b11111111111111111100000100110110;
assign LUT_1[5730] = 32'b11111111111111111110100001001011;
assign LUT_1[5731] = 32'b11111111111111110111110011000111;
assign LUT_1[5732] = 32'b00000000000000001010101100010001;
assign LUT_1[5733] = 32'b00000000000000000011111110001101;
assign LUT_1[5734] = 32'b00000000000000000110011010100010;
assign LUT_1[5735] = 32'b11111111111111111111101100011110;
assign LUT_1[5736] = 32'b00000000000000000010000000101111;
assign LUT_1[5737] = 32'b11111111111111111011010010101011;
assign LUT_1[5738] = 32'b11111111111111111101101111000000;
assign LUT_1[5739] = 32'b11111111111111110111000000111100;
assign LUT_1[5740] = 32'b00000000000000001001111010000110;
assign LUT_1[5741] = 32'b00000000000000000011001100000010;
assign LUT_1[5742] = 32'b00000000000000000101101000010111;
assign LUT_1[5743] = 32'b11111111111111111110111010010011;
assign LUT_1[5744] = 32'b00000000000000000100101110011100;
assign LUT_1[5745] = 32'b11111111111111111110000000011000;
assign LUT_1[5746] = 32'b00000000000000000000011100101101;
assign LUT_1[5747] = 32'b11111111111111111001101110101001;
assign LUT_1[5748] = 32'b00000000000000001100100111110011;
assign LUT_1[5749] = 32'b00000000000000000101111001101111;
assign LUT_1[5750] = 32'b00000000000000001000010110000100;
assign LUT_1[5751] = 32'b00000000000000000001101000000000;
assign LUT_1[5752] = 32'b00000000000000000011111100010001;
assign LUT_1[5753] = 32'b11111111111111111101001110001101;
assign LUT_1[5754] = 32'b11111111111111111111101010100010;
assign LUT_1[5755] = 32'b11111111111111111000111100011110;
assign LUT_1[5756] = 32'b00000000000000001011110101101000;
assign LUT_1[5757] = 32'b00000000000000000101000111100100;
assign LUT_1[5758] = 32'b00000000000000000111100011111001;
assign LUT_1[5759] = 32'b00000000000000000000110101110101;
assign LUT_1[5760] = 32'b00000000000000000010111010010110;
assign LUT_1[5761] = 32'b11111111111111111100001100010010;
assign LUT_1[5762] = 32'b11111111111111111110101000100111;
assign LUT_1[5763] = 32'b11111111111111110111111010100011;
assign LUT_1[5764] = 32'b00000000000000001010110011101101;
assign LUT_1[5765] = 32'b00000000000000000100000101101001;
assign LUT_1[5766] = 32'b00000000000000000110100001111110;
assign LUT_1[5767] = 32'b11111111111111111111110011111010;
assign LUT_1[5768] = 32'b00000000000000000010001000001011;
assign LUT_1[5769] = 32'b11111111111111111011011010000111;
assign LUT_1[5770] = 32'b11111111111111111101110110011100;
assign LUT_1[5771] = 32'b11111111111111110111001000011000;
assign LUT_1[5772] = 32'b00000000000000001010000001100010;
assign LUT_1[5773] = 32'b00000000000000000011010011011110;
assign LUT_1[5774] = 32'b00000000000000000101101111110011;
assign LUT_1[5775] = 32'b11111111111111111111000001101111;
assign LUT_1[5776] = 32'b00000000000000000100110101111000;
assign LUT_1[5777] = 32'b11111111111111111110000111110100;
assign LUT_1[5778] = 32'b00000000000000000000100100001001;
assign LUT_1[5779] = 32'b11111111111111111001110110000101;
assign LUT_1[5780] = 32'b00000000000000001100101111001111;
assign LUT_1[5781] = 32'b00000000000000000110000001001011;
assign LUT_1[5782] = 32'b00000000000000001000011101100000;
assign LUT_1[5783] = 32'b00000000000000000001101111011100;
assign LUT_1[5784] = 32'b00000000000000000100000011101101;
assign LUT_1[5785] = 32'b11111111111111111101010101101001;
assign LUT_1[5786] = 32'b11111111111111111111110001111110;
assign LUT_1[5787] = 32'b11111111111111111001000011111010;
assign LUT_1[5788] = 32'b00000000000000001011111101000100;
assign LUT_1[5789] = 32'b00000000000000000101001111000000;
assign LUT_1[5790] = 32'b00000000000000000111101011010101;
assign LUT_1[5791] = 32'b00000000000000000000111101010001;
assign LUT_1[5792] = 32'b00000000000000000011110101010101;
assign LUT_1[5793] = 32'b11111111111111111101000111010001;
assign LUT_1[5794] = 32'b11111111111111111111100011100110;
assign LUT_1[5795] = 32'b11111111111111111000110101100010;
assign LUT_1[5796] = 32'b00000000000000001011101110101100;
assign LUT_1[5797] = 32'b00000000000000000101000000101000;
assign LUT_1[5798] = 32'b00000000000000000111011100111101;
assign LUT_1[5799] = 32'b00000000000000000000101110111001;
assign LUT_1[5800] = 32'b00000000000000000011000011001010;
assign LUT_1[5801] = 32'b11111111111111111100010101000110;
assign LUT_1[5802] = 32'b11111111111111111110110001011011;
assign LUT_1[5803] = 32'b11111111111111111000000011010111;
assign LUT_1[5804] = 32'b00000000000000001010111100100001;
assign LUT_1[5805] = 32'b00000000000000000100001110011101;
assign LUT_1[5806] = 32'b00000000000000000110101010110010;
assign LUT_1[5807] = 32'b11111111111111111111111100101110;
assign LUT_1[5808] = 32'b00000000000000000101110000110111;
assign LUT_1[5809] = 32'b11111111111111111111000010110011;
assign LUT_1[5810] = 32'b00000000000000000001011111001000;
assign LUT_1[5811] = 32'b11111111111111111010110001000100;
assign LUT_1[5812] = 32'b00000000000000001101101010001110;
assign LUT_1[5813] = 32'b00000000000000000110111100001010;
assign LUT_1[5814] = 32'b00000000000000001001011000011111;
assign LUT_1[5815] = 32'b00000000000000000010101010011011;
assign LUT_1[5816] = 32'b00000000000000000100111110101100;
assign LUT_1[5817] = 32'b11111111111111111110010000101000;
assign LUT_1[5818] = 32'b00000000000000000000101100111101;
assign LUT_1[5819] = 32'b11111111111111111001111110111001;
assign LUT_1[5820] = 32'b00000000000000001100111000000011;
assign LUT_1[5821] = 32'b00000000000000000110001001111111;
assign LUT_1[5822] = 32'b00000000000000001000100110010100;
assign LUT_1[5823] = 32'b00000000000000000001111000010000;
assign LUT_1[5824] = 32'b00000000000000000100110111111110;
assign LUT_1[5825] = 32'b11111111111111111110001001111010;
assign LUT_1[5826] = 32'b00000000000000000000100110001111;
assign LUT_1[5827] = 32'b11111111111111111001111000001011;
assign LUT_1[5828] = 32'b00000000000000001100110001010101;
assign LUT_1[5829] = 32'b00000000000000000110000011010001;
assign LUT_1[5830] = 32'b00000000000000001000011111100110;
assign LUT_1[5831] = 32'b00000000000000000001110001100010;
assign LUT_1[5832] = 32'b00000000000000000100000101110011;
assign LUT_1[5833] = 32'b11111111111111111101010111101111;
assign LUT_1[5834] = 32'b11111111111111111111110100000100;
assign LUT_1[5835] = 32'b11111111111111111001000110000000;
assign LUT_1[5836] = 32'b00000000000000001011111111001010;
assign LUT_1[5837] = 32'b00000000000000000101010001000110;
assign LUT_1[5838] = 32'b00000000000000000111101101011011;
assign LUT_1[5839] = 32'b00000000000000000000111111010111;
assign LUT_1[5840] = 32'b00000000000000000110110011100000;
assign LUT_1[5841] = 32'b00000000000000000000000101011100;
assign LUT_1[5842] = 32'b00000000000000000010100001110001;
assign LUT_1[5843] = 32'b11111111111111111011110011101101;
assign LUT_1[5844] = 32'b00000000000000001110101100110111;
assign LUT_1[5845] = 32'b00000000000000000111111110110011;
assign LUT_1[5846] = 32'b00000000000000001010011011001000;
assign LUT_1[5847] = 32'b00000000000000000011101101000100;
assign LUT_1[5848] = 32'b00000000000000000110000001010101;
assign LUT_1[5849] = 32'b11111111111111111111010011010001;
assign LUT_1[5850] = 32'b00000000000000000001101111100110;
assign LUT_1[5851] = 32'b11111111111111111011000001100010;
assign LUT_1[5852] = 32'b00000000000000001101111010101100;
assign LUT_1[5853] = 32'b00000000000000000111001100101000;
assign LUT_1[5854] = 32'b00000000000000001001101000111101;
assign LUT_1[5855] = 32'b00000000000000000010111010111001;
assign LUT_1[5856] = 32'b00000000000000000101110010111101;
assign LUT_1[5857] = 32'b11111111111111111111000100111001;
assign LUT_1[5858] = 32'b00000000000000000001100001001110;
assign LUT_1[5859] = 32'b11111111111111111010110011001010;
assign LUT_1[5860] = 32'b00000000000000001101101100010100;
assign LUT_1[5861] = 32'b00000000000000000110111110010000;
assign LUT_1[5862] = 32'b00000000000000001001011010100101;
assign LUT_1[5863] = 32'b00000000000000000010101100100001;
assign LUT_1[5864] = 32'b00000000000000000101000000110010;
assign LUT_1[5865] = 32'b11111111111111111110010010101110;
assign LUT_1[5866] = 32'b00000000000000000000101111000011;
assign LUT_1[5867] = 32'b11111111111111111010000000111111;
assign LUT_1[5868] = 32'b00000000000000001100111010001001;
assign LUT_1[5869] = 32'b00000000000000000110001100000101;
assign LUT_1[5870] = 32'b00000000000000001000101000011010;
assign LUT_1[5871] = 32'b00000000000000000001111010010110;
assign LUT_1[5872] = 32'b00000000000000000111101110011111;
assign LUT_1[5873] = 32'b00000000000000000001000000011011;
assign LUT_1[5874] = 32'b00000000000000000011011100110000;
assign LUT_1[5875] = 32'b11111111111111111100101110101100;
assign LUT_1[5876] = 32'b00000000000000001111100111110110;
assign LUT_1[5877] = 32'b00000000000000001000111001110010;
assign LUT_1[5878] = 32'b00000000000000001011010110000111;
assign LUT_1[5879] = 32'b00000000000000000100101000000011;
assign LUT_1[5880] = 32'b00000000000000000110111100010100;
assign LUT_1[5881] = 32'b00000000000000000000001110010000;
assign LUT_1[5882] = 32'b00000000000000000010101010100101;
assign LUT_1[5883] = 32'b11111111111111111011111100100001;
assign LUT_1[5884] = 32'b00000000000000001110110101101011;
assign LUT_1[5885] = 32'b00000000000000001000000111100111;
assign LUT_1[5886] = 32'b00000000000000001010100011111100;
assign LUT_1[5887] = 32'b00000000000000000011110101111000;
assign LUT_1[5888] = 32'b11111111111111111101101110011111;
assign LUT_1[5889] = 32'b11111111111111110111000000011011;
assign LUT_1[5890] = 32'b11111111111111111001011100110000;
assign LUT_1[5891] = 32'b11111111111111110010101110101100;
assign LUT_1[5892] = 32'b00000000000000000101100111110110;
assign LUT_1[5893] = 32'b11111111111111111110111001110010;
assign LUT_1[5894] = 32'b00000000000000000001010110000111;
assign LUT_1[5895] = 32'b11111111111111111010101000000011;
assign LUT_1[5896] = 32'b11111111111111111100111100010100;
assign LUT_1[5897] = 32'b11111111111111110110001110010000;
assign LUT_1[5898] = 32'b11111111111111111000101010100101;
assign LUT_1[5899] = 32'b11111111111111110001111100100001;
assign LUT_1[5900] = 32'b00000000000000000100110101101011;
assign LUT_1[5901] = 32'b11111111111111111110000111100111;
assign LUT_1[5902] = 32'b00000000000000000000100011111100;
assign LUT_1[5903] = 32'b11111111111111111001110101111000;
assign LUT_1[5904] = 32'b11111111111111111111101010000001;
assign LUT_1[5905] = 32'b11111111111111111000111011111101;
assign LUT_1[5906] = 32'b11111111111111111011011000010010;
assign LUT_1[5907] = 32'b11111111111111110100101010001110;
assign LUT_1[5908] = 32'b00000000000000000111100011011000;
assign LUT_1[5909] = 32'b00000000000000000000110101010100;
assign LUT_1[5910] = 32'b00000000000000000011010001101001;
assign LUT_1[5911] = 32'b11111111111111111100100011100101;
assign LUT_1[5912] = 32'b11111111111111111110110111110110;
assign LUT_1[5913] = 32'b11111111111111111000001001110010;
assign LUT_1[5914] = 32'b11111111111111111010100110000111;
assign LUT_1[5915] = 32'b11111111111111110011111000000011;
assign LUT_1[5916] = 32'b00000000000000000110110001001101;
assign LUT_1[5917] = 32'b00000000000000000000000011001001;
assign LUT_1[5918] = 32'b00000000000000000010011111011110;
assign LUT_1[5919] = 32'b11111111111111111011110001011010;
assign LUT_1[5920] = 32'b11111111111111111110101001011110;
assign LUT_1[5921] = 32'b11111111111111110111111011011010;
assign LUT_1[5922] = 32'b11111111111111111010010111101111;
assign LUT_1[5923] = 32'b11111111111111110011101001101011;
assign LUT_1[5924] = 32'b00000000000000000110100010110101;
assign LUT_1[5925] = 32'b11111111111111111111110100110001;
assign LUT_1[5926] = 32'b00000000000000000010010001000110;
assign LUT_1[5927] = 32'b11111111111111111011100011000010;
assign LUT_1[5928] = 32'b11111111111111111101110111010011;
assign LUT_1[5929] = 32'b11111111111111110111001001001111;
assign LUT_1[5930] = 32'b11111111111111111001100101100100;
assign LUT_1[5931] = 32'b11111111111111110010110111100000;
assign LUT_1[5932] = 32'b00000000000000000101110000101010;
assign LUT_1[5933] = 32'b11111111111111111111000010100110;
assign LUT_1[5934] = 32'b00000000000000000001011110111011;
assign LUT_1[5935] = 32'b11111111111111111010110000110111;
assign LUT_1[5936] = 32'b00000000000000000000100101000000;
assign LUT_1[5937] = 32'b11111111111111111001110110111100;
assign LUT_1[5938] = 32'b11111111111111111100010011010001;
assign LUT_1[5939] = 32'b11111111111111110101100101001101;
assign LUT_1[5940] = 32'b00000000000000001000011110010111;
assign LUT_1[5941] = 32'b00000000000000000001110000010011;
assign LUT_1[5942] = 32'b00000000000000000100001100101000;
assign LUT_1[5943] = 32'b11111111111111111101011110100100;
assign LUT_1[5944] = 32'b11111111111111111111110010110101;
assign LUT_1[5945] = 32'b11111111111111111001000100110001;
assign LUT_1[5946] = 32'b11111111111111111011100001000110;
assign LUT_1[5947] = 32'b11111111111111110100110011000010;
assign LUT_1[5948] = 32'b00000000000000000111101100001100;
assign LUT_1[5949] = 32'b00000000000000000000111110001000;
assign LUT_1[5950] = 32'b00000000000000000011011010011101;
assign LUT_1[5951] = 32'b11111111111111111100101100011001;
assign LUT_1[5952] = 32'b11111111111111111111101100000111;
assign LUT_1[5953] = 32'b11111111111111111000111110000011;
assign LUT_1[5954] = 32'b11111111111111111011011010011000;
assign LUT_1[5955] = 32'b11111111111111110100101100010100;
assign LUT_1[5956] = 32'b00000000000000000111100101011110;
assign LUT_1[5957] = 32'b00000000000000000000110111011010;
assign LUT_1[5958] = 32'b00000000000000000011010011101111;
assign LUT_1[5959] = 32'b11111111111111111100100101101011;
assign LUT_1[5960] = 32'b11111111111111111110111001111100;
assign LUT_1[5961] = 32'b11111111111111111000001011111000;
assign LUT_1[5962] = 32'b11111111111111111010101000001101;
assign LUT_1[5963] = 32'b11111111111111110011111010001001;
assign LUT_1[5964] = 32'b00000000000000000110110011010011;
assign LUT_1[5965] = 32'b00000000000000000000000101001111;
assign LUT_1[5966] = 32'b00000000000000000010100001100100;
assign LUT_1[5967] = 32'b11111111111111111011110011100000;
assign LUT_1[5968] = 32'b00000000000000000001100111101001;
assign LUT_1[5969] = 32'b11111111111111111010111001100101;
assign LUT_1[5970] = 32'b11111111111111111101010101111010;
assign LUT_1[5971] = 32'b11111111111111110110100111110110;
assign LUT_1[5972] = 32'b00000000000000001001100001000000;
assign LUT_1[5973] = 32'b00000000000000000010110010111100;
assign LUT_1[5974] = 32'b00000000000000000101001111010001;
assign LUT_1[5975] = 32'b11111111111111111110100001001101;
assign LUT_1[5976] = 32'b00000000000000000000110101011110;
assign LUT_1[5977] = 32'b11111111111111111010000111011010;
assign LUT_1[5978] = 32'b11111111111111111100100011101111;
assign LUT_1[5979] = 32'b11111111111111110101110101101011;
assign LUT_1[5980] = 32'b00000000000000001000101110110101;
assign LUT_1[5981] = 32'b00000000000000000010000000110001;
assign LUT_1[5982] = 32'b00000000000000000100011101000110;
assign LUT_1[5983] = 32'b11111111111111111101101111000010;
assign LUT_1[5984] = 32'b00000000000000000000100111000110;
assign LUT_1[5985] = 32'b11111111111111111001111001000010;
assign LUT_1[5986] = 32'b11111111111111111100010101010111;
assign LUT_1[5987] = 32'b11111111111111110101100111010011;
assign LUT_1[5988] = 32'b00000000000000001000100000011101;
assign LUT_1[5989] = 32'b00000000000000000001110010011001;
assign LUT_1[5990] = 32'b00000000000000000100001110101110;
assign LUT_1[5991] = 32'b11111111111111111101100000101010;
assign LUT_1[5992] = 32'b11111111111111111111110100111011;
assign LUT_1[5993] = 32'b11111111111111111001000110110111;
assign LUT_1[5994] = 32'b11111111111111111011100011001100;
assign LUT_1[5995] = 32'b11111111111111110100110101001000;
assign LUT_1[5996] = 32'b00000000000000000111101110010010;
assign LUT_1[5997] = 32'b00000000000000000001000000001110;
assign LUT_1[5998] = 32'b00000000000000000011011100100011;
assign LUT_1[5999] = 32'b11111111111111111100101110011111;
assign LUT_1[6000] = 32'b00000000000000000010100010101000;
assign LUT_1[6001] = 32'b11111111111111111011110100100100;
assign LUT_1[6002] = 32'b11111111111111111110010000111001;
assign LUT_1[6003] = 32'b11111111111111110111100010110101;
assign LUT_1[6004] = 32'b00000000000000001010011011111111;
assign LUT_1[6005] = 32'b00000000000000000011101101111011;
assign LUT_1[6006] = 32'b00000000000000000110001010010000;
assign LUT_1[6007] = 32'b11111111111111111111011100001100;
assign LUT_1[6008] = 32'b00000000000000000001110000011101;
assign LUT_1[6009] = 32'b11111111111111111011000010011001;
assign LUT_1[6010] = 32'b11111111111111111101011110101110;
assign LUT_1[6011] = 32'b11111111111111110110110000101010;
assign LUT_1[6012] = 32'b00000000000000001001101001110100;
assign LUT_1[6013] = 32'b00000000000000000010111011110000;
assign LUT_1[6014] = 32'b00000000000000000101011000000101;
assign LUT_1[6015] = 32'b11111111111111111110101010000001;
assign LUT_1[6016] = 32'b00000000000000000000101110100010;
assign LUT_1[6017] = 32'b11111111111111111010000000011110;
assign LUT_1[6018] = 32'b11111111111111111100011100110011;
assign LUT_1[6019] = 32'b11111111111111110101101110101111;
assign LUT_1[6020] = 32'b00000000000000001000100111111001;
assign LUT_1[6021] = 32'b00000000000000000001111001110101;
assign LUT_1[6022] = 32'b00000000000000000100010110001010;
assign LUT_1[6023] = 32'b11111111111111111101101000000110;
assign LUT_1[6024] = 32'b11111111111111111111111100010111;
assign LUT_1[6025] = 32'b11111111111111111001001110010011;
assign LUT_1[6026] = 32'b11111111111111111011101010101000;
assign LUT_1[6027] = 32'b11111111111111110100111100100100;
assign LUT_1[6028] = 32'b00000000000000000111110101101110;
assign LUT_1[6029] = 32'b00000000000000000001000111101010;
assign LUT_1[6030] = 32'b00000000000000000011100011111111;
assign LUT_1[6031] = 32'b11111111111111111100110101111011;
assign LUT_1[6032] = 32'b00000000000000000010101010000100;
assign LUT_1[6033] = 32'b11111111111111111011111100000000;
assign LUT_1[6034] = 32'b11111111111111111110011000010101;
assign LUT_1[6035] = 32'b11111111111111110111101010010001;
assign LUT_1[6036] = 32'b00000000000000001010100011011011;
assign LUT_1[6037] = 32'b00000000000000000011110101010111;
assign LUT_1[6038] = 32'b00000000000000000110010001101100;
assign LUT_1[6039] = 32'b11111111111111111111100011101000;
assign LUT_1[6040] = 32'b00000000000000000001110111111001;
assign LUT_1[6041] = 32'b11111111111111111011001001110101;
assign LUT_1[6042] = 32'b11111111111111111101100110001010;
assign LUT_1[6043] = 32'b11111111111111110110111000000110;
assign LUT_1[6044] = 32'b00000000000000001001110001010000;
assign LUT_1[6045] = 32'b00000000000000000011000011001100;
assign LUT_1[6046] = 32'b00000000000000000101011111100001;
assign LUT_1[6047] = 32'b11111111111111111110110001011101;
assign LUT_1[6048] = 32'b00000000000000000001101001100001;
assign LUT_1[6049] = 32'b11111111111111111010111011011101;
assign LUT_1[6050] = 32'b11111111111111111101010111110010;
assign LUT_1[6051] = 32'b11111111111111110110101001101110;
assign LUT_1[6052] = 32'b00000000000000001001100010111000;
assign LUT_1[6053] = 32'b00000000000000000010110100110100;
assign LUT_1[6054] = 32'b00000000000000000101010001001001;
assign LUT_1[6055] = 32'b11111111111111111110100011000101;
assign LUT_1[6056] = 32'b00000000000000000000110111010110;
assign LUT_1[6057] = 32'b11111111111111111010001001010010;
assign LUT_1[6058] = 32'b11111111111111111100100101100111;
assign LUT_1[6059] = 32'b11111111111111110101110111100011;
assign LUT_1[6060] = 32'b00000000000000001000110000101101;
assign LUT_1[6061] = 32'b00000000000000000010000010101001;
assign LUT_1[6062] = 32'b00000000000000000100011110111110;
assign LUT_1[6063] = 32'b11111111111111111101110000111010;
assign LUT_1[6064] = 32'b00000000000000000011100101000011;
assign LUT_1[6065] = 32'b11111111111111111100110110111111;
assign LUT_1[6066] = 32'b11111111111111111111010011010100;
assign LUT_1[6067] = 32'b11111111111111111000100101010000;
assign LUT_1[6068] = 32'b00000000000000001011011110011010;
assign LUT_1[6069] = 32'b00000000000000000100110000010110;
assign LUT_1[6070] = 32'b00000000000000000111001100101011;
assign LUT_1[6071] = 32'b00000000000000000000011110100111;
assign LUT_1[6072] = 32'b00000000000000000010110010111000;
assign LUT_1[6073] = 32'b11111111111111111100000100110100;
assign LUT_1[6074] = 32'b11111111111111111110100001001001;
assign LUT_1[6075] = 32'b11111111111111110111110011000101;
assign LUT_1[6076] = 32'b00000000000000001010101100001111;
assign LUT_1[6077] = 32'b00000000000000000011111110001011;
assign LUT_1[6078] = 32'b00000000000000000110011010100000;
assign LUT_1[6079] = 32'b11111111111111111111101100011100;
assign LUT_1[6080] = 32'b00000000000000000010101100001010;
assign LUT_1[6081] = 32'b11111111111111111011111110000110;
assign LUT_1[6082] = 32'b11111111111111111110011010011011;
assign LUT_1[6083] = 32'b11111111111111110111101100010111;
assign LUT_1[6084] = 32'b00000000000000001010100101100001;
assign LUT_1[6085] = 32'b00000000000000000011110111011101;
assign LUT_1[6086] = 32'b00000000000000000110010011110010;
assign LUT_1[6087] = 32'b11111111111111111111100101101110;
assign LUT_1[6088] = 32'b00000000000000000001111001111111;
assign LUT_1[6089] = 32'b11111111111111111011001011111011;
assign LUT_1[6090] = 32'b11111111111111111101101000010000;
assign LUT_1[6091] = 32'b11111111111111110110111010001100;
assign LUT_1[6092] = 32'b00000000000000001001110011010110;
assign LUT_1[6093] = 32'b00000000000000000011000101010010;
assign LUT_1[6094] = 32'b00000000000000000101100001100111;
assign LUT_1[6095] = 32'b11111111111111111110110011100011;
assign LUT_1[6096] = 32'b00000000000000000100100111101100;
assign LUT_1[6097] = 32'b11111111111111111101111001101000;
assign LUT_1[6098] = 32'b00000000000000000000010101111101;
assign LUT_1[6099] = 32'b11111111111111111001100111111001;
assign LUT_1[6100] = 32'b00000000000000001100100001000011;
assign LUT_1[6101] = 32'b00000000000000000101110010111111;
assign LUT_1[6102] = 32'b00000000000000001000001111010100;
assign LUT_1[6103] = 32'b00000000000000000001100001010000;
assign LUT_1[6104] = 32'b00000000000000000011110101100001;
assign LUT_1[6105] = 32'b11111111111111111101000111011101;
assign LUT_1[6106] = 32'b11111111111111111111100011110010;
assign LUT_1[6107] = 32'b11111111111111111000110101101110;
assign LUT_1[6108] = 32'b00000000000000001011101110111000;
assign LUT_1[6109] = 32'b00000000000000000101000000110100;
assign LUT_1[6110] = 32'b00000000000000000111011101001001;
assign LUT_1[6111] = 32'b00000000000000000000101111000101;
assign LUT_1[6112] = 32'b00000000000000000011100111001001;
assign LUT_1[6113] = 32'b11111111111111111100111001000101;
assign LUT_1[6114] = 32'b11111111111111111111010101011010;
assign LUT_1[6115] = 32'b11111111111111111000100111010110;
assign LUT_1[6116] = 32'b00000000000000001011100000100000;
assign LUT_1[6117] = 32'b00000000000000000100110010011100;
assign LUT_1[6118] = 32'b00000000000000000111001110110001;
assign LUT_1[6119] = 32'b00000000000000000000100000101101;
assign LUT_1[6120] = 32'b00000000000000000010110100111110;
assign LUT_1[6121] = 32'b11111111111111111100000110111010;
assign LUT_1[6122] = 32'b11111111111111111110100011001111;
assign LUT_1[6123] = 32'b11111111111111110111110101001011;
assign LUT_1[6124] = 32'b00000000000000001010101110010101;
assign LUT_1[6125] = 32'b00000000000000000100000000010001;
assign LUT_1[6126] = 32'b00000000000000000110011100100110;
assign LUT_1[6127] = 32'b11111111111111111111101110100010;
assign LUT_1[6128] = 32'b00000000000000000101100010101011;
assign LUT_1[6129] = 32'b11111111111111111110110100100111;
assign LUT_1[6130] = 32'b00000000000000000001010000111100;
assign LUT_1[6131] = 32'b11111111111111111010100010111000;
assign LUT_1[6132] = 32'b00000000000000001101011100000010;
assign LUT_1[6133] = 32'b00000000000000000110101101111110;
assign LUT_1[6134] = 32'b00000000000000001001001010010011;
assign LUT_1[6135] = 32'b00000000000000000010011100001111;
assign LUT_1[6136] = 32'b00000000000000000100110000100000;
assign LUT_1[6137] = 32'b11111111111111111110000010011100;
assign LUT_1[6138] = 32'b00000000000000000000011110110001;
assign LUT_1[6139] = 32'b11111111111111111001110000101101;
assign LUT_1[6140] = 32'b00000000000000001100101001110111;
assign LUT_1[6141] = 32'b00000000000000000101111011110011;
assign LUT_1[6142] = 32'b00000000000000001000011000001000;
assign LUT_1[6143] = 32'b00000000000000000001101010000100;
assign LUT_1[6144] = 32'b00000000000000000000110111000001;
assign LUT_1[6145] = 32'b11111111111111111010001000111101;
assign LUT_1[6146] = 32'b11111111111111111100100101010010;
assign LUT_1[6147] = 32'b11111111111111110101110111001110;
assign LUT_1[6148] = 32'b00000000000000001000110000011000;
assign LUT_1[6149] = 32'b00000000000000000010000010010100;
assign LUT_1[6150] = 32'b00000000000000000100011110101001;
assign LUT_1[6151] = 32'b11111111111111111101110000100101;
assign LUT_1[6152] = 32'b00000000000000000000000100110110;
assign LUT_1[6153] = 32'b11111111111111111001010110110010;
assign LUT_1[6154] = 32'b11111111111111111011110011000111;
assign LUT_1[6155] = 32'b11111111111111110101000101000011;
assign LUT_1[6156] = 32'b00000000000000000111111110001101;
assign LUT_1[6157] = 32'b00000000000000000001010000001001;
assign LUT_1[6158] = 32'b00000000000000000011101100011110;
assign LUT_1[6159] = 32'b11111111111111111100111110011010;
assign LUT_1[6160] = 32'b00000000000000000010110010100011;
assign LUT_1[6161] = 32'b11111111111111111100000100011111;
assign LUT_1[6162] = 32'b11111111111111111110100000110100;
assign LUT_1[6163] = 32'b11111111111111110111110010110000;
assign LUT_1[6164] = 32'b00000000000000001010101011111010;
assign LUT_1[6165] = 32'b00000000000000000011111101110110;
assign LUT_1[6166] = 32'b00000000000000000110011010001011;
assign LUT_1[6167] = 32'b11111111111111111111101100000111;
assign LUT_1[6168] = 32'b00000000000000000010000000011000;
assign LUT_1[6169] = 32'b11111111111111111011010010010100;
assign LUT_1[6170] = 32'b11111111111111111101101110101001;
assign LUT_1[6171] = 32'b11111111111111110111000000100101;
assign LUT_1[6172] = 32'b00000000000000001001111001101111;
assign LUT_1[6173] = 32'b00000000000000000011001011101011;
assign LUT_1[6174] = 32'b00000000000000000101101000000000;
assign LUT_1[6175] = 32'b11111111111111111110111001111100;
assign LUT_1[6176] = 32'b00000000000000000001110010000000;
assign LUT_1[6177] = 32'b11111111111111111011000011111100;
assign LUT_1[6178] = 32'b11111111111111111101100000010001;
assign LUT_1[6179] = 32'b11111111111111110110110010001101;
assign LUT_1[6180] = 32'b00000000000000001001101011010111;
assign LUT_1[6181] = 32'b00000000000000000010111101010011;
assign LUT_1[6182] = 32'b00000000000000000101011001101000;
assign LUT_1[6183] = 32'b11111111111111111110101011100100;
assign LUT_1[6184] = 32'b00000000000000000000111111110101;
assign LUT_1[6185] = 32'b11111111111111111010010001110001;
assign LUT_1[6186] = 32'b11111111111111111100101110000110;
assign LUT_1[6187] = 32'b11111111111111110110000000000010;
assign LUT_1[6188] = 32'b00000000000000001000111001001100;
assign LUT_1[6189] = 32'b00000000000000000010001011001000;
assign LUT_1[6190] = 32'b00000000000000000100100111011101;
assign LUT_1[6191] = 32'b11111111111111111101111001011001;
assign LUT_1[6192] = 32'b00000000000000000011101101100010;
assign LUT_1[6193] = 32'b11111111111111111100111111011110;
assign LUT_1[6194] = 32'b11111111111111111111011011110011;
assign LUT_1[6195] = 32'b11111111111111111000101101101111;
assign LUT_1[6196] = 32'b00000000000000001011100110111001;
assign LUT_1[6197] = 32'b00000000000000000100111000110101;
assign LUT_1[6198] = 32'b00000000000000000111010101001010;
assign LUT_1[6199] = 32'b00000000000000000000100111000110;
assign LUT_1[6200] = 32'b00000000000000000010111011010111;
assign LUT_1[6201] = 32'b11111111111111111100001101010011;
assign LUT_1[6202] = 32'b11111111111111111110101001101000;
assign LUT_1[6203] = 32'b11111111111111110111111011100100;
assign LUT_1[6204] = 32'b00000000000000001010110100101110;
assign LUT_1[6205] = 32'b00000000000000000100000110101010;
assign LUT_1[6206] = 32'b00000000000000000110100010111111;
assign LUT_1[6207] = 32'b11111111111111111111110100111011;
assign LUT_1[6208] = 32'b00000000000000000010110100101001;
assign LUT_1[6209] = 32'b11111111111111111100000110100101;
assign LUT_1[6210] = 32'b11111111111111111110100010111010;
assign LUT_1[6211] = 32'b11111111111111110111110100110110;
assign LUT_1[6212] = 32'b00000000000000001010101110000000;
assign LUT_1[6213] = 32'b00000000000000000011111111111100;
assign LUT_1[6214] = 32'b00000000000000000110011100010001;
assign LUT_1[6215] = 32'b11111111111111111111101110001101;
assign LUT_1[6216] = 32'b00000000000000000010000010011110;
assign LUT_1[6217] = 32'b11111111111111111011010100011010;
assign LUT_1[6218] = 32'b11111111111111111101110000101111;
assign LUT_1[6219] = 32'b11111111111111110111000010101011;
assign LUT_1[6220] = 32'b00000000000000001001111011110101;
assign LUT_1[6221] = 32'b00000000000000000011001101110001;
assign LUT_1[6222] = 32'b00000000000000000101101010000110;
assign LUT_1[6223] = 32'b11111111111111111110111100000010;
assign LUT_1[6224] = 32'b00000000000000000100110000001011;
assign LUT_1[6225] = 32'b11111111111111111110000010000111;
assign LUT_1[6226] = 32'b00000000000000000000011110011100;
assign LUT_1[6227] = 32'b11111111111111111001110000011000;
assign LUT_1[6228] = 32'b00000000000000001100101001100010;
assign LUT_1[6229] = 32'b00000000000000000101111011011110;
assign LUT_1[6230] = 32'b00000000000000001000010111110011;
assign LUT_1[6231] = 32'b00000000000000000001101001101111;
assign LUT_1[6232] = 32'b00000000000000000011111110000000;
assign LUT_1[6233] = 32'b11111111111111111101001111111100;
assign LUT_1[6234] = 32'b11111111111111111111101100010001;
assign LUT_1[6235] = 32'b11111111111111111000111110001101;
assign LUT_1[6236] = 32'b00000000000000001011110111010111;
assign LUT_1[6237] = 32'b00000000000000000101001001010011;
assign LUT_1[6238] = 32'b00000000000000000111100101101000;
assign LUT_1[6239] = 32'b00000000000000000000110111100100;
assign LUT_1[6240] = 32'b00000000000000000011101111101000;
assign LUT_1[6241] = 32'b11111111111111111101000001100100;
assign LUT_1[6242] = 32'b11111111111111111111011101111001;
assign LUT_1[6243] = 32'b11111111111111111000101111110101;
assign LUT_1[6244] = 32'b00000000000000001011101000111111;
assign LUT_1[6245] = 32'b00000000000000000100111010111011;
assign LUT_1[6246] = 32'b00000000000000000111010111010000;
assign LUT_1[6247] = 32'b00000000000000000000101001001100;
assign LUT_1[6248] = 32'b00000000000000000010111101011101;
assign LUT_1[6249] = 32'b11111111111111111100001111011001;
assign LUT_1[6250] = 32'b11111111111111111110101011101110;
assign LUT_1[6251] = 32'b11111111111111110111111101101010;
assign LUT_1[6252] = 32'b00000000000000001010110110110100;
assign LUT_1[6253] = 32'b00000000000000000100001000110000;
assign LUT_1[6254] = 32'b00000000000000000110100101000101;
assign LUT_1[6255] = 32'b11111111111111111111110111000001;
assign LUT_1[6256] = 32'b00000000000000000101101011001010;
assign LUT_1[6257] = 32'b11111111111111111110111101000110;
assign LUT_1[6258] = 32'b00000000000000000001011001011011;
assign LUT_1[6259] = 32'b11111111111111111010101011010111;
assign LUT_1[6260] = 32'b00000000000000001101100100100001;
assign LUT_1[6261] = 32'b00000000000000000110110110011101;
assign LUT_1[6262] = 32'b00000000000000001001010010110010;
assign LUT_1[6263] = 32'b00000000000000000010100100101110;
assign LUT_1[6264] = 32'b00000000000000000100111000111111;
assign LUT_1[6265] = 32'b11111111111111111110001010111011;
assign LUT_1[6266] = 32'b00000000000000000000100111010000;
assign LUT_1[6267] = 32'b11111111111111111001111001001100;
assign LUT_1[6268] = 32'b00000000000000001100110010010110;
assign LUT_1[6269] = 32'b00000000000000000110000100010010;
assign LUT_1[6270] = 32'b00000000000000001000100000100111;
assign LUT_1[6271] = 32'b00000000000000000001110010100011;
assign LUT_1[6272] = 32'b00000000000000000011110111000100;
assign LUT_1[6273] = 32'b11111111111111111101001001000000;
assign LUT_1[6274] = 32'b11111111111111111111100101010101;
assign LUT_1[6275] = 32'b11111111111111111000110111010001;
assign LUT_1[6276] = 32'b00000000000000001011110000011011;
assign LUT_1[6277] = 32'b00000000000000000101000010010111;
assign LUT_1[6278] = 32'b00000000000000000111011110101100;
assign LUT_1[6279] = 32'b00000000000000000000110000101000;
assign LUT_1[6280] = 32'b00000000000000000011000100111001;
assign LUT_1[6281] = 32'b11111111111111111100010110110101;
assign LUT_1[6282] = 32'b11111111111111111110110011001010;
assign LUT_1[6283] = 32'b11111111111111111000000101000110;
assign LUT_1[6284] = 32'b00000000000000001010111110010000;
assign LUT_1[6285] = 32'b00000000000000000100010000001100;
assign LUT_1[6286] = 32'b00000000000000000110101100100001;
assign LUT_1[6287] = 32'b11111111111111111111111110011101;
assign LUT_1[6288] = 32'b00000000000000000101110010100110;
assign LUT_1[6289] = 32'b11111111111111111111000100100010;
assign LUT_1[6290] = 32'b00000000000000000001100000110111;
assign LUT_1[6291] = 32'b11111111111111111010110010110011;
assign LUT_1[6292] = 32'b00000000000000001101101011111101;
assign LUT_1[6293] = 32'b00000000000000000110111101111001;
assign LUT_1[6294] = 32'b00000000000000001001011010001110;
assign LUT_1[6295] = 32'b00000000000000000010101100001010;
assign LUT_1[6296] = 32'b00000000000000000101000000011011;
assign LUT_1[6297] = 32'b11111111111111111110010010010111;
assign LUT_1[6298] = 32'b00000000000000000000101110101100;
assign LUT_1[6299] = 32'b11111111111111111010000000101000;
assign LUT_1[6300] = 32'b00000000000000001100111001110010;
assign LUT_1[6301] = 32'b00000000000000000110001011101110;
assign LUT_1[6302] = 32'b00000000000000001000101000000011;
assign LUT_1[6303] = 32'b00000000000000000001111001111111;
assign LUT_1[6304] = 32'b00000000000000000100110010000011;
assign LUT_1[6305] = 32'b11111111111111111110000011111111;
assign LUT_1[6306] = 32'b00000000000000000000100000010100;
assign LUT_1[6307] = 32'b11111111111111111001110010010000;
assign LUT_1[6308] = 32'b00000000000000001100101011011010;
assign LUT_1[6309] = 32'b00000000000000000101111101010110;
assign LUT_1[6310] = 32'b00000000000000001000011001101011;
assign LUT_1[6311] = 32'b00000000000000000001101011100111;
assign LUT_1[6312] = 32'b00000000000000000011111111111000;
assign LUT_1[6313] = 32'b11111111111111111101010001110100;
assign LUT_1[6314] = 32'b11111111111111111111101110001001;
assign LUT_1[6315] = 32'b11111111111111111001000000000101;
assign LUT_1[6316] = 32'b00000000000000001011111001001111;
assign LUT_1[6317] = 32'b00000000000000000101001011001011;
assign LUT_1[6318] = 32'b00000000000000000111100111100000;
assign LUT_1[6319] = 32'b00000000000000000000111001011100;
assign LUT_1[6320] = 32'b00000000000000000110101101100101;
assign LUT_1[6321] = 32'b11111111111111111111111111100001;
assign LUT_1[6322] = 32'b00000000000000000010011011110110;
assign LUT_1[6323] = 32'b11111111111111111011101101110010;
assign LUT_1[6324] = 32'b00000000000000001110100110111100;
assign LUT_1[6325] = 32'b00000000000000000111111000111000;
assign LUT_1[6326] = 32'b00000000000000001010010101001101;
assign LUT_1[6327] = 32'b00000000000000000011100111001001;
assign LUT_1[6328] = 32'b00000000000000000101111011011010;
assign LUT_1[6329] = 32'b11111111111111111111001101010110;
assign LUT_1[6330] = 32'b00000000000000000001101001101011;
assign LUT_1[6331] = 32'b11111111111111111010111011100111;
assign LUT_1[6332] = 32'b00000000000000001101110100110001;
assign LUT_1[6333] = 32'b00000000000000000111000110101101;
assign LUT_1[6334] = 32'b00000000000000001001100011000010;
assign LUT_1[6335] = 32'b00000000000000000010110100111110;
assign LUT_1[6336] = 32'b00000000000000000101110100101100;
assign LUT_1[6337] = 32'b11111111111111111111000110101000;
assign LUT_1[6338] = 32'b00000000000000000001100010111101;
assign LUT_1[6339] = 32'b11111111111111111010110100111001;
assign LUT_1[6340] = 32'b00000000000000001101101110000011;
assign LUT_1[6341] = 32'b00000000000000000110111111111111;
assign LUT_1[6342] = 32'b00000000000000001001011100010100;
assign LUT_1[6343] = 32'b00000000000000000010101110010000;
assign LUT_1[6344] = 32'b00000000000000000101000010100001;
assign LUT_1[6345] = 32'b11111111111111111110010100011101;
assign LUT_1[6346] = 32'b00000000000000000000110000110010;
assign LUT_1[6347] = 32'b11111111111111111010000010101110;
assign LUT_1[6348] = 32'b00000000000000001100111011111000;
assign LUT_1[6349] = 32'b00000000000000000110001101110100;
assign LUT_1[6350] = 32'b00000000000000001000101010001001;
assign LUT_1[6351] = 32'b00000000000000000001111100000101;
assign LUT_1[6352] = 32'b00000000000000000111110000001110;
assign LUT_1[6353] = 32'b00000000000000000001000010001010;
assign LUT_1[6354] = 32'b00000000000000000011011110011111;
assign LUT_1[6355] = 32'b11111111111111111100110000011011;
assign LUT_1[6356] = 32'b00000000000000001111101001100101;
assign LUT_1[6357] = 32'b00000000000000001000111011100001;
assign LUT_1[6358] = 32'b00000000000000001011010111110110;
assign LUT_1[6359] = 32'b00000000000000000100101001110010;
assign LUT_1[6360] = 32'b00000000000000000110111110000011;
assign LUT_1[6361] = 32'b00000000000000000000001111111111;
assign LUT_1[6362] = 32'b00000000000000000010101100010100;
assign LUT_1[6363] = 32'b11111111111111111011111110010000;
assign LUT_1[6364] = 32'b00000000000000001110110111011010;
assign LUT_1[6365] = 32'b00000000000000001000001001010110;
assign LUT_1[6366] = 32'b00000000000000001010100101101011;
assign LUT_1[6367] = 32'b00000000000000000011110111100111;
assign LUT_1[6368] = 32'b00000000000000000110101111101011;
assign LUT_1[6369] = 32'b00000000000000000000000001100111;
assign LUT_1[6370] = 32'b00000000000000000010011101111100;
assign LUT_1[6371] = 32'b11111111111111111011101111111000;
assign LUT_1[6372] = 32'b00000000000000001110101001000010;
assign LUT_1[6373] = 32'b00000000000000000111111010111110;
assign LUT_1[6374] = 32'b00000000000000001010010111010011;
assign LUT_1[6375] = 32'b00000000000000000011101001001111;
assign LUT_1[6376] = 32'b00000000000000000101111101100000;
assign LUT_1[6377] = 32'b11111111111111111111001111011100;
assign LUT_1[6378] = 32'b00000000000000000001101011110001;
assign LUT_1[6379] = 32'b11111111111111111010111101101101;
assign LUT_1[6380] = 32'b00000000000000001101110110110111;
assign LUT_1[6381] = 32'b00000000000000000111001000110011;
assign LUT_1[6382] = 32'b00000000000000001001100101001000;
assign LUT_1[6383] = 32'b00000000000000000010110111000100;
assign LUT_1[6384] = 32'b00000000000000001000101011001101;
assign LUT_1[6385] = 32'b00000000000000000001111101001001;
assign LUT_1[6386] = 32'b00000000000000000100011001011110;
assign LUT_1[6387] = 32'b11111111111111111101101011011010;
assign LUT_1[6388] = 32'b00000000000000010000100100100100;
assign LUT_1[6389] = 32'b00000000000000001001110110100000;
assign LUT_1[6390] = 32'b00000000000000001100010010110101;
assign LUT_1[6391] = 32'b00000000000000000101100100110001;
assign LUT_1[6392] = 32'b00000000000000000111111001000010;
assign LUT_1[6393] = 32'b00000000000000000001001010111110;
assign LUT_1[6394] = 32'b00000000000000000011100111010011;
assign LUT_1[6395] = 32'b11111111111111111100111001001111;
assign LUT_1[6396] = 32'b00000000000000001111110010011001;
assign LUT_1[6397] = 32'b00000000000000001001000100010101;
assign LUT_1[6398] = 32'b00000000000000001011100000101010;
assign LUT_1[6399] = 32'b00000000000000000100110010100110;
assign LUT_1[6400] = 32'b11111111111111111110101011001101;
assign LUT_1[6401] = 32'b11111111111111110111111101001001;
assign LUT_1[6402] = 32'b11111111111111111010011001011110;
assign LUT_1[6403] = 32'b11111111111111110011101011011010;
assign LUT_1[6404] = 32'b00000000000000000110100100100100;
assign LUT_1[6405] = 32'b11111111111111111111110110100000;
assign LUT_1[6406] = 32'b00000000000000000010010010110101;
assign LUT_1[6407] = 32'b11111111111111111011100100110001;
assign LUT_1[6408] = 32'b11111111111111111101111001000010;
assign LUT_1[6409] = 32'b11111111111111110111001010111110;
assign LUT_1[6410] = 32'b11111111111111111001100111010011;
assign LUT_1[6411] = 32'b11111111111111110010111001001111;
assign LUT_1[6412] = 32'b00000000000000000101110010011001;
assign LUT_1[6413] = 32'b11111111111111111111000100010101;
assign LUT_1[6414] = 32'b00000000000000000001100000101010;
assign LUT_1[6415] = 32'b11111111111111111010110010100110;
assign LUT_1[6416] = 32'b00000000000000000000100110101111;
assign LUT_1[6417] = 32'b11111111111111111001111000101011;
assign LUT_1[6418] = 32'b11111111111111111100010101000000;
assign LUT_1[6419] = 32'b11111111111111110101100110111100;
assign LUT_1[6420] = 32'b00000000000000001000100000000110;
assign LUT_1[6421] = 32'b00000000000000000001110010000010;
assign LUT_1[6422] = 32'b00000000000000000100001110010111;
assign LUT_1[6423] = 32'b11111111111111111101100000010011;
assign LUT_1[6424] = 32'b11111111111111111111110100100100;
assign LUT_1[6425] = 32'b11111111111111111001000110100000;
assign LUT_1[6426] = 32'b11111111111111111011100010110101;
assign LUT_1[6427] = 32'b11111111111111110100110100110001;
assign LUT_1[6428] = 32'b00000000000000000111101101111011;
assign LUT_1[6429] = 32'b00000000000000000000111111110111;
assign LUT_1[6430] = 32'b00000000000000000011011100001100;
assign LUT_1[6431] = 32'b11111111111111111100101110001000;
assign LUT_1[6432] = 32'b11111111111111111111100110001100;
assign LUT_1[6433] = 32'b11111111111111111000111000001000;
assign LUT_1[6434] = 32'b11111111111111111011010100011101;
assign LUT_1[6435] = 32'b11111111111111110100100110011001;
assign LUT_1[6436] = 32'b00000000000000000111011111100011;
assign LUT_1[6437] = 32'b00000000000000000000110001011111;
assign LUT_1[6438] = 32'b00000000000000000011001101110100;
assign LUT_1[6439] = 32'b11111111111111111100011111110000;
assign LUT_1[6440] = 32'b11111111111111111110110100000001;
assign LUT_1[6441] = 32'b11111111111111111000000101111101;
assign LUT_1[6442] = 32'b11111111111111111010100010010010;
assign LUT_1[6443] = 32'b11111111111111110011110100001110;
assign LUT_1[6444] = 32'b00000000000000000110101101011000;
assign LUT_1[6445] = 32'b11111111111111111111111111010100;
assign LUT_1[6446] = 32'b00000000000000000010011011101001;
assign LUT_1[6447] = 32'b11111111111111111011101101100101;
assign LUT_1[6448] = 32'b00000000000000000001100001101110;
assign LUT_1[6449] = 32'b11111111111111111010110011101010;
assign LUT_1[6450] = 32'b11111111111111111101001111111111;
assign LUT_1[6451] = 32'b11111111111111110110100001111011;
assign LUT_1[6452] = 32'b00000000000000001001011011000101;
assign LUT_1[6453] = 32'b00000000000000000010101101000001;
assign LUT_1[6454] = 32'b00000000000000000101001001010110;
assign LUT_1[6455] = 32'b11111111111111111110011011010010;
assign LUT_1[6456] = 32'b00000000000000000000101111100011;
assign LUT_1[6457] = 32'b11111111111111111010000001011111;
assign LUT_1[6458] = 32'b11111111111111111100011101110100;
assign LUT_1[6459] = 32'b11111111111111110101101111110000;
assign LUT_1[6460] = 32'b00000000000000001000101000111010;
assign LUT_1[6461] = 32'b00000000000000000001111010110110;
assign LUT_1[6462] = 32'b00000000000000000100010111001011;
assign LUT_1[6463] = 32'b11111111111111111101101001000111;
assign LUT_1[6464] = 32'b00000000000000000000101000110101;
assign LUT_1[6465] = 32'b11111111111111111001111010110001;
assign LUT_1[6466] = 32'b11111111111111111100010111000110;
assign LUT_1[6467] = 32'b11111111111111110101101001000010;
assign LUT_1[6468] = 32'b00000000000000001000100010001100;
assign LUT_1[6469] = 32'b00000000000000000001110100001000;
assign LUT_1[6470] = 32'b00000000000000000100010000011101;
assign LUT_1[6471] = 32'b11111111111111111101100010011001;
assign LUT_1[6472] = 32'b11111111111111111111110110101010;
assign LUT_1[6473] = 32'b11111111111111111001001000100110;
assign LUT_1[6474] = 32'b11111111111111111011100100111011;
assign LUT_1[6475] = 32'b11111111111111110100110110110111;
assign LUT_1[6476] = 32'b00000000000000000111110000000001;
assign LUT_1[6477] = 32'b00000000000000000001000001111101;
assign LUT_1[6478] = 32'b00000000000000000011011110010010;
assign LUT_1[6479] = 32'b11111111111111111100110000001110;
assign LUT_1[6480] = 32'b00000000000000000010100100010111;
assign LUT_1[6481] = 32'b11111111111111111011110110010011;
assign LUT_1[6482] = 32'b11111111111111111110010010101000;
assign LUT_1[6483] = 32'b11111111111111110111100100100100;
assign LUT_1[6484] = 32'b00000000000000001010011101101110;
assign LUT_1[6485] = 32'b00000000000000000011101111101010;
assign LUT_1[6486] = 32'b00000000000000000110001011111111;
assign LUT_1[6487] = 32'b11111111111111111111011101111011;
assign LUT_1[6488] = 32'b00000000000000000001110010001100;
assign LUT_1[6489] = 32'b11111111111111111011000100001000;
assign LUT_1[6490] = 32'b11111111111111111101100000011101;
assign LUT_1[6491] = 32'b11111111111111110110110010011001;
assign LUT_1[6492] = 32'b00000000000000001001101011100011;
assign LUT_1[6493] = 32'b00000000000000000010111101011111;
assign LUT_1[6494] = 32'b00000000000000000101011001110100;
assign LUT_1[6495] = 32'b11111111111111111110101011110000;
assign LUT_1[6496] = 32'b00000000000000000001100011110100;
assign LUT_1[6497] = 32'b11111111111111111010110101110000;
assign LUT_1[6498] = 32'b11111111111111111101010010000101;
assign LUT_1[6499] = 32'b11111111111111110110100100000001;
assign LUT_1[6500] = 32'b00000000000000001001011101001011;
assign LUT_1[6501] = 32'b00000000000000000010101111000111;
assign LUT_1[6502] = 32'b00000000000000000101001011011100;
assign LUT_1[6503] = 32'b11111111111111111110011101011000;
assign LUT_1[6504] = 32'b00000000000000000000110001101001;
assign LUT_1[6505] = 32'b11111111111111111010000011100101;
assign LUT_1[6506] = 32'b11111111111111111100011111111010;
assign LUT_1[6507] = 32'b11111111111111110101110001110110;
assign LUT_1[6508] = 32'b00000000000000001000101011000000;
assign LUT_1[6509] = 32'b00000000000000000001111100111100;
assign LUT_1[6510] = 32'b00000000000000000100011001010001;
assign LUT_1[6511] = 32'b11111111111111111101101011001101;
assign LUT_1[6512] = 32'b00000000000000000011011111010110;
assign LUT_1[6513] = 32'b11111111111111111100110001010010;
assign LUT_1[6514] = 32'b11111111111111111111001101100111;
assign LUT_1[6515] = 32'b11111111111111111000011111100011;
assign LUT_1[6516] = 32'b00000000000000001011011000101101;
assign LUT_1[6517] = 32'b00000000000000000100101010101001;
assign LUT_1[6518] = 32'b00000000000000000111000110111110;
assign LUT_1[6519] = 32'b00000000000000000000011000111010;
assign LUT_1[6520] = 32'b00000000000000000010101101001011;
assign LUT_1[6521] = 32'b11111111111111111011111111000111;
assign LUT_1[6522] = 32'b11111111111111111110011011011100;
assign LUT_1[6523] = 32'b11111111111111110111101101011000;
assign LUT_1[6524] = 32'b00000000000000001010100110100010;
assign LUT_1[6525] = 32'b00000000000000000011111000011110;
assign LUT_1[6526] = 32'b00000000000000000110010100110011;
assign LUT_1[6527] = 32'b11111111111111111111100110101111;
assign LUT_1[6528] = 32'b00000000000000000001101011010000;
assign LUT_1[6529] = 32'b11111111111111111010111101001100;
assign LUT_1[6530] = 32'b11111111111111111101011001100001;
assign LUT_1[6531] = 32'b11111111111111110110101011011101;
assign LUT_1[6532] = 32'b00000000000000001001100100100111;
assign LUT_1[6533] = 32'b00000000000000000010110110100011;
assign LUT_1[6534] = 32'b00000000000000000101010010111000;
assign LUT_1[6535] = 32'b11111111111111111110100100110100;
assign LUT_1[6536] = 32'b00000000000000000000111001000101;
assign LUT_1[6537] = 32'b11111111111111111010001011000001;
assign LUT_1[6538] = 32'b11111111111111111100100111010110;
assign LUT_1[6539] = 32'b11111111111111110101111001010010;
assign LUT_1[6540] = 32'b00000000000000001000110010011100;
assign LUT_1[6541] = 32'b00000000000000000010000100011000;
assign LUT_1[6542] = 32'b00000000000000000100100000101101;
assign LUT_1[6543] = 32'b11111111111111111101110010101001;
assign LUT_1[6544] = 32'b00000000000000000011100110110010;
assign LUT_1[6545] = 32'b11111111111111111100111000101110;
assign LUT_1[6546] = 32'b11111111111111111111010101000011;
assign LUT_1[6547] = 32'b11111111111111111000100110111111;
assign LUT_1[6548] = 32'b00000000000000001011100000001001;
assign LUT_1[6549] = 32'b00000000000000000100110010000101;
assign LUT_1[6550] = 32'b00000000000000000111001110011010;
assign LUT_1[6551] = 32'b00000000000000000000100000010110;
assign LUT_1[6552] = 32'b00000000000000000010110100100111;
assign LUT_1[6553] = 32'b11111111111111111100000110100011;
assign LUT_1[6554] = 32'b11111111111111111110100010111000;
assign LUT_1[6555] = 32'b11111111111111110111110100110100;
assign LUT_1[6556] = 32'b00000000000000001010101101111110;
assign LUT_1[6557] = 32'b00000000000000000011111111111010;
assign LUT_1[6558] = 32'b00000000000000000110011100001111;
assign LUT_1[6559] = 32'b11111111111111111111101110001011;
assign LUT_1[6560] = 32'b00000000000000000010100110001111;
assign LUT_1[6561] = 32'b11111111111111111011111000001011;
assign LUT_1[6562] = 32'b11111111111111111110010100100000;
assign LUT_1[6563] = 32'b11111111111111110111100110011100;
assign LUT_1[6564] = 32'b00000000000000001010011111100110;
assign LUT_1[6565] = 32'b00000000000000000011110001100010;
assign LUT_1[6566] = 32'b00000000000000000110001101110111;
assign LUT_1[6567] = 32'b11111111111111111111011111110011;
assign LUT_1[6568] = 32'b00000000000000000001110100000100;
assign LUT_1[6569] = 32'b11111111111111111011000110000000;
assign LUT_1[6570] = 32'b11111111111111111101100010010101;
assign LUT_1[6571] = 32'b11111111111111110110110100010001;
assign LUT_1[6572] = 32'b00000000000000001001101101011011;
assign LUT_1[6573] = 32'b00000000000000000010111111010111;
assign LUT_1[6574] = 32'b00000000000000000101011011101100;
assign LUT_1[6575] = 32'b11111111111111111110101101101000;
assign LUT_1[6576] = 32'b00000000000000000100100001110001;
assign LUT_1[6577] = 32'b11111111111111111101110011101101;
assign LUT_1[6578] = 32'b00000000000000000000010000000010;
assign LUT_1[6579] = 32'b11111111111111111001100001111110;
assign LUT_1[6580] = 32'b00000000000000001100011011001000;
assign LUT_1[6581] = 32'b00000000000000000101101101000100;
assign LUT_1[6582] = 32'b00000000000000001000001001011001;
assign LUT_1[6583] = 32'b00000000000000000001011011010101;
assign LUT_1[6584] = 32'b00000000000000000011101111100110;
assign LUT_1[6585] = 32'b11111111111111111101000001100010;
assign LUT_1[6586] = 32'b11111111111111111111011101110111;
assign LUT_1[6587] = 32'b11111111111111111000101111110011;
assign LUT_1[6588] = 32'b00000000000000001011101000111101;
assign LUT_1[6589] = 32'b00000000000000000100111010111001;
assign LUT_1[6590] = 32'b00000000000000000111010111001110;
assign LUT_1[6591] = 32'b00000000000000000000101001001010;
assign LUT_1[6592] = 32'b00000000000000000011101000111000;
assign LUT_1[6593] = 32'b11111111111111111100111010110100;
assign LUT_1[6594] = 32'b11111111111111111111010111001001;
assign LUT_1[6595] = 32'b11111111111111111000101001000101;
assign LUT_1[6596] = 32'b00000000000000001011100010001111;
assign LUT_1[6597] = 32'b00000000000000000100110100001011;
assign LUT_1[6598] = 32'b00000000000000000111010000100000;
assign LUT_1[6599] = 32'b00000000000000000000100010011100;
assign LUT_1[6600] = 32'b00000000000000000010110110101101;
assign LUT_1[6601] = 32'b11111111111111111100001000101001;
assign LUT_1[6602] = 32'b11111111111111111110100100111110;
assign LUT_1[6603] = 32'b11111111111111110111110110111010;
assign LUT_1[6604] = 32'b00000000000000001010110000000100;
assign LUT_1[6605] = 32'b00000000000000000100000010000000;
assign LUT_1[6606] = 32'b00000000000000000110011110010101;
assign LUT_1[6607] = 32'b11111111111111111111110000010001;
assign LUT_1[6608] = 32'b00000000000000000101100100011010;
assign LUT_1[6609] = 32'b11111111111111111110110110010110;
assign LUT_1[6610] = 32'b00000000000000000001010010101011;
assign LUT_1[6611] = 32'b11111111111111111010100100100111;
assign LUT_1[6612] = 32'b00000000000000001101011101110001;
assign LUT_1[6613] = 32'b00000000000000000110101111101101;
assign LUT_1[6614] = 32'b00000000000000001001001100000010;
assign LUT_1[6615] = 32'b00000000000000000010011101111110;
assign LUT_1[6616] = 32'b00000000000000000100110010001111;
assign LUT_1[6617] = 32'b11111111111111111110000100001011;
assign LUT_1[6618] = 32'b00000000000000000000100000100000;
assign LUT_1[6619] = 32'b11111111111111111001110010011100;
assign LUT_1[6620] = 32'b00000000000000001100101011100110;
assign LUT_1[6621] = 32'b00000000000000000101111101100010;
assign LUT_1[6622] = 32'b00000000000000001000011001110111;
assign LUT_1[6623] = 32'b00000000000000000001101011110011;
assign LUT_1[6624] = 32'b00000000000000000100100011110111;
assign LUT_1[6625] = 32'b11111111111111111101110101110011;
assign LUT_1[6626] = 32'b00000000000000000000010010001000;
assign LUT_1[6627] = 32'b11111111111111111001100100000100;
assign LUT_1[6628] = 32'b00000000000000001100011101001110;
assign LUT_1[6629] = 32'b00000000000000000101101111001010;
assign LUT_1[6630] = 32'b00000000000000001000001011011111;
assign LUT_1[6631] = 32'b00000000000000000001011101011011;
assign LUT_1[6632] = 32'b00000000000000000011110001101100;
assign LUT_1[6633] = 32'b11111111111111111101000011101000;
assign LUT_1[6634] = 32'b11111111111111111111011111111101;
assign LUT_1[6635] = 32'b11111111111111111000110001111001;
assign LUT_1[6636] = 32'b00000000000000001011101011000011;
assign LUT_1[6637] = 32'b00000000000000000100111100111111;
assign LUT_1[6638] = 32'b00000000000000000111011001010100;
assign LUT_1[6639] = 32'b00000000000000000000101011010000;
assign LUT_1[6640] = 32'b00000000000000000110011111011001;
assign LUT_1[6641] = 32'b11111111111111111111110001010101;
assign LUT_1[6642] = 32'b00000000000000000010001101101010;
assign LUT_1[6643] = 32'b11111111111111111011011111100110;
assign LUT_1[6644] = 32'b00000000000000001110011000110000;
assign LUT_1[6645] = 32'b00000000000000000111101010101100;
assign LUT_1[6646] = 32'b00000000000000001010000111000001;
assign LUT_1[6647] = 32'b00000000000000000011011000111101;
assign LUT_1[6648] = 32'b00000000000000000101101101001110;
assign LUT_1[6649] = 32'b11111111111111111110111111001010;
assign LUT_1[6650] = 32'b00000000000000000001011011011111;
assign LUT_1[6651] = 32'b11111111111111111010101101011011;
assign LUT_1[6652] = 32'b00000000000000001101100110100101;
assign LUT_1[6653] = 32'b00000000000000000110111000100001;
assign LUT_1[6654] = 32'b00000000000000001001010100110110;
assign LUT_1[6655] = 32'b00000000000000000010100110110010;
assign LUT_1[6656] = 32'b11111111111111111010100101011110;
assign LUT_1[6657] = 32'b11111111111111110011110111011010;
assign LUT_1[6658] = 32'b11111111111111110110010011101111;
assign LUT_1[6659] = 32'b11111111111111101111100101101011;
assign LUT_1[6660] = 32'b00000000000000000010011110110101;
assign LUT_1[6661] = 32'b11111111111111111011110000110001;
assign LUT_1[6662] = 32'b11111111111111111110001101000110;
assign LUT_1[6663] = 32'b11111111111111110111011111000010;
assign LUT_1[6664] = 32'b11111111111111111001110011010011;
assign LUT_1[6665] = 32'b11111111111111110011000101001111;
assign LUT_1[6666] = 32'b11111111111111110101100001100100;
assign LUT_1[6667] = 32'b11111111111111101110110011100000;
assign LUT_1[6668] = 32'b00000000000000000001101100101010;
assign LUT_1[6669] = 32'b11111111111111111010111110100110;
assign LUT_1[6670] = 32'b11111111111111111101011010111011;
assign LUT_1[6671] = 32'b11111111111111110110101100110111;
assign LUT_1[6672] = 32'b11111111111111111100100001000000;
assign LUT_1[6673] = 32'b11111111111111110101110010111100;
assign LUT_1[6674] = 32'b11111111111111111000001111010001;
assign LUT_1[6675] = 32'b11111111111111110001100001001101;
assign LUT_1[6676] = 32'b00000000000000000100011010010111;
assign LUT_1[6677] = 32'b11111111111111111101101100010011;
assign LUT_1[6678] = 32'b00000000000000000000001000101000;
assign LUT_1[6679] = 32'b11111111111111111001011010100100;
assign LUT_1[6680] = 32'b11111111111111111011101110110101;
assign LUT_1[6681] = 32'b11111111111111110101000000110001;
assign LUT_1[6682] = 32'b11111111111111110111011101000110;
assign LUT_1[6683] = 32'b11111111111111110000101111000010;
assign LUT_1[6684] = 32'b00000000000000000011101000001100;
assign LUT_1[6685] = 32'b11111111111111111100111010001000;
assign LUT_1[6686] = 32'b11111111111111111111010110011101;
assign LUT_1[6687] = 32'b11111111111111111000101000011001;
assign LUT_1[6688] = 32'b11111111111111111011100000011101;
assign LUT_1[6689] = 32'b11111111111111110100110010011001;
assign LUT_1[6690] = 32'b11111111111111110111001110101110;
assign LUT_1[6691] = 32'b11111111111111110000100000101010;
assign LUT_1[6692] = 32'b00000000000000000011011001110100;
assign LUT_1[6693] = 32'b11111111111111111100101011110000;
assign LUT_1[6694] = 32'b11111111111111111111001000000101;
assign LUT_1[6695] = 32'b11111111111111111000011010000001;
assign LUT_1[6696] = 32'b11111111111111111010101110010010;
assign LUT_1[6697] = 32'b11111111111111110100000000001110;
assign LUT_1[6698] = 32'b11111111111111110110011100100011;
assign LUT_1[6699] = 32'b11111111111111101111101110011111;
assign LUT_1[6700] = 32'b00000000000000000010100111101001;
assign LUT_1[6701] = 32'b11111111111111111011111001100101;
assign LUT_1[6702] = 32'b11111111111111111110010101111010;
assign LUT_1[6703] = 32'b11111111111111110111100111110110;
assign LUT_1[6704] = 32'b11111111111111111101011011111111;
assign LUT_1[6705] = 32'b11111111111111110110101101111011;
assign LUT_1[6706] = 32'b11111111111111111001001010010000;
assign LUT_1[6707] = 32'b11111111111111110010011100001100;
assign LUT_1[6708] = 32'b00000000000000000101010101010110;
assign LUT_1[6709] = 32'b11111111111111111110100111010010;
assign LUT_1[6710] = 32'b00000000000000000001000011100111;
assign LUT_1[6711] = 32'b11111111111111111010010101100011;
assign LUT_1[6712] = 32'b11111111111111111100101001110100;
assign LUT_1[6713] = 32'b11111111111111110101111011110000;
assign LUT_1[6714] = 32'b11111111111111111000011000000101;
assign LUT_1[6715] = 32'b11111111111111110001101010000001;
assign LUT_1[6716] = 32'b00000000000000000100100011001011;
assign LUT_1[6717] = 32'b11111111111111111101110101000111;
assign LUT_1[6718] = 32'b00000000000000000000010001011100;
assign LUT_1[6719] = 32'b11111111111111111001100011011000;
assign LUT_1[6720] = 32'b11111111111111111100100011000110;
assign LUT_1[6721] = 32'b11111111111111110101110101000010;
assign LUT_1[6722] = 32'b11111111111111111000010001010111;
assign LUT_1[6723] = 32'b11111111111111110001100011010011;
assign LUT_1[6724] = 32'b00000000000000000100011100011101;
assign LUT_1[6725] = 32'b11111111111111111101101110011001;
assign LUT_1[6726] = 32'b00000000000000000000001010101110;
assign LUT_1[6727] = 32'b11111111111111111001011100101010;
assign LUT_1[6728] = 32'b11111111111111111011110000111011;
assign LUT_1[6729] = 32'b11111111111111110101000010110111;
assign LUT_1[6730] = 32'b11111111111111110111011111001100;
assign LUT_1[6731] = 32'b11111111111111110000110001001000;
assign LUT_1[6732] = 32'b00000000000000000011101010010010;
assign LUT_1[6733] = 32'b11111111111111111100111100001110;
assign LUT_1[6734] = 32'b11111111111111111111011000100011;
assign LUT_1[6735] = 32'b11111111111111111000101010011111;
assign LUT_1[6736] = 32'b11111111111111111110011110101000;
assign LUT_1[6737] = 32'b11111111111111110111110000100100;
assign LUT_1[6738] = 32'b11111111111111111010001100111001;
assign LUT_1[6739] = 32'b11111111111111110011011110110101;
assign LUT_1[6740] = 32'b00000000000000000110010111111111;
assign LUT_1[6741] = 32'b11111111111111111111101001111011;
assign LUT_1[6742] = 32'b00000000000000000010000110010000;
assign LUT_1[6743] = 32'b11111111111111111011011000001100;
assign LUT_1[6744] = 32'b11111111111111111101101100011101;
assign LUT_1[6745] = 32'b11111111111111110110111110011001;
assign LUT_1[6746] = 32'b11111111111111111001011010101110;
assign LUT_1[6747] = 32'b11111111111111110010101100101010;
assign LUT_1[6748] = 32'b00000000000000000101100101110100;
assign LUT_1[6749] = 32'b11111111111111111110110111110000;
assign LUT_1[6750] = 32'b00000000000000000001010100000101;
assign LUT_1[6751] = 32'b11111111111111111010100110000001;
assign LUT_1[6752] = 32'b11111111111111111101011110000101;
assign LUT_1[6753] = 32'b11111111111111110110110000000001;
assign LUT_1[6754] = 32'b11111111111111111001001100010110;
assign LUT_1[6755] = 32'b11111111111111110010011110010010;
assign LUT_1[6756] = 32'b00000000000000000101010111011100;
assign LUT_1[6757] = 32'b11111111111111111110101001011000;
assign LUT_1[6758] = 32'b00000000000000000001000101101101;
assign LUT_1[6759] = 32'b11111111111111111010010111101001;
assign LUT_1[6760] = 32'b11111111111111111100101011111010;
assign LUT_1[6761] = 32'b11111111111111110101111101110110;
assign LUT_1[6762] = 32'b11111111111111111000011010001011;
assign LUT_1[6763] = 32'b11111111111111110001101100000111;
assign LUT_1[6764] = 32'b00000000000000000100100101010001;
assign LUT_1[6765] = 32'b11111111111111111101110111001101;
assign LUT_1[6766] = 32'b00000000000000000000010011100010;
assign LUT_1[6767] = 32'b11111111111111111001100101011110;
assign LUT_1[6768] = 32'b11111111111111111111011001100111;
assign LUT_1[6769] = 32'b11111111111111111000101011100011;
assign LUT_1[6770] = 32'b11111111111111111011000111111000;
assign LUT_1[6771] = 32'b11111111111111110100011001110100;
assign LUT_1[6772] = 32'b00000000000000000111010010111110;
assign LUT_1[6773] = 32'b00000000000000000000100100111010;
assign LUT_1[6774] = 32'b00000000000000000011000001001111;
assign LUT_1[6775] = 32'b11111111111111111100010011001011;
assign LUT_1[6776] = 32'b11111111111111111110100111011100;
assign LUT_1[6777] = 32'b11111111111111110111111001011000;
assign LUT_1[6778] = 32'b11111111111111111010010101101101;
assign LUT_1[6779] = 32'b11111111111111110011100111101001;
assign LUT_1[6780] = 32'b00000000000000000110100000110011;
assign LUT_1[6781] = 32'b11111111111111111111110010101111;
assign LUT_1[6782] = 32'b00000000000000000010001111000100;
assign LUT_1[6783] = 32'b11111111111111111011100001000000;
assign LUT_1[6784] = 32'b11111111111111111101100101100001;
assign LUT_1[6785] = 32'b11111111111111110110110111011101;
assign LUT_1[6786] = 32'b11111111111111111001010011110010;
assign LUT_1[6787] = 32'b11111111111111110010100101101110;
assign LUT_1[6788] = 32'b00000000000000000101011110111000;
assign LUT_1[6789] = 32'b11111111111111111110110000110100;
assign LUT_1[6790] = 32'b00000000000000000001001101001001;
assign LUT_1[6791] = 32'b11111111111111111010011111000101;
assign LUT_1[6792] = 32'b11111111111111111100110011010110;
assign LUT_1[6793] = 32'b11111111111111110110000101010010;
assign LUT_1[6794] = 32'b11111111111111111000100001100111;
assign LUT_1[6795] = 32'b11111111111111110001110011100011;
assign LUT_1[6796] = 32'b00000000000000000100101100101101;
assign LUT_1[6797] = 32'b11111111111111111101111110101001;
assign LUT_1[6798] = 32'b00000000000000000000011010111110;
assign LUT_1[6799] = 32'b11111111111111111001101100111010;
assign LUT_1[6800] = 32'b11111111111111111111100001000011;
assign LUT_1[6801] = 32'b11111111111111111000110010111111;
assign LUT_1[6802] = 32'b11111111111111111011001111010100;
assign LUT_1[6803] = 32'b11111111111111110100100001010000;
assign LUT_1[6804] = 32'b00000000000000000111011010011010;
assign LUT_1[6805] = 32'b00000000000000000000101100010110;
assign LUT_1[6806] = 32'b00000000000000000011001000101011;
assign LUT_1[6807] = 32'b11111111111111111100011010100111;
assign LUT_1[6808] = 32'b11111111111111111110101110111000;
assign LUT_1[6809] = 32'b11111111111111111000000000110100;
assign LUT_1[6810] = 32'b11111111111111111010011101001001;
assign LUT_1[6811] = 32'b11111111111111110011101111000101;
assign LUT_1[6812] = 32'b00000000000000000110101000001111;
assign LUT_1[6813] = 32'b11111111111111111111111010001011;
assign LUT_1[6814] = 32'b00000000000000000010010110100000;
assign LUT_1[6815] = 32'b11111111111111111011101000011100;
assign LUT_1[6816] = 32'b11111111111111111110100000100000;
assign LUT_1[6817] = 32'b11111111111111110111110010011100;
assign LUT_1[6818] = 32'b11111111111111111010001110110001;
assign LUT_1[6819] = 32'b11111111111111110011100000101101;
assign LUT_1[6820] = 32'b00000000000000000110011001110111;
assign LUT_1[6821] = 32'b11111111111111111111101011110011;
assign LUT_1[6822] = 32'b00000000000000000010001000001000;
assign LUT_1[6823] = 32'b11111111111111111011011010000100;
assign LUT_1[6824] = 32'b11111111111111111101101110010101;
assign LUT_1[6825] = 32'b11111111111111110111000000010001;
assign LUT_1[6826] = 32'b11111111111111111001011100100110;
assign LUT_1[6827] = 32'b11111111111111110010101110100010;
assign LUT_1[6828] = 32'b00000000000000000101100111101100;
assign LUT_1[6829] = 32'b11111111111111111110111001101000;
assign LUT_1[6830] = 32'b00000000000000000001010101111101;
assign LUT_1[6831] = 32'b11111111111111111010100111111001;
assign LUT_1[6832] = 32'b00000000000000000000011100000010;
assign LUT_1[6833] = 32'b11111111111111111001101101111110;
assign LUT_1[6834] = 32'b11111111111111111100001010010011;
assign LUT_1[6835] = 32'b11111111111111110101011100001111;
assign LUT_1[6836] = 32'b00000000000000001000010101011001;
assign LUT_1[6837] = 32'b00000000000000000001100111010101;
assign LUT_1[6838] = 32'b00000000000000000100000011101010;
assign LUT_1[6839] = 32'b11111111111111111101010101100110;
assign LUT_1[6840] = 32'b11111111111111111111101001110111;
assign LUT_1[6841] = 32'b11111111111111111000111011110011;
assign LUT_1[6842] = 32'b11111111111111111011011000001000;
assign LUT_1[6843] = 32'b11111111111111110100101010000100;
assign LUT_1[6844] = 32'b00000000000000000111100011001110;
assign LUT_1[6845] = 32'b00000000000000000000110101001010;
assign LUT_1[6846] = 32'b00000000000000000011010001011111;
assign LUT_1[6847] = 32'b11111111111111111100100011011011;
assign LUT_1[6848] = 32'b11111111111111111111100011001001;
assign LUT_1[6849] = 32'b11111111111111111000110101000101;
assign LUT_1[6850] = 32'b11111111111111111011010001011010;
assign LUT_1[6851] = 32'b11111111111111110100100011010110;
assign LUT_1[6852] = 32'b00000000000000000111011100100000;
assign LUT_1[6853] = 32'b00000000000000000000101110011100;
assign LUT_1[6854] = 32'b00000000000000000011001010110001;
assign LUT_1[6855] = 32'b11111111111111111100011100101101;
assign LUT_1[6856] = 32'b11111111111111111110110000111110;
assign LUT_1[6857] = 32'b11111111111111111000000010111010;
assign LUT_1[6858] = 32'b11111111111111111010011111001111;
assign LUT_1[6859] = 32'b11111111111111110011110001001011;
assign LUT_1[6860] = 32'b00000000000000000110101010010101;
assign LUT_1[6861] = 32'b11111111111111111111111100010001;
assign LUT_1[6862] = 32'b00000000000000000010011000100110;
assign LUT_1[6863] = 32'b11111111111111111011101010100010;
assign LUT_1[6864] = 32'b00000000000000000001011110101011;
assign LUT_1[6865] = 32'b11111111111111111010110000100111;
assign LUT_1[6866] = 32'b11111111111111111101001100111100;
assign LUT_1[6867] = 32'b11111111111111110110011110111000;
assign LUT_1[6868] = 32'b00000000000000001001011000000010;
assign LUT_1[6869] = 32'b00000000000000000010101001111110;
assign LUT_1[6870] = 32'b00000000000000000101000110010011;
assign LUT_1[6871] = 32'b11111111111111111110011000001111;
assign LUT_1[6872] = 32'b00000000000000000000101100100000;
assign LUT_1[6873] = 32'b11111111111111111001111110011100;
assign LUT_1[6874] = 32'b11111111111111111100011010110001;
assign LUT_1[6875] = 32'b11111111111111110101101100101101;
assign LUT_1[6876] = 32'b00000000000000001000100101110111;
assign LUT_1[6877] = 32'b00000000000000000001110111110011;
assign LUT_1[6878] = 32'b00000000000000000100010100001000;
assign LUT_1[6879] = 32'b11111111111111111101100110000100;
assign LUT_1[6880] = 32'b00000000000000000000011110001000;
assign LUT_1[6881] = 32'b11111111111111111001110000000100;
assign LUT_1[6882] = 32'b11111111111111111100001100011001;
assign LUT_1[6883] = 32'b11111111111111110101011110010101;
assign LUT_1[6884] = 32'b00000000000000001000010111011111;
assign LUT_1[6885] = 32'b00000000000000000001101001011011;
assign LUT_1[6886] = 32'b00000000000000000100000101110000;
assign LUT_1[6887] = 32'b11111111111111111101010111101100;
assign LUT_1[6888] = 32'b11111111111111111111101011111101;
assign LUT_1[6889] = 32'b11111111111111111000111101111001;
assign LUT_1[6890] = 32'b11111111111111111011011010001110;
assign LUT_1[6891] = 32'b11111111111111110100101100001010;
assign LUT_1[6892] = 32'b00000000000000000111100101010100;
assign LUT_1[6893] = 32'b00000000000000000000110111010000;
assign LUT_1[6894] = 32'b00000000000000000011010011100101;
assign LUT_1[6895] = 32'b11111111111111111100100101100001;
assign LUT_1[6896] = 32'b00000000000000000010011001101010;
assign LUT_1[6897] = 32'b11111111111111111011101011100110;
assign LUT_1[6898] = 32'b11111111111111111110000111111011;
assign LUT_1[6899] = 32'b11111111111111110111011001110111;
assign LUT_1[6900] = 32'b00000000000000001010010011000001;
assign LUT_1[6901] = 32'b00000000000000000011100100111101;
assign LUT_1[6902] = 32'b00000000000000000110000001010010;
assign LUT_1[6903] = 32'b11111111111111111111010011001110;
assign LUT_1[6904] = 32'b00000000000000000001100111011111;
assign LUT_1[6905] = 32'b11111111111111111010111001011011;
assign LUT_1[6906] = 32'b11111111111111111101010101110000;
assign LUT_1[6907] = 32'b11111111111111110110100111101100;
assign LUT_1[6908] = 32'b00000000000000001001100000110110;
assign LUT_1[6909] = 32'b00000000000000000010110010110010;
assign LUT_1[6910] = 32'b00000000000000000101001111000111;
assign LUT_1[6911] = 32'b11111111111111111110100001000011;
assign LUT_1[6912] = 32'b11111111111111111000011001101010;
assign LUT_1[6913] = 32'b11111111111111110001101011100110;
assign LUT_1[6914] = 32'b11111111111111110100000111111011;
assign LUT_1[6915] = 32'b11111111111111101101011001110111;
assign LUT_1[6916] = 32'b00000000000000000000010011000001;
assign LUT_1[6917] = 32'b11111111111111111001100100111101;
assign LUT_1[6918] = 32'b11111111111111111100000001010010;
assign LUT_1[6919] = 32'b11111111111111110101010011001110;
assign LUT_1[6920] = 32'b11111111111111110111100111011111;
assign LUT_1[6921] = 32'b11111111111111110000111001011011;
assign LUT_1[6922] = 32'b11111111111111110011010101110000;
assign LUT_1[6923] = 32'b11111111111111101100100111101100;
assign LUT_1[6924] = 32'b11111111111111111111100000110110;
assign LUT_1[6925] = 32'b11111111111111111000110010110010;
assign LUT_1[6926] = 32'b11111111111111111011001111000111;
assign LUT_1[6927] = 32'b11111111111111110100100001000011;
assign LUT_1[6928] = 32'b11111111111111111010010101001100;
assign LUT_1[6929] = 32'b11111111111111110011100111001000;
assign LUT_1[6930] = 32'b11111111111111110110000011011101;
assign LUT_1[6931] = 32'b11111111111111101111010101011001;
assign LUT_1[6932] = 32'b00000000000000000010001110100011;
assign LUT_1[6933] = 32'b11111111111111111011100000011111;
assign LUT_1[6934] = 32'b11111111111111111101111100110100;
assign LUT_1[6935] = 32'b11111111111111110111001110110000;
assign LUT_1[6936] = 32'b11111111111111111001100011000001;
assign LUT_1[6937] = 32'b11111111111111110010110100111101;
assign LUT_1[6938] = 32'b11111111111111110101010001010010;
assign LUT_1[6939] = 32'b11111111111111101110100011001110;
assign LUT_1[6940] = 32'b00000000000000000001011100011000;
assign LUT_1[6941] = 32'b11111111111111111010101110010100;
assign LUT_1[6942] = 32'b11111111111111111101001010101001;
assign LUT_1[6943] = 32'b11111111111111110110011100100101;
assign LUT_1[6944] = 32'b11111111111111111001010100101001;
assign LUT_1[6945] = 32'b11111111111111110010100110100101;
assign LUT_1[6946] = 32'b11111111111111110101000010111010;
assign LUT_1[6947] = 32'b11111111111111101110010100110110;
assign LUT_1[6948] = 32'b00000000000000000001001110000000;
assign LUT_1[6949] = 32'b11111111111111111010011111111100;
assign LUT_1[6950] = 32'b11111111111111111100111100010001;
assign LUT_1[6951] = 32'b11111111111111110110001110001101;
assign LUT_1[6952] = 32'b11111111111111111000100010011110;
assign LUT_1[6953] = 32'b11111111111111110001110100011010;
assign LUT_1[6954] = 32'b11111111111111110100010000101111;
assign LUT_1[6955] = 32'b11111111111111101101100010101011;
assign LUT_1[6956] = 32'b00000000000000000000011011110101;
assign LUT_1[6957] = 32'b11111111111111111001101101110001;
assign LUT_1[6958] = 32'b11111111111111111100001010000110;
assign LUT_1[6959] = 32'b11111111111111110101011100000010;
assign LUT_1[6960] = 32'b11111111111111111011010000001011;
assign LUT_1[6961] = 32'b11111111111111110100100010000111;
assign LUT_1[6962] = 32'b11111111111111110110111110011100;
assign LUT_1[6963] = 32'b11111111111111110000010000011000;
assign LUT_1[6964] = 32'b00000000000000000011001001100010;
assign LUT_1[6965] = 32'b11111111111111111100011011011110;
assign LUT_1[6966] = 32'b11111111111111111110110111110011;
assign LUT_1[6967] = 32'b11111111111111111000001001101111;
assign LUT_1[6968] = 32'b11111111111111111010011110000000;
assign LUT_1[6969] = 32'b11111111111111110011101111111100;
assign LUT_1[6970] = 32'b11111111111111110110001100010001;
assign LUT_1[6971] = 32'b11111111111111101111011110001101;
assign LUT_1[6972] = 32'b00000000000000000010010111010111;
assign LUT_1[6973] = 32'b11111111111111111011101001010011;
assign LUT_1[6974] = 32'b11111111111111111110000101101000;
assign LUT_1[6975] = 32'b11111111111111110111010111100100;
assign LUT_1[6976] = 32'b11111111111111111010010111010010;
assign LUT_1[6977] = 32'b11111111111111110011101001001110;
assign LUT_1[6978] = 32'b11111111111111110110000101100011;
assign LUT_1[6979] = 32'b11111111111111101111010111011111;
assign LUT_1[6980] = 32'b00000000000000000010010000101001;
assign LUT_1[6981] = 32'b11111111111111111011100010100101;
assign LUT_1[6982] = 32'b11111111111111111101111110111010;
assign LUT_1[6983] = 32'b11111111111111110111010000110110;
assign LUT_1[6984] = 32'b11111111111111111001100101000111;
assign LUT_1[6985] = 32'b11111111111111110010110111000011;
assign LUT_1[6986] = 32'b11111111111111110101010011011000;
assign LUT_1[6987] = 32'b11111111111111101110100101010100;
assign LUT_1[6988] = 32'b00000000000000000001011110011110;
assign LUT_1[6989] = 32'b11111111111111111010110000011010;
assign LUT_1[6990] = 32'b11111111111111111101001100101111;
assign LUT_1[6991] = 32'b11111111111111110110011110101011;
assign LUT_1[6992] = 32'b11111111111111111100010010110100;
assign LUT_1[6993] = 32'b11111111111111110101100100110000;
assign LUT_1[6994] = 32'b11111111111111111000000001000101;
assign LUT_1[6995] = 32'b11111111111111110001010011000001;
assign LUT_1[6996] = 32'b00000000000000000100001100001011;
assign LUT_1[6997] = 32'b11111111111111111101011110000111;
assign LUT_1[6998] = 32'b11111111111111111111111010011100;
assign LUT_1[6999] = 32'b11111111111111111001001100011000;
assign LUT_1[7000] = 32'b11111111111111111011100000101001;
assign LUT_1[7001] = 32'b11111111111111110100110010100101;
assign LUT_1[7002] = 32'b11111111111111110111001110111010;
assign LUT_1[7003] = 32'b11111111111111110000100000110110;
assign LUT_1[7004] = 32'b00000000000000000011011010000000;
assign LUT_1[7005] = 32'b11111111111111111100101011111100;
assign LUT_1[7006] = 32'b11111111111111111111001000010001;
assign LUT_1[7007] = 32'b11111111111111111000011010001101;
assign LUT_1[7008] = 32'b11111111111111111011010010010001;
assign LUT_1[7009] = 32'b11111111111111110100100100001101;
assign LUT_1[7010] = 32'b11111111111111110111000000100010;
assign LUT_1[7011] = 32'b11111111111111110000010010011110;
assign LUT_1[7012] = 32'b00000000000000000011001011101000;
assign LUT_1[7013] = 32'b11111111111111111100011101100100;
assign LUT_1[7014] = 32'b11111111111111111110111001111001;
assign LUT_1[7015] = 32'b11111111111111111000001011110101;
assign LUT_1[7016] = 32'b11111111111111111010100000000110;
assign LUT_1[7017] = 32'b11111111111111110011110010000010;
assign LUT_1[7018] = 32'b11111111111111110110001110010111;
assign LUT_1[7019] = 32'b11111111111111101111100000010011;
assign LUT_1[7020] = 32'b00000000000000000010011001011101;
assign LUT_1[7021] = 32'b11111111111111111011101011011001;
assign LUT_1[7022] = 32'b11111111111111111110000111101110;
assign LUT_1[7023] = 32'b11111111111111110111011001101010;
assign LUT_1[7024] = 32'b11111111111111111101001101110011;
assign LUT_1[7025] = 32'b11111111111111110110011111101111;
assign LUT_1[7026] = 32'b11111111111111111000111100000100;
assign LUT_1[7027] = 32'b11111111111111110010001110000000;
assign LUT_1[7028] = 32'b00000000000000000101000111001010;
assign LUT_1[7029] = 32'b11111111111111111110011001000110;
assign LUT_1[7030] = 32'b00000000000000000000110101011011;
assign LUT_1[7031] = 32'b11111111111111111010000111010111;
assign LUT_1[7032] = 32'b11111111111111111100011011101000;
assign LUT_1[7033] = 32'b11111111111111110101101101100100;
assign LUT_1[7034] = 32'b11111111111111111000001001111001;
assign LUT_1[7035] = 32'b11111111111111110001011011110101;
assign LUT_1[7036] = 32'b00000000000000000100010100111111;
assign LUT_1[7037] = 32'b11111111111111111101100110111011;
assign LUT_1[7038] = 32'b00000000000000000000000011010000;
assign LUT_1[7039] = 32'b11111111111111111001010101001100;
assign LUT_1[7040] = 32'b11111111111111111011011001101101;
assign LUT_1[7041] = 32'b11111111111111110100101011101001;
assign LUT_1[7042] = 32'b11111111111111110111000111111110;
assign LUT_1[7043] = 32'b11111111111111110000011001111010;
assign LUT_1[7044] = 32'b00000000000000000011010011000100;
assign LUT_1[7045] = 32'b11111111111111111100100101000000;
assign LUT_1[7046] = 32'b11111111111111111111000001010101;
assign LUT_1[7047] = 32'b11111111111111111000010011010001;
assign LUT_1[7048] = 32'b11111111111111111010100111100010;
assign LUT_1[7049] = 32'b11111111111111110011111001011110;
assign LUT_1[7050] = 32'b11111111111111110110010101110011;
assign LUT_1[7051] = 32'b11111111111111101111100111101111;
assign LUT_1[7052] = 32'b00000000000000000010100000111001;
assign LUT_1[7053] = 32'b11111111111111111011110010110101;
assign LUT_1[7054] = 32'b11111111111111111110001111001010;
assign LUT_1[7055] = 32'b11111111111111110111100001000110;
assign LUT_1[7056] = 32'b11111111111111111101010101001111;
assign LUT_1[7057] = 32'b11111111111111110110100111001011;
assign LUT_1[7058] = 32'b11111111111111111001000011100000;
assign LUT_1[7059] = 32'b11111111111111110010010101011100;
assign LUT_1[7060] = 32'b00000000000000000101001110100110;
assign LUT_1[7061] = 32'b11111111111111111110100000100010;
assign LUT_1[7062] = 32'b00000000000000000000111100110111;
assign LUT_1[7063] = 32'b11111111111111111010001110110011;
assign LUT_1[7064] = 32'b11111111111111111100100011000100;
assign LUT_1[7065] = 32'b11111111111111110101110101000000;
assign LUT_1[7066] = 32'b11111111111111111000010001010101;
assign LUT_1[7067] = 32'b11111111111111110001100011010001;
assign LUT_1[7068] = 32'b00000000000000000100011100011011;
assign LUT_1[7069] = 32'b11111111111111111101101110010111;
assign LUT_1[7070] = 32'b00000000000000000000001010101100;
assign LUT_1[7071] = 32'b11111111111111111001011100101000;
assign LUT_1[7072] = 32'b11111111111111111100010100101100;
assign LUT_1[7073] = 32'b11111111111111110101100110101000;
assign LUT_1[7074] = 32'b11111111111111111000000010111101;
assign LUT_1[7075] = 32'b11111111111111110001010100111001;
assign LUT_1[7076] = 32'b00000000000000000100001110000011;
assign LUT_1[7077] = 32'b11111111111111111101011111111111;
assign LUT_1[7078] = 32'b11111111111111111111111100010100;
assign LUT_1[7079] = 32'b11111111111111111001001110010000;
assign LUT_1[7080] = 32'b11111111111111111011100010100001;
assign LUT_1[7081] = 32'b11111111111111110100110100011101;
assign LUT_1[7082] = 32'b11111111111111110111010000110010;
assign LUT_1[7083] = 32'b11111111111111110000100010101110;
assign LUT_1[7084] = 32'b00000000000000000011011011111000;
assign LUT_1[7085] = 32'b11111111111111111100101101110100;
assign LUT_1[7086] = 32'b11111111111111111111001010001001;
assign LUT_1[7087] = 32'b11111111111111111000011100000101;
assign LUT_1[7088] = 32'b11111111111111111110010000001110;
assign LUT_1[7089] = 32'b11111111111111110111100010001010;
assign LUT_1[7090] = 32'b11111111111111111001111110011111;
assign LUT_1[7091] = 32'b11111111111111110011010000011011;
assign LUT_1[7092] = 32'b00000000000000000110001001100101;
assign LUT_1[7093] = 32'b11111111111111111111011011100001;
assign LUT_1[7094] = 32'b00000000000000000001110111110110;
assign LUT_1[7095] = 32'b11111111111111111011001001110010;
assign LUT_1[7096] = 32'b11111111111111111101011110000011;
assign LUT_1[7097] = 32'b11111111111111110110101111111111;
assign LUT_1[7098] = 32'b11111111111111111001001100010100;
assign LUT_1[7099] = 32'b11111111111111110010011110010000;
assign LUT_1[7100] = 32'b00000000000000000101010111011010;
assign LUT_1[7101] = 32'b11111111111111111110101001010110;
assign LUT_1[7102] = 32'b00000000000000000001000101101011;
assign LUT_1[7103] = 32'b11111111111111111010010111100111;
assign LUT_1[7104] = 32'b11111111111111111101010111010101;
assign LUT_1[7105] = 32'b11111111111111110110101001010001;
assign LUT_1[7106] = 32'b11111111111111111001000101100110;
assign LUT_1[7107] = 32'b11111111111111110010010111100010;
assign LUT_1[7108] = 32'b00000000000000000101010000101100;
assign LUT_1[7109] = 32'b11111111111111111110100010101000;
assign LUT_1[7110] = 32'b00000000000000000000111110111101;
assign LUT_1[7111] = 32'b11111111111111111010010000111001;
assign LUT_1[7112] = 32'b11111111111111111100100101001010;
assign LUT_1[7113] = 32'b11111111111111110101110111000110;
assign LUT_1[7114] = 32'b11111111111111111000010011011011;
assign LUT_1[7115] = 32'b11111111111111110001100101010111;
assign LUT_1[7116] = 32'b00000000000000000100011110100001;
assign LUT_1[7117] = 32'b11111111111111111101110000011101;
assign LUT_1[7118] = 32'b00000000000000000000001100110010;
assign LUT_1[7119] = 32'b11111111111111111001011110101110;
assign LUT_1[7120] = 32'b11111111111111111111010010110111;
assign LUT_1[7121] = 32'b11111111111111111000100100110011;
assign LUT_1[7122] = 32'b11111111111111111011000001001000;
assign LUT_1[7123] = 32'b11111111111111110100010011000100;
assign LUT_1[7124] = 32'b00000000000000000111001100001110;
assign LUT_1[7125] = 32'b00000000000000000000011110001010;
assign LUT_1[7126] = 32'b00000000000000000010111010011111;
assign LUT_1[7127] = 32'b11111111111111111100001100011011;
assign LUT_1[7128] = 32'b11111111111111111110100000101100;
assign LUT_1[7129] = 32'b11111111111111110111110010101000;
assign LUT_1[7130] = 32'b11111111111111111010001110111101;
assign LUT_1[7131] = 32'b11111111111111110011100000111001;
assign LUT_1[7132] = 32'b00000000000000000110011010000011;
assign LUT_1[7133] = 32'b11111111111111111111101011111111;
assign LUT_1[7134] = 32'b00000000000000000010001000010100;
assign LUT_1[7135] = 32'b11111111111111111011011010010000;
assign LUT_1[7136] = 32'b11111111111111111110010010010100;
assign LUT_1[7137] = 32'b11111111111111110111100100010000;
assign LUT_1[7138] = 32'b11111111111111111010000000100101;
assign LUT_1[7139] = 32'b11111111111111110011010010100001;
assign LUT_1[7140] = 32'b00000000000000000110001011101011;
assign LUT_1[7141] = 32'b11111111111111111111011101100111;
assign LUT_1[7142] = 32'b00000000000000000001111001111100;
assign LUT_1[7143] = 32'b11111111111111111011001011111000;
assign LUT_1[7144] = 32'b11111111111111111101100000001001;
assign LUT_1[7145] = 32'b11111111111111110110110010000101;
assign LUT_1[7146] = 32'b11111111111111111001001110011010;
assign LUT_1[7147] = 32'b11111111111111110010100000010110;
assign LUT_1[7148] = 32'b00000000000000000101011001100000;
assign LUT_1[7149] = 32'b11111111111111111110101011011100;
assign LUT_1[7150] = 32'b00000000000000000001000111110001;
assign LUT_1[7151] = 32'b11111111111111111010011001101101;
assign LUT_1[7152] = 32'b00000000000000000000001101110110;
assign LUT_1[7153] = 32'b11111111111111111001011111110010;
assign LUT_1[7154] = 32'b11111111111111111011111100000111;
assign LUT_1[7155] = 32'b11111111111111110101001110000011;
assign LUT_1[7156] = 32'b00000000000000001000000111001101;
assign LUT_1[7157] = 32'b00000000000000000001011001001001;
assign LUT_1[7158] = 32'b00000000000000000011110101011110;
assign LUT_1[7159] = 32'b11111111111111111101000111011010;
assign LUT_1[7160] = 32'b11111111111111111111011011101011;
assign LUT_1[7161] = 32'b11111111111111111000101101100111;
assign LUT_1[7162] = 32'b11111111111111111011001001111100;
assign LUT_1[7163] = 32'b11111111111111110100011011111000;
assign LUT_1[7164] = 32'b00000000000000000111010101000010;
assign LUT_1[7165] = 32'b00000000000000000000100110111110;
assign LUT_1[7166] = 32'b00000000000000000011000011010011;
assign LUT_1[7167] = 32'b11111111111111111100010101001111;
assign LUT_1[7168] = 32'b00000000000000000111001101110001;
assign LUT_1[7169] = 32'b00000000000000000000011111101101;
assign LUT_1[7170] = 32'b00000000000000000010111100000010;
assign LUT_1[7171] = 32'b11111111111111111100001101111110;
assign LUT_1[7172] = 32'b00000000000000001111000111001000;
assign LUT_1[7173] = 32'b00000000000000001000011001000100;
assign LUT_1[7174] = 32'b00000000000000001010110101011001;
assign LUT_1[7175] = 32'b00000000000000000100000111010101;
assign LUT_1[7176] = 32'b00000000000000000110011011100110;
assign LUT_1[7177] = 32'b11111111111111111111101101100010;
assign LUT_1[7178] = 32'b00000000000000000010001001110111;
assign LUT_1[7179] = 32'b11111111111111111011011011110011;
assign LUT_1[7180] = 32'b00000000000000001110010100111101;
assign LUT_1[7181] = 32'b00000000000000000111100110111001;
assign LUT_1[7182] = 32'b00000000000000001010000011001110;
assign LUT_1[7183] = 32'b00000000000000000011010101001010;
assign LUT_1[7184] = 32'b00000000000000001001001001010011;
assign LUT_1[7185] = 32'b00000000000000000010011011001111;
assign LUT_1[7186] = 32'b00000000000000000100110111100100;
assign LUT_1[7187] = 32'b11111111111111111110001001100000;
assign LUT_1[7188] = 32'b00000000000000010001000010101010;
assign LUT_1[7189] = 32'b00000000000000001010010100100110;
assign LUT_1[7190] = 32'b00000000000000001100110000111011;
assign LUT_1[7191] = 32'b00000000000000000110000010110111;
assign LUT_1[7192] = 32'b00000000000000001000010111001000;
assign LUT_1[7193] = 32'b00000000000000000001101001000100;
assign LUT_1[7194] = 32'b00000000000000000100000101011001;
assign LUT_1[7195] = 32'b11111111111111111101010111010101;
assign LUT_1[7196] = 32'b00000000000000010000010000011111;
assign LUT_1[7197] = 32'b00000000000000001001100010011011;
assign LUT_1[7198] = 32'b00000000000000001011111110110000;
assign LUT_1[7199] = 32'b00000000000000000101010000101100;
assign LUT_1[7200] = 32'b00000000000000001000001000110000;
assign LUT_1[7201] = 32'b00000000000000000001011010101100;
assign LUT_1[7202] = 32'b00000000000000000011110111000001;
assign LUT_1[7203] = 32'b11111111111111111101001000111101;
assign LUT_1[7204] = 32'b00000000000000010000000010000111;
assign LUT_1[7205] = 32'b00000000000000001001010100000011;
assign LUT_1[7206] = 32'b00000000000000001011110000011000;
assign LUT_1[7207] = 32'b00000000000000000101000010010100;
assign LUT_1[7208] = 32'b00000000000000000111010110100101;
assign LUT_1[7209] = 32'b00000000000000000000101000100001;
assign LUT_1[7210] = 32'b00000000000000000011000100110110;
assign LUT_1[7211] = 32'b11111111111111111100010110110010;
assign LUT_1[7212] = 32'b00000000000000001111001111111100;
assign LUT_1[7213] = 32'b00000000000000001000100001111000;
assign LUT_1[7214] = 32'b00000000000000001010111110001101;
assign LUT_1[7215] = 32'b00000000000000000100010000001001;
assign LUT_1[7216] = 32'b00000000000000001010000100010010;
assign LUT_1[7217] = 32'b00000000000000000011010110001110;
assign LUT_1[7218] = 32'b00000000000000000101110010100011;
assign LUT_1[7219] = 32'b11111111111111111111000100011111;
assign LUT_1[7220] = 32'b00000000000000010001111101101001;
assign LUT_1[7221] = 32'b00000000000000001011001111100101;
assign LUT_1[7222] = 32'b00000000000000001101101011111010;
assign LUT_1[7223] = 32'b00000000000000000110111101110110;
assign LUT_1[7224] = 32'b00000000000000001001010010000111;
assign LUT_1[7225] = 32'b00000000000000000010100100000011;
assign LUT_1[7226] = 32'b00000000000000000101000000011000;
assign LUT_1[7227] = 32'b11111111111111111110010010010100;
assign LUT_1[7228] = 32'b00000000000000010001001011011110;
assign LUT_1[7229] = 32'b00000000000000001010011101011010;
assign LUT_1[7230] = 32'b00000000000000001100111001101111;
assign LUT_1[7231] = 32'b00000000000000000110001011101011;
assign LUT_1[7232] = 32'b00000000000000001001001011011001;
assign LUT_1[7233] = 32'b00000000000000000010011101010101;
assign LUT_1[7234] = 32'b00000000000000000100111001101010;
assign LUT_1[7235] = 32'b11111111111111111110001011100110;
assign LUT_1[7236] = 32'b00000000000000010001000100110000;
assign LUT_1[7237] = 32'b00000000000000001010010110101100;
assign LUT_1[7238] = 32'b00000000000000001100110011000001;
assign LUT_1[7239] = 32'b00000000000000000110000100111101;
assign LUT_1[7240] = 32'b00000000000000001000011001001110;
assign LUT_1[7241] = 32'b00000000000000000001101011001010;
assign LUT_1[7242] = 32'b00000000000000000100000111011111;
assign LUT_1[7243] = 32'b11111111111111111101011001011011;
assign LUT_1[7244] = 32'b00000000000000010000010010100101;
assign LUT_1[7245] = 32'b00000000000000001001100100100001;
assign LUT_1[7246] = 32'b00000000000000001100000000110110;
assign LUT_1[7247] = 32'b00000000000000000101010010110010;
assign LUT_1[7248] = 32'b00000000000000001011000110111011;
assign LUT_1[7249] = 32'b00000000000000000100011000110111;
assign LUT_1[7250] = 32'b00000000000000000110110101001100;
assign LUT_1[7251] = 32'b00000000000000000000000111001000;
assign LUT_1[7252] = 32'b00000000000000010011000000010010;
assign LUT_1[7253] = 32'b00000000000000001100010010001110;
assign LUT_1[7254] = 32'b00000000000000001110101110100011;
assign LUT_1[7255] = 32'b00000000000000001000000000011111;
assign LUT_1[7256] = 32'b00000000000000001010010100110000;
assign LUT_1[7257] = 32'b00000000000000000011100110101100;
assign LUT_1[7258] = 32'b00000000000000000110000011000001;
assign LUT_1[7259] = 32'b11111111111111111111010100111101;
assign LUT_1[7260] = 32'b00000000000000010010001110000111;
assign LUT_1[7261] = 32'b00000000000000001011100000000011;
assign LUT_1[7262] = 32'b00000000000000001101111100011000;
assign LUT_1[7263] = 32'b00000000000000000111001110010100;
assign LUT_1[7264] = 32'b00000000000000001010000110011000;
assign LUT_1[7265] = 32'b00000000000000000011011000010100;
assign LUT_1[7266] = 32'b00000000000000000101110100101001;
assign LUT_1[7267] = 32'b11111111111111111111000110100101;
assign LUT_1[7268] = 32'b00000000000000010001111111101111;
assign LUT_1[7269] = 32'b00000000000000001011010001101011;
assign LUT_1[7270] = 32'b00000000000000001101101110000000;
assign LUT_1[7271] = 32'b00000000000000000110111111111100;
assign LUT_1[7272] = 32'b00000000000000001001010100001101;
assign LUT_1[7273] = 32'b00000000000000000010100110001001;
assign LUT_1[7274] = 32'b00000000000000000101000010011110;
assign LUT_1[7275] = 32'b11111111111111111110010100011010;
assign LUT_1[7276] = 32'b00000000000000010001001101100100;
assign LUT_1[7277] = 32'b00000000000000001010011111100000;
assign LUT_1[7278] = 32'b00000000000000001100111011110101;
assign LUT_1[7279] = 32'b00000000000000000110001101110001;
assign LUT_1[7280] = 32'b00000000000000001100000001111010;
assign LUT_1[7281] = 32'b00000000000000000101010011110110;
assign LUT_1[7282] = 32'b00000000000000000111110000001011;
assign LUT_1[7283] = 32'b00000000000000000001000010000111;
assign LUT_1[7284] = 32'b00000000000000010011111011010001;
assign LUT_1[7285] = 32'b00000000000000001101001101001101;
assign LUT_1[7286] = 32'b00000000000000001111101001100010;
assign LUT_1[7287] = 32'b00000000000000001000111011011110;
assign LUT_1[7288] = 32'b00000000000000001011001111101111;
assign LUT_1[7289] = 32'b00000000000000000100100001101011;
assign LUT_1[7290] = 32'b00000000000000000110111110000000;
assign LUT_1[7291] = 32'b00000000000000000000001111111100;
assign LUT_1[7292] = 32'b00000000000000010011001001000110;
assign LUT_1[7293] = 32'b00000000000000001100011011000010;
assign LUT_1[7294] = 32'b00000000000000001110110111010111;
assign LUT_1[7295] = 32'b00000000000000001000001001010011;
assign LUT_1[7296] = 32'b00000000000000001010001101110100;
assign LUT_1[7297] = 32'b00000000000000000011011111110000;
assign LUT_1[7298] = 32'b00000000000000000101111100000101;
assign LUT_1[7299] = 32'b11111111111111111111001110000001;
assign LUT_1[7300] = 32'b00000000000000010010000111001011;
assign LUT_1[7301] = 32'b00000000000000001011011001000111;
assign LUT_1[7302] = 32'b00000000000000001101110101011100;
assign LUT_1[7303] = 32'b00000000000000000111000111011000;
assign LUT_1[7304] = 32'b00000000000000001001011011101001;
assign LUT_1[7305] = 32'b00000000000000000010101101100101;
assign LUT_1[7306] = 32'b00000000000000000101001001111010;
assign LUT_1[7307] = 32'b11111111111111111110011011110110;
assign LUT_1[7308] = 32'b00000000000000010001010101000000;
assign LUT_1[7309] = 32'b00000000000000001010100110111100;
assign LUT_1[7310] = 32'b00000000000000001101000011010001;
assign LUT_1[7311] = 32'b00000000000000000110010101001101;
assign LUT_1[7312] = 32'b00000000000000001100001001010110;
assign LUT_1[7313] = 32'b00000000000000000101011011010010;
assign LUT_1[7314] = 32'b00000000000000000111110111100111;
assign LUT_1[7315] = 32'b00000000000000000001001001100011;
assign LUT_1[7316] = 32'b00000000000000010100000010101101;
assign LUT_1[7317] = 32'b00000000000000001101010100101001;
assign LUT_1[7318] = 32'b00000000000000001111110000111110;
assign LUT_1[7319] = 32'b00000000000000001001000010111010;
assign LUT_1[7320] = 32'b00000000000000001011010111001011;
assign LUT_1[7321] = 32'b00000000000000000100101001000111;
assign LUT_1[7322] = 32'b00000000000000000111000101011100;
assign LUT_1[7323] = 32'b00000000000000000000010111011000;
assign LUT_1[7324] = 32'b00000000000000010011010000100010;
assign LUT_1[7325] = 32'b00000000000000001100100010011110;
assign LUT_1[7326] = 32'b00000000000000001110111110110011;
assign LUT_1[7327] = 32'b00000000000000001000010000101111;
assign LUT_1[7328] = 32'b00000000000000001011001000110011;
assign LUT_1[7329] = 32'b00000000000000000100011010101111;
assign LUT_1[7330] = 32'b00000000000000000110110111000100;
assign LUT_1[7331] = 32'b00000000000000000000001001000000;
assign LUT_1[7332] = 32'b00000000000000010011000010001010;
assign LUT_1[7333] = 32'b00000000000000001100010100000110;
assign LUT_1[7334] = 32'b00000000000000001110110000011011;
assign LUT_1[7335] = 32'b00000000000000001000000010010111;
assign LUT_1[7336] = 32'b00000000000000001010010110101000;
assign LUT_1[7337] = 32'b00000000000000000011101000100100;
assign LUT_1[7338] = 32'b00000000000000000110000100111001;
assign LUT_1[7339] = 32'b11111111111111111111010110110101;
assign LUT_1[7340] = 32'b00000000000000010010001111111111;
assign LUT_1[7341] = 32'b00000000000000001011100001111011;
assign LUT_1[7342] = 32'b00000000000000001101111110010000;
assign LUT_1[7343] = 32'b00000000000000000111010000001100;
assign LUT_1[7344] = 32'b00000000000000001101000100010101;
assign LUT_1[7345] = 32'b00000000000000000110010110010001;
assign LUT_1[7346] = 32'b00000000000000001000110010100110;
assign LUT_1[7347] = 32'b00000000000000000010000100100010;
assign LUT_1[7348] = 32'b00000000000000010100111101101100;
assign LUT_1[7349] = 32'b00000000000000001110001111101000;
assign LUT_1[7350] = 32'b00000000000000010000101011111101;
assign LUT_1[7351] = 32'b00000000000000001001111101111001;
assign LUT_1[7352] = 32'b00000000000000001100010010001010;
assign LUT_1[7353] = 32'b00000000000000000101100100000110;
assign LUT_1[7354] = 32'b00000000000000001000000000011011;
assign LUT_1[7355] = 32'b00000000000000000001010010010111;
assign LUT_1[7356] = 32'b00000000000000010100001011100001;
assign LUT_1[7357] = 32'b00000000000000001101011101011101;
assign LUT_1[7358] = 32'b00000000000000001111111001110010;
assign LUT_1[7359] = 32'b00000000000000001001001011101110;
assign LUT_1[7360] = 32'b00000000000000001100001011011100;
assign LUT_1[7361] = 32'b00000000000000000101011101011000;
assign LUT_1[7362] = 32'b00000000000000000111111001101101;
assign LUT_1[7363] = 32'b00000000000000000001001011101001;
assign LUT_1[7364] = 32'b00000000000000010100000100110011;
assign LUT_1[7365] = 32'b00000000000000001101010110101111;
assign LUT_1[7366] = 32'b00000000000000001111110011000100;
assign LUT_1[7367] = 32'b00000000000000001001000101000000;
assign LUT_1[7368] = 32'b00000000000000001011011001010001;
assign LUT_1[7369] = 32'b00000000000000000100101011001101;
assign LUT_1[7370] = 32'b00000000000000000111000111100010;
assign LUT_1[7371] = 32'b00000000000000000000011001011110;
assign LUT_1[7372] = 32'b00000000000000010011010010101000;
assign LUT_1[7373] = 32'b00000000000000001100100100100100;
assign LUT_1[7374] = 32'b00000000000000001111000000111001;
assign LUT_1[7375] = 32'b00000000000000001000010010110101;
assign LUT_1[7376] = 32'b00000000000000001110000110111110;
assign LUT_1[7377] = 32'b00000000000000000111011000111010;
assign LUT_1[7378] = 32'b00000000000000001001110101001111;
assign LUT_1[7379] = 32'b00000000000000000011000111001011;
assign LUT_1[7380] = 32'b00000000000000010110000000010101;
assign LUT_1[7381] = 32'b00000000000000001111010010010001;
assign LUT_1[7382] = 32'b00000000000000010001101110100110;
assign LUT_1[7383] = 32'b00000000000000001011000000100010;
assign LUT_1[7384] = 32'b00000000000000001101010100110011;
assign LUT_1[7385] = 32'b00000000000000000110100110101111;
assign LUT_1[7386] = 32'b00000000000000001001000011000100;
assign LUT_1[7387] = 32'b00000000000000000010010101000000;
assign LUT_1[7388] = 32'b00000000000000010101001110001010;
assign LUT_1[7389] = 32'b00000000000000001110100000000110;
assign LUT_1[7390] = 32'b00000000000000010000111100011011;
assign LUT_1[7391] = 32'b00000000000000001010001110010111;
assign LUT_1[7392] = 32'b00000000000000001101000110011011;
assign LUT_1[7393] = 32'b00000000000000000110011000010111;
assign LUT_1[7394] = 32'b00000000000000001000110100101100;
assign LUT_1[7395] = 32'b00000000000000000010000110101000;
assign LUT_1[7396] = 32'b00000000000000010100111111110010;
assign LUT_1[7397] = 32'b00000000000000001110010001101110;
assign LUT_1[7398] = 32'b00000000000000010000101110000011;
assign LUT_1[7399] = 32'b00000000000000001001111111111111;
assign LUT_1[7400] = 32'b00000000000000001100010100010000;
assign LUT_1[7401] = 32'b00000000000000000101100110001100;
assign LUT_1[7402] = 32'b00000000000000001000000010100001;
assign LUT_1[7403] = 32'b00000000000000000001010100011101;
assign LUT_1[7404] = 32'b00000000000000010100001101100111;
assign LUT_1[7405] = 32'b00000000000000001101011111100011;
assign LUT_1[7406] = 32'b00000000000000001111111011111000;
assign LUT_1[7407] = 32'b00000000000000001001001101110100;
assign LUT_1[7408] = 32'b00000000000000001111000001111101;
assign LUT_1[7409] = 32'b00000000000000001000010011111001;
assign LUT_1[7410] = 32'b00000000000000001010110000001110;
assign LUT_1[7411] = 32'b00000000000000000100000010001010;
assign LUT_1[7412] = 32'b00000000000000010110111011010100;
assign LUT_1[7413] = 32'b00000000000000010000001101010000;
assign LUT_1[7414] = 32'b00000000000000010010101001100101;
assign LUT_1[7415] = 32'b00000000000000001011111011100001;
assign LUT_1[7416] = 32'b00000000000000001110001111110010;
assign LUT_1[7417] = 32'b00000000000000000111100001101110;
assign LUT_1[7418] = 32'b00000000000000001001111110000011;
assign LUT_1[7419] = 32'b00000000000000000011001111111111;
assign LUT_1[7420] = 32'b00000000000000010110001001001001;
assign LUT_1[7421] = 32'b00000000000000001111011011000101;
assign LUT_1[7422] = 32'b00000000000000010001110111011010;
assign LUT_1[7423] = 32'b00000000000000001011001001010110;
assign LUT_1[7424] = 32'b00000000000000000101000001111101;
assign LUT_1[7425] = 32'b11111111111111111110010011111001;
assign LUT_1[7426] = 32'b00000000000000000000110000001110;
assign LUT_1[7427] = 32'b11111111111111111010000010001010;
assign LUT_1[7428] = 32'b00000000000000001100111011010100;
assign LUT_1[7429] = 32'b00000000000000000110001101010000;
assign LUT_1[7430] = 32'b00000000000000001000101001100101;
assign LUT_1[7431] = 32'b00000000000000000001111011100001;
assign LUT_1[7432] = 32'b00000000000000000100001111110010;
assign LUT_1[7433] = 32'b11111111111111111101100001101110;
assign LUT_1[7434] = 32'b11111111111111111111111110000011;
assign LUT_1[7435] = 32'b11111111111111111001001111111111;
assign LUT_1[7436] = 32'b00000000000000001100001001001001;
assign LUT_1[7437] = 32'b00000000000000000101011011000101;
assign LUT_1[7438] = 32'b00000000000000000111110111011010;
assign LUT_1[7439] = 32'b00000000000000000001001001010110;
assign LUT_1[7440] = 32'b00000000000000000110111101011111;
assign LUT_1[7441] = 32'b00000000000000000000001111011011;
assign LUT_1[7442] = 32'b00000000000000000010101011110000;
assign LUT_1[7443] = 32'b11111111111111111011111101101100;
assign LUT_1[7444] = 32'b00000000000000001110110110110110;
assign LUT_1[7445] = 32'b00000000000000001000001000110010;
assign LUT_1[7446] = 32'b00000000000000001010100101000111;
assign LUT_1[7447] = 32'b00000000000000000011110111000011;
assign LUT_1[7448] = 32'b00000000000000000110001011010100;
assign LUT_1[7449] = 32'b11111111111111111111011101010000;
assign LUT_1[7450] = 32'b00000000000000000001111001100101;
assign LUT_1[7451] = 32'b11111111111111111011001011100001;
assign LUT_1[7452] = 32'b00000000000000001110000100101011;
assign LUT_1[7453] = 32'b00000000000000000111010110100111;
assign LUT_1[7454] = 32'b00000000000000001001110010111100;
assign LUT_1[7455] = 32'b00000000000000000011000100111000;
assign LUT_1[7456] = 32'b00000000000000000101111100111100;
assign LUT_1[7457] = 32'b11111111111111111111001110111000;
assign LUT_1[7458] = 32'b00000000000000000001101011001101;
assign LUT_1[7459] = 32'b11111111111111111010111101001001;
assign LUT_1[7460] = 32'b00000000000000001101110110010011;
assign LUT_1[7461] = 32'b00000000000000000111001000001111;
assign LUT_1[7462] = 32'b00000000000000001001100100100100;
assign LUT_1[7463] = 32'b00000000000000000010110110100000;
assign LUT_1[7464] = 32'b00000000000000000101001010110001;
assign LUT_1[7465] = 32'b11111111111111111110011100101101;
assign LUT_1[7466] = 32'b00000000000000000000111001000010;
assign LUT_1[7467] = 32'b11111111111111111010001010111110;
assign LUT_1[7468] = 32'b00000000000000001101000100001000;
assign LUT_1[7469] = 32'b00000000000000000110010110000100;
assign LUT_1[7470] = 32'b00000000000000001000110010011001;
assign LUT_1[7471] = 32'b00000000000000000010000100010101;
assign LUT_1[7472] = 32'b00000000000000000111111000011110;
assign LUT_1[7473] = 32'b00000000000000000001001010011010;
assign LUT_1[7474] = 32'b00000000000000000011100110101111;
assign LUT_1[7475] = 32'b11111111111111111100111000101011;
assign LUT_1[7476] = 32'b00000000000000001111110001110101;
assign LUT_1[7477] = 32'b00000000000000001001000011110001;
assign LUT_1[7478] = 32'b00000000000000001011100000000110;
assign LUT_1[7479] = 32'b00000000000000000100110010000010;
assign LUT_1[7480] = 32'b00000000000000000111000110010011;
assign LUT_1[7481] = 32'b00000000000000000000011000001111;
assign LUT_1[7482] = 32'b00000000000000000010110100100100;
assign LUT_1[7483] = 32'b11111111111111111100000110100000;
assign LUT_1[7484] = 32'b00000000000000001110111111101010;
assign LUT_1[7485] = 32'b00000000000000001000010001100110;
assign LUT_1[7486] = 32'b00000000000000001010101101111011;
assign LUT_1[7487] = 32'b00000000000000000011111111110111;
assign LUT_1[7488] = 32'b00000000000000000110111111100101;
assign LUT_1[7489] = 32'b00000000000000000000010001100001;
assign LUT_1[7490] = 32'b00000000000000000010101101110110;
assign LUT_1[7491] = 32'b11111111111111111011111111110010;
assign LUT_1[7492] = 32'b00000000000000001110111000111100;
assign LUT_1[7493] = 32'b00000000000000001000001010111000;
assign LUT_1[7494] = 32'b00000000000000001010100111001101;
assign LUT_1[7495] = 32'b00000000000000000011111001001001;
assign LUT_1[7496] = 32'b00000000000000000110001101011010;
assign LUT_1[7497] = 32'b11111111111111111111011111010110;
assign LUT_1[7498] = 32'b00000000000000000001111011101011;
assign LUT_1[7499] = 32'b11111111111111111011001101100111;
assign LUT_1[7500] = 32'b00000000000000001110000110110001;
assign LUT_1[7501] = 32'b00000000000000000111011000101101;
assign LUT_1[7502] = 32'b00000000000000001001110101000010;
assign LUT_1[7503] = 32'b00000000000000000011000110111110;
assign LUT_1[7504] = 32'b00000000000000001000111011000111;
assign LUT_1[7505] = 32'b00000000000000000010001101000011;
assign LUT_1[7506] = 32'b00000000000000000100101001011000;
assign LUT_1[7507] = 32'b11111111111111111101111011010100;
assign LUT_1[7508] = 32'b00000000000000010000110100011110;
assign LUT_1[7509] = 32'b00000000000000001010000110011010;
assign LUT_1[7510] = 32'b00000000000000001100100010101111;
assign LUT_1[7511] = 32'b00000000000000000101110100101011;
assign LUT_1[7512] = 32'b00000000000000001000001000111100;
assign LUT_1[7513] = 32'b00000000000000000001011010111000;
assign LUT_1[7514] = 32'b00000000000000000011110111001101;
assign LUT_1[7515] = 32'b11111111111111111101001001001001;
assign LUT_1[7516] = 32'b00000000000000010000000010010011;
assign LUT_1[7517] = 32'b00000000000000001001010100001111;
assign LUT_1[7518] = 32'b00000000000000001011110000100100;
assign LUT_1[7519] = 32'b00000000000000000101000010100000;
assign LUT_1[7520] = 32'b00000000000000000111111010100100;
assign LUT_1[7521] = 32'b00000000000000000001001100100000;
assign LUT_1[7522] = 32'b00000000000000000011101000110101;
assign LUT_1[7523] = 32'b11111111111111111100111010110001;
assign LUT_1[7524] = 32'b00000000000000001111110011111011;
assign LUT_1[7525] = 32'b00000000000000001001000101110111;
assign LUT_1[7526] = 32'b00000000000000001011100010001100;
assign LUT_1[7527] = 32'b00000000000000000100110100001000;
assign LUT_1[7528] = 32'b00000000000000000111001000011001;
assign LUT_1[7529] = 32'b00000000000000000000011010010101;
assign LUT_1[7530] = 32'b00000000000000000010110110101010;
assign LUT_1[7531] = 32'b11111111111111111100001000100110;
assign LUT_1[7532] = 32'b00000000000000001111000001110000;
assign LUT_1[7533] = 32'b00000000000000001000010011101100;
assign LUT_1[7534] = 32'b00000000000000001010110000000001;
assign LUT_1[7535] = 32'b00000000000000000100000001111101;
assign LUT_1[7536] = 32'b00000000000000001001110110000110;
assign LUT_1[7537] = 32'b00000000000000000011001000000010;
assign LUT_1[7538] = 32'b00000000000000000101100100010111;
assign LUT_1[7539] = 32'b11111111111111111110110110010011;
assign LUT_1[7540] = 32'b00000000000000010001101111011101;
assign LUT_1[7541] = 32'b00000000000000001011000001011001;
assign LUT_1[7542] = 32'b00000000000000001101011101101110;
assign LUT_1[7543] = 32'b00000000000000000110101111101010;
assign LUT_1[7544] = 32'b00000000000000001001000011111011;
assign LUT_1[7545] = 32'b00000000000000000010010101110111;
assign LUT_1[7546] = 32'b00000000000000000100110010001100;
assign LUT_1[7547] = 32'b11111111111111111110000100001000;
assign LUT_1[7548] = 32'b00000000000000010000111101010010;
assign LUT_1[7549] = 32'b00000000000000001010001111001110;
assign LUT_1[7550] = 32'b00000000000000001100101011100011;
assign LUT_1[7551] = 32'b00000000000000000101111101011111;
assign LUT_1[7552] = 32'b00000000000000001000000010000000;
assign LUT_1[7553] = 32'b00000000000000000001010011111100;
assign LUT_1[7554] = 32'b00000000000000000011110000010001;
assign LUT_1[7555] = 32'b11111111111111111101000010001101;
assign LUT_1[7556] = 32'b00000000000000001111111011010111;
assign LUT_1[7557] = 32'b00000000000000001001001101010011;
assign LUT_1[7558] = 32'b00000000000000001011101001101000;
assign LUT_1[7559] = 32'b00000000000000000100111011100100;
assign LUT_1[7560] = 32'b00000000000000000111001111110101;
assign LUT_1[7561] = 32'b00000000000000000000100001110001;
assign LUT_1[7562] = 32'b00000000000000000010111110000110;
assign LUT_1[7563] = 32'b11111111111111111100010000000010;
assign LUT_1[7564] = 32'b00000000000000001111001001001100;
assign LUT_1[7565] = 32'b00000000000000001000011011001000;
assign LUT_1[7566] = 32'b00000000000000001010110111011101;
assign LUT_1[7567] = 32'b00000000000000000100001001011001;
assign LUT_1[7568] = 32'b00000000000000001001111101100010;
assign LUT_1[7569] = 32'b00000000000000000011001111011110;
assign LUT_1[7570] = 32'b00000000000000000101101011110011;
assign LUT_1[7571] = 32'b11111111111111111110111101101111;
assign LUT_1[7572] = 32'b00000000000000010001110110111001;
assign LUT_1[7573] = 32'b00000000000000001011001000110101;
assign LUT_1[7574] = 32'b00000000000000001101100101001010;
assign LUT_1[7575] = 32'b00000000000000000110110111000110;
assign LUT_1[7576] = 32'b00000000000000001001001011010111;
assign LUT_1[7577] = 32'b00000000000000000010011101010011;
assign LUT_1[7578] = 32'b00000000000000000100111001101000;
assign LUT_1[7579] = 32'b11111111111111111110001011100100;
assign LUT_1[7580] = 32'b00000000000000010001000100101110;
assign LUT_1[7581] = 32'b00000000000000001010010110101010;
assign LUT_1[7582] = 32'b00000000000000001100110010111111;
assign LUT_1[7583] = 32'b00000000000000000110000100111011;
assign LUT_1[7584] = 32'b00000000000000001000111100111111;
assign LUT_1[7585] = 32'b00000000000000000010001110111011;
assign LUT_1[7586] = 32'b00000000000000000100101011010000;
assign LUT_1[7587] = 32'b11111111111111111101111101001100;
assign LUT_1[7588] = 32'b00000000000000010000110110010110;
assign LUT_1[7589] = 32'b00000000000000001010001000010010;
assign LUT_1[7590] = 32'b00000000000000001100100100100111;
assign LUT_1[7591] = 32'b00000000000000000101110110100011;
assign LUT_1[7592] = 32'b00000000000000001000001010110100;
assign LUT_1[7593] = 32'b00000000000000000001011100110000;
assign LUT_1[7594] = 32'b00000000000000000011111001000101;
assign LUT_1[7595] = 32'b11111111111111111101001011000001;
assign LUT_1[7596] = 32'b00000000000000010000000100001011;
assign LUT_1[7597] = 32'b00000000000000001001010110000111;
assign LUT_1[7598] = 32'b00000000000000001011110010011100;
assign LUT_1[7599] = 32'b00000000000000000101000100011000;
assign LUT_1[7600] = 32'b00000000000000001010111000100001;
assign LUT_1[7601] = 32'b00000000000000000100001010011101;
assign LUT_1[7602] = 32'b00000000000000000110100110110010;
assign LUT_1[7603] = 32'b11111111111111111111111000101110;
assign LUT_1[7604] = 32'b00000000000000010010110001111000;
assign LUT_1[7605] = 32'b00000000000000001100000011110100;
assign LUT_1[7606] = 32'b00000000000000001110100000001001;
assign LUT_1[7607] = 32'b00000000000000000111110010000101;
assign LUT_1[7608] = 32'b00000000000000001010000110010110;
assign LUT_1[7609] = 32'b00000000000000000011011000010010;
assign LUT_1[7610] = 32'b00000000000000000101110100100111;
assign LUT_1[7611] = 32'b11111111111111111111000110100011;
assign LUT_1[7612] = 32'b00000000000000010001111111101101;
assign LUT_1[7613] = 32'b00000000000000001011010001101001;
assign LUT_1[7614] = 32'b00000000000000001101101101111110;
assign LUT_1[7615] = 32'b00000000000000000110111111111010;
assign LUT_1[7616] = 32'b00000000000000001001111111101000;
assign LUT_1[7617] = 32'b00000000000000000011010001100100;
assign LUT_1[7618] = 32'b00000000000000000101101101111001;
assign LUT_1[7619] = 32'b11111111111111111110111111110101;
assign LUT_1[7620] = 32'b00000000000000010001111000111111;
assign LUT_1[7621] = 32'b00000000000000001011001010111011;
assign LUT_1[7622] = 32'b00000000000000001101100111010000;
assign LUT_1[7623] = 32'b00000000000000000110111001001100;
assign LUT_1[7624] = 32'b00000000000000001001001101011101;
assign LUT_1[7625] = 32'b00000000000000000010011111011001;
assign LUT_1[7626] = 32'b00000000000000000100111011101110;
assign LUT_1[7627] = 32'b11111111111111111110001101101010;
assign LUT_1[7628] = 32'b00000000000000010001000110110100;
assign LUT_1[7629] = 32'b00000000000000001010011000110000;
assign LUT_1[7630] = 32'b00000000000000001100110101000101;
assign LUT_1[7631] = 32'b00000000000000000110000111000001;
assign LUT_1[7632] = 32'b00000000000000001011111011001010;
assign LUT_1[7633] = 32'b00000000000000000101001101000110;
assign LUT_1[7634] = 32'b00000000000000000111101001011011;
assign LUT_1[7635] = 32'b00000000000000000000111011010111;
assign LUT_1[7636] = 32'b00000000000000010011110100100001;
assign LUT_1[7637] = 32'b00000000000000001101000110011101;
assign LUT_1[7638] = 32'b00000000000000001111100010110010;
assign LUT_1[7639] = 32'b00000000000000001000110100101110;
assign LUT_1[7640] = 32'b00000000000000001011001000111111;
assign LUT_1[7641] = 32'b00000000000000000100011010111011;
assign LUT_1[7642] = 32'b00000000000000000110110111010000;
assign LUT_1[7643] = 32'b00000000000000000000001001001100;
assign LUT_1[7644] = 32'b00000000000000010011000010010110;
assign LUT_1[7645] = 32'b00000000000000001100010100010010;
assign LUT_1[7646] = 32'b00000000000000001110110000100111;
assign LUT_1[7647] = 32'b00000000000000001000000010100011;
assign LUT_1[7648] = 32'b00000000000000001010111010100111;
assign LUT_1[7649] = 32'b00000000000000000100001100100011;
assign LUT_1[7650] = 32'b00000000000000000110101000111000;
assign LUT_1[7651] = 32'b11111111111111111111111010110100;
assign LUT_1[7652] = 32'b00000000000000010010110011111110;
assign LUT_1[7653] = 32'b00000000000000001100000101111010;
assign LUT_1[7654] = 32'b00000000000000001110100010001111;
assign LUT_1[7655] = 32'b00000000000000000111110100001011;
assign LUT_1[7656] = 32'b00000000000000001010001000011100;
assign LUT_1[7657] = 32'b00000000000000000011011010011000;
assign LUT_1[7658] = 32'b00000000000000000101110110101101;
assign LUT_1[7659] = 32'b11111111111111111111001000101001;
assign LUT_1[7660] = 32'b00000000000000010010000001110011;
assign LUT_1[7661] = 32'b00000000000000001011010011101111;
assign LUT_1[7662] = 32'b00000000000000001101110000000100;
assign LUT_1[7663] = 32'b00000000000000000111000010000000;
assign LUT_1[7664] = 32'b00000000000000001100110110001001;
assign LUT_1[7665] = 32'b00000000000000000110001000000101;
assign LUT_1[7666] = 32'b00000000000000001000100100011010;
assign LUT_1[7667] = 32'b00000000000000000001110110010110;
assign LUT_1[7668] = 32'b00000000000000010100101111100000;
assign LUT_1[7669] = 32'b00000000000000001110000001011100;
assign LUT_1[7670] = 32'b00000000000000010000011101110001;
assign LUT_1[7671] = 32'b00000000000000001001101111101101;
assign LUT_1[7672] = 32'b00000000000000001100000011111110;
assign LUT_1[7673] = 32'b00000000000000000101010101111010;
assign LUT_1[7674] = 32'b00000000000000000111110010001111;
assign LUT_1[7675] = 32'b00000000000000000001000100001011;
assign LUT_1[7676] = 32'b00000000000000010011111101010101;
assign LUT_1[7677] = 32'b00000000000000001101001111010001;
assign LUT_1[7678] = 32'b00000000000000001111101011100110;
assign LUT_1[7679] = 32'b00000000000000001000111101100010;
assign LUT_1[7680] = 32'b00000000000000000000111100001110;
assign LUT_1[7681] = 32'b11111111111111111010001110001010;
assign LUT_1[7682] = 32'b11111111111111111100101010011111;
assign LUT_1[7683] = 32'b11111111111111110101111100011011;
assign LUT_1[7684] = 32'b00000000000000001000110101100101;
assign LUT_1[7685] = 32'b00000000000000000010000111100001;
assign LUT_1[7686] = 32'b00000000000000000100100011110110;
assign LUT_1[7687] = 32'b11111111111111111101110101110010;
assign LUT_1[7688] = 32'b00000000000000000000001010000011;
assign LUT_1[7689] = 32'b11111111111111111001011011111111;
assign LUT_1[7690] = 32'b11111111111111111011111000010100;
assign LUT_1[7691] = 32'b11111111111111110101001010010000;
assign LUT_1[7692] = 32'b00000000000000001000000011011010;
assign LUT_1[7693] = 32'b00000000000000000001010101010110;
assign LUT_1[7694] = 32'b00000000000000000011110001101011;
assign LUT_1[7695] = 32'b11111111111111111101000011100111;
assign LUT_1[7696] = 32'b00000000000000000010110111110000;
assign LUT_1[7697] = 32'b11111111111111111100001001101100;
assign LUT_1[7698] = 32'b11111111111111111110100110000001;
assign LUT_1[7699] = 32'b11111111111111110111110111111101;
assign LUT_1[7700] = 32'b00000000000000001010110001000111;
assign LUT_1[7701] = 32'b00000000000000000100000011000011;
assign LUT_1[7702] = 32'b00000000000000000110011111011000;
assign LUT_1[7703] = 32'b11111111111111111111110001010100;
assign LUT_1[7704] = 32'b00000000000000000010000101100101;
assign LUT_1[7705] = 32'b11111111111111111011010111100001;
assign LUT_1[7706] = 32'b11111111111111111101110011110110;
assign LUT_1[7707] = 32'b11111111111111110111000101110010;
assign LUT_1[7708] = 32'b00000000000000001001111110111100;
assign LUT_1[7709] = 32'b00000000000000000011010000111000;
assign LUT_1[7710] = 32'b00000000000000000101101101001101;
assign LUT_1[7711] = 32'b11111111111111111110111111001001;
assign LUT_1[7712] = 32'b00000000000000000001110111001101;
assign LUT_1[7713] = 32'b11111111111111111011001001001001;
assign LUT_1[7714] = 32'b11111111111111111101100101011110;
assign LUT_1[7715] = 32'b11111111111111110110110111011010;
assign LUT_1[7716] = 32'b00000000000000001001110000100100;
assign LUT_1[7717] = 32'b00000000000000000011000010100000;
assign LUT_1[7718] = 32'b00000000000000000101011110110101;
assign LUT_1[7719] = 32'b11111111111111111110110000110001;
assign LUT_1[7720] = 32'b00000000000000000001000101000010;
assign LUT_1[7721] = 32'b11111111111111111010010110111110;
assign LUT_1[7722] = 32'b11111111111111111100110011010011;
assign LUT_1[7723] = 32'b11111111111111110110000101001111;
assign LUT_1[7724] = 32'b00000000000000001000111110011001;
assign LUT_1[7725] = 32'b00000000000000000010010000010101;
assign LUT_1[7726] = 32'b00000000000000000100101100101010;
assign LUT_1[7727] = 32'b11111111111111111101111110100110;
assign LUT_1[7728] = 32'b00000000000000000011110010101111;
assign LUT_1[7729] = 32'b11111111111111111101000100101011;
assign LUT_1[7730] = 32'b11111111111111111111100001000000;
assign LUT_1[7731] = 32'b11111111111111111000110010111100;
assign LUT_1[7732] = 32'b00000000000000001011101100000110;
assign LUT_1[7733] = 32'b00000000000000000100111110000010;
assign LUT_1[7734] = 32'b00000000000000000111011010010111;
assign LUT_1[7735] = 32'b00000000000000000000101100010011;
assign LUT_1[7736] = 32'b00000000000000000011000000100100;
assign LUT_1[7737] = 32'b11111111111111111100010010100000;
assign LUT_1[7738] = 32'b11111111111111111110101110110101;
assign LUT_1[7739] = 32'b11111111111111111000000000110001;
assign LUT_1[7740] = 32'b00000000000000001010111001111011;
assign LUT_1[7741] = 32'b00000000000000000100001011110111;
assign LUT_1[7742] = 32'b00000000000000000110101000001100;
assign LUT_1[7743] = 32'b11111111111111111111111010001000;
assign LUT_1[7744] = 32'b00000000000000000010111001110110;
assign LUT_1[7745] = 32'b11111111111111111100001011110010;
assign LUT_1[7746] = 32'b11111111111111111110101000000111;
assign LUT_1[7747] = 32'b11111111111111110111111010000011;
assign LUT_1[7748] = 32'b00000000000000001010110011001101;
assign LUT_1[7749] = 32'b00000000000000000100000101001001;
assign LUT_1[7750] = 32'b00000000000000000110100001011110;
assign LUT_1[7751] = 32'b11111111111111111111110011011010;
assign LUT_1[7752] = 32'b00000000000000000010000111101011;
assign LUT_1[7753] = 32'b11111111111111111011011001100111;
assign LUT_1[7754] = 32'b11111111111111111101110101111100;
assign LUT_1[7755] = 32'b11111111111111110111000111111000;
assign LUT_1[7756] = 32'b00000000000000001010000001000010;
assign LUT_1[7757] = 32'b00000000000000000011010010111110;
assign LUT_1[7758] = 32'b00000000000000000101101111010011;
assign LUT_1[7759] = 32'b11111111111111111111000001001111;
assign LUT_1[7760] = 32'b00000000000000000100110101011000;
assign LUT_1[7761] = 32'b11111111111111111110000111010100;
assign LUT_1[7762] = 32'b00000000000000000000100011101001;
assign LUT_1[7763] = 32'b11111111111111111001110101100101;
assign LUT_1[7764] = 32'b00000000000000001100101110101111;
assign LUT_1[7765] = 32'b00000000000000000110000000101011;
assign LUT_1[7766] = 32'b00000000000000001000011101000000;
assign LUT_1[7767] = 32'b00000000000000000001101110111100;
assign LUT_1[7768] = 32'b00000000000000000100000011001101;
assign LUT_1[7769] = 32'b11111111111111111101010101001001;
assign LUT_1[7770] = 32'b11111111111111111111110001011110;
assign LUT_1[7771] = 32'b11111111111111111001000011011010;
assign LUT_1[7772] = 32'b00000000000000001011111100100100;
assign LUT_1[7773] = 32'b00000000000000000101001110100000;
assign LUT_1[7774] = 32'b00000000000000000111101010110101;
assign LUT_1[7775] = 32'b00000000000000000000111100110001;
assign LUT_1[7776] = 32'b00000000000000000011110100110101;
assign LUT_1[7777] = 32'b11111111111111111101000110110001;
assign LUT_1[7778] = 32'b11111111111111111111100011000110;
assign LUT_1[7779] = 32'b11111111111111111000110101000010;
assign LUT_1[7780] = 32'b00000000000000001011101110001100;
assign LUT_1[7781] = 32'b00000000000000000101000000001000;
assign LUT_1[7782] = 32'b00000000000000000111011100011101;
assign LUT_1[7783] = 32'b00000000000000000000101110011001;
assign LUT_1[7784] = 32'b00000000000000000011000010101010;
assign LUT_1[7785] = 32'b11111111111111111100010100100110;
assign LUT_1[7786] = 32'b11111111111111111110110000111011;
assign LUT_1[7787] = 32'b11111111111111111000000010110111;
assign LUT_1[7788] = 32'b00000000000000001010111100000001;
assign LUT_1[7789] = 32'b00000000000000000100001101111101;
assign LUT_1[7790] = 32'b00000000000000000110101010010010;
assign LUT_1[7791] = 32'b11111111111111111111111100001110;
assign LUT_1[7792] = 32'b00000000000000000101110000010111;
assign LUT_1[7793] = 32'b11111111111111111111000010010011;
assign LUT_1[7794] = 32'b00000000000000000001011110101000;
assign LUT_1[7795] = 32'b11111111111111111010110000100100;
assign LUT_1[7796] = 32'b00000000000000001101101001101110;
assign LUT_1[7797] = 32'b00000000000000000110111011101010;
assign LUT_1[7798] = 32'b00000000000000001001010111111111;
assign LUT_1[7799] = 32'b00000000000000000010101001111011;
assign LUT_1[7800] = 32'b00000000000000000100111110001100;
assign LUT_1[7801] = 32'b11111111111111111110010000001000;
assign LUT_1[7802] = 32'b00000000000000000000101100011101;
assign LUT_1[7803] = 32'b11111111111111111001111110011001;
assign LUT_1[7804] = 32'b00000000000000001100110111100011;
assign LUT_1[7805] = 32'b00000000000000000110001001011111;
assign LUT_1[7806] = 32'b00000000000000001000100101110100;
assign LUT_1[7807] = 32'b00000000000000000001110111110000;
assign LUT_1[7808] = 32'b00000000000000000011111100010001;
assign LUT_1[7809] = 32'b11111111111111111101001110001101;
assign LUT_1[7810] = 32'b11111111111111111111101010100010;
assign LUT_1[7811] = 32'b11111111111111111000111100011110;
assign LUT_1[7812] = 32'b00000000000000001011110101101000;
assign LUT_1[7813] = 32'b00000000000000000101000111100100;
assign LUT_1[7814] = 32'b00000000000000000111100011111001;
assign LUT_1[7815] = 32'b00000000000000000000110101110101;
assign LUT_1[7816] = 32'b00000000000000000011001010000110;
assign LUT_1[7817] = 32'b11111111111111111100011100000010;
assign LUT_1[7818] = 32'b11111111111111111110111000010111;
assign LUT_1[7819] = 32'b11111111111111111000001010010011;
assign LUT_1[7820] = 32'b00000000000000001011000011011101;
assign LUT_1[7821] = 32'b00000000000000000100010101011001;
assign LUT_1[7822] = 32'b00000000000000000110110001101110;
assign LUT_1[7823] = 32'b00000000000000000000000011101010;
assign LUT_1[7824] = 32'b00000000000000000101110111110011;
assign LUT_1[7825] = 32'b11111111111111111111001001101111;
assign LUT_1[7826] = 32'b00000000000000000001100110000100;
assign LUT_1[7827] = 32'b11111111111111111010111000000000;
assign LUT_1[7828] = 32'b00000000000000001101110001001010;
assign LUT_1[7829] = 32'b00000000000000000111000011000110;
assign LUT_1[7830] = 32'b00000000000000001001011111011011;
assign LUT_1[7831] = 32'b00000000000000000010110001010111;
assign LUT_1[7832] = 32'b00000000000000000101000101101000;
assign LUT_1[7833] = 32'b11111111111111111110010111100100;
assign LUT_1[7834] = 32'b00000000000000000000110011111001;
assign LUT_1[7835] = 32'b11111111111111111010000101110101;
assign LUT_1[7836] = 32'b00000000000000001100111110111111;
assign LUT_1[7837] = 32'b00000000000000000110010000111011;
assign LUT_1[7838] = 32'b00000000000000001000101101010000;
assign LUT_1[7839] = 32'b00000000000000000001111111001100;
assign LUT_1[7840] = 32'b00000000000000000100110111010000;
assign LUT_1[7841] = 32'b11111111111111111110001001001100;
assign LUT_1[7842] = 32'b00000000000000000000100101100001;
assign LUT_1[7843] = 32'b11111111111111111001110111011101;
assign LUT_1[7844] = 32'b00000000000000001100110000100111;
assign LUT_1[7845] = 32'b00000000000000000110000010100011;
assign LUT_1[7846] = 32'b00000000000000001000011110111000;
assign LUT_1[7847] = 32'b00000000000000000001110000110100;
assign LUT_1[7848] = 32'b00000000000000000100000101000101;
assign LUT_1[7849] = 32'b11111111111111111101010111000001;
assign LUT_1[7850] = 32'b11111111111111111111110011010110;
assign LUT_1[7851] = 32'b11111111111111111001000101010010;
assign LUT_1[7852] = 32'b00000000000000001011111110011100;
assign LUT_1[7853] = 32'b00000000000000000101010000011000;
assign LUT_1[7854] = 32'b00000000000000000111101100101101;
assign LUT_1[7855] = 32'b00000000000000000000111110101001;
assign LUT_1[7856] = 32'b00000000000000000110110010110010;
assign LUT_1[7857] = 32'b00000000000000000000000100101110;
assign LUT_1[7858] = 32'b00000000000000000010100001000011;
assign LUT_1[7859] = 32'b11111111111111111011110010111111;
assign LUT_1[7860] = 32'b00000000000000001110101100001001;
assign LUT_1[7861] = 32'b00000000000000000111111110000101;
assign LUT_1[7862] = 32'b00000000000000001010011010011010;
assign LUT_1[7863] = 32'b00000000000000000011101100010110;
assign LUT_1[7864] = 32'b00000000000000000110000000100111;
assign LUT_1[7865] = 32'b11111111111111111111010010100011;
assign LUT_1[7866] = 32'b00000000000000000001101110111000;
assign LUT_1[7867] = 32'b11111111111111111011000000110100;
assign LUT_1[7868] = 32'b00000000000000001101111001111110;
assign LUT_1[7869] = 32'b00000000000000000111001011111010;
assign LUT_1[7870] = 32'b00000000000000001001101000001111;
assign LUT_1[7871] = 32'b00000000000000000010111010001011;
assign LUT_1[7872] = 32'b00000000000000000101111001111001;
assign LUT_1[7873] = 32'b11111111111111111111001011110101;
assign LUT_1[7874] = 32'b00000000000000000001101000001010;
assign LUT_1[7875] = 32'b11111111111111111010111010000110;
assign LUT_1[7876] = 32'b00000000000000001101110011010000;
assign LUT_1[7877] = 32'b00000000000000000111000101001100;
assign LUT_1[7878] = 32'b00000000000000001001100001100001;
assign LUT_1[7879] = 32'b00000000000000000010110011011101;
assign LUT_1[7880] = 32'b00000000000000000101000111101110;
assign LUT_1[7881] = 32'b11111111111111111110011001101010;
assign LUT_1[7882] = 32'b00000000000000000000110101111111;
assign LUT_1[7883] = 32'b11111111111111111010000111111011;
assign LUT_1[7884] = 32'b00000000000000001101000001000101;
assign LUT_1[7885] = 32'b00000000000000000110010011000001;
assign LUT_1[7886] = 32'b00000000000000001000101111010110;
assign LUT_1[7887] = 32'b00000000000000000010000001010010;
assign LUT_1[7888] = 32'b00000000000000000111110101011011;
assign LUT_1[7889] = 32'b00000000000000000001000111010111;
assign LUT_1[7890] = 32'b00000000000000000011100011101100;
assign LUT_1[7891] = 32'b11111111111111111100110101101000;
assign LUT_1[7892] = 32'b00000000000000001111101110110010;
assign LUT_1[7893] = 32'b00000000000000001001000000101110;
assign LUT_1[7894] = 32'b00000000000000001011011101000011;
assign LUT_1[7895] = 32'b00000000000000000100101110111111;
assign LUT_1[7896] = 32'b00000000000000000111000011010000;
assign LUT_1[7897] = 32'b00000000000000000000010101001100;
assign LUT_1[7898] = 32'b00000000000000000010110001100001;
assign LUT_1[7899] = 32'b11111111111111111100000011011101;
assign LUT_1[7900] = 32'b00000000000000001110111100100111;
assign LUT_1[7901] = 32'b00000000000000001000001110100011;
assign LUT_1[7902] = 32'b00000000000000001010101010111000;
assign LUT_1[7903] = 32'b00000000000000000011111100110100;
assign LUT_1[7904] = 32'b00000000000000000110110100111000;
assign LUT_1[7905] = 32'b00000000000000000000000110110100;
assign LUT_1[7906] = 32'b00000000000000000010100011001001;
assign LUT_1[7907] = 32'b11111111111111111011110101000101;
assign LUT_1[7908] = 32'b00000000000000001110101110001111;
assign LUT_1[7909] = 32'b00000000000000001000000000001011;
assign LUT_1[7910] = 32'b00000000000000001010011100100000;
assign LUT_1[7911] = 32'b00000000000000000011101110011100;
assign LUT_1[7912] = 32'b00000000000000000110000010101101;
assign LUT_1[7913] = 32'b11111111111111111111010100101001;
assign LUT_1[7914] = 32'b00000000000000000001110000111110;
assign LUT_1[7915] = 32'b11111111111111111011000010111010;
assign LUT_1[7916] = 32'b00000000000000001101111100000100;
assign LUT_1[7917] = 32'b00000000000000000111001110000000;
assign LUT_1[7918] = 32'b00000000000000001001101010010101;
assign LUT_1[7919] = 32'b00000000000000000010111100010001;
assign LUT_1[7920] = 32'b00000000000000001000110000011010;
assign LUT_1[7921] = 32'b00000000000000000010000010010110;
assign LUT_1[7922] = 32'b00000000000000000100011110101011;
assign LUT_1[7923] = 32'b11111111111111111101110000100111;
assign LUT_1[7924] = 32'b00000000000000010000101001110001;
assign LUT_1[7925] = 32'b00000000000000001001111011101101;
assign LUT_1[7926] = 32'b00000000000000001100011000000010;
assign LUT_1[7927] = 32'b00000000000000000101101001111110;
assign LUT_1[7928] = 32'b00000000000000000111111110001111;
assign LUT_1[7929] = 32'b00000000000000000001010000001011;
assign LUT_1[7930] = 32'b00000000000000000011101100100000;
assign LUT_1[7931] = 32'b11111111111111111100111110011100;
assign LUT_1[7932] = 32'b00000000000000001111110111100110;
assign LUT_1[7933] = 32'b00000000000000001001001001100010;
assign LUT_1[7934] = 32'b00000000000000001011100101110111;
assign LUT_1[7935] = 32'b00000000000000000100110111110011;
assign LUT_1[7936] = 32'b11111111111111111110110000011010;
assign LUT_1[7937] = 32'b11111111111111111000000010010110;
assign LUT_1[7938] = 32'b11111111111111111010011110101011;
assign LUT_1[7939] = 32'b11111111111111110011110000100111;
assign LUT_1[7940] = 32'b00000000000000000110101001110001;
assign LUT_1[7941] = 32'b11111111111111111111111011101101;
assign LUT_1[7942] = 32'b00000000000000000010011000000010;
assign LUT_1[7943] = 32'b11111111111111111011101001111110;
assign LUT_1[7944] = 32'b11111111111111111101111110001111;
assign LUT_1[7945] = 32'b11111111111111110111010000001011;
assign LUT_1[7946] = 32'b11111111111111111001101100100000;
assign LUT_1[7947] = 32'b11111111111111110010111110011100;
assign LUT_1[7948] = 32'b00000000000000000101110111100110;
assign LUT_1[7949] = 32'b11111111111111111111001001100010;
assign LUT_1[7950] = 32'b00000000000000000001100101110111;
assign LUT_1[7951] = 32'b11111111111111111010110111110011;
assign LUT_1[7952] = 32'b00000000000000000000101011111100;
assign LUT_1[7953] = 32'b11111111111111111001111101111000;
assign LUT_1[7954] = 32'b11111111111111111100011010001101;
assign LUT_1[7955] = 32'b11111111111111110101101100001001;
assign LUT_1[7956] = 32'b00000000000000001000100101010011;
assign LUT_1[7957] = 32'b00000000000000000001110111001111;
assign LUT_1[7958] = 32'b00000000000000000100010011100100;
assign LUT_1[7959] = 32'b11111111111111111101100101100000;
assign LUT_1[7960] = 32'b11111111111111111111111001110001;
assign LUT_1[7961] = 32'b11111111111111111001001011101101;
assign LUT_1[7962] = 32'b11111111111111111011101000000010;
assign LUT_1[7963] = 32'b11111111111111110100111001111110;
assign LUT_1[7964] = 32'b00000000000000000111110011001000;
assign LUT_1[7965] = 32'b00000000000000000001000101000100;
assign LUT_1[7966] = 32'b00000000000000000011100001011001;
assign LUT_1[7967] = 32'b11111111111111111100110011010101;
assign LUT_1[7968] = 32'b11111111111111111111101011011001;
assign LUT_1[7969] = 32'b11111111111111111000111101010101;
assign LUT_1[7970] = 32'b11111111111111111011011001101010;
assign LUT_1[7971] = 32'b11111111111111110100101011100110;
assign LUT_1[7972] = 32'b00000000000000000111100100110000;
assign LUT_1[7973] = 32'b00000000000000000000110110101100;
assign LUT_1[7974] = 32'b00000000000000000011010011000001;
assign LUT_1[7975] = 32'b11111111111111111100100100111101;
assign LUT_1[7976] = 32'b11111111111111111110111001001110;
assign LUT_1[7977] = 32'b11111111111111111000001011001010;
assign LUT_1[7978] = 32'b11111111111111111010100111011111;
assign LUT_1[7979] = 32'b11111111111111110011111001011011;
assign LUT_1[7980] = 32'b00000000000000000110110010100101;
assign LUT_1[7981] = 32'b00000000000000000000000100100001;
assign LUT_1[7982] = 32'b00000000000000000010100000110110;
assign LUT_1[7983] = 32'b11111111111111111011110010110010;
assign LUT_1[7984] = 32'b00000000000000000001100110111011;
assign LUT_1[7985] = 32'b11111111111111111010111000110111;
assign LUT_1[7986] = 32'b11111111111111111101010101001100;
assign LUT_1[7987] = 32'b11111111111111110110100111001000;
assign LUT_1[7988] = 32'b00000000000000001001100000010010;
assign LUT_1[7989] = 32'b00000000000000000010110010001110;
assign LUT_1[7990] = 32'b00000000000000000101001110100011;
assign LUT_1[7991] = 32'b11111111111111111110100000011111;
assign LUT_1[7992] = 32'b00000000000000000000110100110000;
assign LUT_1[7993] = 32'b11111111111111111010000110101100;
assign LUT_1[7994] = 32'b11111111111111111100100011000001;
assign LUT_1[7995] = 32'b11111111111111110101110100111101;
assign LUT_1[7996] = 32'b00000000000000001000101110000111;
assign LUT_1[7997] = 32'b00000000000000000010000000000011;
assign LUT_1[7998] = 32'b00000000000000000100011100011000;
assign LUT_1[7999] = 32'b11111111111111111101101110010100;
assign LUT_1[8000] = 32'b00000000000000000000101110000010;
assign LUT_1[8001] = 32'b11111111111111111001111111111110;
assign LUT_1[8002] = 32'b11111111111111111100011100010011;
assign LUT_1[8003] = 32'b11111111111111110101101110001111;
assign LUT_1[8004] = 32'b00000000000000001000100111011001;
assign LUT_1[8005] = 32'b00000000000000000001111001010101;
assign LUT_1[8006] = 32'b00000000000000000100010101101010;
assign LUT_1[8007] = 32'b11111111111111111101100111100110;
assign LUT_1[8008] = 32'b11111111111111111111111011110111;
assign LUT_1[8009] = 32'b11111111111111111001001101110011;
assign LUT_1[8010] = 32'b11111111111111111011101010001000;
assign LUT_1[8011] = 32'b11111111111111110100111100000100;
assign LUT_1[8012] = 32'b00000000000000000111110101001110;
assign LUT_1[8013] = 32'b00000000000000000001000111001010;
assign LUT_1[8014] = 32'b00000000000000000011100011011111;
assign LUT_1[8015] = 32'b11111111111111111100110101011011;
assign LUT_1[8016] = 32'b00000000000000000010101001100100;
assign LUT_1[8017] = 32'b11111111111111111011111011100000;
assign LUT_1[8018] = 32'b11111111111111111110010111110101;
assign LUT_1[8019] = 32'b11111111111111110111101001110001;
assign LUT_1[8020] = 32'b00000000000000001010100010111011;
assign LUT_1[8021] = 32'b00000000000000000011110100110111;
assign LUT_1[8022] = 32'b00000000000000000110010001001100;
assign LUT_1[8023] = 32'b11111111111111111111100011001000;
assign LUT_1[8024] = 32'b00000000000000000001110111011001;
assign LUT_1[8025] = 32'b11111111111111111011001001010101;
assign LUT_1[8026] = 32'b11111111111111111101100101101010;
assign LUT_1[8027] = 32'b11111111111111110110110111100110;
assign LUT_1[8028] = 32'b00000000000000001001110000110000;
assign LUT_1[8029] = 32'b00000000000000000011000010101100;
assign LUT_1[8030] = 32'b00000000000000000101011111000001;
assign LUT_1[8031] = 32'b11111111111111111110110000111101;
assign LUT_1[8032] = 32'b00000000000000000001101001000001;
assign LUT_1[8033] = 32'b11111111111111111010111010111101;
assign LUT_1[8034] = 32'b11111111111111111101010111010010;
assign LUT_1[8035] = 32'b11111111111111110110101001001110;
assign LUT_1[8036] = 32'b00000000000000001001100010011000;
assign LUT_1[8037] = 32'b00000000000000000010110100010100;
assign LUT_1[8038] = 32'b00000000000000000101010000101001;
assign LUT_1[8039] = 32'b11111111111111111110100010100101;
assign LUT_1[8040] = 32'b00000000000000000000110110110110;
assign LUT_1[8041] = 32'b11111111111111111010001000110010;
assign LUT_1[8042] = 32'b11111111111111111100100101000111;
assign LUT_1[8043] = 32'b11111111111111110101110111000011;
assign LUT_1[8044] = 32'b00000000000000001000110000001101;
assign LUT_1[8045] = 32'b00000000000000000010000010001001;
assign LUT_1[8046] = 32'b00000000000000000100011110011110;
assign LUT_1[8047] = 32'b11111111111111111101110000011010;
assign LUT_1[8048] = 32'b00000000000000000011100100100011;
assign LUT_1[8049] = 32'b11111111111111111100110110011111;
assign LUT_1[8050] = 32'b11111111111111111111010010110100;
assign LUT_1[8051] = 32'b11111111111111111000100100110000;
assign LUT_1[8052] = 32'b00000000000000001011011101111010;
assign LUT_1[8053] = 32'b00000000000000000100101111110110;
assign LUT_1[8054] = 32'b00000000000000000111001100001011;
assign LUT_1[8055] = 32'b00000000000000000000011110000111;
assign LUT_1[8056] = 32'b00000000000000000010110010011000;
assign LUT_1[8057] = 32'b11111111111111111100000100010100;
assign LUT_1[8058] = 32'b11111111111111111110100000101001;
assign LUT_1[8059] = 32'b11111111111111110111110010100101;
assign LUT_1[8060] = 32'b00000000000000001010101011101111;
assign LUT_1[8061] = 32'b00000000000000000011111101101011;
assign LUT_1[8062] = 32'b00000000000000000110011010000000;
assign LUT_1[8063] = 32'b11111111111111111111101011111100;
assign LUT_1[8064] = 32'b00000000000000000001110000011101;
assign LUT_1[8065] = 32'b11111111111111111011000010011001;
assign LUT_1[8066] = 32'b11111111111111111101011110101110;
assign LUT_1[8067] = 32'b11111111111111110110110000101010;
assign LUT_1[8068] = 32'b00000000000000001001101001110100;
assign LUT_1[8069] = 32'b00000000000000000010111011110000;
assign LUT_1[8070] = 32'b00000000000000000101011000000101;
assign LUT_1[8071] = 32'b11111111111111111110101010000001;
assign LUT_1[8072] = 32'b00000000000000000000111110010010;
assign LUT_1[8073] = 32'b11111111111111111010010000001110;
assign LUT_1[8074] = 32'b11111111111111111100101100100011;
assign LUT_1[8075] = 32'b11111111111111110101111110011111;
assign LUT_1[8076] = 32'b00000000000000001000110111101001;
assign LUT_1[8077] = 32'b00000000000000000010001001100101;
assign LUT_1[8078] = 32'b00000000000000000100100101111010;
assign LUT_1[8079] = 32'b11111111111111111101110111110110;
assign LUT_1[8080] = 32'b00000000000000000011101011111111;
assign LUT_1[8081] = 32'b11111111111111111100111101111011;
assign LUT_1[8082] = 32'b11111111111111111111011010010000;
assign LUT_1[8083] = 32'b11111111111111111000101100001100;
assign LUT_1[8084] = 32'b00000000000000001011100101010110;
assign LUT_1[8085] = 32'b00000000000000000100110111010010;
assign LUT_1[8086] = 32'b00000000000000000111010011100111;
assign LUT_1[8087] = 32'b00000000000000000000100101100011;
assign LUT_1[8088] = 32'b00000000000000000010111001110100;
assign LUT_1[8089] = 32'b11111111111111111100001011110000;
assign LUT_1[8090] = 32'b11111111111111111110101000000101;
assign LUT_1[8091] = 32'b11111111111111110111111010000001;
assign LUT_1[8092] = 32'b00000000000000001010110011001011;
assign LUT_1[8093] = 32'b00000000000000000100000101000111;
assign LUT_1[8094] = 32'b00000000000000000110100001011100;
assign LUT_1[8095] = 32'b11111111111111111111110011011000;
assign LUT_1[8096] = 32'b00000000000000000010101011011100;
assign LUT_1[8097] = 32'b11111111111111111011111101011000;
assign LUT_1[8098] = 32'b11111111111111111110011001101101;
assign LUT_1[8099] = 32'b11111111111111110111101011101001;
assign LUT_1[8100] = 32'b00000000000000001010100100110011;
assign LUT_1[8101] = 32'b00000000000000000011110110101111;
assign LUT_1[8102] = 32'b00000000000000000110010011000100;
assign LUT_1[8103] = 32'b11111111111111111111100101000000;
assign LUT_1[8104] = 32'b00000000000000000001111001010001;
assign LUT_1[8105] = 32'b11111111111111111011001011001101;
assign LUT_1[8106] = 32'b11111111111111111101100111100010;
assign LUT_1[8107] = 32'b11111111111111110110111001011110;
assign LUT_1[8108] = 32'b00000000000000001001110010101000;
assign LUT_1[8109] = 32'b00000000000000000011000100100100;
assign LUT_1[8110] = 32'b00000000000000000101100000111001;
assign LUT_1[8111] = 32'b11111111111111111110110010110101;
assign LUT_1[8112] = 32'b00000000000000000100100110111110;
assign LUT_1[8113] = 32'b11111111111111111101111000111010;
assign LUT_1[8114] = 32'b00000000000000000000010101001111;
assign LUT_1[8115] = 32'b11111111111111111001100111001011;
assign LUT_1[8116] = 32'b00000000000000001100100000010101;
assign LUT_1[8117] = 32'b00000000000000000101110010010001;
assign LUT_1[8118] = 32'b00000000000000001000001110100110;
assign LUT_1[8119] = 32'b00000000000000000001100000100010;
assign LUT_1[8120] = 32'b00000000000000000011110100110011;
assign LUT_1[8121] = 32'b11111111111111111101000110101111;
assign LUT_1[8122] = 32'b11111111111111111111100011000100;
assign LUT_1[8123] = 32'b11111111111111111000110101000000;
assign LUT_1[8124] = 32'b00000000000000001011101110001010;
assign LUT_1[8125] = 32'b00000000000000000101000000000110;
assign LUT_1[8126] = 32'b00000000000000000111011100011011;
assign LUT_1[8127] = 32'b00000000000000000000101110010111;
assign LUT_1[8128] = 32'b00000000000000000011101110000101;
assign LUT_1[8129] = 32'b11111111111111111101000000000001;
assign LUT_1[8130] = 32'b11111111111111111111011100010110;
assign LUT_1[8131] = 32'b11111111111111111000101110010010;
assign LUT_1[8132] = 32'b00000000000000001011100111011100;
assign LUT_1[8133] = 32'b00000000000000000100111001011000;
assign LUT_1[8134] = 32'b00000000000000000111010101101101;
assign LUT_1[8135] = 32'b00000000000000000000100111101001;
assign LUT_1[8136] = 32'b00000000000000000010111011111010;
assign LUT_1[8137] = 32'b11111111111111111100001101110110;
assign LUT_1[8138] = 32'b11111111111111111110101010001011;
assign LUT_1[8139] = 32'b11111111111111110111111100000111;
assign LUT_1[8140] = 32'b00000000000000001010110101010001;
assign LUT_1[8141] = 32'b00000000000000000100000111001101;
assign LUT_1[8142] = 32'b00000000000000000110100011100010;
assign LUT_1[8143] = 32'b11111111111111111111110101011110;
assign LUT_1[8144] = 32'b00000000000000000101101001100111;
assign LUT_1[8145] = 32'b11111111111111111110111011100011;
assign LUT_1[8146] = 32'b00000000000000000001010111111000;
assign LUT_1[8147] = 32'b11111111111111111010101001110100;
assign LUT_1[8148] = 32'b00000000000000001101100010111110;
assign LUT_1[8149] = 32'b00000000000000000110110100111010;
assign LUT_1[8150] = 32'b00000000000000001001010001001111;
assign LUT_1[8151] = 32'b00000000000000000010100011001011;
assign LUT_1[8152] = 32'b00000000000000000100110111011100;
assign LUT_1[8153] = 32'b11111111111111111110001001011000;
assign LUT_1[8154] = 32'b00000000000000000000100101101101;
assign LUT_1[8155] = 32'b11111111111111111001110111101001;
assign LUT_1[8156] = 32'b00000000000000001100110000110011;
assign LUT_1[8157] = 32'b00000000000000000110000010101111;
assign LUT_1[8158] = 32'b00000000000000001000011111000100;
assign LUT_1[8159] = 32'b00000000000000000001110001000000;
assign LUT_1[8160] = 32'b00000000000000000100101001000100;
assign LUT_1[8161] = 32'b11111111111111111101111011000000;
assign LUT_1[8162] = 32'b00000000000000000000010111010101;
assign LUT_1[8163] = 32'b11111111111111111001101001010001;
assign LUT_1[8164] = 32'b00000000000000001100100010011011;
assign LUT_1[8165] = 32'b00000000000000000101110100010111;
assign LUT_1[8166] = 32'b00000000000000001000010000101100;
assign LUT_1[8167] = 32'b00000000000000000001100010101000;
assign LUT_1[8168] = 32'b00000000000000000011110110111001;
assign LUT_1[8169] = 32'b11111111111111111101001000110101;
assign LUT_1[8170] = 32'b11111111111111111111100101001010;
assign LUT_1[8171] = 32'b11111111111111111000110111000110;
assign LUT_1[8172] = 32'b00000000000000001011110000010000;
assign LUT_1[8173] = 32'b00000000000000000101000010001100;
assign LUT_1[8174] = 32'b00000000000000000111011110100001;
assign LUT_1[8175] = 32'b00000000000000000000110000011101;
assign LUT_1[8176] = 32'b00000000000000000110100100100110;
assign LUT_1[8177] = 32'b11111111111111111111110110100010;
assign LUT_1[8178] = 32'b00000000000000000010010010110111;
assign LUT_1[8179] = 32'b11111111111111111011100100110011;
assign LUT_1[8180] = 32'b00000000000000001110011101111101;
assign LUT_1[8181] = 32'b00000000000000000111101111111001;
assign LUT_1[8182] = 32'b00000000000000001010001100001110;
assign LUT_1[8183] = 32'b00000000000000000011011110001010;
assign LUT_1[8184] = 32'b00000000000000000101110010011011;
assign LUT_1[8185] = 32'b11111111111111111111000100010111;
assign LUT_1[8186] = 32'b00000000000000000001100000101100;
assign LUT_1[8187] = 32'b11111111111111111010110010101000;
assign LUT_1[8188] = 32'b00000000000000001101101011110010;
assign LUT_1[8189] = 32'b00000000000000000110111101101110;
assign LUT_1[8190] = 32'b00000000000000001001011010000011;
assign LUT_1[8191] = 32'b00000000000000000010101011111111;
assign LUT_1[8192] = 32'b00000000000000000011001000100011;
assign LUT_1[8193] = 32'b11111111111111111100011010011111;
assign LUT_1[8194] = 32'b11111111111111111110110110110100;
assign LUT_1[8195] = 32'b11111111111111111000001000110000;
assign LUT_1[8196] = 32'b00000000000000001011000001111010;
assign LUT_1[8197] = 32'b00000000000000000100010011110110;
assign LUT_1[8198] = 32'b00000000000000000110110000001011;
assign LUT_1[8199] = 32'b00000000000000000000000010000111;
assign LUT_1[8200] = 32'b00000000000000000010010110011000;
assign LUT_1[8201] = 32'b11111111111111111011101000010100;
assign LUT_1[8202] = 32'b11111111111111111110000100101001;
assign LUT_1[8203] = 32'b11111111111111110111010110100101;
assign LUT_1[8204] = 32'b00000000000000001010001111101111;
assign LUT_1[8205] = 32'b00000000000000000011100001101011;
assign LUT_1[8206] = 32'b00000000000000000101111110000000;
assign LUT_1[8207] = 32'b11111111111111111111001111111100;
assign LUT_1[8208] = 32'b00000000000000000101000100000101;
assign LUT_1[8209] = 32'b11111111111111111110010110000001;
assign LUT_1[8210] = 32'b00000000000000000000110010010110;
assign LUT_1[8211] = 32'b11111111111111111010000100010010;
assign LUT_1[8212] = 32'b00000000000000001100111101011100;
assign LUT_1[8213] = 32'b00000000000000000110001111011000;
assign LUT_1[8214] = 32'b00000000000000001000101011101101;
assign LUT_1[8215] = 32'b00000000000000000001111101101001;
assign LUT_1[8216] = 32'b00000000000000000100010001111010;
assign LUT_1[8217] = 32'b11111111111111111101100011110110;
assign LUT_1[8218] = 32'b00000000000000000000000000001011;
assign LUT_1[8219] = 32'b11111111111111111001010010000111;
assign LUT_1[8220] = 32'b00000000000000001100001011010001;
assign LUT_1[8221] = 32'b00000000000000000101011101001101;
assign LUT_1[8222] = 32'b00000000000000000111111001100010;
assign LUT_1[8223] = 32'b00000000000000000001001011011110;
assign LUT_1[8224] = 32'b00000000000000000100000011100010;
assign LUT_1[8225] = 32'b11111111111111111101010101011110;
assign LUT_1[8226] = 32'b11111111111111111111110001110011;
assign LUT_1[8227] = 32'b11111111111111111001000011101111;
assign LUT_1[8228] = 32'b00000000000000001011111100111001;
assign LUT_1[8229] = 32'b00000000000000000101001110110101;
assign LUT_1[8230] = 32'b00000000000000000111101011001010;
assign LUT_1[8231] = 32'b00000000000000000000111101000110;
assign LUT_1[8232] = 32'b00000000000000000011010001010111;
assign LUT_1[8233] = 32'b11111111111111111100100011010011;
assign LUT_1[8234] = 32'b11111111111111111110111111101000;
assign LUT_1[8235] = 32'b11111111111111111000010001100100;
assign LUT_1[8236] = 32'b00000000000000001011001010101110;
assign LUT_1[8237] = 32'b00000000000000000100011100101010;
assign LUT_1[8238] = 32'b00000000000000000110111000111111;
assign LUT_1[8239] = 32'b00000000000000000000001010111011;
assign LUT_1[8240] = 32'b00000000000000000101111111000100;
assign LUT_1[8241] = 32'b11111111111111111111010001000000;
assign LUT_1[8242] = 32'b00000000000000000001101101010101;
assign LUT_1[8243] = 32'b11111111111111111010111111010001;
assign LUT_1[8244] = 32'b00000000000000001101111000011011;
assign LUT_1[8245] = 32'b00000000000000000111001010010111;
assign LUT_1[8246] = 32'b00000000000000001001100110101100;
assign LUT_1[8247] = 32'b00000000000000000010111000101000;
assign LUT_1[8248] = 32'b00000000000000000101001100111001;
assign LUT_1[8249] = 32'b11111111111111111110011110110101;
assign LUT_1[8250] = 32'b00000000000000000000111011001010;
assign LUT_1[8251] = 32'b11111111111111111010001101000110;
assign LUT_1[8252] = 32'b00000000000000001101000110010000;
assign LUT_1[8253] = 32'b00000000000000000110011000001100;
assign LUT_1[8254] = 32'b00000000000000001000110100100001;
assign LUT_1[8255] = 32'b00000000000000000010000110011101;
assign LUT_1[8256] = 32'b00000000000000000101000110001011;
assign LUT_1[8257] = 32'b11111111111111111110011000000111;
assign LUT_1[8258] = 32'b00000000000000000000110100011100;
assign LUT_1[8259] = 32'b11111111111111111010000110011000;
assign LUT_1[8260] = 32'b00000000000000001100111111100010;
assign LUT_1[8261] = 32'b00000000000000000110010001011110;
assign LUT_1[8262] = 32'b00000000000000001000101101110011;
assign LUT_1[8263] = 32'b00000000000000000001111111101111;
assign LUT_1[8264] = 32'b00000000000000000100010100000000;
assign LUT_1[8265] = 32'b11111111111111111101100101111100;
assign LUT_1[8266] = 32'b00000000000000000000000010010001;
assign LUT_1[8267] = 32'b11111111111111111001010100001101;
assign LUT_1[8268] = 32'b00000000000000001100001101010111;
assign LUT_1[8269] = 32'b00000000000000000101011111010011;
assign LUT_1[8270] = 32'b00000000000000000111111011101000;
assign LUT_1[8271] = 32'b00000000000000000001001101100100;
assign LUT_1[8272] = 32'b00000000000000000111000001101101;
assign LUT_1[8273] = 32'b00000000000000000000010011101001;
assign LUT_1[8274] = 32'b00000000000000000010101111111110;
assign LUT_1[8275] = 32'b11111111111111111100000001111010;
assign LUT_1[8276] = 32'b00000000000000001110111011000100;
assign LUT_1[8277] = 32'b00000000000000001000001101000000;
assign LUT_1[8278] = 32'b00000000000000001010101001010101;
assign LUT_1[8279] = 32'b00000000000000000011111011010001;
assign LUT_1[8280] = 32'b00000000000000000110001111100010;
assign LUT_1[8281] = 32'b11111111111111111111100001011110;
assign LUT_1[8282] = 32'b00000000000000000001111101110011;
assign LUT_1[8283] = 32'b11111111111111111011001111101111;
assign LUT_1[8284] = 32'b00000000000000001110001000111001;
assign LUT_1[8285] = 32'b00000000000000000111011010110101;
assign LUT_1[8286] = 32'b00000000000000001001110111001010;
assign LUT_1[8287] = 32'b00000000000000000011001001000110;
assign LUT_1[8288] = 32'b00000000000000000110000001001010;
assign LUT_1[8289] = 32'b11111111111111111111010011000110;
assign LUT_1[8290] = 32'b00000000000000000001101111011011;
assign LUT_1[8291] = 32'b11111111111111111011000001010111;
assign LUT_1[8292] = 32'b00000000000000001101111010100001;
assign LUT_1[8293] = 32'b00000000000000000111001100011101;
assign LUT_1[8294] = 32'b00000000000000001001101000110010;
assign LUT_1[8295] = 32'b00000000000000000010111010101110;
assign LUT_1[8296] = 32'b00000000000000000101001110111111;
assign LUT_1[8297] = 32'b11111111111111111110100000111011;
assign LUT_1[8298] = 32'b00000000000000000000111101010000;
assign LUT_1[8299] = 32'b11111111111111111010001111001100;
assign LUT_1[8300] = 32'b00000000000000001101001000010110;
assign LUT_1[8301] = 32'b00000000000000000110011010010010;
assign LUT_1[8302] = 32'b00000000000000001000110110100111;
assign LUT_1[8303] = 32'b00000000000000000010001000100011;
assign LUT_1[8304] = 32'b00000000000000000111111100101100;
assign LUT_1[8305] = 32'b00000000000000000001001110101000;
assign LUT_1[8306] = 32'b00000000000000000011101010111101;
assign LUT_1[8307] = 32'b11111111111111111100111100111001;
assign LUT_1[8308] = 32'b00000000000000001111110110000011;
assign LUT_1[8309] = 32'b00000000000000001001000111111111;
assign LUT_1[8310] = 32'b00000000000000001011100100010100;
assign LUT_1[8311] = 32'b00000000000000000100110110010000;
assign LUT_1[8312] = 32'b00000000000000000111001010100001;
assign LUT_1[8313] = 32'b00000000000000000000011100011101;
assign LUT_1[8314] = 32'b00000000000000000010111000110010;
assign LUT_1[8315] = 32'b11111111111111111100001010101110;
assign LUT_1[8316] = 32'b00000000000000001111000011111000;
assign LUT_1[8317] = 32'b00000000000000001000010101110100;
assign LUT_1[8318] = 32'b00000000000000001010110010001001;
assign LUT_1[8319] = 32'b00000000000000000100000100000101;
assign LUT_1[8320] = 32'b00000000000000000110001000100110;
assign LUT_1[8321] = 32'b11111111111111111111011010100010;
assign LUT_1[8322] = 32'b00000000000000000001110110110111;
assign LUT_1[8323] = 32'b11111111111111111011001000110011;
assign LUT_1[8324] = 32'b00000000000000001110000001111101;
assign LUT_1[8325] = 32'b00000000000000000111010011111001;
assign LUT_1[8326] = 32'b00000000000000001001110000001110;
assign LUT_1[8327] = 32'b00000000000000000011000010001010;
assign LUT_1[8328] = 32'b00000000000000000101010110011011;
assign LUT_1[8329] = 32'b11111111111111111110101000010111;
assign LUT_1[8330] = 32'b00000000000000000001000100101100;
assign LUT_1[8331] = 32'b11111111111111111010010110101000;
assign LUT_1[8332] = 32'b00000000000000001101001111110010;
assign LUT_1[8333] = 32'b00000000000000000110100001101110;
assign LUT_1[8334] = 32'b00000000000000001000111110000011;
assign LUT_1[8335] = 32'b00000000000000000010001111111111;
assign LUT_1[8336] = 32'b00000000000000001000000100001000;
assign LUT_1[8337] = 32'b00000000000000000001010110000100;
assign LUT_1[8338] = 32'b00000000000000000011110010011001;
assign LUT_1[8339] = 32'b11111111111111111101000100010101;
assign LUT_1[8340] = 32'b00000000000000001111111101011111;
assign LUT_1[8341] = 32'b00000000000000001001001111011011;
assign LUT_1[8342] = 32'b00000000000000001011101011110000;
assign LUT_1[8343] = 32'b00000000000000000100111101101100;
assign LUT_1[8344] = 32'b00000000000000000111010001111101;
assign LUT_1[8345] = 32'b00000000000000000000100011111001;
assign LUT_1[8346] = 32'b00000000000000000011000000001110;
assign LUT_1[8347] = 32'b11111111111111111100010010001010;
assign LUT_1[8348] = 32'b00000000000000001111001011010100;
assign LUT_1[8349] = 32'b00000000000000001000011101010000;
assign LUT_1[8350] = 32'b00000000000000001010111001100101;
assign LUT_1[8351] = 32'b00000000000000000100001011100001;
assign LUT_1[8352] = 32'b00000000000000000111000011100101;
assign LUT_1[8353] = 32'b00000000000000000000010101100001;
assign LUT_1[8354] = 32'b00000000000000000010110001110110;
assign LUT_1[8355] = 32'b11111111111111111100000011110010;
assign LUT_1[8356] = 32'b00000000000000001110111100111100;
assign LUT_1[8357] = 32'b00000000000000001000001110111000;
assign LUT_1[8358] = 32'b00000000000000001010101011001101;
assign LUT_1[8359] = 32'b00000000000000000011111101001001;
assign LUT_1[8360] = 32'b00000000000000000110010001011010;
assign LUT_1[8361] = 32'b11111111111111111111100011010110;
assign LUT_1[8362] = 32'b00000000000000000001111111101011;
assign LUT_1[8363] = 32'b11111111111111111011010001100111;
assign LUT_1[8364] = 32'b00000000000000001110001010110001;
assign LUT_1[8365] = 32'b00000000000000000111011100101101;
assign LUT_1[8366] = 32'b00000000000000001001111001000010;
assign LUT_1[8367] = 32'b00000000000000000011001010111110;
assign LUT_1[8368] = 32'b00000000000000001000111111000111;
assign LUT_1[8369] = 32'b00000000000000000010010001000011;
assign LUT_1[8370] = 32'b00000000000000000100101101011000;
assign LUT_1[8371] = 32'b11111111111111111101111111010100;
assign LUT_1[8372] = 32'b00000000000000010000111000011110;
assign LUT_1[8373] = 32'b00000000000000001010001010011010;
assign LUT_1[8374] = 32'b00000000000000001100100110101111;
assign LUT_1[8375] = 32'b00000000000000000101111000101011;
assign LUT_1[8376] = 32'b00000000000000001000001100111100;
assign LUT_1[8377] = 32'b00000000000000000001011110111000;
assign LUT_1[8378] = 32'b00000000000000000011111011001101;
assign LUT_1[8379] = 32'b11111111111111111101001101001001;
assign LUT_1[8380] = 32'b00000000000000010000000110010011;
assign LUT_1[8381] = 32'b00000000000000001001011000001111;
assign LUT_1[8382] = 32'b00000000000000001011110100100100;
assign LUT_1[8383] = 32'b00000000000000000101000110100000;
assign LUT_1[8384] = 32'b00000000000000001000000110001110;
assign LUT_1[8385] = 32'b00000000000000000001011000001010;
assign LUT_1[8386] = 32'b00000000000000000011110100011111;
assign LUT_1[8387] = 32'b11111111111111111101000110011011;
assign LUT_1[8388] = 32'b00000000000000001111111111100101;
assign LUT_1[8389] = 32'b00000000000000001001010001100001;
assign LUT_1[8390] = 32'b00000000000000001011101101110110;
assign LUT_1[8391] = 32'b00000000000000000100111111110010;
assign LUT_1[8392] = 32'b00000000000000000111010100000011;
assign LUT_1[8393] = 32'b00000000000000000000100101111111;
assign LUT_1[8394] = 32'b00000000000000000011000010010100;
assign LUT_1[8395] = 32'b11111111111111111100010100010000;
assign LUT_1[8396] = 32'b00000000000000001111001101011010;
assign LUT_1[8397] = 32'b00000000000000001000011111010110;
assign LUT_1[8398] = 32'b00000000000000001010111011101011;
assign LUT_1[8399] = 32'b00000000000000000100001101100111;
assign LUT_1[8400] = 32'b00000000000000001010000001110000;
assign LUT_1[8401] = 32'b00000000000000000011010011101100;
assign LUT_1[8402] = 32'b00000000000000000101110000000001;
assign LUT_1[8403] = 32'b11111111111111111111000001111101;
assign LUT_1[8404] = 32'b00000000000000010001111011000111;
assign LUT_1[8405] = 32'b00000000000000001011001101000011;
assign LUT_1[8406] = 32'b00000000000000001101101001011000;
assign LUT_1[8407] = 32'b00000000000000000110111011010100;
assign LUT_1[8408] = 32'b00000000000000001001001111100101;
assign LUT_1[8409] = 32'b00000000000000000010100001100001;
assign LUT_1[8410] = 32'b00000000000000000100111101110110;
assign LUT_1[8411] = 32'b11111111111111111110001111110010;
assign LUT_1[8412] = 32'b00000000000000010001001000111100;
assign LUT_1[8413] = 32'b00000000000000001010011010111000;
assign LUT_1[8414] = 32'b00000000000000001100110111001101;
assign LUT_1[8415] = 32'b00000000000000000110001001001001;
assign LUT_1[8416] = 32'b00000000000000001001000001001101;
assign LUT_1[8417] = 32'b00000000000000000010010011001001;
assign LUT_1[8418] = 32'b00000000000000000100101111011110;
assign LUT_1[8419] = 32'b11111111111111111110000001011010;
assign LUT_1[8420] = 32'b00000000000000010000111010100100;
assign LUT_1[8421] = 32'b00000000000000001010001100100000;
assign LUT_1[8422] = 32'b00000000000000001100101000110101;
assign LUT_1[8423] = 32'b00000000000000000101111010110001;
assign LUT_1[8424] = 32'b00000000000000001000001111000010;
assign LUT_1[8425] = 32'b00000000000000000001100000111110;
assign LUT_1[8426] = 32'b00000000000000000011111101010011;
assign LUT_1[8427] = 32'b11111111111111111101001111001111;
assign LUT_1[8428] = 32'b00000000000000010000001000011001;
assign LUT_1[8429] = 32'b00000000000000001001011010010101;
assign LUT_1[8430] = 32'b00000000000000001011110110101010;
assign LUT_1[8431] = 32'b00000000000000000101001000100110;
assign LUT_1[8432] = 32'b00000000000000001010111100101111;
assign LUT_1[8433] = 32'b00000000000000000100001110101011;
assign LUT_1[8434] = 32'b00000000000000000110101011000000;
assign LUT_1[8435] = 32'b11111111111111111111111100111100;
assign LUT_1[8436] = 32'b00000000000000010010110110000110;
assign LUT_1[8437] = 32'b00000000000000001100001000000010;
assign LUT_1[8438] = 32'b00000000000000001110100100010111;
assign LUT_1[8439] = 32'b00000000000000000111110110010011;
assign LUT_1[8440] = 32'b00000000000000001010001010100100;
assign LUT_1[8441] = 32'b00000000000000000011011100100000;
assign LUT_1[8442] = 32'b00000000000000000101111000110101;
assign LUT_1[8443] = 32'b11111111111111111111001010110001;
assign LUT_1[8444] = 32'b00000000000000010010000011111011;
assign LUT_1[8445] = 32'b00000000000000001011010101110111;
assign LUT_1[8446] = 32'b00000000000000001101110010001100;
assign LUT_1[8447] = 32'b00000000000000000111000100001000;
assign LUT_1[8448] = 32'b00000000000000000000111100101111;
assign LUT_1[8449] = 32'b11111111111111111010001110101011;
assign LUT_1[8450] = 32'b11111111111111111100101011000000;
assign LUT_1[8451] = 32'b11111111111111110101111100111100;
assign LUT_1[8452] = 32'b00000000000000001000110110000110;
assign LUT_1[8453] = 32'b00000000000000000010001000000010;
assign LUT_1[8454] = 32'b00000000000000000100100100010111;
assign LUT_1[8455] = 32'b11111111111111111101110110010011;
assign LUT_1[8456] = 32'b00000000000000000000001010100100;
assign LUT_1[8457] = 32'b11111111111111111001011100100000;
assign LUT_1[8458] = 32'b11111111111111111011111000110101;
assign LUT_1[8459] = 32'b11111111111111110101001010110001;
assign LUT_1[8460] = 32'b00000000000000001000000011111011;
assign LUT_1[8461] = 32'b00000000000000000001010101110111;
assign LUT_1[8462] = 32'b00000000000000000011110010001100;
assign LUT_1[8463] = 32'b11111111111111111101000100001000;
assign LUT_1[8464] = 32'b00000000000000000010111000010001;
assign LUT_1[8465] = 32'b11111111111111111100001010001101;
assign LUT_1[8466] = 32'b11111111111111111110100110100010;
assign LUT_1[8467] = 32'b11111111111111110111111000011110;
assign LUT_1[8468] = 32'b00000000000000001010110001101000;
assign LUT_1[8469] = 32'b00000000000000000100000011100100;
assign LUT_1[8470] = 32'b00000000000000000110011111111001;
assign LUT_1[8471] = 32'b11111111111111111111110001110101;
assign LUT_1[8472] = 32'b00000000000000000010000110000110;
assign LUT_1[8473] = 32'b11111111111111111011011000000010;
assign LUT_1[8474] = 32'b11111111111111111101110100010111;
assign LUT_1[8475] = 32'b11111111111111110111000110010011;
assign LUT_1[8476] = 32'b00000000000000001001111111011101;
assign LUT_1[8477] = 32'b00000000000000000011010001011001;
assign LUT_1[8478] = 32'b00000000000000000101101101101110;
assign LUT_1[8479] = 32'b11111111111111111110111111101010;
assign LUT_1[8480] = 32'b00000000000000000001110111101110;
assign LUT_1[8481] = 32'b11111111111111111011001001101010;
assign LUT_1[8482] = 32'b11111111111111111101100101111111;
assign LUT_1[8483] = 32'b11111111111111110110110111111011;
assign LUT_1[8484] = 32'b00000000000000001001110001000101;
assign LUT_1[8485] = 32'b00000000000000000011000011000001;
assign LUT_1[8486] = 32'b00000000000000000101011111010110;
assign LUT_1[8487] = 32'b11111111111111111110110001010010;
assign LUT_1[8488] = 32'b00000000000000000001000101100011;
assign LUT_1[8489] = 32'b11111111111111111010010111011111;
assign LUT_1[8490] = 32'b11111111111111111100110011110100;
assign LUT_1[8491] = 32'b11111111111111110110000101110000;
assign LUT_1[8492] = 32'b00000000000000001000111110111010;
assign LUT_1[8493] = 32'b00000000000000000010010000110110;
assign LUT_1[8494] = 32'b00000000000000000100101101001011;
assign LUT_1[8495] = 32'b11111111111111111101111111000111;
assign LUT_1[8496] = 32'b00000000000000000011110011010000;
assign LUT_1[8497] = 32'b11111111111111111101000101001100;
assign LUT_1[8498] = 32'b11111111111111111111100001100001;
assign LUT_1[8499] = 32'b11111111111111111000110011011101;
assign LUT_1[8500] = 32'b00000000000000001011101100100111;
assign LUT_1[8501] = 32'b00000000000000000100111110100011;
assign LUT_1[8502] = 32'b00000000000000000111011010111000;
assign LUT_1[8503] = 32'b00000000000000000000101100110100;
assign LUT_1[8504] = 32'b00000000000000000011000001000101;
assign LUT_1[8505] = 32'b11111111111111111100010011000001;
assign LUT_1[8506] = 32'b11111111111111111110101111010110;
assign LUT_1[8507] = 32'b11111111111111111000000001010010;
assign LUT_1[8508] = 32'b00000000000000001010111010011100;
assign LUT_1[8509] = 32'b00000000000000000100001100011000;
assign LUT_1[8510] = 32'b00000000000000000110101000101101;
assign LUT_1[8511] = 32'b11111111111111111111111010101001;
assign LUT_1[8512] = 32'b00000000000000000010111010010111;
assign LUT_1[8513] = 32'b11111111111111111100001100010011;
assign LUT_1[8514] = 32'b11111111111111111110101000101000;
assign LUT_1[8515] = 32'b11111111111111110111111010100100;
assign LUT_1[8516] = 32'b00000000000000001010110011101110;
assign LUT_1[8517] = 32'b00000000000000000100000101101010;
assign LUT_1[8518] = 32'b00000000000000000110100001111111;
assign LUT_1[8519] = 32'b11111111111111111111110011111011;
assign LUT_1[8520] = 32'b00000000000000000010001000001100;
assign LUT_1[8521] = 32'b11111111111111111011011010001000;
assign LUT_1[8522] = 32'b11111111111111111101110110011101;
assign LUT_1[8523] = 32'b11111111111111110111001000011001;
assign LUT_1[8524] = 32'b00000000000000001010000001100011;
assign LUT_1[8525] = 32'b00000000000000000011010011011111;
assign LUT_1[8526] = 32'b00000000000000000101101111110100;
assign LUT_1[8527] = 32'b11111111111111111111000001110000;
assign LUT_1[8528] = 32'b00000000000000000100110101111001;
assign LUT_1[8529] = 32'b11111111111111111110000111110101;
assign LUT_1[8530] = 32'b00000000000000000000100100001010;
assign LUT_1[8531] = 32'b11111111111111111001110110000110;
assign LUT_1[8532] = 32'b00000000000000001100101111010000;
assign LUT_1[8533] = 32'b00000000000000000110000001001100;
assign LUT_1[8534] = 32'b00000000000000001000011101100001;
assign LUT_1[8535] = 32'b00000000000000000001101111011101;
assign LUT_1[8536] = 32'b00000000000000000100000011101110;
assign LUT_1[8537] = 32'b11111111111111111101010101101010;
assign LUT_1[8538] = 32'b11111111111111111111110001111111;
assign LUT_1[8539] = 32'b11111111111111111001000011111011;
assign LUT_1[8540] = 32'b00000000000000001011111101000101;
assign LUT_1[8541] = 32'b00000000000000000101001111000001;
assign LUT_1[8542] = 32'b00000000000000000111101011010110;
assign LUT_1[8543] = 32'b00000000000000000000111101010010;
assign LUT_1[8544] = 32'b00000000000000000011110101010110;
assign LUT_1[8545] = 32'b11111111111111111101000111010010;
assign LUT_1[8546] = 32'b11111111111111111111100011100111;
assign LUT_1[8547] = 32'b11111111111111111000110101100011;
assign LUT_1[8548] = 32'b00000000000000001011101110101101;
assign LUT_1[8549] = 32'b00000000000000000101000000101001;
assign LUT_1[8550] = 32'b00000000000000000111011100111110;
assign LUT_1[8551] = 32'b00000000000000000000101110111010;
assign LUT_1[8552] = 32'b00000000000000000011000011001011;
assign LUT_1[8553] = 32'b11111111111111111100010101000111;
assign LUT_1[8554] = 32'b11111111111111111110110001011100;
assign LUT_1[8555] = 32'b11111111111111111000000011011000;
assign LUT_1[8556] = 32'b00000000000000001010111100100010;
assign LUT_1[8557] = 32'b00000000000000000100001110011110;
assign LUT_1[8558] = 32'b00000000000000000110101010110011;
assign LUT_1[8559] = 32'b11111111111111111111111100101111;
assign LUT_1[8560] = 32'b00000000000000000101110000111000;
assign LUT_1[8561] = 32'b11111111111111111111000010110100;
assign LUT_1[8562] = 32'b00000000000000000001011111001001;
assign LUT_1[8563] = 32'b11111111111111111010110001000101;
assign LUT_1[8564] = 32'b00000000000000001101101010001111;
assign LUT_1[8565] = 32'b00000000000000000110111100001011;
assign LUT_1[8566] = 32'b00000000000000001001011000100000;
assign LUT_1[8567] = 32'b00000000000000000010101010011100;
assign LUT_1[8568] = 32'b00000000000000000100111110101101;
assign LUT_1[8569] = 32'b11111111111111111110010000101001;
assign LUT_1[8570] = 32'b00000000000000000000101100111110;
assign LUT_1[8571] = 32'b11111111111111111001111110111010;
assign LUT_1[8572] = 32'b00000000000000001100111000000100;
assign LUT_1[8573] = 32'b00000000000000000110001010000000;
assign LUT_1[8574] = 32'b00000000000000001000100110010101;
assign LUT_1[8575] = 32'b00000000000000000001111000010001;
assign LUT_1[8576] = 32'b00000000000000000011111100110010;
assign LUT_1[8577] = 32'b11111111111111111101001110101110;
assign LUT_1[8578] = 32'b11111111111111111111101011000011;
assign LUT_1[8579] = 32'b11111111111111111000111100111111;
assign LUT_1[8580] = 32'b00000000000000001011110110001001;
assign LUT_1[8581] = 32'b00000000000000000101001000000101;
assign LUT_1[8582] = 32'b00000000000000000111100100011010;
assign LUT_1[8583] = 32'b00000000000000000000110110010110;
assign LUT_1[8584] = 32'b00000000000000000011001010100111;
assign LUT_1[8585] = 32'b11111111111111111100011100100011;
assign LUT_1[8586] = 32'b11111111111111111110111000111000;
assign LUT_1[8587] = 32'b11111111111111111000001010110100;
assign LUT_1[8588] = 32'b00000000000000001011000011111110;
assign LUT_1[8589] = 32'b00000000000000000100010101111010;
assign LUT_1[8590] = 32'b00000000000000000110110010001111;
assign LUT_1[8591] = 32'b00000000000000000000000100001011;
assign LUT_1[8592] = 32'b00000000000000000101111000010100;
assign LUT_1[8593] = 32'b11111111111111111111001010010000;
assign LUT_1[8594] = 32'b00000000000000000001100110100101;
assign LUT_1[8595] = 32'b11111111111111111010111000100001;
assign LUT_1[8596] = 32'b00000000000000001101110001101011;
assign LUT_1[8597] = 32'b00000000000000000111000011100111;
assign LUT_1[8598] = 32'b00000000000000001001011111111100;
assign LUT_1[8599] = 32'b00000000000000000010110001111000;
assign LUT_1[8600] = 32'b00000000000000000101000110001001;
assign LUT_1[8601] = 32'b11111111111111111110011000000101;
assign LUT_1[8602] = 32'b00000000000000000000110100011010;
assign LUT_1[8603] = 32'b11111111111111111010000110010110;
assign LUT_1[8604] = 32'b00000000000000001100111111100000;
assign LUT_1[8605] = 32'b00000000000000000110010001011100;
assign LUT_1[8606] = 32'b00000000000000001000101101110001;
assign LUT_1[8607] = 32'b00000000000000000001111111101101;
assign LUT_1[8608] = 32'b00000000000000000100110111110001;
assign LUT_1[8609] = 32'b11111111111111111110001001101101;
assign LUT_1[8610] = 32'b00000000000000000000100110000010;
assign LUT_1[8611] = 32'b11111111111111111001110111111110;
assign LUT_1[8612] = 32'b00000000000000001100110001001000;
assign LUT_1[8613] = 32'b00000000000000000110000011000100;
assign LUT_1[8614] = 32'b00000000000000001000011111011001;
assign LUT_1[8615] = 32'b00000000000000000001110001010101;
assign LUT_1[8616] = 32'b00000000000000000100000101100110;
assign LUT_1[8617] = 32'b11111111111111111101010111100010;
assign LUT_1[8618] = 32'b11111111111111111111110011110111;
assign LUT_1[8619] = 32'b11111111111111111001000101110011;
assign LUT_1[8620] = 32'b00000000000000001011111110111101;
assign LUT_1[8621] = 32'b00000000000000000101010000111001;
assign LUT_1[8622] = 32'b00000000000000000111101101001110;
assign LUT_1[8623] = 32'b00000000000000000000111111001010;
assign LUT_1[8624] = 32'b00000000000000000110110011010011;
assign LUT_1[8625] = 32'b00000000000000000000000101001111;
assign LUT_1[8626] = 32'b00000000000000000010100001100100;
assign LUT_1[8627] = 32'b11111111111111111011110011100000;
assign LUT_1[8628] = 32'b00000000000000001110101100101010;
assign LUT_1[8629] = 32'b00000000000000000111111110100110;
assign LUT_1[8630] = 32'b00000000000000001010011010111011;
assign LUT_1[8631] = 32'b00000000000000000011101100110111;
assign LUT_1[8632] = 32'b00000000000000000110000001001000;
assign LUT_1[8633] = 32'b11111111111111111111010011000100;
assign LUT_1[8634] = 32'b00000000000000000001101111011001;
assign LUT_1[8635] = 32'b11111111111111111011000001010101;
assign LUT_1[8636] = 32'b00000000000000001101111010011111;
assign LUT_1[8637] = 32'b00000000000000000111001100011011;
assign LUT_1[8638] = 32'b00000000000000001001101000110000;
assign LUT_1[8639] = 32'b00000000000000000010111010101100;
assign LUT_1[8640] = 32'b00000000000000000101111010011010;
assign LUT_1[8641] = 32'b11111111111111111111001100010110;
assign LUT_1[8642] = 32'b00000000000000000001101000101011;
assign LUT_1[8643] = 32'b11111111111111111010111010100111;
assign LUT_1[8644] = 32'b00000000000000001101110011110001;
assign LUT_1[8645] = 32'b00000000000000000111000101101101;
assign LUT_1[8646] = 32'b00000000000000001001100010000010;
assign LUT_1[8647] = 32'b00000000000000000010110011111110;
assign LUT_1[8648] = 32'b00000000000000000101001000001111;
assign LUT_1[8649] = 32'b11111111111111111110011010001011;
assign LUT_1[8650] = 32'b00000000000000000000110110100000;
assign LUT_1[8651] = 32'b11111111111111111010001000011100;
assign LUT_1[8652] = 32'b00000000000000001101000001100110;
assign LUT_1[8653] = 32'b00000000000000000110010011100010;
assign LUT_1[8654] = 32'b00000000000000001000101111110111;
assign LUT_1[8655] = 32'b00000000000000000010000001110011;
assign LUT_1[8656] = 32'b00000000000000000111110101111100;
assign LUT_1[8657] = 32'b00000000000000000001000111111000;
assign LUT_1[8658] = 32'b00000000000000000011100100001101;
assign LUT_1[8659] = 32'b11111111111111111100110110001001;
assign LUT_1[8660] = 32'b00000000000000001111101111010011;
assign LUT_1[8661] = 32'b00000000000000001001000001001111;
assign LUT_1[8662] = 32'b00000000000000001011011101100100;
assign LUT_1[8663] = 32'b00000000000000000100101111100000;
assign LUT_1[8664] = 32'b00000000000000000111000011110001;
assign LUT_1[8665] = 32'b00000000000000000000010101101101;
assign LUT_1[8666] = 32'b00000000000000000010110010000010;
assign LUT_1[8667] = 32'b11111111111111111100000011111110;
assign LUT_1[8668] = 32'b00000000000000001110111101001000;
assign LUT_1[8669] = 32'b00000000000000001000001111000100;
assign LUT_1[8670] = 32'b00000000000000001010101011011001;
assign LUT_1[8671] = 32'b00000000000000000011111101010101;
assign LUT_1[8672] = 32'b00000000000000000110110101011001;
assign LUT_1[8673] = 32'b00000000000000000000000111010101;
assign LUT_1[8674] = 32'b00000000000000000010100011101010;
assign LUT_1[8675] = 32'b11111111111111111011110101100110;
assign LUT_1[8676] = 32'b00000000000000001110101110110000;
assign LUT_1[8677] = 32'b00000000000000001000000000101100;
assign LUT_1[8678] = 32'b00000000000000001010011101000001;
assign LUT_1[8679] = 32'b00000000000000000011101110111101;
assign LUT_1[8680] = 32'b00000000000000000110000011001110;
assign LUT_1[8681] = 32'b11111111111111111111010101001010;
assign LUT_1[8682] = 32'b00000000000000000001110001011111;
assign LUT_1[8683] = 32'b11111111111111111011000011011011;
assign LUT_1[8684] = 32'b00000000000000001101111100100101;
assign LUT_1[8685] = 32'b00000000000000000111001110100001;
assign LUT_1[8686] = 32'b00000000000000001001101010110110;
assign LUT_1[8687] = 32'b00000000000000000010111100110010;
assign LUT_1[8688] = 32'b00000000000000001000110000111011;
assign LUT_1[8689] = 32'b00000000000000000010000010110111;
assign LUT_1[8690] = 32'b00000000000000000100011111001100;
assign LUT_1[8691] = 32'b11111111111111111101110001001000;
assign LUT_1[8692] = 32'b00000000000000010000101010010010;
assign LUT_1[8693] = 32'b00000000000000001001111100001110;
assign LUT_1[8694] = 32'b00000000000000001100011000100011;
assign LUT_1[8695] = 32'b00000000000000000101101010011111;
assign LUT_1[8696] = 32'b00000000000000000111111110110000;
assign LUT_1[8697] = 32'b00000000000000000001010000101100;
assign LUT_1[8698] = 32'b00000000000000000011101101000001;
assign LUT_1[8699] = 32'b11111111111111111100111110111101;
assign LUT_1[8700] = 32'b00000000000000001111111000000111;
assign LUT_1[8701] = 32'b00000000000000001001001010000011;
assign LUT_1[8702] = 32'b00000000000000001011100110011000;
assign LUT_1[8703] = 32'b00000000000000000100111000010100;
assign LUT_1[8704] = 32'b11111111111111111100110111000000;
assign LUT_1[8705] = 32'b11111111111111110110001000111100;
assign LUT_1[8706] = 32'b11111111111111111000100101010001;
assign LUT_1[8707] = 32'b11111111111111110001110111001101;
assign LUT_1[8708] = 32'b00000000000000000100110000010111;
assign LUT_1[8709] = 32'b11111111111111111110000010010011;
assign LUT_1[8710] = 32'b00000000000000000000011110101000;
assign LUT_1[8711] = 32'b11111111111111111001110000100100;
assign LUT_1[8712] = 32'b11111111111111111100000100110101;
assign LUT_1[8713] = 32'b11111111111111110101010110110001;
assign LUT_1[8714] = 32'b11111111111111110111110011000110;
assign LUT_1[8715] = 32'b11111111111111110001000101000010;
assign LUT_1[8716] = 32'b00000000000000000011111110001100;
assign LUT_1[8717] = 32'b11111111111111111101010000001000;
assign LUT_1[8718] = 32'b11111111111111111111101100011101;
assign LUT_1[8719] = 32'b11111111111111111000111110011001;
assign LUT_1[8720] = 32'b11111111111111111110110010100010;
assign LUT_1[8721] = 32'b11111111111111111000000100011110;
assign LUT_1[8722] = 32'b11111111111111111010100000110011;
assign LUT_1[8723] = 32'b11111111111111110011110010101111;
assign LUT_1[8724] = 32'b00000000000000000110101011111001;
assign LUT_1[8725] = 32'b11111111111111111111111101110101;
assign LUT_1[8726] = 32'b00000000000000000010011010001010;
assign LUT_1[8727] = 32'b11111111111111111011101100000110;
assign LUT_1[8728] = 32'b11111111111111111110000000010111;
assign LUT_1[8729] = 32'b11111111111111110111010010010011;
assign LUT_1[8730] = 32'b11111111111111111001101110101000;
assign LUT_1[8731] = 32'b11111111111111110011000000100100;
assign LUT_1[8732] = 32'b00000000000000000101111001101110;
assign LUT_1[8733] = 32'b11111111111111111111001011101010;
assign LUT_1[8734] = 32'b00000000000000000001100111111111;
assign LUT_1[8735] = 32'b11111111111111111010111001111011;
assign LUT_1[8736] = 32'b11111111111111111101110001111111;
assign LUT_1[8737] = 32'b11111111111111110111000011111011;
assign LUT_1[8738] = 32'b11111111111111111001100000010000;
assign LUT_1[8739] = 32'b11111111111111110010110010001100;
assign LUT_1[8740] = 32'b00000000000000000101101011010110;
assign LUT_1[8741] = 32'b11111111111111111110111101010010;
assign LUT_1[8742] = 32'b00000000000000000001011001100111;
assign LUT_1[8743] = 32'b11111111111111111010101011100011;
assign LUT_1[8744] = 32'b11111111111111111100111111110100;
assign LUT_1[8745] = 32'b11111111111111110110010001110000;
assign LUT_1[8746] = 32'b11111111111111111000101110000101;
assign LUT_1[8747] = 32'b11111111111111110010000000000001;
assign LUT_1[8748] = 32'b00000000000000000100111001001011;
assign LUT_1[8749] = 32'b11111111111111111110001011000111;
assign LUT_1[8750] = 32'b00000000000000000000100111011100;
assign LUT_1[8751] = 32'b11111111111111111001111001011000;
assign LUT_1[8752] = 32'b11111111111111111111101101100001;
assign LUT_1[8753] = 32'b11111111111111111000111111011101;
assign LUT_1[8754] = 32'b11111111111111111011011011110010;
assign LUT_1[8755] = 32'b11111111111111110100101101101110;
assign LUT_1[8756] = 32'b00000000000000000111100110111000;
assign LUT_1[8757] = 32'b00000000000000000000111000110100;
assign LUT_1[8758] = 32'b00000000000000000011010101001001;
assign LUT_1[8759] = 32'b11111111111111111100100111000101;
assign LUT_1[8760] = 32'b11111111111111111110111011010110;
assign LUT_1[8761] = 32'b11111111111111111000001101010010;
assign LUT_1[8762] = 32'b11111111111111111010101001100111;
assign LUT_1[8763] = 32'b11111111111111110011111011100011;
assign LUT_1[8764] = 32'b00000000000000000110110100101101;
assign LUT_1[8765] = 32'b00000000000000000000000110101001;
assign LUT_1[8766] = 32'b00000000000000000010100010111110;
assign LUT_1[8767] = 32'b11111111111111111011110100111010;
assign LUT_1[8768] = 32'b11111111111111111110110100101000;
assign LUT_1[8769] = 32'b11111111111111111000000110100100;
assign LUT_1[8770] = 32'b11111111111111111010100010111001;
assign LUT_1[8771] = 32'b11111111111111110011110100110101;
assign LUT_1[8772] = 32'b00000000000000000110101101111111;
assign LUT_1[8773] = 32'b11111111111111111111111111111011;
assign LUT_1[8774] = 32'b00000000000000000010011100010000;
assign LUT_1[8775] = 32'b11111111111111111011101110001100;
assign LUT_1[8776] = 32'b11111111111111111110000010011101;
assign LUT_1[8777] = 32'b11111111111111110111010100011001;
assign LUT_1[8778] = 32'b11111111111111111001110000101110;
assign LUT_1[8779] = 32'b11111111111111110011000010101010;
assign LUT_1[8780] = 32'b00000000000000000101111011110100;
assign LUT_1[8781] = 32'b11111111111111111111001101110000;
assign LUT_1[8782] = 32'b00000000000000000001101010000101;
assign LUT_1[8783] = 32'b11111111111111111010111100000001;
assign LUT_1[8784] = 32'b00000000000000000000110000001010;
assign LUT_1[8785] = 32'b11111111111111111010000010000110;
assign LUT_1[8786] = 32'b11111111111111111100011110011011;
assign LUT_1[8787] = 32'b11111111111111110101110000010111;
assign LUT_1[8788] = 32'b00000000000000001000101001100001;
assign LUT_1[8789] = 32'b00000000000000000001111011011101;
assign LUT_1[8790] = 32'b00000000000000000100010111110010;
assign LUT_1[8791] = 32'b11111111111111111101101001101110;
assign LUT_1[8792] = 32'b11111111111111111111111101111111;
assign LUT_1[8793] = 32'b11111111111111111001001111111011;
assign LUT_1[8794] = 32'b11111111111111111011101100010000;
assign LUT_1[8795] = 32'b11111111111111110100111110001100;
assign LUT_1[8796] = 32'b00000000000000000111110111010110;
assign LUT_1[8797] = 32'b00000000000000000001001001010010;
assign LUT_1[8798] = 32'b00000000000000000011100101100111;
assign LUT_1[8799] = 32'b11111111111111111100110111100011;
assign LUT_1[8800] = 32'b11111111111111111111101111100111;
assign LUT_1[8801] = 32'b11111111111111111001000001100011;
assign LUT_1[8802] = 32'b11111111111111111011011101111000;
assign LUT_1[8803] = 32'b11111111111111110100101111110100;
assign LUT_1[8804] = 32'b00000000000000000111101000111110;
assign LUT_1[8805] = 32'b00000000000000000000111010111010;
assign LUT_1[8806] = 32'b00000000000000000011010111001111;
assign LUT_1[8807] = 32'b11111111111111111100101001001011;
assign LUT_1[8808] = 32'b11111111111111111110111101011100;
assign LUT_1[8809] = 32'b11111111111111111000001111011000;
assign LUT_1[8810] = 32'b11111111111111111010101011101101;
assign LUT_1[8811] = 32'b11111111111111110011111101101001;
assign LUT_1[8812] = 32'b00000000000000000110110110110011;
assign LUT_1[8813] = 32'b00000000000000000000001000101111;
assign LUT_1[8814] = 32'b00000000000000000010100101000100;
assign LUT_1[8815] = 32'b11111111111111111011110111000000;
assign LUT_1[8816] = 32'b00000000000000000001101011001001;
assign LUT_1[8817] = 32'b11111111111111111010111101000101;
assign LUT_1[8818] = 32'b11111111111111111101011001011010;
assign LUT_1[8819] = 32'b11111111111111110110101011010110;
assign LUT_1[8820] = 32'b00000000000000001001100100100000;
assign LUT_1[8821] = 32'b00000000000000000010110110011100;
assign LUT_1[8822] = 32'b00000000000000000101010010110001;
assign LUT_1[8823] = 32'b11111111111111111110100100101101;
assign LUT_1[8824] = 32'b00000000000000000000111000111110;
assign LUT_1[8825] = 32'b11111111111111111010001010111010;
assign LUT_1[8826] = 32'b11111111111111111100100111001111;
assign LUT_1[8827] = 32'b11111111111111110101111001001011;
assign LUT_1[8828] = 32'b00000000000000001000110010010101;
assign LUT_1[8829] = 32'b00000000000000000010000100010001;
assign LUT_1[8830] = 32'b00000000000000000100100000100110;
assign LUT_1[8831] = 32'b11111111111111111101110010100010;
assign LUT_1[8832] = 32'b11111111111111111111110111000011;
assign LUT_1[8833] = 32'b11111111111111111001001000111111;
assign LUT_1[8834] = 32'b11111111111111111011100101010100;
assign LUT_1[8835] = 32'b11111111111111110100110111010000;
assign LUT_1[8836] = 32'b00000000000000000111110000011010;
assign LUT_1[8837] = 32'b00000000000000000001000010010110;
assign LUT_1[8838] = 32'b00000000000000000011011110101011;
assign LUT_1[8839] = 32'b11111111111111111100110000100111;
assign LUT_1[8840] = 32'b11111111111111111111000100111000;
assign LUT_1[8841] = 32'b11111111111111111000010110110100;
assign LUT_1[8842] = 32'b11111111111111111010110011001001;
assign LUT_1[8843] = 32'b11111111111111110100000101000101;
assign LUT_1[8844] = 32'b00000000000000000110111110001111;
assign LUT_1[8845] = 32'b00000000000000000000010000001011;
assign LUT_1[8846] = 32'b00000000000000000010101100100000;
assign LUT_1[8847] = 32'b11111111111111111011111110011100;
assign LUT_1[8848] = 32'b00000000000000000001110010100101;
assign LUT_1[8849] = 32'b11111111111111111011000100100001;
assign LUT_1[8850] = 32'b11111111111111111101100000110110;
assign LUT_1[8851] = 32'b11111111111111110110110010110010;
assign LUT_1[8852] = 32'b00000000000000001001101011111100;
assign LUT_1[8853] = 32'b00000000000000000010111101111000;
assign LUT_1[8854] = 32'b00000000000000000101011010001101;
assign LUT_1[8855] = 32'b11111111111111111110101100001001;
assign LUT_1[8856] = 32'b00000000000000000001000000011010;
assign LUT_1[8857] = 32'b11111111111111111010010010010110;
assign LUT_1[8858] = 32'b11111111111111111100101110101011;
assign LUT_1[8859] = 32'b11111111111111110110000000100111;
assign LUT_1[8860] = 32'b00000000000000001000111001110001;
assign LUT_1[8861] = 32'b00000000000000000010001011101101;
assign LUT_1[8862] = 32'b00000000000000000100101000000010;
assign LUT_1[8863] = 32'b11111111111111111101111001111110;
assign LUT_1[8864] = 32'b00000000000000000000110010000010;
assign LUT_1[8865] = 32'b11111111111111111010000011111110;
assign LUT_1[8866] = 32'b11111111111111111100100000010011;
assign LUT_1[8867] = 32'b11111111111111110101110010001111;
assign LUT_1[8868] = 32'b00000000000000001000101011011001;
assign LUT_1[8869] = 32'b00000000000000000001111101010101;
assign LUT_1[8870] = 32'b00000000000000000100011001101010;
assign LUT_1[8871] = 32'b11111111111111111101101011100110;
assign LUT_1[8872] = 32'b11111111111111111111111111110111;
assign LUT_1[8873] = 32'b11111111111111111001010001110011;
assign LUT_1[8874] = 32'b11111111111111111011101110001000;
assign LUT_1[8875] = 32'b11111111111111110101000000000100;
assign LUT_1[8876] = 32'b00000000000000000111111001001110;
assign LUT_1[8877] = 32'b00000000000000000001001011001010;
assign LUT_1[8878] = 32'b00000000000000000011100111011111;
assign LUT_1[8879] = 32'b11111111111111111100111001011011;
assign LUT_1[8880] = 32'b00000000000000000010101101100100;
assign LUT_1[8881] = 32'b11111111111111111011111111100000;
assign LUT_1[8882] = 32'b11111111111111111110011011110101;
assign LUT_1[8883] = 32'b11111111111111110111101101110001;
assign LUT_1[8884] = 32'b00000000000000001010100110111011;
assign LUT_1[8885] = 32'b00000000000000000011111000110111;
assign LUT_1[8886] = 32'b00000000000000000110010101001100;
assign LUT_1[8887] = 32'b11111111111111111111100111001000;
assign LUT_1[8888] = 32'b00000000000000000001111011011001;
assign LUT_1[8889] = 32'b11111111111111111011001101010101;
assign LUT_1[8890] = 32'b11111111111111111101101001101010;
assign LUT_1[8891] = 32'b11111111111111110110111011100110;
assign LUT_1[8892] = 32'b00000000000000001001110100110000;
assign LUT_1[8893] = 32'b00000000000000000011000110101100;
assign LUT_1[8894] = 32'b00000000000000000101100011000001;
assign LUT_1[8895] = 32'b11111111111111111110110100111101;
assign LUT_1[8896] = 32'b00000000000000000001110100101011;
assign LUT_1[8897] = 32'b11111111111111111011000110100111;
assign LUT_1[8898] = 32'b11111111111111111101100010111100;
assign LUT_1[8899] = 32'b11111111111111110110110100111000;
assign LUT_1[8900] = 32'b00000000000000001001101110000010;
assign LUT_1[8901] = 32'b00000000000000000010111111111110;
assign LUT_1[8902] = 32'b00000000000000000101011100010011;
assign LUT_1[8903] = 32'b11111111111111111110101110001111;
assign LUT_1[8904] = 32'b00000000000000000001000010100000;
assign LUT_1[8905] = 32'b11111111111111111010010100011100;
assign LUT_1[8906] = 32'b11111111111111111100110000110001;
assign LUT_1[8907] = 32'b11111111111111110110000010101101;
assign LUT_1[8908] = 32'b00000000000000001000111011110111;
assign LUT_1[8909] = 32'b00000000000000000010001101110011;
assign LUT_1[8910] = 32'b00000000000000000100101010001000;
assign LUT_1[8911] = 32'b11111111111111111101111100000100;
assign LUT_1[8912] = 32'b00000000000000000011110000001101;
assign LUT_1[8913] = 32'b11111111111111111101000010001001;
assign LUT_1[8914] = 32'b11111111111111111111011110011110;
assign LUT_1[8915] = 32'b11111111111111111000110000011010;
assign LUT_1[8916] = 32'b00000000000000001011101001100100;
assign LUT_1[8917] = 32'b00000000000000000100111011100000;
assign LUT_1[8918] = 32'b00000000000000000111010111110101;
assign LUT_1[8919] = 32'b00000000000000000000101001110001;
assign LUT_1[8920] = 32'b00000000000000000010111110000010;
assign LUT_1[8921] = 32'b11111111111111111100001111111110;
assign LUT_1[8922] = 32'b11111111111111111110101100010011;
assign LUT_1[8923] = 32'b11111111111111110111111110001111;
assign LUT_1[8924] = 32'b00000000000000001010110111011001;
assign LUT_1[8925] = 32'b00000000000000000100001001010101;
assign LUT_1[8926] = 32'b00000000000000000110100101101010;
assign LUT_1[8927] = 32'b11111111111111111111110111100110;
assign LUT_1[8928] = 32'b00000000000000000010101111101010;
assign LUT_1[8929] = 32'b11111111111111111100000001100110;
assign LUT_1[8930] = 32'b11111111111111111110011101111011;
assign LUT_1[8931] = 32'b11111111111111110111101111110111;
assign LUT_1[8932] = 32'b00000000000000001010101001000001;
assign LUT_1[8933] = 32'b00000000000000000011111010111101;
assign LUT_1[8934] = 32'b00000000000000000110010111010010;
assign LUT_1[8935] = 32'b11111111111111111111101001001110;
assign LUT_1[8936] = 32'b00000000000000000001111101011111;
assign LUT_1[8937] = 32'b11111111111111111011001111011011;
assign LUT_1[8938] = 32'b11111111111111111101101011110000;
assign LUT_1[8939] = 32'b11111111111111110110111101101100;
assign LUT_1[8940] = 32'b00000000000000001001110110110110;
assign LUT_1[8941] = 32'b00000000000000000011001000110010;
assign LUT_1[8942] = 32'b00000000000000000101100101000111;
assign LUT_1[8943] = 32'b11111111111111111110110111000011;
assign LUT_1[8944] = 32'b00000000000000000100101011001100;
assign LUT_1[8945] = 32'b11111111111111111101111101001000;
assign LUT_1[8946] = 32'b00000000000000000000011001011101;
assign LUT_1[8947] = 32'b11111111111111111001101011011001;
assign LUT_1[8948] = 32'b00000000000000001100100100100011;
assign LUT_1[8949] = 32'b00000000000000000101110110011111;
assign LUT_1[8950] = 32'b00000000000000001000010010110100;
assign LUT_1[8951] = 32'b00000000000000000001100100110000;
assign LUT_1[8952] = 32'b00000000000000000011111001000001;
assign LUT_1[8953] = 32'b11111111111111111101001010111101;
assign LUT_1[8954] = 32'b11111111111111111111100111010010;
assign LUT_1[8955] = 32'b11111111111111111000111001001110;
assign LUT_1[8956] = 32'b00000000000000001011110010011000;
assign LUT_1[8957] = 32'b00000000000000000101000100010100;
assign LUT_1[8958] = 32'b00000000000000000111100000101001;
assign LUT_1[8959] = 32'b00000000000000000000110010100101;
assign LUT_1[8960] = 32'b11111111111111111010101011001100;
assign LUT_1[8961] = 32'b11111111111111110011111101001000;
assign LUT_1[8962] = 32'b11111111111111110110011001011101;
assign LUT_1[8963] = 32'b11111111111111101111101011011001;
assign LUT_1[8964] = 32'b00000000000000000010100100100011;
assign LUT_1[8965] = 32'b11111111111111111011110110011111;
assign LUT_1[8966] = 32'b11111111111111111110010010110100;
assign LUT_1[8967] = 32'b11111111111111110111100100110000;
assign LUT_1[8968] = 32'b11111111111111111001111001000001;
assign LUT_1[8969] = 32'b11111111111111110011001010111101;
assign LUT_1[8970] = 32'b11111111111111110101100111010010;
assign LUT_1[8971] = 32'b11111111111111101110111001001110;
assign LUT_1[8972] = 32'b00000000000000000001110010011000;
assign LUT_1[8973] = 32'b11111111111111111011000100010100;
assign LUT_1[8974] = 32'b11111111111111111101100000101001;
assign LUT_1[8975] = 32'b11111111111111110110110010100101;
assign LUT_1[8976] = 32'b11111111111111111100100110101110;
assign LUT_1[8977] = 32'b11111111111111110101111000101010;
assign LUT_1[8978] = 32'b11111111111111111000010100111111;
assign LUT_1[8979] = 32'b11111111111111110001100110111011;
assign LUT_1[8980] = 32'b00000000000000000100100000000101;
assign LUT_1[8981] = 32'b11111111111111111101110010000001;
assign LUT_1[8982] = 32'b00000000000000000000001110010110;
assign LUT_1[8983] = 32'b11111111111111111001100000010010;
assign LUT_1[8984] = 32'b11111111111111111011110100100011;
assign LUT_1[8985] = 32'b11111111111111110101000110011111;
assign LUT_1[8986] = 32'b11111111111111110111100010110100;
assign LUT_1[8987] = 32'b11111111111111110000110100110000;
assign LUT_1[8988] = 32'b00000000000000000011101101111010;
assign LUT_1[8989] = 32'b11111111111111111100111111110110;
assign LUT_1[8990] = 32'b11111111111111111111011100001011;
assign LUT_1[8991] = 32'b11111111111111111000101110000111;
assign LUT_1[8992] = 32'b11111111111111111011100110001011;
assign LUT_1[8993] = 32'b11111111111111110100111000000111;
assign LUT_1[8994] = 32'b11111111111111110111010100011100;
assign LUT_1[8995] = 32'b11111111111111110000100110011000;
assign LUT_1[8996] = 32'b00000000000000000011011111100010;
assign LUT_1[8997] = 32'b11111111111111111100110001011110;
assign LUT_1[8998] = 32'b11111111111111111111001101110011;
assign LUT_1[8999] = 32'b11111111111111111000011111101111;
assign LUT_1[9000] = 32'b11111111111111111010110100000000;
assign LUT_1[9001] = 32'b11111111111111110100000101111100;
assign LUT_1[9002] = 32'b11111111111111110110100010010001;
assign LUT_1[9003] = 32'b11111111111111101111110100001101;
assign LUT_1[9004] = 32'b00000000000000000010101101010111;
assign LUT_1[9005] = 32'b11111111111111111011111111010011;
assign LUT_1[9006] = 32'b11111111111111111110011011101000;
assign LUT_1[9007] = 32'b11111111111111110111101101100100;
assign LUT_1[9008] = 32'b11111111111111111101100001101101;
assign LUT_1[9009] = 32'b11111111111111110110110011101001;
assign LUT_1[9010] = 32'b11111111111111111001001111111110;
assign LUT_1[9011] = 32'b11111111111111110010100001111010;
assign LUT_1[9012] = 32'b00000000000000000101011011000100;
assign LUT_1[9013] = 32'b11111111111111111110101101000000;
assign LUT_1[9014] = 32'b00000000000000000001001001010101;
assign LUT_1[9015] = 32'b11111111111111111010011011010001;
assign LUT_1[9016] = 32'b11111111111111111100101111100010;
assign LUT_1[9017] = 32'b11111111111111110110000001011110;
assign LUT_1[9018] = 32'b11111111111111111000011101110011;
assign LUT_1[9019] = 32'b11111111111111110001101111101111;
assign LUT_1[9020] = 32'b00000000000000000100101000111001;
assign LUT_1[9021] = 32'b11111111111111111101111010110101;
assign LUT_1[9022] = 32'b00000000000000000000010111001010;
assign LUT_1[9023] = 32'b11111111111111111001101001000110;
assign LUT_1[9024] = 32'b11111111111111111100101000110100;
assign LUT_1[9025] = 32'b11111111111111110101111010110000;
assign LUT_1[9026] = 32'b11111111111111111000010111000101;
assign LUT_1[9027] = 32'b11111111111111110001101001000001;
assign LUT_1[9028] = 32'b00000000000000000100100010001011;
assign LUT_1[9029] = 32'b11111111111111111101110100000111;
assign LUT_1[9030] = 32'b00000000000000000000010000011100;
assign LUT_1[9031] = 32'b11111111111111111001100010011000;
assign LUT_1[9032] = 32'b11111111111111111011110110101001;
assign LUT_1[9033] = 32'b11111111111111110101001000100101;
assign LUT_1[9034] = 32'b11111111111111110111100100111010;
assign LUT_1[9035] = 32'b11111111111111110000110110110110;
assign LUT_1[9036] = 32'b00000000000000000011110000000000;
assign LUT_1[9037] = 32'b11111111111111111101000001111100;
assign LUT_1[9038] = 32'b11111111111111111111011110010001;
assign LUT_1[9039] = 32'b11111111111111111000110000001101;
assign LUT_1[9040] = 32'b11111111111111111110100100010110;
assign LUT_1[9041] = 32'b11111111111111110111110110010010;
assign LUT_1[9042] = 32'b11111111111111111010010010100111;
assign LUT_1[9043] = 32'b11111111111111110011100100100011;
assign LUT_1[9044] = 32'b00000000000000000110011101101101;
assign LUT_1[9045] = 32'b11111111111111111111101111101001;
assign LUT_1[9046] = 32'b00000000000000000010001011111110;
assign LUT_1[9047] = 32'b11111111111111111011011101111010;
assign LUT_1[9048] = 32'b11111111111111111101110010001011;
assign LUT_1[9049] = 32'b11111111111111110111000100000111;
assign LUT_1[9050] = 32'b11111111111111111001100000011100;
assign LUT_1[9051] = 32'b11111111111111110010110010011000;
assign LUT_1[9052] = 32'b00000000000000000101101011100010;
assign LUT_1[9053] = 32'b11111111111111111110111101011110;
assign LUT_1[9054] = 32'b00000000000000000001011001110011;
assign LUT_1[9055] = 32'b11111111111111111010101011101111;
assign LUT_1[9056] = 32'b11111111111111111101100011110011;
assign LUT_1[9057] = 32'b11111111111111110110110101101111;
assign LUT_1[9058] = 32'b11111111111111111001010010000100;
assign LUT_1[9059] = 32'b11111111111111110010100100000000;
assign LUT_1[9060] = 32'b00000000000000000101011101001010;
assign LUT_1[9061] = 32'b11111111111111111110101111000110;
assign LUT_1[9062] = 32'b00000000000000000001001011011011;
assign LUT_1[9063] = 32'b11111111111111111010011101010111;
assign LUT_1[9064] = 32'b11111111111111111100110001101000;
assign LUT_1[9065] = 32'b11111111111111110110000011100100;
assign LUT_1[9066] = 32'b11111111111111111000011111111001;
assign LUT_1[9067] = 32'b11111111111111110001110001110101;
assign LUT_1[9068] = 32'b00000000000000000100101010111111;
assign LUT_1[9069] = 32'b11111111111111111101111100111011;
assign LUT_1[9070] = 32'b00000000000000000000011001010000;
assign LUT_1[9071] = 32'b11111111111111111001101011001100;
assign LUT_1[9072] = 32'b11111111111111111111011111010101;
assign LUT_1[9073] = 32'b11111111111111111000110001010001;
assign LUT_1[9074] = 32'b11111111111111111011001101100110;
assign LUT_1[9075] = 32'b11111111111111110100011111100010;
assign LUT_1[9076] = 32'b00000000000000000111011000101100;
assign LUT_1[9077] = 32'b00000000000000000000101010101000;
assign LUT_1[9078] = 32'b00000000000000000011000110111101;
assign LUT_1[9079] = 32'b11111111111111111100011000111001;
assign LUT_1[9080] = 32'b11111111111111111110101101001010;
assign LUT_1[9081] = 32'b11111111111111110111111111000110;
assign LUT_1[9082] = 32'b11111111111111111010011011011011;
assign LUT_1[9083] = 32'b11111111111111110011101101010111;
assign LUT_1[9084] = 32'b00000000000000000110100110100001;
assign LUT_1[9085] = 32'b11111111111111111111111000011101;
assign LUT_1[9086] = 32'b00000000000000000010010100110010;
assign LUT_1[9087] = 32'b11111111111111111011100110101110;
assign LUT_1[9088] = 32'b11111111111111111101101011001111;
assign LUT_1[9089] = 32'b11111111111111110110111101001011;
assign LUT_1[9090] = 32'b11111111111111111001011001100000;
assign LUT_1[9091] = 32'b11111111111111110010101011011100;
assign LUT_1[9092] = 32'b00000000000000000101100100100110;
assign LUT_1[9093] = 32'b11111111111111111110110110100010;
assign LUT_1[9094] = 32'b00000000000000000001010010110111;
assign LUT_1[9095] = 32'b11111111111111111010100100110011;
assign LUT_1[9096] = 32'b11111111111111111100111001000100;
assign LUT_1[9097] = 32'b11111111111111110110001011000000;
assign LUT_1[9098] = 32'b11111111111111111000100111010101;
assign LUT_1[9099] = 32'b11111111111111110001111001010001;
assign LUT_1[9100] = 32'b00000000000000000100110010011011;
assign LUT_1[9101] = 32'b11111111111111111110000100010111;
assign LUT_1[9102] = 32'b00000000000000000000100000101100;
assign LUT_1[9103] = 32'b11111111111111111001110010101000;
assign LUT_1[9104] = 32'b11111111111111111111100110110001;
assign LUT_1[9105] = 32'b11111111111111111000111000101101;
assign LUT_1[9106] = 32'b11111111111111111011010101000010;
assign LUT_1[9107] = 32'b11111111111111110100100110111110;
assign LUT_1[9108] = 32'b00000000000000000111100000001000;
assign LUT_1[9109] = 32'b00000000000000000000110010000100;
assign LUT_1[9110] = 32'b00000000000000000011001110011001;
assign LUT_1[9111] = 32'b11111111111111111100100000010101;
assign LUT_1[9112] = 32'b11111111111111111110110100100110;
assign LUT_1[9113] = 32'b11111111111111111000000110100010;
assign LUT_1[9114] = 32'b11111111111111111010100010110111;
assign LUT_1[9115] = 32'b11111111111111110011110100110011;
assign LUT_1[9116] = 32'b00000000000000000110101101111101;
assign LUT_1[9117] = 32'b11111111111111111111111111111001;
assign LUT_1[9118] = 32'b00000000000000000010011100001110;
assign LUT_1[9119] = 32'b11111111111111111011101110001010;
assign LUT_1[9120] = 32'b11111111111111111110100110001110;
assign LUT_1[9121] = 32'b11111111111111110111111000001010;
assign LUT_1[9122] = 32'b11111111111111111010010100011111;
assign LUT_1[9123] = 32'b11111111111111110011100110011011;
assign LUT_1[9124] = 32'b00000000000000000110011111100101;
assign LUT_1[9125] = 32'b11111111111111111111110001100001;
assign LUT_1[9126] = 32'b00000000000000000010001101110110;
assign LUT_1[9127] = 32'b11111111111111111011011111110010;
assign LUT_1[9128] = 32'b11111111111111111101110100000011;
assign LUT_1[9129] = 32'b11111111111111110111000101111111;
assign LUT_1[9130] = 32'b11111111111111111001100010010100;
assign LUT_1[9131] = 32'b11111111111111110010110100010000;
assign LUT_1[9132] = 32'b00000000000000000101101101011010;
assign LUT_1[9133] = 32'b11111111111111111110111111010110;
assign LUT_1[9134] = 32'b00000000000000000001011011101011;
assign LUT_1[9135] = 32'b11111111111111111010101101100111;
assign LUT_1[9136] = 32'b00000000000000000000100001110000;
assign LUT_1[9137] = 32'b11111111111111111001110011101100;
assign LUT_1[9138] = 32'b11111111111111111100010000000001;
assign LUT_1[9139] = 32'b11111111111111110101100001111101;
assign LUT_1[9140] = 32'b00000000000000001000011011000111;
assign LUT_1[9141] = 32'b00000000000000000001101101000011;
assign LUT_1[9142] = 32'b00000000000000000100001001011000;
assign LUT_1[9143] = 32'b11111111111111111101011011010100;
assign LUT_1[9144] = 32'b11111111111111111111101111100101;
assign LUT_1[9145] = 32'b11111111111111111001000001100001;
assign LUT_1[9146] = 32'b11111111111111111011011101110110;
assign LUT_1[9147] = 32'b11111111111111110100101111110010;
assign LUT_1[9148] = 32'b00000000000000000111101000111100;
assign LUT_1[9149] = 32'b00000000000000000000111010111000;
assign LUT_1[9150] = 32'b00000000000000000011010111001101;
assign LUT_1[9151] = 32'b11111111111111111100101001001001;
assign LUT_1[9152] = 32'b11111111111111111111101000110111;
assign LUT_1[9153] = 32'b11111111111111111000111010110011;
assign LUT_1[9154] = 32'b11111111111111111011010111001000;
assign LUT_1[9155] = 32'b11111111111111110100101001000100;
assign LUT_1[9156] = 32'b00000000000000000111100010001110;
assign LUT_1[9157] = 32'b00000000000000000000110100001010;
assign LUT_1[9158] = 32'b00000000000000000011010000011111;
assign LUT_1[9159] = 32'b11111111111111111100100010011011;
assign LUT_1[9160] = 32'b11111111111111111110110110101100;
assign LUT_1[9161] = 32'b11111111111111111000001000101000;
assign LUT_1[9162] = 32'b11111111111111111010100100111101;
assign LUT_1[9163] = 32'b11111111111111110011110110111001;
assign LUT_1[9164] = 32'b00000000000000000110110000000011;
assign LUT_1[9165] = 32'b00000000000000000000000001111111;
assign LUT_1[9166] = 32'b00000000000000000010011110010100;
assign LUT_1[9167] = 32'b11111111111111111011110000010000;
assign LUT_1[9168] = 32'b00000000000000000001100100011001;
assign LUT_1[9169] = 32'b11111111111111111010110110010101;
assign LUT_1[9170] = 32'b11111111111111111101010010101010;
assign LUT_1[9171] = 32'b11111111111111110110100100100110;
assign LUT_1[9172] = 32'b00000000000000001001011101110000;
assign LUT_1[9173] = 32'b00000000000000000010101111101100;
assign LUT_1[9174] = 32'b00000000000000000101001100000001;
assign LUT_1[9175] = 32'b11111111111111111110011101111101;
assign LUT_1[9176] = 32'b00000000000000000000110010001110;
assign LUT_1[9177] = 32'b11111111111111111010000100001010;
assign LUT_1[9178] = 32'b11111111111111111100100000011111;
assign LUT_1[9179] = 32'b11111111111111110101110010011011;
assign LUT_1[9180] = 32'b00000000000000001000101011100101;
assign LUT_1[9181] = 32'b00000000000000000001111101100001;
assign LUT_1[9182] = 32'b00000000000000000100011001110110;
assign LUT_1[9183] = 32'b11111111111111111101101011110010;
assign LUT_1[9184] = 32'b00000000000000000000100011110110;
assign LUT_1[9185] = 32'b11111111111111111001110101110010;
assign LUT_1[9186] = 32'b11111111111111111100010010000111;
assign LUT_1[9187] = 32'b11111111111111110101100100000011;
assign LUT_1[9188] = 32'b00000000000000001000011101001101;
assign LUT_1[9189] = 32'b00000000000000000001101111001001;
assign LUT_1[9190] = 32'b00000000000000000100001011011110;
assign LUT_1[9191] = 32'b11111111111111111101011101011010;
assign LUT_1[9192] = 32'b11111111111111111111110001101011;
assign LUT_1[9193] = 32'b11111111111111111001000011100111;
assign LUT_1[9194] = 32'b11111111111111111011011111111100;
assign LUT_1[9195] = 32'b11111111111111110100110001111000;
assign LUT_1[9196] = 32'b00000000000000000111101011000010;
assign LUT_1[9197] = 32'b00000000000000000000111100111110;
assign LUT_1[9198] = 32'b00000000000000000011011001010011;
assign LUT_1[9199] = 32'b11111111111111111100101011001111;
assign LUT_1[9200] = 32'b00000000000000000010011111011000;
assign LUT_1[9201] = 32'b11111111111111111011110001010100;
assign LUT_1[9202] = 32'b11111111111111111110001101101001;
assign LUT_1[9203] = 32'b11111111111111110111011111100101;
assign LUT_1[9204] = 32'b00000000000000001010011000101111;
assign LUT_1[9205] = 32'b00000000000000000011101010101011;
assign LUT_1[9206] = 32'b00000000000000000110000111000000;
assign LUT_1[9207] = 32'b11111111111111111111011000111100;
assign LUT_1[9208] = 32'b00000000000000000001101101001101;
assign LUT_1[9209] = 32'b11111111111111111010111111001001;
assign LUT_1[9210] = 32'b11111111111111111101011011011110;
assign LUT_1[9211] = 32'b11111111111111110110101101011010;
assign LUT_1[9212] = 32'b00000000000000001001100110100100;
assign LUT_1[9213] = 32'b00000000000000000010111000100000;
assign LUT_1[9214] = 32'b00000000000000000101010100110101;
assign LUT_1[9215] = 32'b11111111111111111110100110110001;
assign LUT_1[9216] = 32'b00000000000000001001011111010011;
assign LUT_1[9217] = 32'b00000000000000000010110001001111;
assign LUT_1[9218] = 32'b00000000000000000101001101100100;
assign LUT_1[9219] = 32'b11111111111111111110011111100000;
assign LUT_1[9220] = 32'b00000000000000010001011000101010;
assign LUT_1[9221] = 32'b00000000000000001010101010100110;
assign LUT_1[9222] = 32'b00000000000000001101000110111011;
assign LUT_1[9223] = 32'b00000000000000000110011000110111;
assign LUT_1[9224] = 32'b00000000000000001000101101001000;
assign LUT_1[9225] = 32'b00000000000000000001111111000100;
assign LUT_1[9226] = 32'b00000000000000000100011011011001;
assign LUT_1[9227] = 32'b11111111111111111101101101010101;
assign LUT_1[9228] = 32'b00000000000000010000100110011111;
assign LUT_1[9229] = 32'b00000000000000001001111000011011;
assign LUT_1[9230] = 32'b00000000000000001100010100110000;
assign LUT_1[9231] = 32'b00000000000000000101100110101100;
assign LUT_1[9232] = 32'b00000000000000001011011010110101;
assign LUT_1[9233] = 32'b00000000000000000100101100110001;
assign LUT_1[9234] = 32'b00000000000000000111001001000110;
assign LUT_1[9235] = 32'b00000000000000000000011011000010;
assign LUT_1[9236] = 32'b00000000000000010011010100001100;
assign LUT_1[9237] = 32'b00000000000000001100100110001000;
assign LUT_1[9238] = 32'b00000000000000001111000010011101;
assign LUT_1[9239] = 32'b00000000000000001000010100011001;
assign LUT_1[9240] = 32'b00000000000000001010101000101010;
assign LUT_1[9241] = 32'b00000000000000000011111010100110;
assign LUT_1[9242] = 32'b00000000000000000110010110111011;
assign LUT_1[9243] = 32'b11111111111111111111101000110111;
assign LUT_1[9244] = 32'b00000000000000010010100010000001;
assign LUT_1[9245] = 32'b00000000000000001011110011111101;
assign LUT_1[9246] = 32'b00000000000000001110010000010010;
assign LUT_1[9247] = 32'b00000000000000000111100010001110;
assign LUT_1[9248] = 32'b00000000000000001010011010010010;
assign LUT_1[9249] = 32'b00000000000000000011101100001110;
assign LUT_1[9250] = 32'b00000000000000000110001000100011;
assign LUT_1[9251] = 32'b11111111111111111111011010011111;
assign LUT_1[9252] = 32'b00000000000000010010010011101001;
assign LUT_1[9253] = 32'b00000000000000001011100101100101;
assign LUT_1[9254] = 32'b00000000000000001110000001111010;
assign LUT_1[9255] = 32'b00000000000000000111010011110110;
assign LUT_1[9256] = 32'b00000000000000001001101000000111;
assign LUT_1[9257] = 32'b00000000000000000010111010000011;
assign LUT_1[9258] = 32'b00000000000000000101010110011000;
assign LUT_1[9259] = 32'b11111111111111111110101000010100;
assign LUT_1[9260] = 32'b00000000000000010001100001011110;
assign LUT_1[9261] = 32'b00000000000000001010110011011010;
assign LUT_1[9262] = 32'b00000000000000001101001111101111;
assign LUT_1[9263] = 32'b00000000000000000110100001101011;
assign LUT_1[9264] = 32'b00000000000000001100010101110100;
assign LUT_1[9265] = 32'b00000000000000000101100111110000;
assign LUT_1[9266] = 32'b00000000000000001000000100000101;
assign LUT_1[9267] = 32'b00000000000000000001010110000001;
assign LUT_1[9268] = 32'b00000000000000010100001111001011;
assign LUT_1[9269] = 32'b00000000000000001101100001000111;
assign LUT_1[9270] = 32'b00000000000000001111111101011100;
assign LUT_1[9271] = 32'b00000000000000001001001111011000;
assign LUT_1[9272] = 32'b00000000000000001011100011101001;
assign LUT_1[9273] = 32'b00000000000000000100110101100101;
assign LUT_1[9274] = 32'b00000000000000000111010001111010;
assign LUT_1[9275] = 32'b00000000000000000000100011110110;
assign LUT_1[9276] = 32'b00000000000000010011011101000000;
assign LUT_1[9277] = 32'b00000000000000001100101110111100;
assign LUT_1[9278] = 32'b00000000000000001111001011010001;
assign LUT_1[9279] = 32'b00000000000000001000011101001101;
assign LUT_1[9280] = 32'b00000000000000001011011100111011;
assign LUT_1[9281] = 32'b00000000000000000100101110110111;
assign LUT_1[9282] = 32'b00000000000000000111001011001100;
assign LUT_1[9283] = 32'b00000000000000000000011101001000;
assign LUT_1[9284] = 32'b00000000000000010011010110010010;
assign LUT_1[9285] = 32'b00000000000000001100101000001110;
assign LUT_1[9286] = 32'b00000000000000001111000100100011;
assign LUT_1[9287] = 32'b00000000000000001000010110011111;
assign LUT_1[9288] = 32'b00000000000000001010101010110000;
assign LUT_1[9289] = 32'b00000000000000000011111100101100;
assign LUT_1[9290] = 32'b00000000000000000110011001000001;
assign LUT_1[9291] = 32'b11111111111111111111101010111101;
assign LUT_1[9292] = 32'b00000000000000010010100100000111;
assign LUT_1[9293] = 32'b00000000000000001011110110000011;
assign LUT_1[9294] = 32'b00000000000000001110010010011000;
assign LUT_1[9295] = 32'b00000000000000000111100100010100;
assign LUT_1[9296] = 32'b00000000000000001101011000011101;
assign LUT_1[9297] = 32'b00000000000000000110101010011001;
assign LUT_1[9298] = 32'b00000000000000001001000110101110;
assign LUT_1[9299] = 32'b00000000000000000010011000101010;
assign LUT_1[9300] = 32'b00000000000000010101010001110100;
assign LUT_1[9301] = 32'b00000000000000001110100011110000;
assign LUT_1[9302] = 32'b00000000000000010001000000000101;
assign LUT_1[9303] = 32'b00000000000000001010010010000001;
assign LUT_1[9304] = 32'b00000000000000001100100110010010;
assign LUT_1[9305] = 32'b00000000000000000101111000001110;
assign LUT_1[9306] = 32'b00000000000000001000010100100011;
assign LUT_1[9307] = 32'b00000000000000000001100110011111;
assign LUT_1[9308] = 32'b00000000000000010100011111101001;
assign LUT_1[9309] = 32'b00000000000000001101110001100101;
assign LUT_1[9310] = 32'b00000000000000010000001101111010;
assign LUT_1[9311] = 32'b00000000000000001001011111110110;
assign LUT_1[9312] = 32'b00000000000000001100010111111010;
assign LUT_1[9313] = 32'b00000000000000000101101001110110;
assign LUT_1[9314] = 32'b00000000000000001000000110001011;
assign LUT_1[9315] = 32'b00000000000000000001011000000111;
assign LUT_1[9316] = 32'b00000000000000010100010001010001;
assign LUT_1[9317] = 32'b00000000000000001101100011001101;
assign LUT_1[9318] = 32'b00000000000000001111111111100010;
assign LUT_1[9319] = 32'b00000000000000001001010001011110;
assign LUT_1[9320] = 32'b00000000000000001011100101101111;
assign LUT_1[9321] = 32'b00000000000000000100110111101011;
assign LUT_1[9322] = 32'b00000000000000000111010100000000;
assign LUT_1[9323] = 32'b00000000000000000000100101111100;
assign LUT_1[9324] = 32'b00000000000000010011011111000110;
assign LUT_1[9325] = 32'b00000000000000001100110001000010;
assign LUT_1[9326] = 32'b00000000000000001111001101010111;
assign LUT_1[9327] = 32'b00000000000000001000011111010011;
assign LUT_1[9328] = 32'b00000000000000001110010011011100;
assign LUT_1[9329] = 32'b00000000000000000111100101011000;
assign LUT_1[9330] = 32'b00000000000000001010000001101101;
assign LUT_1[9331] = 32'b00000000000000000011010011101001;
assign LUT_1[9332] = 32'b00000000000000010110001100110011;
assign LUT_1[9333] = 32'b00000000000000001111011110101111;
assign LUT_1[9334] = 32'b00000000000000010001111011000100;
assign LUT_1[9335] = 32'b00000000000000001011001101000000;
assign LUT_1[9336] = 32'b00000000000000001101100001010001;
assign LUT_1[9337] = 32'b00000000000000000110110011001101;
assign LUT_1[9338] = 32'b00000000000000001001001111100010;
assign LUT_1[9339] = 32'b00000000000000000010100001011110;
assign LUT_1[9340] = 32'b00000000000000010101011010101000;
assign LUT_1[9341] = 32'b00000000000000001110101100100100;
assign LUT_1[9342] = 32'b00000000000000010001001000111001;
assign LUT_1[9343] = 32'b00000000000000001010011010110101;
assign LUT_1[9344] = 32'b00000000000000001100011111010110;
assign LUT_1[9345] = 32'b00000000000000000101110001010010;
assign LUT_1[9346] = 32'b00000000000000001000001101100111;
assign LUT_1[9347] = 32'b00000000000000000001011111100011;
assign LUT_1[9348] = 32'b00000000000000010100011000101101;
assign LUT_1[9349] = 32'b00000000000000001101101010101001;
assign LUT_1[9350] = 32'b00000000000000010000000110111110;
assign LUT_1[9351] = 32'b00000000000000001001011000111010;
assign LUT_1[9352] = 32'b00000000000000001011101101001011;
assign LUT_1[9353] = 32'b00000000000000000100111111000111;
assign LUT_1[9354] = 32'b00000000000000000111011011011100;
assign LUT_1[9355] = 32'b00000000000000000000101101011000;
assign LUT_1[9356] = 32'b00000000000000010011100110100010;
assign LUT_1[9357] = 32'b00000000000000001100111000011110;
assign LUT_1[9358] = 32'b00000000000000001111010100110011;
assign LUT_1[9359] = 32'b00000000000000001000100110101111;
assign LUT_1[9360] = 32'b00000000000000001110011010111000;
assign LUT_1[9361] = 32'b00000000000000000111101100110100;
assign LUT_1[9362] = 32'b00000000000000001010001001001001;
assign LUT_1[9363] = 32'b00000000000000000011011011000101;
assign LUT_1[9364] = 32'b00000000000000010110010100001111;
assign LUT_1[9365] = 32'b00000000000000001111100110001011;
assign LUT_1[9366] = 32'b00000000000000010010000010100000;
assign LUT_1[9367] = 32'b00000000000000001011010100011100;
assign LUT_1[9368] = 32'b00000000000000001101101000101101;
assign LUT_1[9369] = 32'b00000000000000000110111010101001;
assign LUT_1[9370] = 32'b00000000000000001001010110111110;
assign LUT_1[9371] = 32'b00000000000000000010101000111010;
assign LUT_1[9372] = 32'b00000000000000010101100010000100;
assign LUT_1[9373] = 32'b00000000000000001110110100000000;
assign LUT_1[9374] = 32'b00000000000000010001010000010101;
assign LUT_1[9375] = 32'b00000000000000001010100010010001;
assign LUT_1[9376] = 32'b00000000000000001101011010010101;
assign LUT_1[9377] = 32'b00000000000000000110101100010001;
assign LUT_1[9378] = 32'b00000000000000001001001000100110;
assign LUT_1[9379] = 32'b00000000000000000010011010100010;
assign LUT_1[9380] = 32'b00000000000000010101010011101100;
assign LUT_1[9381] = 32'b00000000000000001110100101101000;
assign LUT_1[9382] = 32'b00000000000000010001000001111101;
assign LUT_1[9383] = 32'b00000000000000001010010011111001;
assign LUT_1[9384] = 32'b00000000000000001100101000001010;
assign LUT_1[9385] = 32'b00000000000000000101111010000110;
assign LUT_1[9386] = 32'b00000000000000001000010110011011;
assign LUT_1[9387] = 32'b00000000000000000001101000010111;
assign LUT_1[9388] = 32'b00000000000000010100100001100001;
assign LUT_1[9389] = 32'b00000000000000001101110011011101;
assign LUT_1[9390] = 32'b00000000000000010000001111110010;
assign LUT_1[9391] = 32'b00000000000000001001100001101110;
assign LUT_1[9392] = 32'b00000000000000001111010101110111;
assign LUT_1[9393] = 32'b00000000000000001000100111110011;
assign LUT_1[9394] = 32'b00000000000000001011000100001000;
assign LUT_1[9395] = 32'b00000000000000000100010110000100;
assign LUT_1[9396] = 32'b00000000000000010111001111001110;
assign LUT_1[9397] = 32'b00000000000000010000100001001010;
assign LUT_1[9398] = 32'b00000000000000010010111101011111;
assign LUT_1[9399] = 32'b00000000000000001100001111011011;
assign LUT_1[9400] = 32'b00000000000000001110100011101100;
assign LUT_1[9401] = 32'b00000000000000000111110101101000;
assign LUT_1[9402] = 32'b00000000000000001010010001111101;
assign LUT_1[9403] = 32'b00000000000000000011100011111001;
assign LUT_1[9404] = 32'b00000000000000010110011101000011;
assign LUT_1[9405] = 32'b00000000000000001111101110111111;
assign LUT_1[9406] = 32'b00000000000000010010001011010100;
assign LUT_1[9407] = 32'b00000000000000001011011101010000;
assign LUT_1[9408] = 32'b00000000000000001110011100111110;
assign LUT_1[9409] = 32'b00000000000000000111101110111010;
assign LUT_1[9410] = 32'b00000000000000001010001011001111;
assign LUT_1[9411] = 32'b00000000000000000011011101001011;
assign LUT_1[9412] = 32'b00000000000000010110010110010101;
assign LUT_1[9413] = 32'b00000000000000001111101000010001;
assign LUT_1[9414] = 32'b00000000000000010010000100100110;
assign LUT_1[9415] = 32'b00000000000000001011010110100010;
assign LUT_1[9416] = 32'b00000000000000001101101010110011;
assign LUT_1[9417] = 32'b00000000000000000110111100101111;
assign LUT_1[9418] = 32'b00000000000000001001011001000100;
assign LUT_1[9419] = 32'b00000000000000000010101011000000;
assign LUT_1[9420] = 32'b00000000000000010101100100001010;
assign LUT_1[9421] = 32'b00000000000000001110110110000110;
assign LUT_1[9422] = 32'b00000000000000010001010010011011;
assign LUT_1[9423] = 32'b00000000000000001010100100010111;
assign LUT_1[9424] = 32'b00000000000000010000011000100000;
assign LUT_1[9425] = 32'b00000000000000001001101010011100;
assign LUT_1[9426] = 32'b00000000000000001100000110110001;
assign LUT_1[9427] = 32'b00000000000000000101011000101101;
assign LUT_1[9428] = 32'b00000000000000011000010001110111;
assign LUT_1[9429] = 32'b00000000000000010001100011110011;
assign LUT_1[9430] = 32'b00000000000000010100000000001000;
assign LUT_1[9431] = 32'b00000000000000001101010010000100;
assign LUT_1[9432] = 32'b00000000000000001111100110010101;
assign LUT_1[9433] = 32'b00000000000000001000111000010001;
assign LUT_1[9434] = 32'b00000000000000001011010100100110;
assign LUT_1[9435] = 32'b00000000000000000100100110100010;
assign LUT_1[9436] = 32'b00000000000000010111011111101100;
assign LUT_1[9437] = 32'b00000000000000010000110001101000;
assign LUT_1[9438] = 32'b00000000000000010011001101111101;
assign LUT_1[9439] = 32'b00000000000000001100011111111001;
assign LUT_1[9440] = 32'b00000000000000001111010111111101;
assign LUT_1[9441] = 32'b00000000000000001000101001111001;
assign LUT_1[9442] = 32'b00000000000000001011000110001110;
assign LUT_1[9443] = 32'b00000000000000000100011000001010;
assign LUT_1[9444] = 32'b00000000000000010111010001010100;
assign LUT_1[9445] = 32'b00000000000000010000100011010000;
assign LUT_1[9446] = 32'b00000000000000010010111111100101;
assign LUT_1[9447] = 32'b00000000000000001100010001100001;
assign LUT_1[9448] = 32'b00000000000000001110100101110010;
assign LUT_1[9449] = 32'b00000000000000000111110111101110;
assign LUT_1[9450] = 32'b00000000000000001010010100000011;
assign LUT_1[9451] = 32'b00000000000000000011100101111111;
assign LUT_1[9452] = 32'b00000000000000010110011111001001;
assign LUT_1[9453] = 32'b00000000000000001111110001000101;
assign LUT_1[9454] = 32'b00000000000000010010001101011010;
assign LUT_1[9455] = 32'b00000000000000001011011111010110;
assign LUT_1[9456] = 32'b00000000000000010001010011011111;
assign LUT_1[9457] = 32'b00000000000000001010100101011011;
assign LUT_1[9458] = 32'b00000000000000001101000001110000;
assign LUT_1[9459] = 32'b00000000000000000110010011101100;
assign LUT_1[9460] = 32'b00000000000000011001001100110110;
assign LUT_1[9461] = 32'b00000000000000010010011110110010;
assign LUT_1[9462] = 32'b00000000000000010100111011000111;
assign LUT_1[9463] = 32'b00000000000000001110001101000011;
assign LUT_1[9464] = 32'b00000000000000010000100001010100;
assign LUT_1[9465] = 32'b00000000000000001001110011010000;
assign LUT_1[9466] = 32'b00000000000000001100001111100101;
assign LUT_1[9467] = 32'b00000000000000000101100001100001;
assign LUT_1[9468] = 32'b00000000000000011000011010101011;
assign LUT_1[9469] = 32'b00000000000000010001101100100111;
assign LUT_1[9470] = 32'b00000000000000010100001000111100;
assign LUT_1[9471] = 32'b00000000000000001101011010111000;
assign LUT_1[9472] = 32'b00000000000000000111010011011111;
assign LUT_1[9473] = 32'b00000000000000000000100101011011;
assign LUT_1[9474] = 32'b00000000000000000011000001110000;
assign LUT_1[9475] = 32'b11111111111111111100010011101100;
assign LUT_1[9476] = 32'b00000000000000001111001100110110;
assign LUT_1[9477] = 32'b00000000000000001000011110110010;
assign LUT_1[9478] = 32'b00000000000000001010111011000111;
assign LUT_1[9479] = 32'b00000000000000000100001101000011;
assign LUT_1[9480] = 32'b00000000000000000110100001010100;
assign LUT_1[9481] = 32'b11111111111111111111110011010000;
assign LUT_1[9482] = 32'b00000000000000000010001111100101;
assign LUT_1[9483] = 32'b11111111111111111011100001100001;
assign LUT_1[9484] = 32'b00000000000000001110011010101011;
assign LUT_1[9485] = 32'b00000000000000000111101100100111;
assign LUT_1[9486] = 32'b00000000000000001010001000111100;
assign LUT_1[9487] = 32'b00000000000000000011011010111000;
assign LUT_1[9488] = 32'b00000000000000001001001111000001;
assign LUT_1[9489] = 32'b00000000000000000010100000111101;
assign LUT_1[9490] = 32'b00000000000000000100111101010010;
assign LUT_1[9491] = 32'b11111111111111111110001111001110;
assign LUT_1[9492] = 32'b00000000000000010001001000011000;
assign LUT_1[9493] = 32'b00000000000000001010011010010100;
assign LUT_1[9494] = 32'b00000000000000001100110110101001;
assign LUT_1[9495] = 32'b00000000000000000110001000100101;
assign LUT_1[9496] = 32'b00000000000000001000011100110110;
assign LUT_1[9497] = 32'b00000000000000000001101110110010;
assign LUT_1[9498] = 32'b00000000000000000100001011000111;
assign LUT_1[9499] = 32'b11111111111111111101011101000011;
assign LUT_1[9500] = 32'b00000000000000010000010110001101;
assign LUT_1[9501] = 32'b00000000000000001001101000001001;
assign LUT_1[9502] = 32'b00000000000000001100000100011110;
assign LUT_1[9503] = 32'b00000000000000000101010110011010;
assign LUT_1[9504] = 32'b00000000000000001000001110011110;
assign LUT_1[9505] = 32'b00000000000000000001100000011010;
assign LUT_1[9506] = 32'b00000000000000000011111100101111;
assign LUT_1[9507] = 32'b11111111111111111101001110101011;
assign LUT_1[9508] = 32'b00000000000000010000000111110101;
assign LUT_1[9509] = 32'b00000000000000001001011001110001;
assign LUT_1[9510] = 32'b00000000000000001011110110000110;
assign LUT_1[9511] = 32'b00000000000000000101001000000010;
assign LUT_1[9512] = 32'b00000000000000000111011100010011;
assign LUT_1[9513] = 32'b00000000000000000000101110001111;
assign LUT_1[9514] = 32'b00000000000000000011001010100100;
assign LUT_1[9515] = 32'b11111111111111111100011100100000;
assign LUT_1[9516] = 32'b00000000000000001111010101101010;
assign LUT_1[9517] = 32'b00000000000000001000100111100110;
assign LUT_1[9518] = 32'b00000000000000001011000011111011;
assign LUT_1[9519] = 32'b00000000000000000100010101110111;
assign LUT_1[9520] = 32'b00000000000000001010001010000000;
assign LUT_1[9521] = 32'b00000000000000000011011011111100;
assign LUT_1[9522] = 32'b00000000000000000101111000010001;
assign LUT_1[9523] = 32'b11111111111111111111001010001101;
assign LUT_1[9524] = 32'b00000000000000010010000011010111;
assign LUT_1[9525] = 32'b00000000000000001011010101010011;
assign LUT_1[9526] = 32'b00000000000000001101110001101000;
assign LUT_1[9527] = 32'b00000000000000000111000011100100;
assign LUT_1[9528] = 32'b00000000000000001001010111110101;
assign LUT_1[9529] = 32'b00000000000000000010101001110001;
assign LUT_1[9530] = 32'b00000000000000000101000110000110;
assign LUT_1[9531] = 32'b11111111111111111110011000000010;
assign LUT_1[9532] = 32'b00000000000000010001010001001100;
assign LUT_1[9533] = 32'b00000000000000001010100011001000;
assign LUT_1[9534] = 32'b00000000000000001100111111011101;
assign LUT_1[9535] = 32'b00000000000000000110010001011001;
assign LUT_1[9536] = 32'b00000000000000001001010001000111;
assign LUT_1[9537] = 32'b00000000000000000010100011000011;
assign LUT_1[9538] = 32'b00000000000000000100111111011000;
assign LUT_1[9539] = 32'b11111111111111111110010001010100;
assign LUT_1[9540] = 32'b00000000000000010001001010011110;
assign LUT_1[9541] = 32'b00000000000000001010011100011010;
assign LUT_1[9542] = 32'b00000000000000001100111000101111;
assign LUT_1[9543] = 32'b00000000000000000110001010101011;
assign LUT_1[9544] = 32'b00000000000000001000011110111100;
assign LUT_1[9545] = 32'b00000000000000000001110000111000;
assign LUT_1[9546] = 32'b00000000000000000100001101001101;
assign LUT_1[9547] = 32'b11111111111111111101011111001001;
assign LUT_1[9548] = 32'b00000000000000010000011000010011;
assign LUT_1[9549] = 32'b00000000000000001001101010001111;
assign LUT_1[9550] = 32'b00000000000000001100000110100100;
assign LUT_1[9551] = 32'b00000000000000000101011000100000;
assign LUT_1[9552] = 32'b00000000000000001011001100101001;
assign LUT_1[9553] = 32'b00000000000000000100011110100101;
assign LUT_1[9554] = 32'b00000000000000000110111010111010;
assign LUT_1[9555] = 32'b00000000000000000000001100110110;
assign LUT_1[9556] = 32'b00000000000000010011000110000000;
assign LUT_1[9557] = 32'b00000000000000001100010111111100;
assign LUT_1[9558] = 32'b00000000000000001110110100010001;
assign LUT_1[9559] = 32'b00000000000000001000000110001101;
assign LUT_1[9560] = 32'b00000000000000001010011010011110;
assign LUT_1[9561] = 32'b00000000000000000011101100011010;
assign LUT_1[9562] = 32'b00000000000000000110001000101111;
assign LUT_1[9563] = 32'b11111111111111111111011010101011;
assign LUT_1[9564] = 32'b00000000000000010010010011110101;
assign LUT_1[9565] = 32'b00000000000000001011100101110001;
assign LUT_1[9566] = 32'b00000000000000001110000010000110;
assign LUT_1[9567] = 32'b00000000000000000111010100000010;
assign LUT_1[9568] = 32'b00000000000000001010001100000110;
assign LUT_1[9569] = 32'b00000000000000000011011110000010;
assign LUT_1[9570] = 32'b00000000000000000101111010010111;
assign LUT_1[9571] = 32'b11111111111111111111001100010011;
assign LUT_1[9572] = 32'b00000000000000010010000101011101;
assign LUT_1[9573] = 32'b00000000000000001011010111011001;
assign LUT_1[9574] = 32'b00000000000000001101110011101110;
assign LUT_1[9575] = 32'b00000000000000000111000101101010;
assign LUT_1[9576] = 32'b00000000000000001001011001111011;
assign LUT_1[9577] = 32'b00000000000000000010101011110111;
assign LUT_1[9578] = 32'b00000000000000000101001000001100;
assign LUT_1[9579] = 32'b11111111111111111110011010001000;
assign LUT_1[9580] = 32'b00000000000000010001010011010010;
assign LUT_1[9581] = 32'b00000000000000001010100101001110;
assign LUT_1[9582] = 32'b00000000000000001101000001100011;
assign LUT_1[9583] = 32'b00000000000000000110010011011111;
assign LUT_1[9584] = 32'b00000000000000001100000111101000;
assign LUT_1[9585] = 32'b00000000000000000101011001100100;
assign LUT_1[9586] = 32'b00000000000000000111110101111001;
assign LUT_1[9587] = 32'b00000000000000000001000111110101;
assign LUT_1[9588] = 32'b00000000000000010100000000111111;
assign LUT_1[9589] = 32'b00000000000000001101010010111011;
assign LUT_1[9590] = 32'b00000000000000001111101111010000;
assign LUT_1[9591] = 32'b00000000000000001001000001001100;
assign LUT_1[9592] = 32'b00000000000000001011010101011101;
assign LUT_1[9593] = 32'b00000000000000000100100111011001;
assign LUT_1[9594] = 32'b00000000000000000111000011101110;
assign LUT_1[9595] = 32'b00000000000000000000010101101010;
assign LUT_1[9596] = 32'b00000000000000010011001110110100;
assign LUT_1[9597] = 32'b00000000000000001100100000110000;
assign LUT_1[9598] = 32'b00000000000000001110111101000101;
assign LUT_1[9599] = 32'b00000000000000001000001111000001;
assign LUT_1[9600] = 32'b00000000000000001010010011100010;
assign LUT_1[9601] = 32'b00000000000000000011100101011110;
assign LUT_1[9602] = 32'b00000000000000000110000001110011;
assign LUT_1[9603] = 32'b11111111111111111111010011101111;
assign LUT_1[9604] = 32'b00000000000000010010001100111001;
assign LUT_1[9605] = 32'b00000000000000001011011110110101;
assign LUT_1[9606] = 32'b00000000000000001101111011001010;
assign LUT_1[9607] = 32'b00000000000000000111001101000110;
assign LUT_1[9608] = 32'b00000000000000001001100001010111;
assign LUT_1[9609] = 32'b00000000000000000010110011010011;
assign LUT_1[9610] = 32'b00000000000000000101001111101000;
assign LUT_1[9611] = 32'b11111111111111111110100001100100;
assign LUT_1[9612] = 32'b00000000000000010001011010101110;
assign LUT_1[9613] = 32'b00000000000000001010101100101010;
assign LUT_1[9614] = 32'b00000000000000001101001000111111;
assign LUT_1[9615] = 32'b00000000000000000110011010111011;
assign LUT_1[9616] = 32'b00000000000000001100001111000100;
assign LUT_1[9617] = 32'b00000000000000000101100001000000;
assign LUT_1[9618] = 32'b00000000000000000111111101010101;
assign LUT_1[9619] = 32'b00000000000000000001001111010001;
assign LUT_1[9620] = 32'b00000000000000010100001000011011;
assign LUT_1[9621] = 32'b00000000000000001101011010010111;
assign LUT_1[9622] = 32'b00000000000000001111110110101100;
assign LUT_1[9623] = 32'b00000000000000001001001000101000;
assign LUT_1[9624] = 32'b00000000000000001011011100111001;
assign LUT_1[9625] = 32'b00000000000000000100101110110101;
assign LUT_1[9626] = 32'b00000000000000000111001011001010;
assign LUT_1[9627] = 32'b00000000000000000000011101000110;
assign LUT_1[9628] = 32'b00000000000000010011010110010000;
assign LUT_1[9629] = 32'b00000000000000001100101000001100;
assign LUT_1[9630] = 32'b00000000000000001111000100100001;
assign LUT_1[9631] = 32'b00000000000000001000010110011101;
assign LUT_1[9632] = 32'b00000000000000001011001110100001;
assign LUT_1[9633] = 32'b00000000000000000100100000011101;
assign LUT_1[9634] = 32'b00000000000000000110111100110010;
assign LUT_1[9635] = 32'b00000000000000000000001110101110;
assign LUT_1[9636] = 32'b00000000000000010011000111111000;
assign LUT_1[9637] = 32'b00000000000000001100011001110100;
assign LUT_1[9638] = 32'b00000000000000001110110110001001;
assign LUT_1[9639] = 32'b00000000000000001000001000000101;
assign LUT_1[9640] = 32'b00000000000000001010011100010110;
assign LUT_1[9641] = 32'b00000000000000000011101110010010;
assign LUT_1[9642] = 32'b00000000000000000110001010100111;
assign LUT_1[9643] = 32'b11111111111111111111011100100011;
assign LUT_1[9644] = 32'b00000000000000010010010101101101;
assign LUT_1[9645] = 32'b00000000000000001011100111101001;
assign LUT_1[9646] = 32'b00000000000000001110000011111110;
assign LUT_1[9647] = 32'b00000000000000000111010101111010;
assign LUT_1[9648] = 32'b00000000000000001101001010000011;
assign LUT_1[9649] = 32'b00000000000000000110011011111111;
assign LUT_1[9650] = 32'b00000000000000001000111000010100;
assign LUT_1[9651] = 32'b00000000000000000010001010010000;
assign LUT_1[9652] = 32'b00000000000000010101000011011010;
assign LUT_1[9653] = 32'b00000000000000001110010101010110;
assign LUT_1[9654] = 32'b00000000000000010000110001101011;
assign LUT_1[9655] = 32'b00000000000000001010000011100111;
assign LUT_1[9656] = 32'b00000000000000001100010111111000;
assign LUT_1[9657] = 32'b00000000000000000101101001110100;
assign LUT_1[9658] = 32'b00000000000000001000000110001001;
assign LUT_1[9659] = 32'b00000000000000000001011000000101;
assign LUT_1[9660] = 32'b00000000000000010100010001001111;
assign LUT_1[9661] = 32'b00000000000000001101100011001011;
assign LUT_1[9662] = 32'b00000000000000001111111111100000;
assign LUT_1[9663] = 32'b00000000000000001001010001011100;
assign LUT_1[9664] = 32'b00000000000000001100010001001010;
assign LUT_1[9665] = 32'b00000000000000000101100011000110;
assign LUT_1[9666] = 32'b00000000000000000111111111011011;
assign LUT_1[9667] = 32'b00000000000000000001010001010111;
assign LUT_1[9668] = 32'b00000000000000010100001010100001;
assign LUT_1[9669] = 32'b00000000000000001101011100011101;
assign LUT_1[9670] = 32'b00000000000000001111111000110010;
assign LUT_1[9671] = 32'b00000000000000001001001010101110;
assign LUT_1[9672] = 32'b00000000000000001011011110111111;
assign LUT_1[9673] = 32'b00000000000000000100110000111011;
assign LUT_1[9674] = 32'b00000000000000000111001101010000;
assign LUT_1[9675] = 32'b00000000000000000000011111001100;
assign LUT_1[9676] = 32'b00000000000000010011011000010110;
assign LUT_1[9677] = 32'b00000000000000001100101010010010;
assign LUT_1[9678] = 32'b00000000000000001111000110100111;
assign LUT_1[9679] = 32'b00000000000000001000011000100011;
assign LUT_1[9680] = 32'b00000000000000001110001100101100;
assign LUT_1[9681] = 32'b00000000000000000111011110101000;
assign LUT_1[9682] = 32'b00000000000000001001111010111101;
assign LUT_1[9683] = 32'b00000000000000000011001100111001;
assign LUT_1[9684] = 32'b00000000000000010110000110000011;
assign LUT_1[9685] = 32'b00000000000000001111010111111111;
assign LUT_1[9686] = 32'b00000000000000010001110100010100;
assign LUT_1[9687] = 32'b00000000000000001011000110010000;
assign LUT_1[9688] = 32'b00000000000000001101011010100001;
assign LUT_1[9689] = 32'b00000000000000000110101100011101;
assign LUT_1[9690] = 32'b00000000000000001001001000110010;
assign LUT_1[9691] = 32'b00000000000000000010011010101110;
assign LUT_1[9692] = 32'b00000000000000010101010011111000;
assign LUT_1[9693] = 32'b00000000000000001110100101110100;
assign LUT_1[9694] = 32'b00000000000000010001000010001001;
assign LUT_1[9695] = 32'b00000000000000001010010100000101;
assign LUT_1[9696] = 32'b00000000000000001101001100001001;
assign LUT_1[9697] = 32'b00000000000000000110011110000101;
assign LUT_1[9698] = 32'b00000000000000001000111010011010;
assign LUT_1[9699] = 32'b00000000000000000010001100010110;
assign LUT_1[9700] = 32'b00000000000000010101000101100000;
assign LUT_1[9701] = 32'b00000000000000001110010111011100;
assign LUT_1[9702] = 32'b00000000000000010000110011110001;
assign LUT_1[9703] = 32'b00000000000000001010000101101101;
assign LUT_1[9704] = 32'b00000000000000001100011001111110;
assign LUT_1[9705] = 32'b00000000000000000101101011111010;
assign LUT_1[9706] = 32'b00000000000000001000001000001111;
assign LUT_1[9707] = 32'b00000000000000000001011010001011;
assign LUT_1[9708] = 32'b00000000000000010100010011010101;
assign LUT_1[9709] = 32'b00000000000000001101100101010001;
assign LUT_1[9710] = 32'b00000000000000010000000001100110;
assign LUT_1[9711] = 32'b00000000000000001001010011100010;
assign LUT_1[9712] = 32'b00000000000000001111000111101011;
assign LUT_1[9713] = 32'b00000000000000001000011001100111;
assign LUT_1[9714] = 32'b00000000000000001010110101111100;
assign LUT_1[9715] = 32'b00000000000000000100000111111000;
assign LUT_1[9716] = 32'b00000000000000010111000001000010;
assign LUT_1[9717] = 32'b00000000000000010000010010111110;
assign LUT_1[9718] = 32'b00000000000000010010101111010011;
assign LUT_1[9719] = 32'b00000000000000001100000001001111;
assign LUT_1[9720] = 32'b00000000000000001110010101100000;
assign LUT_1[9721] = 32'b00000000000000000111100111011100;
assign LUT_1[9722] = 32'b00000000000000001010000011110001;
assign LUT_1[9723] = 32'b00000000000000000011010101101101;
assign LUT_1[9724] = 32'b00000000000000010110001110110111;
assign LUT_1[9725] = 32'b00000000000000001111100000110011;
assign LUT_1[9726] = 32'b00000000000000010001111101001000;
assign LUT_1[9727] = 32'b00000000000000001011001111000100;
assign LUT_1[9728] = 32'b00000000000000000011001101110000;
assign LUT_1[9729] = 32'b11111111111111111100011111101100;
assign LUT_1[9730] = 32'b11111111111111111110111100000001;
assign LUT_1[9731] = 32'b11111111111111111000001101111101;
assign LUT_1[9732] = 32'b00000000000000001011000111000111;
assign LUT_1[9733] = 32'b00000000000000000100011001000011;
assign LUT_1[9734] = 32'b00000000000000000110110101011000;
assign LUT_1[9735] = 32'b00000000000000000000000111010100;
assign LUT_1[9736] = 32'b00000000000000000010011011100101;
assign LUT_1[9737] = 32'b11111111111111111011101101100001;
assign LUT_1[9738] = 32'b11111111111111111110001001110110;
assign LUT_1[9739] = 32'b11111111111111110111011011110010;
assign LUT_1[9740] = 32'b00000000000000001010010100111100;
assign LUT_1[9741] = 32'b00000000000000000011100110111000;
assign LUT_1[9742] = 32'b00000000000000000110000011001101;
assign LUT_1[9743] = 32'b11111111111111111111010101001001;
assign LUT_1[9744] = 32'b00000000000000000101001001010010;
assign LUT_1[9745] = 32'b11111111111111111110011011001110;
assign LUT_1[9746] = 32'b00000000000000000000110111100011;
assign LUT_1[9747] = 32'b11111111111111111010001001011111;
assign LUT_1[9748] = 32'b00000000000000001101000010101001;
assign LUT_1[9749] = 32'b00000000000000000110010100100101;
assign LUT_1[9750] = 32'b00000000000000001000110000111010;
assign LUT_1[9751] = 32'b00000000000000000010000010110110;
assign LUT_1[9752] = 32'b00000000000000000100010111000111;
assign LUT_1[9753] = 32'b11111111111111111101101001000011;
assign LUT_1[9754] = 32'b00000000000000000000000101011000;
assign LUT_1[9755] = 32'b11111111111111111001010111010100;
assign LUT_1[9756] = 32'b00000000000000001100010000011110;
assign LUT_1[9757] = 32'b00000000000000000101100010011010;
assign LUT_1[9758] = 32'b00000000000000000111111110101111;
assign LUT_1[9759] = 32'b00000000000000000001010000101011;
assign LUT_1[9760] = 32'b00000000000000000100001000101111;
assign LUT_1[9761] = 32'b11111111111111111101011010101011;
assign LUT_1[9762] = 32'b11111111111111111111110111000000;
assign LUT_1[9763] = 32'b11111111111111111001001000111100;
assign LUT_1[9764] = 32'b00000000000000001100000010000110;
assign LUT_1[9765] = 32'b00000000000000000101010100000010;
assign LUT_1[9766] = 32'b00000000000000000111110000010111;
assign LUT_1[9767] = 32'b00000000000000000001000010010011;
assign LUT_1[9768] = 32'b00000000000000000011010110100100;
assign LUT_1[9769] = 32'b11111111111111111100101000100000;
assign LUT_1[9770] = 32'b11111111111111111111000100110101;
assign LUT_1[9771] = 32'b11111111111111111000010110110001;
assign LUT_1[9772] = 32'b00000000000000001011001111111011;
assign LUT_1[9773] = 32'b00000000000000000100100001110111;
assign LUT_1[9774] = 32'b00000000000000000110111110001100;
assign LUT_1[9775] = 32'b00000000000000000000010000001000;
assign LUT_1[9776] = 32'b00000000000000000110000100010001;
assign LUT_1[9777] = 32'b11111111111111111111010110001101;
assign LUT_1[9778] = 32'b00000000000000000001110010100010;
assign LUT_1[9779] = 32'b11111111111111111011000100011110;
assign LUT_1[9780] = 32'b00000000000000001101111101101000;
assign LUT_1[9781] = 32'b00000000000000000111001111100100;
assign LUT_1[9782] = 32'b00000000000000001001101011111001;
assign LUT_1[9783] = 32'b00000000000000000010111101110101;
assign LUT_1[9784] = 32'b00000000000000000101010010000110;
assign LUT_1[9785] = 32'b11111111111111111110100100000010;
assign LUT_1[9786] = 32'b00000000000000000001000000010111;
assign LUT_1[9787] = 32'b11111111111111111010010010010011;
assign LUT_1[9788] = 32'b00000000000000001101001011011101;
assign LUT_1[9789] = 32'b00000000000000000110011101011001;
assign LUT_1[9790] = 32'b00000000000000001000111001101110;
assign LUT_1[9791] = 32'b00000000000000000010001011101010;
assign LUT_1[9792] = 32'b00000000000000000101001011011000;
assign LUT_1[9793] = 32'b11111111111111111110011101010100;
assign LUT_1[9794] = 32'b00000000000000000000111001101001;
assign LUT_1[9795] = 32'b11111111111111111010001011100101;
assign LUT_1[9796] = 32'b00000000000000001101000100101111;
assign LUT_1[9797] = 32'b00000000000000000110010110101011;
assign LUT_1[9798] = 32'b00000000000000001000110011000000;
assign LUT_1[9799] = 32'b00000000000000000010000100111100;
assign LUT_1[9800] = 32'b00000000000000000100011001001101;
assign LUT_1[9801] = 32'b11111111111111111101101011001001;
assign LUT_1[9802] = 32'b00000000000000000000000111011110;
assign LUT_1[9803] = 32'b11111111111111111001011001011010;
assign LUT_1[9804] = 32'b00000000000000001100010010100100;
assign LUT_1[9805] = 32'b00000000000000000101100100100000;
assign LUT_1[9806] = 32'b00000000000000001000000000110101;
assign LUT_1[9807] = 32'b00000000000000000001010010110001;
assign LUT_1[9808] = 32'b00000000000000000111000110111010;
assign LUT_1[9809] = 32'b00000000000000000000011000110110;
assign LUT_1[9810] = 32'b00000000000000000010110101001011;
assign LUT_1[9811] = 32'b11111111111111111100000111000111;
assign LUT_1[9812] = 32'b00000000000000001111000000010001;
assign LUT_1[9813] = 32'b00000000000000001000010010001101;
assign LUT_1[9814] = 32'b00000000000000001010101110100010;
assign LUT_1[9815] = 32'b00000000000000000100000000011110;
assign LUT_1[9816] = 32'b00000000000000000110010100101111;
assign LUT_1[9817] = 32'b11111111111111111111100110101011;
assign LUT_1[9818] = 32'b00000000000000000010000011000000;
assign LUT_1[9819] = 32'b11111111111111111011010100111100;
assign LUT_1[9820] = 32'b00000000000000001110001110000110;
assign LUT_1[9821] = 32'b00000000000000000111100000000010;
assign LUT_1[9822] = 32'b00000000000000001001111100010111;
assign LUT_1[9823] = 32'b00000000000000000011001110010011;
assign LUT_1[9824] = 32'b00000000000000000110000110010111;
assign LUT_1[9825] = 32'b11111111111111111111011000010011;
assign LUT_1[9826] = 32'b00000000000000000001110100101000;
assign LUT_1[9827] = 32'b11111111111111111011000110100100;
assign LUT_1[9828] = 32'b00000000000000001101111111101110;
assign LUT_1[9829] = 32'b00000000000000000111010001101010;
assign LUT_1[9830] = 32'b00000000000000001001101101111111;
assign LUT_1[9831] = 32'b00000000000000000010111111111011;
assign LUT_1[9832] = 32'b00000000000000000101010100001100;
assign LUT_1[9833] = 32'b11111111111111111110100110001000;
assign LUT_1[9834] = 32'b00000000000000000001000010011101;
assign LUT_1[9835] = 32'b11111111111111111010010100011001;
assign LUT_1[9836] = 32'b00000000000000001101001101100011;
assign LUT_1[9837] = 32'b00000000000000000110011111011111;
assign LUT_1[9838] = 32'b00000000000000001000111011110100;
assign LUT_1[9839] = 32'b00000000000000000010001101110000;
assign LUT_1[9840] = 32'b00000000000000001000000001111001;
assign LUT_1[9841] = 32'b00000000000000000001010011110101;
assign LUT_1[9842] = 32'b00000000000000000011110000001010;
assign LUT_1[9843] = 32'b11111111111111111101000010000110;
assign LUT_1[9844] = 32'b00000000000000001111111011010000;
assign LUT_1[9845] = 32'b00000000000000001001001101001100;
assign LUT_1[9846] = 32'b00000000000000001011101001100001;
assign LUT_1[9847] = 32'b00000000000000000100111011011101;
assign LUT_1[9848] = 32'b00000000000000000111001111101110;
assign LUT_1[9849] = 32'b00000000000000000000100001101010;
assign LUT_1[9850] = 32'b00000000000000000010111101111111;
assign LUT_1[9851] = 32'b11111111111111111100001111111011;
assign LUT_1[9852] = 32'b00000000000000001111001001000101;
assign LUT_1[9853] = 32'b00000000000000001000011011000001;
assign LUT_1[9854] = 32'b00000000000000001010110111010110;
assign LUT_1[9855] = 32'b00000000000000000100001001010010;
assign LUT_1[9856] = 32'b00000000000000000110001101110011;
assign LUT_1[9857] = 32'b11111111111111111111011111101111;
assign LUT_1[9858] = 32'b00000000000000000001111100000100;
assign LUT_1[9859] = 32'b11111111111111111011001110000000;
assign LUT_1[9860] = 32'b00000000000000001110000111001010;
assign LUT_1[9861] = 32'b00000000000000000111011001000110;
assign LUT_1[9862] = 32'b00000000000000001001110101011011;
assign LUT_1[9863] = 32'b00000000000000000011000111010111;
assign LUT_1[9864] = 32'b00000000000000000101011011101000;
assign LUT_1[9865] = 32'b11111111111111111110101101100100;
assign LUT_1[9866] = 32'b00000000000000000001001001111001;
assign LUT_1[9867] = 32'b11111111111111111010011011110101;
assign LUT_1[9868] = 32'b00000000000000001101010100111111;
assign LUT_1[9869] = 32'b00000000000000000110100110111011;
assign LUT_1[9870] = 32'b00000000000000001001000011010000;
assign LUT_1[9871] = 32'b00000000000000000010010101001100;
assign LUT_1[9872] = 32'b00000000000000001000001001010101;
assign LUT_1[9873] = 32'b00000000000000000001011011010001;
assign LUT_1[9874] = 32'b00000000000000000011110111100110;
assign LUT_1[9875] = 32'b11111111111111111101001001100010;
assign LUT_1[9876] = 32'b00000000000000010000000010101100;
assign LUT_1[9877] = 32'b00000000000000001001010100101000;
assign LUT_1[9878] = 32'b00000000000000001011110000111101;
assign LUT_1[9879] = 32'b00000000000000000101000010111001;
assign LUT_1[9880] = 32'b00000000000000000111010111001010;
assign LUT_1[9881] = 32'b00000000000000000000101001000110;
assign LUT_1[9882] = 32'b00000000000000000011000101011011;
assign LUT_1[9883] = 32'b11111111111111111100010111010111;
assign LUT_1[9884] = 32'b00000000000000001111010000100001;
assign LUT_1[9885] = 32'b00000000000000001000100010011101;
assign LUT_1[9886] = 32'b00000000000000001010111110110010;
assign LUT_1[9887] = 32'b00000000000000000100010000101110;
assign LUT_1[9888] = 32'b00000000000000000111001000110010;
assign LUT_1[9889] = 32'b00000000000000000000011010101110;
assign LUT_1[9890] = 32'b00000000000000000010110111000011;
assign LUT_1[9891] = 32'b11111111111111111100001000111111;
assign LUT_1[9892] = 32'b00000000000000001111000010001001;
assign LUT_1[9893] = 32'b00000000000000001000010100000101;
assign LUT_1[9894] = 32'b00000000000000001010110000011010;
assign LUT_1[9895] = 32'b00000000000000000100000010010110;
assign LUT_1[9896] = 32'b00000000000000000110010110100111;
assign LUT_1[9897] = 32'b11111111111111111111101000100011;
assign LUT_1[9898] = 32'b00000000000000000010000100111000;
assign LUT_1[9899] = 32'b11111111111111111011010110110100;
assign LUT_1[9900] = 32'b00000000000000001110001111111110;
assign LUT_1[9901] = 32'b00000000000000000111100001111010;
assign LUT_1[9902] = 32'b00000000000000001001111110001111;
assign LUT_1[9903] = 32'b00000000000000000011010000001011;
assign LUT_1[9904] = 32'b00000000000000001001000100010100;
assign LUT_1[9905] = 32'b00000000000000000010010110010000;
assign LUT_1[9906] = 32'b00000000000000000100110010100101;
assign LUT_1[9907] = 32'b11111111111111111110000100100001;
assign LUT_1[9908] = 32'b00000000000000010000111101101011;
assign LUT_1[9909] = 32'b00000000000000001010001111100111;
assign LUT_1[9910] = 32'b00000000000000001100101011111100;
assign LUT_1[9911] = 32'b00000000000000000101111101111000;
assign LUT_1[9912] = 32'b00000000000000001000010010001001;
assign LUT_1[9913] = 32'b00000000000000000001100100000101;
assign LUT_1[9914] = 32'b00000000000000000100000000011010;
assign LUT_1[9915] = 32'b11111111111111111101010010010110;
assign LUT_1[9916] = 32'b00000000000000010000001011100000;
assign LUT_1[9917] = 32'b00000000000000001001011101011100;
assign LUT_1[9918] = 32'b00000000000000001011111001110001;
assign LUT_1[9919] = 32'b00000000000000000101001011101101;
assign LUT_1[9920] = 32'b00000000000000001000001011011011;
assign LUT_1[9921] = 32'b00000000000000000001011101010111;
assign LUT_1[9922] = 32'b00000000000000000011111001101100;
assign LUT_1[9923] = 32'b11111111111111111101001011101000;
assign LUT_1[9924] = 32'b00000000000000010000000100110010;
assign LUT_1[9925] = 32'b00000000000000001001010110101110;
assign LUT_1[9926] = 32'b00000000000000001011110011000011;
assign LUT_1[9927] = 32'b00000000000000000101000100111111;
assign LUT_1[9928] = 32'b00000000000000000111011001010000;
assign LUT_1[9929] = 32'b00000000000000000000101011001100;
assign LUT_1[9930] = 32'b00000000000000000011000111100001;
assign LUT_1[9931] = 32'b11111111111111111100011001011101;
assign LUT_1[9932] = 32'b00000000000000001111010010100111;
assign LUT_1[9933] = 32'b00000000000000001000100100100011;
assign LUT_1[9934] = 32'b00000000000000001011000000111000;
assign LUT_1[9935] = 32'b00000000000000000100010010110100;
assign LUT_1[9936] = 32'b00000000000000001010000110111101;
assign LUT_1[9937] = 32'b00000000000000000011011000111001;
assign LUT_1[9938] = 32'b00000000000000000101110101001110;
assign LUT_1[9939] = 32'b11111111111111111111000111001010;
assign LUT_1[9940] = 32'b00000000000000010010000000010100;
assign LUT_1[9941] = 32'b00000000000000001011010010010000;
assign LUT_1[9942] = 32'b00000000000000001101101110100101;
assign LUT_1[9943] = 32'b00000000000000000111000000100001;
assign LUT_1[9944] = 32'b00000000000000001001010100110010;
assign LUT_1[9945] = 32'b00000000000000000010100110101110;
assign LUT_1[9946] = 32'b00000000000000000101000011000011;
assign LUT_1[9947] = 32'b11111111111111111110010100111111;
assign LUT_1[9948] = 32'b00000000000000010001001110001001;
assign LUT_1[9949] = 32'b00000000000000001010100000000101;
assign LUT_1[9950] = 32'b00000000000000001100111100011010;
assign LUT_1[9951] = 32'b00000000000000000110001110010110;
assign LUT_1[9952] = 32'b00000000000000001001000110011010;
assign LUT_1[9953] = 32'b00000000000000000010011000010110;
assign LUT_1[9954] = 32'b00000000000000000100110100101011;
assign LUT_1[9955] = 32'b11111111111111111110000110100111;
assign LUT_1[9956] = 32'b00000000000000010000111111110001;
assign LUT_1[9957] = 32'b00000000000000001010010001101101;
assign LUT_1[9958] = 32'b00000000000000001100101110000010;
assign LUT_1[9959] = 32'b00000000000000000101111111111110;
assign LUT_1[9960] = 32'b00000000000000001000010100001111;
assign LUT_1[9961] = 32'b00000000000000000001100110001011;
assign LUT_1[9962] = 32'b00000000000000000100000010100000;
assign LUT_1[9963] = 32'b11111111111111111101010100011100;
assign LUT_1[9964] = 32'b00000000000000010000001101100110;
assign LUT_1[9965] = 32'b00000000000000001001011111100010;
assign LUT_1[9966] = 32'b00000000000000001011111011110111;
assign LUT_1[9967] = 32'b00000000000000000101001101110011;
assign LUT_1[9968] = 32'b00000000000000001011000001111100;
assign LUT_1[9969] = 32'b00000000000000000100010011111000;
assign LUT_1[9970] = 32'b00000000000000000110110000001101;
assign LUT_1[9971] = 32'b00000000000000000000000010001001;
assign LUT_1[9972] = 32'b00000000000000010010111011010011;
assign LUT_1[9973] = 32'b00000000000000001100001101001111;
assign LUT_1[9974] = 32'b00000000000000001110101001100100;
assign LUT_1[9975] = 32'b00000000000000000111111011100000;
assign LUT_1[9976] = 32'b00000000000000001010001111110001;
assign LUT_1[9977] = 32'b00000000000000000011100001101101;
assign LUT_1[9978] = 32'b00000000000000000101111110000010;
assign LUT_1[9979] = 32'b11111111111111111111001111111110;
assign LUT_1[9980] = 32'b00000000000000010010001001001000;
assign LUT_1[9981] = 32'b00000000000000001011011011000100;
assign LUT_1[9982] = 32'b00000000000000001101110111011001;
assign LUT_1[9983] = 32'b00000000000000000111001001010101;
assign LUT_1[9984] = 32'b00000000000000000001000001111100;
assign LUT_1[9985] = 32'b11111111111111111010010011111000;
assign LUT_1[9986] = 32'b11111111111111111100110000001101;
assign LUT_1[9987] = 32'b11111111111111110110000010001001;
assign LUT_1[9988] = 32'b00000000000000001000111011010011;
assign LUT_1[9989] = 32'b00000000000000000010001101001111;
assign LUT_1[9990] = 32'b00000000000000000100101001100100;
assign LUT_1[9991] = 32'b11111111111111111101111011100000;
assign LUT_1[9992] = 32'b00000000000000000000001111110001;
assign LUT_1[9993] = 32'b11111111111111111001100001101101;
assign LUT_1[9994] = 32'b11111111111111111011111110000010;
assign LUT_1[9995] = 32'b11111111111111110101001111111110;
assign LUT_1[9996] = 32'b00000000000000001000001001001000;
assign LUT_1[9997] = 32'b00000000000000000001011011000100;
assign LUT_1[9998] = 32'b00000000000000000011110111011001;
assign LUT_1[9999] = 32'b11111111111111111101001001010101;
assign LUT_1[10000] = 32'b00000000000000000010111101011110;
assign LUT_1[10001] = 32'b11111111111111111100001111011010;
assign LUT_1[10002] = 32'b11111111111111111110101011101111;
assign LUT_1[10003] = 32'b11111111111111110111111101101011;
assign LUT_1[10004] = 32'b00000000000000001010110110110101;
assign LUT_1[10005] = 32'b00000000000000000100001000110001;
assign LUT_1[10006] = 32'b00000000000000000110100101000110;
assign LUT_1[10007] = 32'b11111111111111111111110111000010;
assign LUT_1[10008] = 32'b00000000000000000010001011010011;
assign LUT_1[10009] = 32'b11111111111111111011011101001111;
assign LUT_1[10010] = 32'b11111111111111111101111001100100;
assign LUT_1[10011] = 32'b11111111111111110111001011100000;
assign LUT_1[10012] = 32'b00000000000000001010000100101010;
assign LUT_1[10013] = 32'b00000000000000000011010110100110;
assign LUT_1[10014] = 32'b00000000000000000101110010111011;
assign LUT_1[10015] = 32'b11111111111111111111000100110111;
assign LUT_1[10016] = 32'b00000000000000000001111100111011;
assign LUT_1[10017] = 32'b11111111111111111011001110110111;
assign LUT_1[10018] = 32'b11111111111111111101101011001100;
assign LUT_1[10019] = 32'b11111111111111110110111101001000;
assign LUT_1[10020] = 32'b00000000000000001001110110010010;
assign LUT_1[10021] = 32'b00000000000000000011001000001110;
assign LUT_1[10022] = 32'b00000000000000000101100100100011;
assign LUT_1[10023] = 32'b11111111111111111110110110011111;
assign LUT_1[10024] = 32'b00000000000000000001001010110000;
assign LUT_1[10025] = 32'b11111111111111111010011100101100;
assign LUT_1[10026] = 32'b11111111111111111100111001000001;
assign LUT_1[10027] = 32'b11111111111111110110001010111101;
assign LUT_1[10028] = 32'b00000000000000001001000100000111;
assign LUT_1[10029] = 32'b00000000000000000010010110000011;
assign LUT_1[10030] = 32'b00000000000000000100110010011000;
assign LUT_1[10031] = 32'b11111111111111111110000100010100;
assign LUT_1[10032] = 32'b00000000000000000011111000011101;
assign LUT_1[10033] = 32'b11111111111111111101001010011001;
assign LUT_1[10034] = 32'b11111111111111111111100110101110;
assign LUT_1[10035] = 32'b11111111111111111000111000101010;
assign LUT_1[10036] = 32'b00000000000000001011110001110100;
assign LUT_1[10037] = 32'b00000000000000000101000011110000;
assign LUT_1[10038] = 32'b00000000000000000111100000000101;
assign LUT_1[10039] = 32'b00000000000000000000110010000001;
assign LUT_1[10040] = 32'b00000000000000000011000110010010;
assign LUT_1[10041] = 32'b11111111111111111100011000001110;
assign LUT_1[10042] = 32'b11111111111111111110110100100011;
assign LUT_1[10043] = 32'b11111111111111111000000110011111;
assign LUT_1[10044] = 32'b00000000000000001010111111101001;
assign LUT_1[10045] = 32'b00000000000000000100010001100101;
assign LUT_1[10046] = 32'b00000000000000000110101101111010;
assign LUT_1[10047] = 32'b11111111111111111111111111110110;
assign LUT_1[10048] = 32'b00000000000000000010111111100100;
assign LUT_1[10049] = 32'b11111111111111111100010001100000;
assign LUT_1[10050] = 32'b11111111111111111110101101110101;
assign LUT_1[10051] = 32'b11111111111111110111111111110001;
assign LUT_1[10052] = 32'b00000000000000001010111000111011;
assign LUT_1[10053] = 32'b00000000000000000100001010110111;
assign LUT_1[10054] = 32'b00000000000000000110100111001100;
assign LUT_1[10055] = 32'b11111111111111111111111001001000;
assign LUT_1[10056] = 32'b00000000000000000010001101011001;
assign LUT_1[10057] = 32'b11111111111111111011011111010101;
assign LUT_1[10058] = 32'b11111111111111111101111011101010;
assign LUT_1[10059] = 32'b11111111111111110111001101100110;
assign LUT_1[10060] = 32'b00000000000000001010000110110000;
assign LUT_1[10061] = 32'b00000000000000000011011000101100;
assign LUT_1[10062] = 32'b00000000000000000101110101000001;
assign LUT_1[10063] = 32'b11111111111111111111000110111101;
assign LUT_1[10064] = 32'b00000000000000000100111011000110;
assign LUT_1[10065] = 32'b11111111111111111110001101000010;
assign LUT_1[10066] = 32'b00000000000000000000101001010111;
assign LUT_1[10067] = 32'b11111111111111111001111011010011;
assign LUT_1[10068] = 32'b00000000000000001100110100011101;
assign LUT_1[10069] = 32'b00000000000000000110000110011001;
assign LUT_1[10070] = 32'b00000000000000001000100010101110;
assign LUT_1[10071] = 32'b00000000000000000001110100101010;
assign LUT_1[10072] = 32'b00000000000000000100001000111011;
assign LUT_1[10073] = 32'b11111111111111111101011010110111;
assign LUT_1[10074] = 32'b11111111111111111111110111001100;
assign LUT_1[10075] = 32'b11111111111111111001001001001000;
assign LUT_1[10076] = 32'b00000000000000001100000010010010;
assign LUT_1[10077] = 32'b00000000000000000101010100001110;
assign LUT_1[10078] = 32'b00000000000000000111110000100011;
assign LUT_1[10079] = 32'b00000000000000000001000010011111;
assign LUT_1[10080] = 32'b00000000000000000011111010100011;
assign LUT_1[10081] = 32'b11111111111111111101001100011111;
assign LUT_1[10082] = 32'b11111111111111111111101000110100;
assign LUT_1[10083] = 32'b11111111111111111000111010110000;
assign LUT_1[10084] = 32'b00000000000000001011110011111010;
assign LUT_1[10085] = 32'b00000000000000000101000101110110;
assign LUT_1[10086] = 32'b00000000000000000111100010001011;
assign LUT_1[10087] = 32'b00000000000000000000110100000111;
assign LUT_1[10088] = 32'b00000000000000000011001000011000;
assign LUT_1[10089] = 32'b11111111111111111100011010010100;
assign LUT_1[10090] = 32'b11111111111111111110110110101001;
assign LUT_1[10091] = 32'b11111111111111111000001000100101;
assign LUT_1[10092] = 32'b00000000000000001011000001101111;
assign LUT_1[10093] = 32'b00000000000000000100010011101011;
assign LUT_1[10094] = 32'b00000000000000000110110000000000;
assign LUT_1[10095] = 32'b00000000000000000000000001111100;
assign LUT_1[10096] = 32'b00000000000000000101110110000101;
assign LUT_1[10097] = 32'b11111111111111111111001000000001;
assign LUT_1[10098] = 32'b00000000000000000001100100010110;
assign LUT_1[10099] = 32'b11111111111111111010110110010010;
assign LUT_1[10100] = 32'b00000000000000001101101111011100;
assign LUT_1[10101] = 32'b00000000000000000111000001011000;
assign LUT_1[10102] = 32'b00000000000000001001011101101101;
assign LUT_1[10103] = 32'b00000000000000000010101111101001;
assign LUT_1[10104] = 32'b00000000000000000101000011111010;
assign LUT_1[10105] = 32'b11111111111111111110010101110110;
assign LUT_1[10106] = 32'b00000000000000000000110010001011;
assign LUT_1[10107] = 32'b11111111111111111010000100000111;
assign LUT_1[10108] = 32'b00000000000000001100111101010001;
assign LUT_1[10109] = 32'b00000000000000000110001111001101;
assign LUT_1[10110] = 32'b00000000000000001000101011100010;
assign LUT_1[10111] = 32'b00000000000000000001111101011110;
assign LUT_1[10112] = 32'b00000000000000000100000001111111;
assign LUT_1[10113] = 32'b11111111111111111101010011111011;
assign LUT_1[10114] = 32'b11111111111111111111110000010000;
assign LUT_1[10115] = 32'b11111111111111111001000010001100;
assign LUT_1[10116] = 32'b00000000000000001011111011010110;
assign LUT_1[10117] = 32'b00000000000000000101001101010010;
assign LUT_1[10118] = 32'b00000000000000000111101001100111;
assign LUT_1[10119] = 32'b00000000000000000000111011100011;
assign LUT_1[10120] = 32'b00000000000000000011001111110100;
assign LUT_1[10121] = 32'b11111111111111111100100001110000;
assign LUT_1[10122] = 32'b11111111111111111110111110000101;
assign LUT_1[10123] = 32'b11111111111111111000010000000001;
assign LUT_1[10124] = 32'b00000000000000001011001001001011;
assign LUT_1[10125] = 32'b00000000000000000100011011000111;
assign LUT_1[10126] = 32'b00000000000000000110110111011100;
assign LUT_1[10127] = 32'b00000000000000000000001001011000;
assign LUT_1[10128] = 32'b00000000000000000101111101100001;
assign LUT_1[10129] = 32'b11111111111111111111001111011101;
assign LUT_1[10130] = 32'b00000000000000000001101011110010;
assign LUT_1[10131] = 32'b11111111111111111010111101101110;
assign LUT_1[10132] = 32'b00000000000000001101110110111000;
assign LUT_1[10133] = 32'b00000000000000000111001000110100;
assign LUT_1[10134] = 32'b00000000000000001001100101001001;
assign LUT_1[10135] = 32'b00000000000000000010110111000101;
assign LUT_1[10136] = 32'b00000000000000000101001011010110;
assign LUT_1[10137] = 32'b11111111111111111110011101010010;
assign LUT_1[10138] = 32'b00000000000000000000111001100111;
assign LUT_1[10139] = 32'b11111111111111111010001011100011;
assign LUT_1[10140] = 32'b00000000000000001101000100101101;
assign LUT_1[10141] = 32'b00000000000000000110010110101001;
assign LUT_1[10142] = 32'b00000000000000001000110010111110;
assign LUT_1[10143] = 32'b00000000000000000010000100111010;
assign LUT_1[10144] = 32'b00000000000000000100111100111110;
assign LUT_1[10145] = 32'b11111111111111111110001110111010;
assign LUT_1[10146] = 32'b00000000000000000000101011001111;
assign LUT_1[10147] = 32'b11111111111111111001111101001011;
assign LUT_1[10148] = 32'b00000000000000001100110110010101;
assign LUT_1[10149] = 32'b00000000000000000110001000010001;
assign LUT_1[10150] = 32'b00000000000000001000100100100110;
assign LUT_1[10151] = 32'b00000000000000000001110110100010;
assign LUT_1[10152] = 32'b00000000000000000100001010110011;
assign LUT_1[10153] = 32'b11111111111111111101011100101111;
assign LUT_1[10154] = 32'b11111111111111111111111001000100;
assign LUT_1[10155] = 32'b11111111111111111001001011000000;
assign LUT_1[10156] = 32'b00000000000000001100000100001010;
assign LUT_1[10157] = 32'b00000000000000000101010110000110;
assign LUT_1[10158] = 32'b00000000000000000111110010011011;
assign LUT_1[10159] = 32'b00000000000000000001000100010111;
assign LUT_1[10160] = 32'b00000000000000000110111000100000;
assign LUT_1[10161] = 32'b00000000000000000000001010011100;
assign LUT_1[10162] = 32'b00000000000000000010100110110001;
assign LUT_1[10163] = 32'b11111111111111111011111000101101;
assign LUT_1[10164] = 32'b00000000000000001110110001110111;
assign LUT_1[10165] = 32'b00000000000000001000000011110011;
assign LUT_1[10166] = 32'b00000000000000001010100000001000;
assign LUT_1[10167] = 32'b00000000000000000011110010000100;
assign LUT_1[10168] = 32'b00000000000000000110000110010101;
assign LUT_1[10169] = 32'b11111111111111111111011000010001;
assign LUT_1[10170] = 32'b00000000000000000001110100100110;
assign LUT_1[10171] = 32'b11111111111111111011000110100010;
assign LUT_1[10172] = 32'b00000000000000001101111111101100;
assign LUT_1[10173] = 32'b00000000000000000111010001101000;
assign LUT_1[10174] = 32'b00000000000000001001101101111101;
assign LUT_1[10175] = 32'b00000000000000000010111111111001;
assign LUT_1[10176] = 32'b00000000000000000101111111100111;
assign LUT_1[10177] = 32'b11111111111111111111010001100011;
assign LUT_1[10178] = 32'b00000000000000000001101101111000;
assign LUT_1[10179] = 32'b11111111111111111010111111110100;
assign LUT_1[10180] = 32'b00000000000000001101111000111110;
assign LUT_1[10181] = 32'b00000000000000000111001010111010;
assign LUT_1[10182] = 32'b00000000000000001001100111001111;
assign LUT_1[10183] = 32'b00000000000000000010111001001011;
assign LUT_1[10184] = 32'b00000000000000000101001101011100;
assign LUT_1[10185] = 32'b11111111111111111110011111011000;
assign LUT_1[10186] = 32'b00000000000000000000111011101101;
assign LUT_1[10187] = 32'b11111111111111111010001101101001;
assign LUT_1[10188] = 32'b00000000000000001101000110110011;
assign LUT_1[10189] = 32'b00000000000000000110011000101111;
assign LUT_1[10190] = 32'b00000000000000001000110101000100;
assign LUT_1[10191] = 32'b00000000000000000010000111000000;
assign LUT_1[10192] = 32'b00000000000000000111111011001001;
assign LUT_1[10193] = 32'b00000000000000000001001101000101;
assign LUT_1[10194] = 32'b00000000000000000011101001011010;
assign LUT_1[10195] = 32'b11111111111111111100111011010110;
assign LUT_1[10196] = 32'b00000000000000001111110100100000;
assign LUT_1[10197] = 32'b00000000000000001001000110011100;
assign LUT_1[10198] = 32'b00000000000000001011100010110001;
assign LUT_1[10199] = 32'b00000000000000000100110100101101;
assign LUT_1[10200] = 32'b00000000000000000111001000111110;
assign LUT_1[10201] = 32'b00000000000000000000011010111010;
assign LUT_1[10202] = 32'b00000000000000000010110111001111;
assign LUT_1[10203] = 32'b11111111111111111100001001001011;
assign LUT_1[10204] = 32'b00000000000000001111000010010101;
assign LUT_1[10205] = 32'b00000000000000001000010100010001;
assign LUT_1[10206] = 32'b00000000000000001010110000100110;
assign LUT_1[10207] = 32'b00000000000000000100000010100010;
assign LUT_1[10208] = 32'b00000000000000000110111010100110;
assign LUT_1[10209] = 32'b00000000000000000000001100100010;
assign LUT_1[10210] = 32'b00000000000000000010101000110111;
assign LUT_1[10211] = 32'b11111111111111111011111010110011;
assign LUT_1[10212] = 32'b00000000000000001110110011111101;
assign LUT_1[10213] = 32'b00000000000000001000000101111001;
assign LUT_1[10214] = 32'b00000000000000001010100010001110;
assign LUT_1[10215] = 32'b00000000000000000011110100001010;
assign LUT_1[10216] = 32'b00000000000000000110001000011011;
assign LUT_1[10217] = 32'b11111111111111111111011010010111;
assign LUT_1[10218] = 32'b00000000000000000001110110101100;
assign LUT_1[10219] = 32'b11111111111111111011001000101000;
assign LUT_1[10220] = 32'b00000000000000001110000001110010;
assign LUT_1[10221] = 32'b00000000000000000111010011101110;
assign LUT_1[10222] = 32'b00000000000000001001110000000011;
assign LUT_1[10223] = 32'b00000000000000000011000001111111;
assign LUT_1[10224] = 32'b00000000000000001000110110001000;
assign LUT_1[10225] = 32'b00000000000000000010001000000100;
assign LUT_1[10226] = 32'b00000000000000000100100100011001;
assign LUT_1[10227] = 32'b11111111111111111101110110010101;
assign LUT_1[10228] = 32'b00000000000000010000101111011111;
assign LUT_1[10229] = 32'b00000000000000001010000001011011;
assign LUT_1[10230] = 32'b00000000000000001100011101110000;
assign LUT_1[10231] = 32'b00000000000000000101101111101100;
assign LUT_1[10232] = 32'b00000000000000001000000011111101;
assign LUT_1[10233] = 32'b00000000000000000001010101111001;
assign LUT_1[10234] = 32'b00000000000000000011110010001110;
assign LUT_1[10235] = 32'b11111111111111111101000100001010;
assign LUT_1[10236] = 32'b00000000000000001111111101010100;
assign LUT_1[10237] = 32'b00000000000000001001001111010000;
assign LUT_1[10238] = 32'b00000000000000001011101011100101;
assign LUT_1[10239] = 32'b00000000000000000100111101100001;
assign LUT_1[10240] = 32'b00000000000000000100001010011110;
assign LUT_1[10241] = 32'b11111111111111111101011100011010;
assign LUT_1[10242] = 32'b11111111111111111111111000101111;
assign LUT_1[10243] = 32'b11111111111111111001001010101011;
assign LUT_1[10244] = 32'b00000000000000001100000011110101;
assign LUT_1[10245] = 32'b00000000000000000101010101110001;
assign LUT_1[10246] = 32'b00000000000000000111110010000110;
assign LUT_1[10247] = 32'b00000000000000000001000100000010;
assign LUT_1[10248] = 32'b00000000000000000011011000010011;
assign LUT_1[10249] = 32'b11111111111111111100101010001111;
assign LUT_1[10250] = 32'b11111111111111111111000110100100;
assign LUT_1[10251] = 32'b11111111111111111000011000100000;
assign LUT_1[10252] = 32'b00000000000000001011010001101010;
assign LUT_1[10253] = 32'b00000000000000000100100011100110;
assign LUT_1[10254] = 32'b00000000000000000110111111111011;
assign LUT_1[10255] = 32'b00000000000000000000010001110111;
assign LUT_1[10256] = 32'b00000000000000000110000110000000;
assign LUT_1[10257] = 32'b11111111111111111111010111111100;
assign LUT_1[10258] = 32'b00000000000000000001110100010001;
assign LUT_1[10259] = 32'b11111111111111111011000110001101;
assign LUT_1[10260] = 32'b00000000000000001101111111010111;
assign LUT_1[10261] = 32'b00000000000000000111010001010011;
assign LUT_1[10262] = 32'b00000000000000001001101101101000;
assign LUT_1[10263] = 32'b00000000000000000010111111100100;
assign LUT_1[10264] = 32'b00000000000000000101010011110101;
assign LUT_1[10265] = 32'b11111111111111111110100101110001;
assign LUT_1[10266] = 32'b00000000000000000001000010000110;
assign LUT_1[10267] = 32'b11111111111111111010010100000010;
assign LUT_1[10268] = 32'b00000000000000001101001101001100;
assign LUT_1[10269] = 32'b00000000000000000110011111001000;
assign LUT_1[10270] = 32'b00000000000000001000111011011101;
assign LUT_1[10271] = 32'b00000000000000000010001101011001;
assign LUT_1[10272] = 32'b00000000000000000101000101011101;
assign LUT_1[10273] = 32'b11111111111111111110010111011001;
assign LUT_1[10274] = 32'b00000000000000000000110011101110;
assign LUT_1[10275] = 32'b11111111111111111010000101101010;
assign LUT_1[10276] = 32'b00000000000000001100111110110100;
assign LUT_1[10277] = 32'b00000000000000000110010000110000;
assign LUT_1[10278] = 32'b00000000000000001000101101000101;
assign LUT_1[10279] = 32'b00000000000000000001111111000001;
assign LUT_1[10280] = 32'b00000000000000000100010011010010;
assign LUT_1[10281] = 32'b11111111111111111101100101001110;
assign LUT_1[10282] = 32'b00000000000000000000000001100011;
assign LUT_1[10283] = 32'b11111111111111111001010011011111;
assign LUT_1[10284] = 32'b00000000000000001100001100101001;
assign LUT_1[10285] = 32'b00000000000000000101011110100101;
assign LUT_1[10286] = 32'b00000000000000000111111010111010;
assign LUT_1[10287] = 32'b00000000000000000001001100110110;
assign LUT_1[10288] = 32'b00000000000000000111000000111111;
assign LUT_1[10289] = 32'b00000000000000000000010010111011;
assign LUT_1[10290] = 32'b00000000000000000010101111010000;
assign LUT_1[10291] = 32'b11111111111111111100000001001100;
assign LUT_1[10292] = 32'b00000000000000001110111010010110;
assign LUT_1[10293] = 32'b00000000000000001000001100010010;
assign LUT_1[10294] = 32'b00000000000000001010101000100111;
assign LUT_1[10295] = 32'b00000000000000000011111010100011;
assign LUT_1[10296] = 32'b00000000000000000110001110110100;
assign LUT_1[10297] = 32'b11111111111111111111100000110000;
assign LUT_1[10298] = 32'b00000000000000000001111101000101;
assign LUT_1[10299] = 32'b11111111111111111011001111000001;
assign LUT_1[10300] = 32'b00000000000000001110001000001011;
assign LUT_1[10301] = 32'b00000000000000000111011010000111;
assign LUT_1[10302] = 32'b00000000000000001001110110011100;
assign LUT_1[10303] = 32'b00000000000000000011001000011000;
assign LUT_1[10304] = 32'b00000000000000000110001000000110;
assign LUT_1[10305] = 32'b11111111111111111111011010000010;
assign LUT_1[10306] = 32'b00000000000000000001110110010111;
assign LUT_1[10307] = 32'b11111111111111111011001000010011;
assign LUT_1[10308] = 32'b00000000000000001110000001011101;
assign LUT_1[10309] = 32'b00000000000000000111010011011001;
assign LUT_1[10310] = 32'b00000000000000001001101111101110;
assign LUT_1[10311] = 32'b00000000000000000011000001101010;
assign LUT_1[10312] = 32'b00000000000000000101010101111011;
assign LUT_1[10313] = 32'b11111111111111111110100111110111;
assign LUT_1[10314] = 32'b00000000000000000001000100001100;
assign LUT_1[10315] = 32'b11111111111111111010010110001000;
assign LUT_1[10316] = 32'b00000000000000001101001111010010;
assign LUT_1[10317] = 32'b00000000000000000110100001001110;
assign LUT_1[10318] = 32'b00000000000000001000111101100011;
assign LUT_1[10319] = 32'b00000000000000000010001111011111;
assign LUT_1[10320] = 32'b00000000000000001000000011101000;
assign LUT_1[10321] = 32'b00000000000000000001010101100100;
assign LUT_1[10322] = 32'b00000000000000000011110001111001;
assign LUT_1[10323] = 32'b11111111111111111101000011110101;
assign LUT_1[10324] = 32'b00000000000000001111111100111111;
assign LUT_1[10325] = 32'b00000000000000001001001110111011;
assign LUT_1[10326] = 32'b00000000000000001011101011010000;
assign LUT_1[10327] = 32'b00000000000000000100111101001100;
assign LUT_1[10328] = 32'b00000000000000000111010001011101;
assign LUT_1[10329] = 32'b00000000000000000000100011011001;
assign LUT_1[10330] = 32'b00000000000000000010111111101110;
assign LUT_1[10331] = 32'b11111111111111111100010001101010;
assign LUT_1[10332] = 32'b00000000000000001111001010110100;
assign LUT_1[10333] = 32'b00000000000000001000011100110000;
assign LUT_1[10334] = 32'b00000000000000001010111001000101;
assign LUT_1[10335] = 32'b00000000000000000100001011000001;
assign LUT_1[10336] = 32'b00000000000000000111000011000101;
assign LUT_1[10337] = 32'b00000000000000000000010101000001;
assign LUT_1[10338] = 32'b00000000000000000010110001010110;
assign LUT_1[10339] = 32'b11111111111111111100000011010010;
assign LUT_1[10340] = 32'b00000000000000001110111100011100;
assign LUT_1[10341] = 32'b00000000000000001000001110011000;
assign LUT_1[10342] = 32'b00000000000000001010101010101101;
assign LUT_1[10343] = 32'b00000000000000000011111100101001;
assign LUT_1[10344] = 32'b00000000000000000110010000111010;
assign LUT_1[10345] = 32'b11111111111111111111100010110110;
assign LUT_1[10346] = 32'b00000000000000000001111111001011;
assign LUT_1[10347] = 32'b11111111111111111011010001000111;
assign LUT_1[10348] = 32'b00000000000000001110001010010001;
assign LUT_1[10349] = 32'b00000000000000000111011100001101;
assign LUT_1[10350] = 32'b00000000000000001001111000100010;
assign LUT_1[10351] = 32'b00000000000000000011001010011110;
assign LUT_1[10352] = 32'b00000000000000001000111110100111;
assign LUT_1[10353] = 32'b00000000000000000010010000100011;
assign LUT_1[10354] = 32'b00000000000000000100101100111000;
assign LUT_1[10355] = 32'b11111111111111111101111110110100;
assign LUT_1[10356] = 32'b00000000000000010000110111111110;
assign LUT_1[10357] = 32'b00000000000000001010001001111010;
assign LUT_1[10358] = 32'b00000000000000001100100110001111;
assign LUT_1[10359] = 32'b00000000000000000101111000001011;
assign LUT_1[10360] = 32'b00000000000000001000001100011100;
assign LUT_1[10361] = 32'b00000000000000000001011110011000;
assign LUT_1[10362] = 32'b00000000000000000011111010101101;
assign LUT_1[10363] = 32'b11111111111111111101001100101001;
assign LUT_1[10364] = 32'b00000000000000010000000101110011;
assign LUT_1[10365] = 32'b00000000000000001001010111101111;
assign LUT_1[10366] = 32'b00000000000000001011110100000100;
assign LUT_1[10367] = 32'b00000000000000000101000110000000;
assign LUT_1[10368] = 32'b00000000000000000111001010100001;
assign LUT_1[10369] = 32'b00000000000000000000011100011101;
assign LUT_1[10370] = 32'b00000000000000000010111000110010;
assign LUT_1[10371] = 32'b11111111111111111100001010101110;
assign LUT_1[10372] = 32'b00000000000000001111000011111000;
assign LUT_1[10373] = 32'b00000000000000001000010101110100;
assign LUT_1[10374] = 32'b00000000000000001010110010001001;
assign LUT_1[10375] = 32'b00000000000000000100000100000101;
assign LUT_1[10376] = 32'b00000000000000000110011000010110;
assign LUT_1[10377] = 32'b11111111111111111111101010010010;
assign LUT_1[10378] = 32'b00000000000000000010000110100111;
assign LUT_1[10379] = 32'b11111111111111111011011000100011;
assign LUT_1[10380] = 32'b00000000000000001110010001101101;
assign LUT_1[10381] = 32'b00000000000000000111100011101001;
assign LUT_1[10382] = 32'b00000000000000001001111111111110;
assign LUT_1[10383] = 32'b00000000000000000011010001111010;
assign LUT_1[10384] = 32'b00000000000000001001000110000011;
assign LUT_1[10385] = 32'b00000000000000000010010111111111;
assign LUT_1[10386] = 32'b00000000000000000100110100010100;
assign LUT_1[10387] = 32'b11111111111111111110000110010000;
assign LUT_1[10388] = 32'b00000000000000010000111111011010;
assign LUT_1[10389] = 32'b00000000000000001010010001010110;
assign LUT_1[10390] = 32'b00000000000000001100101101101011;
assign LUT_1[10391] = 32'b00000000000000000101111111100111;
assign LUT_1[10392] = 32'b00000000000000001000010011111000;
assign LUT_1[10393] = 32'b00000000000000000001100101110100;
assign LUT_1[10394] = 32'b00000000000000000100000010001001;
assign LUT_1[10395] = 32'b11111111111111111101010100000101;
assign LUT_1[10396] = 32'b00000000000000010000001101001111;
assign LUT_1[10397] = 32'b00000000000000001001011111001011;
assign LUT_1[10398] = 32'b00000000000000001011111011100000;
assign LUT_1[10399] = 32'b00000000000000000101001101011100;
assign LUT_1[10400] = 32'b00000000000000001000000101100000;
assign LUT_1[10401] = 32'b00000000000000000001010111011100;
assign LUT_1[10402] = 32'b00000000000000000011110011110001;
assign LUT_1[10403] = 32'b11111111111111111101000101101101;
assign LUT_1[10404] = 32'b00000000000000001111111110110111;
assign LUT_1[10405] = 32'b00000000000000001001010000110011;
assign LUT_1[10406] = 32'b00000000000000001011101101001000;
assign LUT_1[10407] = 32'b00000000000000000100111111000100;
assign LUT_1[10408] = 32'b00000000000000000111010011010101;
assign LUT_1[10409] = 32'b00000000000000000000100101010001;
assign LUT_1[10410] = 32'b00000000000000000011000001100110;
assign LUT_1[10411] = 32'b11111111111111111100010011100010;
assign LUT_1[10412] = 32'b00000000000000001111001100101100;
assign LUT_1[10413] = 32'b00000000000000001000011110101000;
assign LUT_1[10414] = 32'b00000000000000001010111010111101;
assign LUT_1[10415] = 32'b00000000000000000100001100111001;
assign LUT_1[10416] = 32'b00000000000000001010000001000010;
assign LUT_1[10417] = 32'b00000000000000000011010010111110;
assign LUT_1[10418] = 32'b00000000000000000101101111010011;
assign LUT_1[10419] = 32'b11111111111111111111000001001111;
assign LUT_1[10420] = 32'b00000000000000010001111010011001;
assign LUT_1[10421] = 32'b00000000000000001011001100010101;
assign LUT_1[10422] = 32'b00000000000000001101101000101010;
assign LUT_1[10423] = 32'b00000000000000000110111010100110;
assign LUT_1[10424] = 32'b00000000000000001001001110110111;
assign LUT_1[10425] = 32'b00000000000000000010100000110011;
assign LUT_1[10426] = 32'b00000000000000000100111101001000;
assign LUT_1[10427] = 32'b11111111111111111110001111000100;
assign LUT_1[10428] = 32'b00000000000000010001001000001110;
assign LUT_1[10429] = 32'b00000000000000001010011010001010;
assign LUT_1[10430] = 32'b00000000000000001100110110011111;
assign LUT_1[10431] = 32'b00000000000000000110001000011011;
assign LUT_1[10432] = 32'b00000000000000001001001000001001;
assign LUT_1[10433] = 32'b00000000000000000010011010000101;
assign LUT_1[10434] = 32'b00000000000000000100110110011010;
assign LUT_1[10435] = 32'b11111111111111111110001000010110;
assign LUT_1[10436] = 32'b00000000000000010001000001100000;
assign LUT_1[10437] = 32'b00000000000000001010010011011100;
assign LUT_1[10438] = 32'b00000000000000001100101111110001;
assign LUT_1[10439] = 32'b00000000000000000110000001101101;
assign LUT_1[10440] = 32'b00000000000000001000010101111110;
assign LUT_1[10441] = 32'b00000000000000000001100111111010;
assign LUT_1[10442] = 32'b00000000000000000100000100001111;
assign LUT_1[10443] = 32'b11111111111111111101010110001011;
assign LUT_1[10444] = 32'b00000000000000010000001111010101;
assign LUT_1[10445] = 32'b00000000000000001001100001010001;
assign LUT_1[10446] = 32'b00000000000000001011111101100110;
assign LUT_1[10447] = 32'b00000000000000000101001111100010;
assign LUT_1[10448] = 32'b00000000000000001011000011101011;
assign LUT_1[10449] = 32'b00000000000000000100010101100111;
assign LUT_1[10450] = 32'b00000000000000000110110001111100;
assign LUT_1[10451] = 32'b00000000000000000000000011111000;
assign LUT_1[10452] = 32'b00000000000000010010111101000010;
assign LUT_1[10453] = 32'b00000000000000001100001110111110;
assign LUT_1[10454] = 32'b00000000000000001110101011010011;
assign LUT_1[10455] = 32'b00000000000000000111111101001111;
assign LUT_1[10456] = 32'b00000000000000001010010001100000;
assign LUT_1[10457] = 32'b00000000000000000011100011011100;
assign LUT_1[10458] = 32'b00000000000000000101111111110001;
assign LUT_1[10459] = 32'b11111111111111111111010001101101;
assign LUT_1[10460] = 32'b00000000000000010010001010110111;
assign LUT_1[10461] = 32'b00000000000000001011011100110011;
assign LUT_1[10462] = 32'b00000000000000001101111001001000;
assign LUT_1[10463] = 32'b00000000000000000111001011000100;
assign LUT_1[10464] = 32'b00000000000000001010000011001000;
assign LUT_1[10465] = 32'b00000000000000000011010101000100;
assign LUT_1[10466] = 32'b00000000000000000101110001011001;
assign LUT_1[10467] = 32'b11111111111111111111000011010101;
assign LUT_1[10468] = 32'b00000000000000010001111100011111;
assign LUT_1[10469] = 32'b00000000000000001011001110011011;
assign LUT_1[10470] = 32'b00000000000000001101101010110000;
assign LUT_1[10471] = 32'b00000000000000000110111100101100;
assign LUT_1[10472] = 32'b00000000000000001001010000111101;
assign LUT_1[10473] = 32'b00000000000000000010100010111001;
assign LUT_1[10474] = 32'b00000000000000000100111111001110;
assign LUT_1[10475] = 32'b11111111111111111110010001001010;
assign LUT_1[10476] = 32'b00000000000000010001001010010100;
assign LUT_1[10477] = 32'b00000000000000001010011100010000;
assign LUT_1[10478] = 32'b00000000000000001100111000100101;
assign LUT_1[10479] = 32'b00000000000000000110001010100001;
assign LUT_1[10480] = 32'b00000000000000001011111110101010;
assign LUT_1[10481] = 32'b00000000000000000101010000100110;
assign LUT_1[10482] = 32'b00000000000000000111101100111011;
assign LUT_1[10483] = 32'b00000000000000000000111110110111;
assign LUT_1[10484] = 32'b00000000000000010011111000000001;
assign LUT_1[10485] = 32'b00000000000000001101001001111101;
assign LUT_1[10486] = 32'b00000000000000001111100110010010;
assign LUT_1[10487] = 32'b00000000000000001000111000001110;
assign LUT_1[10488] = 32'b00000000000000001011001100011111;
assign LUT_1[10489] = 32'b00000000000000000100011110011011;
assign LUT_1[10490] = 32'b00000000000000000110111010110000;
assign LUT_1[10491] = 32'b00000000000000000000001100101100;
assign LUT_1[10492] = 32'b00000000000000010011000101110110;
assign LUT_1[10493] = 32'b00000000000000001100010111110010;
assign LUT_1[10494] = 32'b00000000000000001110110100000111;
assign LUT_1[10495] = 32'b00000000000000001000000110000011;
assign LUT_1[10496] = 32'b00000000000000000001111110101010;
assign LUT_1[10497] = 32'b11111111111111111011010000100110;
assign LUT_1[10498] = 32'b11111111111111111101101100111011;
assign LUT_1[10499] = 32'b11111111111111110110111110110111;
assign LUT_1[10500] = 32'b00000000000000001001111000000001;
assign LUT_1[10501] = 32'b00000000000000000011001001111101;
assign LUT_1[10502] = 32'b00000000000000000101100110010010;
assign LUT_1[10503] = 32'b11111111111111111110111000001110;
assign LUT_1[10504] = 32'b00000000000000000001001100011111;
assign LUT_1[10505] = 32'b11111111111111111010011110011011;
assign LUT_1[10506] = 32'b11111111111111111100111010110000;
assign LUT_1[10507] = 32'b11111111111111110110001100101100;
assign LUT_1[10508] = 32'b00000000000000001001000101110110;
assign LUT_1[10509] = 32'b00000000000000000010010111110010;
assign LUT_1[10510] = 32'b00000000000000000100110100000111;
assign LUT_1[10511] = 32'b11111111111111111110000110000011;
assign LUT_1[10512] = 32'b00000000000000000011111010001100;
assign LUT_1[10513] = 32'b11111111111111111101001100001000;
assign LUT_1[10514] = 32'b11111111111111111111101000011101;
assign LUT_1[10515] = 32'b11111111111111111000111010011001;
assign LUT_1[10516] = 32'b00000000000000001011110011100011;
assign LUT_1[10517] = 32'b00000000000000000101000101011111;
assign LUT_1[10518] = 32'b00000000000000000111100001110100;
assign LUT_1[10519] = 32'b00000000000000000000110011110000;
assign LUT_1[10520] = 32'b00000000000000000011001000000001;
assign LUT_1[10521] = 32'b11111111111111111100011001111101;
assign LUT_1[10522] = 32'b11111111111111111110110110010010;
assign LUT_1[10523] = 32'b11111111111111111000001000001110;
assign LUT_1[10524] = 32'b00000000000000001011000001011000;
assign LUT_1[10525] = 32'b00000000000000000100010011010100;
assign LUT_1[10526] = 32'b00000000000000000110101111101001;
assign LUT_1[10527] = 32'b00000000000000000000000001100101;
assign LUT_1[10528] = 32'b00000000000000000010111001101001;
assign LUT_1[10529] = 32'b11111111111111111100001011100101;
assign LUT_1[10530] = 32'b11111111111111111110100111111010;
assign LUT_1[10531] = 32'b11111111111111110111111001110110;
assign LUT_1[10532] = 32'b00000000000000001010110011000000;
assign LUT_1[10533] = 32'b00000000000000000100000100111100;
assign LUT_1[10534] = 32'b00000000000000000110100001010001;
assign LUT_1[10535] = 32'b11111111111111111111110011001101;
assign LUT_1[10536] = 32'b00000000000000000010000111011110;
assign LUT_1[10537] = 32'b11111111111111111011011001011010;
assign LUT_1[10538] = 32'b11111111111111111101110101101111;
assign LUT_1[10539] = 32'b11111111111111110111000111101011;
assign LUT_1[10540] = 32'b00000000000000001010000000110101;
assign LUT_1[10541] = 32'b00000000000000000011010010110001;
assign LUT_1[10542] = 32'b00000000000000000101101111000110;
assign LUT_1[10543] = 32'b11111111111111111111000001000010;
assign LUT_1[10544] = 32'b00000000000000000100110101001011;
assign LUT_1[10545] = 32'b11111111111111111110000111000111;
assign LUT_1[10546] = 32'b00000000000000000000100011011100;
assign LUT_1[10547] = 32'b11111111111111111001110101011000;
assign LUT_1[10548] = 32'b00000000000000001100101110100010;
assign LUT_1[10549] = 32'b00000000000000000110000000011110;
assign LUT_1[10550] = 32'b00000000000000001000011100110011;
assign LUT_1[10551] = 32'b00000000000000000001101110101111;
assign LUT_1[10552] = 32'b00000000000000000100000011000000;
assign LUT_1[10553] = 32'b11111111111111111101010100111100;
assign LUT_1[10554] = 32'b11111111111111111111110001010001;
assign LUT_1[10555] = 32'b11111111111111111001000011001101;
assign LUT_1[10556] = 32'b00000000000000001011111100010111;
assign LUT_1[10557] = 32'b00000000000000000101001110010011;
assign LUT_1[10558] = 32'b00000000000000000111101010101000;
assign LUT_1[10559] = 32'b00000000000000000000111100100100;
assign LUT_1[10560] = 32'b00000000000000000011111100010010;
assign LUT_1[10561] = 32'b11111111111111111101001110001110;
assign LUT_1[10562] = 32'b11111111111111111111101010100011;
assign LUT_1[10563] = 32'b11111111111111111000111100011111;
assign LUT_1[10564] = 32'b00000000000000001011110101101001;
assign LUT_1[10565] = 32'b00000000000000000101000111100101;
assign LUT_1[10566] = 32'b00000000000000000111100011111010;
assign LUT_1[10567] = 32'b00000000000000000000110101110110;
assign LUT_1[10568] = 32'b00000000000000000011001010000111;
assign LUT_1[10569] = 32'b11111111111111111100011100000011;
assign LUT_1[10570] = 32'b11111111111111111110111000011000;
assign LUT_1[10571] = 32'b11111111111111111000001010010100;
assign LUT_1[10572] = 32'b00000000000000001011000011011110;
assign LUT_1[10573] = 32'b00000000000000000100010101011010;
assign LUT_1[10574] = 32'b00000000000000000110110001101111;
assign LUT_1[10575] = 32'b00000000000000000000000011101011;
assign LUT_1[10576] = 32'b00000000000000000101110111110100;
assign LUT_1[10577] = 32'b11111111111111111111001001110000;
assign LUT_1[10578] = 32'b00000000000000000001100110000101;
assign LUT_1[10579] = 32'b11111111111111111010111000000001;
assign LUT_1[10580] = 32'b00000000000000001101110001001011;
assign LUT_1[10581] = 32'b00000000000000000111000011000111;
assign LUT_1[10582] = 32'b00000000000000001001011111011100;
assign LUT_1[10583] = 32'b00000000000000000010110001011000;
assign LUT_1[10584] = 32'b00000000000000000101000101101001;
assign LUT_1[10585] = 32'b11111111111111111110010111100101;
assign LUT_1[10586] = 32'b00000000000000000000110011111010;
assign LUT_1[10587] = 32'b11111111111111111010000101110110;
assign LUT_1[10588] = 32'b00000000000000001100111111000000;
assign LUT_1[10589] = 32'b00000000000000000110010000111100;
assign LUT_1[10590] = 32'b00000000000000001000101101010001;
assign LUT_1[10591] = 32'b00000000000000000001111111001101;
assign LUT_1[10592] = 32'b00000000000000000100110111010001;
assign LUT_1[10593] = 32'b11111111111111111110001001001101;
assign LUT_1[10594] = 32'b00000000000000000000100101100010;
assign LUT_1[10595] = 32'b11111111111111111001110111011110;
assign LUT_1[10596] = 32'b00000000000000001100110000101000;
assign LUT_1[10597] = 32'b00000000000000000110000010100100;
assign LUT_1[10598] = 32'b00000000000000001000011110111001;
assign LUT_1[10599] = 32'b00000000000000000001110000110101;
assign LUT_1[10600] = 32'b00000000000000000100000101000110;
assign LUT_1[10601] = 32'b11111111111111111101010111000010;
assign LUT_1[10602] = 32'b11111111111111111111110011010111;
assign LUT_1[10603] = 32'b11111111111111111001000101010011;
assign LUT_1[10604] = 32'b00000000000000001011111110011101;
assign LUT_1[10605] = 32'b00000000000000000101010000011001;
assign LUT_1[10606] = 32'b00000000000000000111101100101110;
assign LUT_1[10607] = 32'b00000000000000000000111110101010;
assign LUT_1[10608] = 32'b00000000000000000110110010110011;
assign LUT_1[10609] = 32'b00000000000000000000000100101111;
assign LUT_1[10610] = 32'b00000000000000000010100001000100;
assign LUT_1[10611] = 32'b11111111111111111011110011000000;
assign LUT_1[10612] = 32'b00000000000000001110101100001010;
assign LUT_1[10613] = 32'b00000000000000000111111110000110;
assign LUT_1[10614] = 32'b00000000000000001010011010011011;
assign LUT_1[10615] = 32'b00000000000000000011101100010111;
assign LUT_1[10616] = 32'b00000000000000000110000000101000;
assign LUT_1[10617] = 32'b11111111111111111111010010100100;
assign LUT_1[10618] = 32'b00000000000000000001101110111001;
assign LUT_1[10619] = 32'b11111111111111111011000000110101;
assign LUT_1[10620] = 32'b00000000000000001101111001111111;
assign LUT_1[10621] = 32'b00000000000000000111001011111011;
assign LUT_1[10622] = 32'b00000000000000001001101000010000;
assign LUT_1[10623] = 32'b00000000000000000010111010001100;
assign LUT_1[10624] = 32'b00000000000000000100111110101101;
assign LUT_1[10625] = 32'b11111111111111111110010000101001;
assign LUT_1[10626] = 32'b00000000000000000000101100111110;
assign LUT_1[10627] = 32'b11111111111111111001111110111010;
assign LUT_1[10628] = 32'b00000000000000001100111000000100;
assign LUT_1[10629] = 32'b00000000000000000110001010000000;
assign LUT_1[10630] = 32'b00000000000000001000100110010101;
assign LUT_1[10631] = 32'b00000000000000000001111000010001;
assign LUT_1[10632] = 32'b00000000000000000100001100100010;
assign LUT_1[10633] = 32'b11111111111111111101011110011110;
assign LUT_1[10634] = 32'b11111111111111111111111010110011;
assign LUT_1[10635] = 32'b11111111111111111001001100101111;
assign LUT_1[10636] = 32'b00000000000000001100000101111001;
assign LUT_1[10637] = 32'b00000000000000000101010111110101;
assign LUT_1[10638] = 32'b00000000000000000111110100001010;
assign LUT_1[10639] = 32'b00000000000000000001000110000110;
assign LUT_1[10640] = 32'b00000000000000000110111010001111;
assign LUT_1[10641] = 32'b00000000000000000000001100001011;
assign LUT_1[10642] = 32'b00000000000000000010101000100000;
assign LUT_1[10643] = 32'b11111111111111111011111010011100;
assign LUT_1[10644] = 32'b00000000000000001110110011100110;
assign LUT_1[10645] = 32'b00000000000000001000000101100010;
assign LUT_1[10646] = 32'b00000000000000001010100001110111;
assign LUT_1[10647] = 32'b00000000000000000011110011110011;
assign LUT_1[10648] = 32'b00000000000000000110001000000100;
assign LUT_1[10649] = 32'b11111111111111111111011010000000;
assign LUT_1[10650] = 32'b00000000000000000001110110010101;
assign LUT_1[10651] = 32'b11111111111111111011001000010001;
assign LUT_1[10652] = 32'b00000000000000001110000001011011;
assign LUT_1[10653] = 32'b00000000000000000111010011010111;
assign LUT_1[10654] = 32'b00000000000000001001101111101100;
assign LUT_1[10655] = 32'b00000000000000000011000001101000;
assign LUT_1[10656] = 32'b00000000000000000101111001101100;
assign LUT_1[10657] = 32'b11111111111111111111001011101000;
assign LUT_1[10658] = 32'b00000000000000000001100111111101;
assign LUT_1[10659] = 32'b11111111111111111010111001111001;
assign LUT_1[10660] = 32'b00000000000000001101110011000011;
assign LUT_1[10661] = 32'b00000000000000000111000100111111;
assign LUT_1[10662] = 32'b00000000000000001001100001010100;
assign LUT_1[10663] = 32'b00000000000000000010110011010000;
assign LUT_1[10664] = 32'b00000000000000000101000111100001;
assign LUT_1[10665] = 32'b11111111111111111110011001011101;
assign LUT_1[10666] = 32'b00000000000000000000110101110010;
assign LUT_1[10667] = 32'b11111111111111111010000111101110;
assign LUT_1[10668] = 32'b00000000000000001101000000111000;
assign LUT_1[10669] = 32'b00000000000000000110010010110100;
assign LUT_1[10670] = 32'b00000000000000001000101111001001;
assign LUT_1[10671] = 32'b00000000000000000010000001000101;
assign LUT_1[10672] = 32'b00000000000000000111110101001110;
assign LUT_1[10673] = 32'b00000000000000000001000111001010;
assign LUT_1[10674] = 32'b00000000000000000011100011011111;
assign LUT_1[10675] = 32'b11111111111111111100110101011011;
assign LUT_1[10676] = 32'b00000000000000001111101110100101;
assign LUT_1[10677] = 32'b00000000000000001001000000100001;
assign LUT_1[10678] = 32'b00000000000000001011011100110110;
assign LUT_1[10679] = 32'b00000000000000000100101110110010;
assign LUT_1[10680] = 32'b00000000000000000111000011000011;
assign LUT_1[10681] = 32'b00000000000000000000010100111111;
assign LUT_1[10682] = 32'b00000000000000000010110001010100;
assign LUT_1[10683] = 32'b11111111111111111100000011010000;
assign LUT_1[10684] = 32'b00000000000000001110111100011010;
assign LUT_1[10685] = 32'b00000000000000001000001110010110;
assign LUT_1[10686] = 32'b00000000000000001010101010101011;
assign LUT_1[10687] = 32'b00000000000000000011111100100111;
assign LUT_1[10688] = 32'b00000000000000000110111100010101;
assign LUT_1[10689] = 32'b00000000000000000000001110010001;
assign LUT_1[10690] = 32'b00000000000000000010101010100110;
assign LUT_1[10691] = 32'b11111111111111111011111100100010;
assign LUT_1[10692] = 32'b00000000000000001110110101101100;
assign LUT_1[10693] = 32'b00000000000000001000000111101000;
assign LUT_1[10694] = 32'b00000000000000001010100011111101;
assign LUT_1[10695] = 32'b00000000000000000011110101111001;
assign LUT_1[10696] = 32'b00000000000000000110001010001010;
assign LUT_1[10697] = 32'b11111111111111111111011100000110;
assign LUT_1[10698] = 32'b00000000000000000001111000011011;
assign LUT_1[10699] = 32'b11111111111111111011001010010111;
assign LUT_1[10700] = 32'b00000000000000001110000011100001;
assign LUT_1[10701] = 32'b00000000000000000111010101011101;
assign LUT_1[10702] = 32'b00000000000000001001110001110010;
assign LUT_1[10703] = 32'b00000000000000000011000011101110;
assign LUT_1[10704] = 32'b00000000000000001000110111110111;
assign LUT_1[10705] = 32'b00000000000000000010001001110011;
assign LUT_1[10706] = 32'b00000000000000000100100110001000;
assign LUT_1[10707] = 32'b11111111111111111101111000000100;
assign LUT_1[10708] = 32'b00000000000000010000110001001110;
assign LUT_1[10709] = 32'b00000000000000001010000011001010;
assign LUT_1[10710] = 32'b00000000000000001100011111011111;
assign LUT_1[10711] = 32'b00000000000000000101110001011011;
assign LUT_1[10712] = 32'b00000000000000001000000101101100;
assign LUT_1[10713] = 32'b00000000000000000001010111101000;
assign LUT_1[10714] = 32'b00000000000000000011110011111101;
assign LUT_1[10715] = 32'b11111111111111111101000101111001;
assign LUT_1[10716] = 32'b00000000000000001111111111000011;
assign LUT_1[10717] = 32'b00000000000000001001010000111111;
assign LUT_1[10718] = 32'b00000000000000001011101101010100;
assign LUT_1[10719] = 32'b00000000000000000100111111010000;
assign LUT_1[10720] = 32'b00000000000000000111110111010100;
assign LUT_1[10721] = 32'b00000000000000000001001001010000;
assign LUT_1[10722] = 32'b00000000000000000011100101100101;
assign LUT_1[10723] = 32'b11111111111111111100110111100001;
assign LUT_1[10724] = 32'b00000000000000001111110000101011;
assign LUT_1[10725] = 32'b00000000000000001001000010100111;
assign LUT_1[10726] = 32'b00000000000000001011011110111100;
assign LUT_1[10727] = 32'b00000000000000000100110000111000;
assign LUT_1[10728] = 32'b00000000000000000111000101001001;
assign LUT_1[10729] = 32'b00000000000000000000010111000101;
assign LUT_1[10730] = 32'b00000000000000000010110011011010;
assign LUT_1[10731] = 32'b11111111111111111100000101010110;
assign LUT_1[10732] = 32'b00000000000000001110111110100000;
assign LUT_1[10733] = 32'b00000000000000001000010000011100;
assign LUT_1[10734] = 32'b00000000000000001010101100110001;
assign LUT_1[10735] = 32'b00000000000000000011111110101101;
assign LUT_1[10736] = 32'b00000000000000001001110010110110;
assign LUT_1[10737] = 32'b00000000000000000011000100110010;
assign LUT_1[10738] = 32'b00000000000000000101100001000111;
assign LUT_1[10739] = 32'b11111111111111111110110011000011;
assign LUT_1[10740] = 32'b00000000000000010001101100001101;
assign LUT_1[10741] = 32'b00000000000000001010111110001001;
assign LUT_1[10742] = 32'b00000000000000001101011010011110;
assign LUT_1[10743] = 32'b00000000000000000110101100011010;
assign LUT_1[10744] = 32'b00000000000000001001000000101011;
assign LUT_1[10745] = 32'b00000000000000000010010010100111;
assign LUT_1[10746] = 32'b00000000000000000100101110111100;
assign LUT_1[10747] = 32'b11111111111111111110000000111000;
assign LUT_1[10748] = 32'b00000000000000010000111010000010;
assign LUT_1[10749] = 32'b00000000000000001010001011111110;
assign LUT_1[10750] = 32'b00000000000000001100101000010011;
assign LUT_1[10751] = 32'b00000000000000000101111010001111;
assign LUT_1[10752] = 32'b11111111111111111101111000111011;
assign LUT_1[10753] = 32'b11111111111111110111001010110111;
assign LUT_1[10754] = 32'b11111111111111111001100111001100;
assign LUT_1[10755] = 32'b11111111111111110010111001001000;
assign LUT_1[10756] = 32'b00000000000000000101110010010010;
assign LUT_1[10757] = 32'b11111111111111111111000100001110;
assign LUT_1[10758] = 32'b00000000000000000001100000100011;
assign LUT_1[10759] = 32'b11111111111111111010110010011111;
assign LUT_1[10760] = 32'b11111111111111111101000110110000;
assign LUT_1[10761] = 32'b11111111111111110110011000101100;
assign LUT_1[10762] = 32'b11111111111111111000110101000001;
assign LUT_1[10763] = 32'b11111111111111110010000110111101;
assign LUT_1[10764] = 32'b00000000000000000101000000000111;
assign LUT_1[10765] = 32'b11111111111111111110010010000011;
assign LUT_1[10766] = 32'b00000000000000000000101110011000;
assign LUT_1[10767] = 32'b11111111111111111010000000010100;
assign LUT_1[10768] = 32'b11111111111111111111110100011101;
assign LUT_1[10769] = 32'b11111111111111111001000110011001;
assign LUT_1[10770] = 32'b11111111111111111011100010101110;
assign LUT_1[10771] = 32'b11111111111111110100110100101010;
assign LUT_1[10772] = 32'b00000000000000000111101101110100;
assign LUT_1[10773] = 32'b00000000000000000000111111110000;
assign LUT_1[10774] = 32'b00000000000000000011011100000101;
assign LUT_1[10775] = 32'b11111111111111111100101110000001;
assign LUT_1[10776] = 32'b11111111111111111111000010010010;
assign LUT_1[10777] = 32'b11111111111111111000010100001110;
assign LUT_1[10778] = 32'b11111111111111111010110000100011;
assign LUT_1[10779] = 32'b11111111111111110100000010011111;
assign LUT_1[10780] = 32'b00000000000000000110111011101001;
assign LUT_1[10781] = 32'b00000000000000000000001101100101;
assign LUT_1[10782] = 32'b00000000000000000010101001111010;
assign LUT_1[10783] = 32'b11111111111111111011111011110110;
assign LUT_1[10784] = 32'b11111111111111111110110011111010;
assign LUT_1[10785] = 32'b11111111111111111000000101110110;
assign LUT_1[10786] = 32'b11111111111111111010100010001011;
assign LUT_1[10787] = 32'b11111111111111110011110100000111;
assign LUT_1[10788] = 32'b00000000000000000110101101010001;
assign LUT_1[10789] = 32'b11111111111111111111111111001101;
assign LUT_1[10790] = 32'b00000000000000000010011011100010;
assign LUT_1[10791] = 32'b11111111111111111011101101011110;
assign LUT_1[10792] = 32'b11111111111111111110000001101111;
assign LUT_1[10793] = 32'b11111111111111110111010011101011;
assign LUT_1[10794] = 32'b11111111111111111001110000000000;
assign LUT_1[10795] = 32'b11111111111111110011000001111100;
assign LUT_1[10796] = 32'b00000000000000000101111011000110;
assign LUT_1[10797] = 32'b11111111111111111111001101000010;
assign LUT_1[10798] = 32'b00000000000000000001101001010111;
assign LUT_1[10799] = 32'b11111111111111111010111011010011;
assign LUT_1[10800] = 32'b00000000000000000000101111011100;
assign LUT_1[10801] = 32'b11111111111111111010000001011000;
assign LUT_1[10802] = 32'b11111111111111111100011101101101;
assign LUT_1[10803] = 32'b11111111111111110101101111101001;
assign LUT_1[10804] = 32'b00000000000000001000101000110011;
assign LUT_1[10805] = 32'b00000000000000000001111010101111;
assign LUT_1[10806] = 32'b00000000000000000100010111000100;
assign LUT_1[10807] = 32'b11111111111111111101101001000000;
assign LUT_1[10808] = 32'b11111111111111111111111101010001;
assign LUT_1[10809] = 32'b11111111111111111001001111001101;
assign LUT_1[10810] = 32'b11111111111111111011101011100010;
assign LUT_1[10811] = 32'b11111111111111110100111101011110;
assign LUT_1[10812] = 32'b00000000000000000111110110101000;
assign LUT_1[10813] = 32'b00000000000000000001001000100100;
assign LUT_1[10814] = 32'b00000000000000000011100100111001;
assign LUT_1[10815] = 32'b11111111111111111100110110110101;
assign LUT_1[10816] = 32'b11111111111111111111110110100011;
assign LUT_1[10817] = 32'b11111111111111111001001000011111;
assign LUT_1[10818] = 32'b11111111111111111011100100110100;
assign LUT_1[10819] = 32'b11111111111111110100110110110000;
assign LUT_1[10820] = 32'b00000000000000000111101111111010;
assign LUT_1[10821] = 32'b00000000000000000001000001110110;
assign LUT_1[10822] = 32'b00000000000000000011011110001011;
assign LUT_1[10823] = 32'b11111111111111111100110000000111;
assign LUT_1[10824] = 32'b11111111111111111111000100011000;
assign LUT_1[10825] = 32'b11111111111111111000010110010100;
assign LUT_1[10826] = 32'b11111111111111111010110010101001;
assign LUT_1[10827] = 32'b11111111111111110100000100100101;
assign LUT_1[10828] = 32'b00000000000000000110111101101111;
assign LUT_1[10829] = 32'b00000000000000000000001111101011;
assign LUT_1[10830] = 32'b00000000000000000010101100000000;
assign LUT_1[10831] = 32'b11111111111111111011111101111100;
assign LUT_1[10832] = 32'b00000000000000000001110010000101;
assign LUT_1[10833] = 32'b11111111111111111011000100000001;
assign LUT_1[10834] = 32'b11111111111111111101100000010110;
assign LUT_1[10835] = 32'b11111111111111110110110010010010;
assign LUT_1[10836] = 32'b00000000000000001001101011011100;
assign LUT_1[10837] = 32'b00000000000000000010111101011000;
assign LUT_1[10838] = 32'b00000000000000000101011001101101;
assign LUT_1[10839] = 32'b11111111111111111110101011101001;
assign LUT_1[10840] = 32'b00000000000000000000111111111010;
assign LUT_1[10841] = 32'b11111111111111111010010001110110;
assign LUT_1[10842] = 32'b11111111111111111100101110001011;
assign LUT_1[10843] = 32'b11111111111111110110000000000111;
assign LUT_1[10844] = 32'b00000000000000001000111001010001;
assign LUT_1[10845] = 32'b00000000000000000010001011001101;
assign LUT_1[10846] = 32'b00000000000000000100100111100010;
assign LUT_1[10847] = 32'b11111111111111111101111001011110;
assign LUT_1[10848] = 32'b00000000000000000000110001100010;
assign LUT_1[10849] = 32'b11111111111111111010000011011110;
assign LUT_1[10850] = 32'b11111111111111111100011111110011;
assign LUT_1[10851] = 32'b11111111111111110101110001101111;
assign LUT_1[10852] = 32'b00000000000000001000101010111001;
assign LUT_1[10853] = 32'b00000000000000000001111100110101;
assign LUT_1[10854] = 32'b00000000000000000100011001001010;
assign LUT_1[10855] = 32'b11111111111111111101101011000110;
assign LUT_1[10856] = 32'b11111111111111111111111111010111;
assign LUT_1[10857] = 32'b11111111111111111001010001010011;
assign LUT_1[10858] = 32'b11111111111111111011101101101000;
assign LUT_1[10859] = 32'b11111111111111110100111111100100;
assign LUT_1[10860] = 32'b00000000000000000111111000101110;
assign LUT_1[10861] = 32'b00000000000000000001001010101010;
assign LUT_1[10862] = 32'b00000000000000000011100110111111;
assign LUT_1[10863] = 32'b11111111111111111100111000111011;
assign LUT_1[10864] = 32'b00000000000000000010101101000100;
assign LUT_1[10865] = 32'b11111111111111111011111111000000;
assign LUT_1[10866] = 32'b11111111111111111110011011010101;
assign LUT_1[10867] = 32'b11111111111111110111101101010001;
assign LUT_1[10868] = 32'b00000000000000001010100110011011;
assign LUT_1[10869] = 32'b00000000000000000011111000010111;
assign LUT_1[10870] = 32'b00000000000000000110010100101100;
assign LUT_1[10871] = 32'b11111111111111111111100110101000;
assign LUT_1[10872] = 32'b00000000000000000001111010111001;
assign LUT_1[10873] = 32'b11111111111111111011001100110101;
assign LUT_1[10874] = 32'b11111111111111111101101001001010;
assign LUT_1[10875] = 32'b11111111111111110110111011000110;
assign LUT_1[10876] = 32'b00000000000000001001110100010000;
assign LUT_1[10877] = 32'b00000000000000000011000110001100;
assign LUT_1[10878] = 32'b00000000000000000101100010100001;
assign LUT_1[10879] = 32'b11111111111111111110110100011101;
assign LUT_1[10880] = 32'b00000000000000000000111000111110;
assign LUT_1[10881] = 32'b11111111111111111010001010111010;
assign LUT_1[10882] = 32'b11111111111111111100100111001111;
assign LUT_1[10883] = 32'b11111111111111110101111001001011;
assign LUT_1[10884] = 32'b00000000000000001000110010010101;
assign LUT_1[10885] = 32'b00000000000000000010000100010001;
assign LUT_1[10886] = 32'b00000000000000000100100000100110;
assign LUT_1[10887] = 32'b11111111111111111101110010100010;
assign LUT_1[10888] = 32'b00000000000000000000000110110011;
assign LUT_1[10889] = 32'b11111111111111111001011000101111;
assign LUT_1[10890] = 32'b11111111111111111011110101000100;
assign LUT_1[10891] = 32'b11111111111111110101000111000000;
assign LUT_1[10892] = 32'b00000000000000001000000000001010;
assign LUT_1[10893] = 32'b00000000000000000001010010000110;
assign LUT_1[10894] = 32'b00000000000000000011101110011011;
assign LUT_1[10895] = 32'b11111111111111111101000000010111;
assign LUT_1[10896] = 32'b00000000000000000010110100100000;
assign LUT_1[10897] = 32'b11111111111111111100000110011100;
assign LUT_1[10898] = 32'b11111111111111111110100010110001;
assign LUT_1[10899] = 32'b11111111111111110111110100101101;
assign LUT_1[10900] = 32'b00000000000000001010101101110111;
assign LUT_1[10901] = 32'b00000000000000000011111111110011;
assign LUT_1[10902] = 32'b00000000000000000110011100001000;
assign LUT_1[10903] = 32'b11111111111111111111101110000100;
assign LUT_1[10904] = 32'b00000000000000000010000010010101;
assign LUT_1[10905] = 32'b11111111111111111011010100010001;
assign LUT_1[10906] = 32'b11111111111111111101110000100110;
assign LUT_1[10907] = 32'b11111111111111110111000010100010;
assign LUT_1[10908] = 32'b00000000000000001001111011101100;
assign LUT_1[10909] = 32'b00000000000000000011001101101000;
assign LUT_1[10910] = 32'b00000000000000000101101001111101;
assign LUT_1[10911] = 32'b11111111111111111110111011111001;
assign LUT_1[10912] = 32'b00000000000000000001110011111101;
assign LUT_1[10913] = 32'b11111111111111111011000101111001;
assign LUT_1[10914] = 32'b11111111111111111101100010001110;
assign LUT_1[10915] = 32'b11111111111111110110110100001010;
assign LUT_1[10916] = 32'b00000000000000001001101101010100;
assign LUT_1[10917] = 32'b00000000000000000010111111010000;
assign LUT_1[10918] = 32'b00000000000000000101011011100101;
assign LUT_1[10919] = 32'b11111111111111111110101101100001;
assign LUT_1[10920] = 32'b00000000000000000001000001110010;
assign LUT_1[10921] = 32'b11111111111111111010010011101110;
assign LUT_1[10922] = 32'b11111111111111111100110000000011;
assign LUT_1[10923] = 32'b11111111111111110110000001111111;
assign LUT_1[10924] = 32'b00000000000000001000111011001001;
assign LUT_1[10925] = 32'b00000000000000000010001101000101;
assign LUT_1[10926] = 32'b00000000000000000100101001011010;
assign LUT_1[10927] = 32'b11111111111111111101111011010110;
assign LUT_1[10928] = 32'b00000000000000000011101111011111;
assign LUT_1[10929] = 32'b11111111111111111101000001011011;
assign LUT_1[10930] = 32'b11111111111111111111011101110000;
assign LUT_1[10931] = 32'b11111111111111111000101111101100;
assign LUT_1[10932] = 32'b00000000000000001011101000110110;
assign LUT_1[10933] = 32'b00000000000000000100111010110010;
assign LUT_1[10934] = 32'b00000000000000000111010111000111;
assign LUT_1[10935] = 32'b00000000000000000000101001000011;
assign LUT_1[10936] = 32'b00000000000000000010111101010100;
assign LUT_1[10937] = 32'b11111111111111111100001111010000;
assign LUT_1[10938] = 32'b11111111111111111110101011100101;
assign LUT_1[10939] = 32'b11111111111111110111111101100001;
assign LUT_1[10940] = 32'b00000000000000001010110110101011;
assign LUT_1[10941] = 32'b00000000000000000100001000100111;
assign LUT_1[10942] = 32'b00000000000000000110100100111100;
assign LUT_1[10943] = 32'b11111111111111111111110110111000;
assign LUT_1[10944] = 32'b00000000000000000010110110100110;
assign LUT_1[10945] = 32'b11111111111111111100001000100010;
assign LUT_1[10946] = 32'b11111111111111111110100100110111;
assign LUT_1[10947] = 32'b11111111111111110111110110110011;
assign LUT_1[10948] = 32'b00000000000000001010101111111101;
assign LUT_1[10949] = 32'b00000000000000000100000001111001;
assign LUT_1[10950] = 32'b00000000000000000110011110001110;
assign LUT_1[10951] = 32'b11111111111111111111110000001010;
assign LUT_1[10952] = 32'b00000000000000000010000100011011;
assign LUT_1[10953] = 32'b11111111111111111011010110010111;
assign LUT_1[10954] = 32'b11111111111111111101110010101100;
assign LUT_1[10955] = 32'b11111111111111110111000100101000;
assign LUT_1[10956] = 32'b00000000000000001001111101110010;
assign LUT_1[10957] = 32'b00000000000000000011001111101110;
assign LUT_1[10958] = 32'b00000000000000000101101100000011;
assign LUT_1[10959] = 32'b11111111111111111110111101111111;
assign LUT_1[10960] = 32'b00000000000000000100110010001000;
assign LUT_1[10961] = 32'b11111111111111111110000100000100;
assign LUT_1[10962] = 32'b00000000000000000000100000011001;
assign LUT_1[10963] = 32'b11111111111111111001110010010101;
assign LUT_1[10964] = 32'b00000000000000001100101011011111;
assign LUT_1[10965] = 32'b00000000000000000101111101011011;
assign LUT_1[10966] = 32'b00000000000000001000011001110000;
assign LUT_1[10967] = 32'b00000000000000000001101011101100;
assign LUT_1[10968] = 32'b00000000000000000011111111111101;
assign LUT_1[10969] = 32'b11111111111111111101010001111001;
assign LUT_1[10970] = 32'b11111111111111111111101110001110;
assign LUT_1[10971] = 32'b11111111111111111001000000001010;
assign LUT_1[10972] = 32'b00000000000000001011111001010100;
assign LUT_1[10973] = 32'b00000000000000000101001011010000;
assign LUT_1[10974] = 32'b00000000000000000111100111100101;
assign LUT_1[10975] = 32'b00000000000000000000111001100001;
assign LUT_1[10976] = 32'b00000000000000000011110001100101;
assign LUT_1[10977] = 32'b11111111111111111101000011100001;
assign LUT_1[10978] = 32'b11111111111111111111011111110110;
assign LUT_1[10979] = 32'b11111111111111111000110001110010;
assign LUT_1[10980] = 32'b00000000000000001011101010111100;
assign LUT_1[10981] = 32'b00000000000000000100111100111000;
assign LUT_1[10982] = 32'b00000000000000000111011001001101;
assign LUT_1[10983] = 32'b00000000000000000000101011001001;
assign LUT_1[10984] = 32'b00000000000000000010111111011010;
assign LUT_1[10985] = 32'b11111111111111111100010001010110;
assign LUT_1[10986] = 32'b11111111111111111110101101101011;
assign LUT_1[10987] = 32'b11111111111111110111111111100111;
assign LUT_1[10988] = 32'b00000000000000001010111000110001;
assign LUT_1[10989] = 32'b00000000000000000100001010101101;
assign LUT_1[10990] = 32'b00000000000000000110100111000010;
assign LUT_1[10991] = 32'b11111111111111111111111000111110;
assign LUT_1[10992] = 32'b00000000000000000101101101000111;
assign LUT_1[10993] = 32'b11111111111111111110111111000011;
assign LUT_1[10994] = 32'b00000000000000000001011011011000;
assign LUT_1[10995] = 32'b11111111111111111010101101010100;
assign LUT_1[10996] = 32'b00000000000000001101100110011110;
assign LUT_1[10997] = 32'b00000000000000000110111000011010;
assign LUT_1[10998] = 32'b00000000000000001001010100101111;
assign LUT_1[10999] = 32'b00000000000000000010100110101011;
assign LUT_1[11000] = 32'b00000000000000000100111010111100;
assign LUT_1[11001] = 32'b11111111111111111110001100111000;
assign LUT_1[11002] = 32'b00000000000000000000101001001101;
assign LUT_1[11003] = 32'b11111111111111111001111011001001;
assign LUT_1[11004] = 32'b00000000000000001100110100010011;
assign LUT_1[11005] = 32'b00000000000000000110000110001111;
assign LUT_1[11006] = 32'b00000000000000001000100010100100;
assign LUT_1[11007] = 32'b00000000000000000001110100100000;
assign LUT_1[11008] = 32'b11111111111111111011101101000111;
assign LUT_1[11009] = 32'b11111111111111110100111111000011;
assign LUT_1[11010] = 32'b11111111111111110111011011011000;
assign LUT_1[11011] = 32'b11111111111111110000101101010100;
assign LUT_1[11012] = 32'b00000000000000000011100110011110;
assign LUT_1[11013] = 32'b11111111111111111100111000011010;
assign LUT_1[11014] = 32'b11111111111111111111010100101111;
assign LUT_1[11015] = 32'b11111111111111111000100110101011;
assign LUT_1[11016] = 32'b11111111111111111010111010111100;
assign LUT_1[11017] = 32'b11111111111111110100001100111000;
assign LUT_1[11018] = 32'b11111111111111110110101001001101;
assign LUT_1[11019] = 32'b11111111111111101111111011001001;
assign LUT_1[11020] = 32'b00000000000000000010110100010011;
assign LUT_1[11021] = 32'b11111111111111111100000110001111;
assign LUT_1[11022] = 32'b11111111111111111110100010100100;
assign LUT_1[11023] = 32'b11111111111111110111110100100000;
assign LUT_1[11024] = 32'b11111111111111111101101000101001;
assign LUT_1[11025] = 32'b11111111111111110110111010100101;
assign LUT_1[11026] = 32'b11111111111111111001010110111010;
assign LUT_1[11027] = 32'b11111111111111110010101000110110;
assign LUT_1[11028] = 32'b00000000000000000101100010000000;
assign LUT_1[11029] = 32'b11111111111111111110110011111100;
assign LUT_1[11030] = 32'b00000000000000000001010000010001;
assign LUT_1[11031] = 32'b11111111111111111010100010001101;
assign LUT_1[11032] = 32'b11111111111111111100110110011110;
assign LUT_1[11033] = 32'b11111111111111110110001000011010;
assign LUT_1[11034] = 32'b11111111111111111000100100101111;
assign LUT_1[11035] = 32'b11111111111111110001110110101011;
assign LUT_1[11036] = 32'b00000000000000000100101111110101;
assign LUT_1[11037] = 32'b11111111111111111110000001110001;
assign LUT_1[11038] = 32'b00000000000000000000011110000110;
assign LUT_1[11039] = 32'b11111111111111111001110000000010;
assign LUT_1[11040] = 32'b11111111111111111100101000000110;
assign LUT_1[11041] = 32'b11111111111111110101111010000010;
assign LUT_1[11042] = 32'b11111111111111111000010110010111;
assign LUT_1[11043] = 32'b11111111111111110001101000010011;
assign LUT_1[11044] = 32'b00000000000000000100100001011101;
assign LUT_1[11045] = 32'b11111111111111111101110011011001;
assign LUT_1[11046] = 32'b00000000000000000000001111101110;
assign LUT_1[11047] = 32'b11111111111111111001100001101010;
assign LUT_1[11048] = 32'b11111111111111111011110101111011;
assign LUT_1[11049] = 32'b11111111111111110101000111110111;
assign LUT_1[11050] = 32'b11111111111111110111100100001100;
assign LUT_1[11051] = 32'b11111111111111110000110110001000;
assign LUT_1[11052] = 32'b00000000000000000011101111010010;
assign LUT_1[11053] = 32'b11111111111111111101000001001110;
assign LUT_1[11054] = 32'b11111111111111111111011101100011;
assign LUT_1[11055] = 32'b11111111111111111000101111011111;
assign LUT_1[11056] = 32'b11111111111111111110100011101000;
assign LUT_1[11057] = 32'b11111111111111110111110101100100;
assign LUT_1[11058] = 32'b11111111111111111010010001111001;
assign LUT_1[11059] = 32'b11111111111111110011100011110101;
assign LUT_1[11060] = 32'b00000000000000000110011100111111;
assign LUT_1[11061] = 32'b11111111111111111111101110111011;
assign LUT_1[11062] = 32'b00000000000000000010001011010000;
assign LUT_1[11063] = 32'b11111111111111111011011101001100;
assign LUT_1[11064] = 32'b11111111111111111101110001011101;
assign LUT_1[11065] = 32'b11111111111111110111000011011001;
assign LUT_1[11066] = 32'b11111111111111111001011111101110;
assign LUT_1[11067] = 32'b11111111111111110010110001101010;
assign LUT_1[11068] = 32'b00000000000000000101101010110100;
assign LUT_1[11069] = 32'b11111111111111111110111100110000;
assign LUT_1[11070] = 32'b00000000000000000001011001000101;
assign LUT_1[11071] = 32'b11111111111111111010101011000001;
assign LUT_1[11072] = 32'b11111111111111111101101010101111;
assign LUT_1[11073] = 32'b11111111111111110110111100101011;
assign LUT_1[11074] = 32'b11111111111111111001011001000000;
assign LUT_1[11075] = 32'b11111111111111110010101010111100;
assign LUT_1[11076] = 32'b00000000000000000101100100000110;
assign LUT_1[11077] = 32'b11111111111111111110110110000010;
assign LUT_1[11078] = 32'b00000000000000000001010010010111;
assign LUT_1[11079] = 32'b11111111111111111010100100010011;
assign LUT_1[11080] = 32'b11111111111111111100111000100100;
assign LUT_1[11081] = 32'b11111111111111110110001010100000;
assign LUT_1[11082] = 32'b11111111111111111000100110110101;
assign LUT_1[11083] = 32'b11111111111111110001111000110001;
assign LUT_1[11084] = 32'b00000000000000000100110001111011;
assign LUT_1[11085] = 32'b11111111111111111110000011110111;
assign LUT_1[11086] = 32'b00000000000000000000100000001100;
assign LUT_1[11087] = 32'b11111111111111111001110010001000;
assign LUT_1[11088] = 32'b11111111111111111111100110010001;
assign LUT_1[11089] = 32'b11111111111111111000111000001101;
assign LUT_1[11090] = 32'b11111111111111111011010100100010;
assign LUT_1[11091] = 32'b11111111111111110100100110011110;
assign LUT_1[11092] = 32'b00000000000000000111011111101000;
assign LUT_1[11093] = 32'b00000000000000000000110001100100;
assign LUT_1[11094] = 32'b00000000000000000011001101111001;
assign LUT_1[11095] = 32'b11111111111111111100011111110101;
assign LUT_1[11096] = 32'b11111111111111111110110100000110;
assign LUT_1[11097] = 32'b11111111111111111000000110000010;
assign LUT_1[11098] = 32'b11111111111111111010100010010111;
assign LUT_1[11099] = 32'b11111111111111110011110100010011;
assign LUT_1[11100] = 32'b00000000000000000110101101011101;
assign LUT_1[11101] = 32'b11111111111111111111111111011001;
assign LUT_1[11102] = 32'b00000000000000000010011011101110;
assign LUT_1[11103] = 32'b11111111111111111011101101101010;
assign LUT_1[11104] = 32'b11111111111111111110100101101110;
assign LUT_1[11105] = 32'b11111111111111110111110111101010;
assign LUT_1[11106] = 32'b11111111111111111010010011111111;
assign LUT_1[11107] = 32'b11111111111111110011100101111011;
assign LUT_1[11108] = 32'b00000000000000000110011111000101;
assign LUT_1[11109] = 32'b11111111111111111111110001000001;
assign LUT_1[11110] = 32'b00000000000000000010001101010110;
assign LUT_1[11111] = 32'b11111111111111111011011111010010;
assign LUT_1[11112] = 32'b11111111111111111101110011100011;
assign LUT_1[11113] = 32'b11111111111111110111000101011111;
assign LUT_1[11114] = 32'b11111111111111111001100001110100;
assign LUT_1[11115] = 32'b11111111111111110010110011110000;
assign LUT_1[11116] = 32'b00000000000000000101101100111010;
assign LUT_1[11117] = 32'b11111111111111111110111110110110;
assign LUT_1[11118] = 32'b00000000000000000001011011001011;
assign LUT_1[11119] = 32'b11111111111111111010101101000111;
assign LUT_1[11120] = 32'b00000000000000000000100001010000;
assign LUT_1[11121] = 32'b11111111111111111001110011001100;
assign LUT_1[11122] = 32'b11111111111111111100001111100001;
assign LUT_1[11123] = 32'b11111111111111110101100001011101;
assign LUT_1[11124] = 32'b00000000000000001000011010100111;
assign LUT_1[11125] = 32'b00000000000000000001101100100011;
assign LUT_1[11126] = 32'b00000000000000000100001000111000;
assign LUT_1[11127] = 32'b11111111111111111101011010110100;
assign LUT_1[11128] = 32'b11111111111111111111101111000101;
assign LUT_1[11129] = 32'b11111111111111111001000001000001;
assign LUT_1[11130] = 32'b11111111111111111011011101010110;
assign LUT_1[11131] = 32'b11111111111111110100101111010010;
assign LUT_1[11132] = 32'b00000000000000000111101000011100;
assign LUT_1[11133] = 32'b00000000000000000000111010011000;
assign LUT_1[11134] = 32'b00000000000000000011010110101101;
assign LUT_1[11135] = 32'b11111111111111111100101000101001;
assign LUT_1[11136] = 32'b11111111111111111110101101001010;
assign LUT_1[11137] = 32'b11111111111111110111111111000110;
assign LUT_1[11138] = 32'b11111111111111111010011011011011;
assign LUT_1[11139] = 32'b11111111111111110011101101010111;
assign LUT_1[11140] = 32'b00000000000000000110100110100001;
assign LUT_1[11141] = 32'b11111111111111111111111000011101;
assign LUT_1[11142] = 32'b00000000000000000010010100110010;
assign LUT_1[11143] = 32'b11111111111111111011100110101110;
assign LUT_1[11144] = 32'b11111111111111111101111010111111;
assign LUT_1[11145] = 32'b11111111111111110111001100111011;
assign LUT_1[11146] = 32'b11111111111111111001101001010000;
assign LUT_1[11147] = 32'b11111111111111110010111011001100;
assign LUT_1[11148] = 32'b00000000000000000101110100010110;
assign LUT_1[11149] = 32'b11111111111111111111000110010010;
assign LUT_1[11150] = 32'b00000000000000000001100010100111;
assign LUT_1[11151] = 32'b11111111111111111010110100100011;
assign LUT_1[11152] = 32'b00000000000000000000101000101100;
assign LUT_1[11153] = 32'b11111111111111111001111010101000;
assign LUT_1[11154] = 32'b11111111111111111100010110111101;
assign LUT_1[11155] = 32'b11111111111111110101101000111001;
assign LUT_1[11156] = 32'b00000000000000001000100010000011;
assign LUT_1[11157] = 32'b00000000000000000001110011111111;
assign LUT_1[11158] = 32'b00000000000000000100010000010100;
assign LUT_1[11159] = 32'b11111111111111111101100010010000;
assign LUT_1[11160] = 32'b11111111111111111111110110100001;
assign LUT_1[11161] = 32'b11111111111111111001001000011101;
assign LUT_1[11162] = 32'b11111111111111111011100100110010;
assign LUT_1[11163] = 32'b11111111111111110100110110101110;
assign LUT_1[11164] = 32'b00000000000000000111101111111000;
assign LUT_1[11165] = 32'b00000000000000000001000001110100;
assign LUT_1[11166] = 32'b00000000000000000011011110001001;
assign LUT_1[11167] = 32'b11111111111111111100110000000101;
assign LUT_1[11168] = 32'b11111111111111111111101000001001;
assign LUT_1[11169] = 32'b11111111111111111000111010000101;
assign LUT_1[11170] = 32'b11111111111111111011010110011010;
assign LUT_1[11171] = 32'b11111111111111110100101000010110;
assign LUT_1[11172] = 32'b00000000000000000111100001100000;
assign LUT_1[11173] = 32'b00000000000000000000110011011100;
assign LUT_1[11174] = 32'b00000000000000000011001111110001;
assign LUT_1[11175] = 32'b11111111111111111100100001101101;
assign LUT_1[11176] = 32'b11111111111111111110110101111110;
assign LUT_1[11177] = 32'b11111111111111111000000111111010;
assign LUT_1[11178] = 32'b11111111111111111010100100001111;
assign LUT_1[11179] = 32'b11111111111111110011110110001011;
assign LUT_1[11180] = 32'b00000000000000000110101111010101;
assign LUT_1[11181] = 32'b00000000000000000000000001010001;
assign LUT_1[11182] = 32'b00000000000000000010011101100110;
assign LUT_1[11183] = 32'b11111111111111111011101111100010;
assign LUT_1[11184] = 32'b00000000000000000001100011101011;
assign LUT_1[11185] = 32'b11111111111111111010110101100111;
assign LUT_1[11186] = 32'b11111111111111111101010001111100;
assign LUT_1[11187] = 32'b11111111111111110110100011111000;
assign LUT_1[11188] = 32'b00000000000000001001011101000010;
assign LUT_1[11189] = 32'b00000000000000000010101110111110;
assign LUT_1[11190] = 32'b00000000000000000101001011010011;
assign LUT_1[11191] = 32'b11111111111111111110011101001111;
assign LUT_1[11192] = 32'b00000000000000000000110001100000;
assign LUT_1[11193] = 32'b11111111111111111010000011011100;
assign LUT_1[11194] = 32'b11111111111111111100011111110001;
assign LUT_1[11195] = 32'b11111111111111110101110001101101;
assign LUT_1[11196] = 32'b00000000000000001000101010110111;
assign LUT_1[11197] = 32'b00000000000000000001111100110011;
assign LUT_1[11198] = 32'b00000000000000000100011001001000;
assign LUT_1[11199] = 32'b11111111111111111101101011000100;
assign LUT_1[11200] = 32'b00000000000000000000101010110010;
assign LUT_1[11201] = 32'b11111111111111111001111100101110;
assign LUT_1[11202] = 32'b11111111111111111100011001000011;
assign LUT_1[11203] = 32'b11111111111111110101101010111111;
assign LUT_1[11204] = 32'b00000000000000001000100100001001;
assign LUT_1[11205] = 32'b00000000000000000001110110000101;
assign LUT_1[11206] = 32'b00000000000000000100010010011010;
assign LUT_1[11207] = 32'b11111111111111111101100100010110;
assign LUT_1[11208] = 32'b11111111111111111111111000100111;
assign LUT_1[11209] = 32'b11111111111111111001001010100011;
assign LUT_1[11210] = 32'b11111111111111111011100110111000;
assign LUT_1[11211] = 32'b11111111111111110100111000110100;
assign LUT_1[11212] = 32'b00000000000000000111110001111110;
assign LUT_1[11213] = 32'b00000000000000000001000011111010;
assign LUT_1[11214] = 32'b00000000000000000011100000001111;
assign LUT_1[11215] = 32'b11111111111111111100110010001011;
assign LUT_1[11216] = 32'b00000000000000000010100110010100;
assign LUT_1[11217] = 32'b11111111111111111011111000010000;
assign LUT_1[11218] = 32'b11111111111111111110010100100101;
assign LUT_1[11219] = 32'b11111111111111110111100110100001;
assign LUT_1[11220] = 32'b00000000000000001010011111101011;
assign LUT_1[11221] = 32'b00000000000000000011110001100111;
assign LUT_1[11222] = 32'b00000000000000000110001101111100;
assign LUT_1[11223] = 32'b11111111111111111111011111111000;
assign LUT_1[11224] = 32'b00000000000000000001110100001001;
assign LUT_1[11225] = 32'b11111111111111111011000110000101;
assign LUT_1[11226] = 32'b11111111111111111101100010011010;
assign LUT_1[11227] = 32'b11111111111111110110110100010110;
assign LUT_1[11228] = 32'b00000000000000001001101101100000;
assign LUT_1[11229] = 32'b00000000000000000010111111011100;
assign LUT_1[11230] = 32'b00000000000000000101011011110001;
assign LUT_1[11231] = 32'b11111111111111111110101101101101;
assign LUT_1[11232] = 32'b00000000000000000001100101110001;
assign LUT_1[11233] = 32'b11111111111111111010110111101101;
assign LUT_1[11234] = 32'b11111111111111111101010100000010;
assign LUT_1[11235] = 32'b11111111111111110110100101111110;
assign LUT_1[11236] = 32'b00000000000000001001011111001000;
assign LUT_1[11237] = 32'b00000000000000000010110001000100;
assign LUT_1[11238] = 32'b00000000000000000101001101011001;
assign LUT_1[11239] = 32'b11111111111111111110011111010101;
assign LUT_1[11240] = 32'b00000000000000000000110011100110;
assign LUT_1[11241] = 32'b11111111111111111010000101100010;
assign LUT_1[11242] = 32'b11111111111111111100100001110111;
assign LUT_1[11243] = 32'b11111111111111110101110011110011;
assign LUT_1[11244] = 32'b00000000000000001000101100111101;
assign LUT_1[11245] = 32'b00000000000000000001111110111001;
assign LUT_1[11246] = 32'b00000000000000000100011011001110;
assign LUT_1[11247] = 32'b11111111111111111101101101001010;
assign LUT_1[11248] = 32'b00000000000000000011100001010011;
assign LUT_1[11249] = 32'b11111111111111111100110011001111;
assign LUT_1[11250] = 32'b11111111111111111111001111100100;
assign LUT_1[11251] = 32'b11111111111111111000100001100000;
assign LUT_1[11252] = 32'b00000000000000001011011010101010;
assign LUT_1[11253] = 32'b00000000000000000100101100100110;
assign LUT_1[11254] = 32'b00000000000000000111001000111011;
assign LUT_1[11255] = 32'b00000000000000000000011010110111;
assign LUT_1[11256] = 32'b00000000000000000010101111001000;
assign LUT_1[11257] = 32'b11111111111111111100000001000100;
assign LUT_1[11258] = 32'b11111111111111111110011101011001;
assign LUT_1[11259] = 32'b11111111111111110111101111010101;
assign LUT_1[11260] = 32'b00000000000000001010101000011111;
assign LUT_1[11261] = 32'b00000000000000000011111010011011;
assign LUT_1[11262] = 32'b00000000000000000110010110110000;
assign LUT_1[11263] = 32'b11111111111111111111101000101100;
assign LUT_1[11264] = 32'b00000000000000001010100001001110;
assign LUT_1[11265] = 32'b00000000000000000011110011001010;
assign LUT_1[11266] = 32'b00000000000000000110001111011111;
assign LUT_1[11267] = 32'b11111111111111111111100001011011;
assign LUT_1[11268] = 32'b00000000000000010010011010100101;
assign LUT_1[11269] = 32'b00000000000000001011101100100001;
assign LUT_1[11270] = 32'b00000000000000001110001000110110;
assign LUT_1[11271] = 32'b00000000000000000111011010110010;
assign LUT_1[11272] = 32'b00000000000000001001101111000011;
assign LUT_1[11273] = 32'b00000000000000000011000000111111;
assign LUT_1[11274] = 32'b00000000000000000101011101010100;
assign LUT_1[11275] = 32'b11111111111111111110101111010000;
assign LUT_1[11276] = 32'b00000000000000010001101000011010;
assign LUT_1[11277] = 32'b00000000000000001010111010010110;
assign LUT_1[11278] = 32'b00000000000000001101010110101011;
assign LUT_1[11279] = 32'b00000000000000000110101000100111;
assign LUT_1[11280] = 32'b00000000000000001100011100110000;
assign LUT_1[11281] = 32'b00000000000000000101101110101100;
assign LUT_1[11282] = 32'b00000000000000001000001011000001;
assign LUT_1[11283] = 32'b00000000000000000001011100111101;
assign LUT_1[11284] = 32'b00000000000000010100010110000111;
assign LUT_1[11285] = 32'b00000000000000001101101000000011;
assign LUT_1[11286] = 32'b00000000000000010000000100011000;
assign LUT_1[11287] = 32'b00000000000000001001010110010100;
assign LUT_1[11288] = 32'b00000000000000001011101010100101;
assign LUT_1[11289] = 32'b00000000000000000100111100100001;
assign LUT_1[11290] = 32'b00000000000000000111011000110110;
assign LUT_1[11291] = 32'b00000000000000000000101010110010;
assign LUT_1[11292] = 32'b00000000000000010011100011111100;
assign LUT_1[11293] = 32'b00000000000000001100110101111000;
assign LUT_1[11294] = 32'b00000000000000001111010010001101;
assign LUT_1[11295] = 32'b00000000000000001000100100001001;
assign LUT_1[11296] = 32'b00000000000000001011011100001101;
assign LUT_1[11297] = 32'b00000000000000000100101110001001;
assign LUT_1[11298] = 32'b00000000000000000111001010011110;
assign LUT_1[11299] = 32'b00000000000000000000011100011010;
assign LUT_1[11300] = 32'b00000000000000010011010101100100;
assign LUT_1[11301] = 32'b00000000000000001100100111100000;
assign LUT_1[11302] = 32'b00000000000000001111000011110101;
assign LUT_1[11303] = 32'b00000000000000001000010101110001;
assign LUT_1[11304] = 32'b00000000000000001010101010000010;
assign LUT_1[11305] = 32'b00000000000000000011111011111110;
assign LUT_1[11306] = 32'b00000000000000000110011000010011;
assign LUT_1[11307] = 32'b11111111111111111111101010001111;
assign LUT_1[11308] = 32'b00000000000000010010100011011001;
assign LUT_1[11309] = 32'b00000000000000001011110101010101;
assign LUT_1[11310] = 32'b00000000000000001110010001101010;
assign LUT_1[11311] = 32'b00000000000000000111100011100110;
assign LUT_1[11312] = 32'b00000000000000001101010111101111;
assign LUT_1[11313] = 32'b00000000000000000110101001101011;
assign LUT_1[11314] = 32'b00000000000000001001000110000000;
assign LUT_1[11315] = 32'b00000000000000000010010111111100;
assign LUT_1[11316] = 32'b00000000000000010101010001000110;
assign LUT_1[11317] = 32'b00000000000000001110100011000010;
assign LUT_1[11318] = 32'b00000000000000010000111111010111;
assign LUT_1[11319] = 32'b00000000000000001010010001010011;
assign LUT_1[11320] = 32'b00000000000000001100100101100100;
assign LUT_1[11321] = 32'b00000000000000000101110111100000;
assign LUT_1[11322] = 32'b00000000000000001000010011110101;
assign LUT_1[11323] = 32'b00000000000000000001100101110001;
assign LUT_1[11324] = 32'b00000000000000010100011110111011;
assign LUT_1[11325] = 32'b00000000000000001101110000110111;
assign LUT_1[11326] = 32'b00000000000000010000001101001100;
assign LUT_1[11327] = 32'b00000000000000001001011111001000;
assign LUT_1[11328] = 32'b00000000000000001100011110110110;
assign LUT_1[11329] = 32'b00000000000000000101110000110010;
assign LUT_1[11330] = 32'b00000000000000001000001101000111;
assign LUT_1[11331] = 32'b00000000000000000001011111000011;
assign LUT_1[11332] = 32'b00000000000000010100011000001101;
assign LUT_1[11333] = 32'b00000000000000001101101010001001;
assign LUT_1[11334] = 32'b00000000000000010000000110011110;
assign LUT_1[11335] = 32'b00000000000000001001011000011010;
assign LUT_1[11336] = 32'b00000000000000001011101100101011;
assign LUT_1[11337] = 32'b00000000000000000100111110100111;
assign LUT_1[11338] = 32'b00000000000000000111011010111100;
assign LUT_1[11339] = 32'b00000000000000000000101100111000;
assign LUT_1[11340] = 32'b00000000000000010011100110000010;
assign LUT_1[11341] = 32'b00000000000000001100110111111110;
assign LUT_1[11342] = 32'b00000000000000001111010100010011;
assign LUT_1[11343] = 32'b00000000000000001000100110001111;
assign LUT_1[11344] = 32'b00000000000000001110011010011000;
assign LUT_1[11345] = 32'b00000000000000000111101100010100;
assign LUT_1[11346] = 32'b00000000000000001010001000101001;
assign LUT_1[11347] = 32'b00000000000000000011011010100101;
assign LUT_1[11348] = 32'b00000000000000010110010011101111;
assign LUT_1[11349] = 32'b00000000000000001111100101101011;
assign LUT_1[11350] = 32'b00000000000000010010000010000000;
assign LUT_1[11351] = 32'b00000000000000001011010011111100;
assign LUT_1[11352] = 32'b00000000000000001101101000001101;
assign LUT_1[11353] = 32'b00000000000000000110111010001001;
assign LUT_1[11354] = 32'b00000000000000001001010110011110;
assign LUT_1[11355] = 32'b00000000000000000010101000011010;
assign LUT_1[11356] = 32'b00000000000000010101100001100100;
assign LUT_1[11357] = 32'b00000000000000001110110011100000;
assign LUT_1[11358] = 32'b00000000000000010001001111110101;
assign LUT_1[11359] = 32'b00000000000000001010100001110001;
assign LUT_1[11360] = 32'b00000000000000001101011001110101;
assign LUT_1[11361] = 32'b00000000000000000110101011110001;
assign LUT_1[11362] = 32'b00000000000000001001001000000110;
assign LUT_1[11363] = 32'b00000000000000000010011010000010;
assign LUT_1[11364] = 32'b00000000000000010101010011001100;
assign LUT_1[11365] = 32'b00000000000000001110100101001000;
assign LUT_1[11366] = 32'b00000000000000010001000001011101;
assign LUT_1[11367] = 32'b00000000000000001010010011011001;
assign LUT_1[11368] = 32'b00000000000000001100100111101010;
assign LUT_1[11369] = 32'b00000000000000000101111001100110;
assign LUT_1[11370] = 32'b00000000000000001000010101111011;
assign LUT_1[11371] = 32'b00000000000000000001100111110111;
assign LUT_1[11372] = 32'b00000000000000010100100001000001;
assign LUT_1[11373] = 32'b00000000000000001101110010111101;
assign LUT_1[11374] = 32'b00000000000000010000001111010010;
assign LUT_1[11375] = 32'b00000000000000001001100001001110;
assign LUT_1[11376] = 32'b00000000000000001111010101010111;
assign LUT_1[11377] = 32'b00000000000000001000100111010011;
assign LUT_1[11378] = 32'b00000000000000001011000011101000;
assign LUT_1[11379] = 32'b00000000000000000100010101100100;
assign LUT_1[11380] = 32'b00000000000000010111001110101110;
assign LUT_1[11381] = 32'b00000000000000010000100000101010;
assign LUT_1[11382] = 32'b00000000000000010010111100111111;
assign LUT_1[11383] = 32'b00000000000000001100001110111011;
assign LUT_1[11384] = 32'b00000000000000001110100011001100;
assign LUT_1[11385] = 32'b00000000000000000111110101001000;
assign LUT_1[11386] = 32'b00000000000000001010010001011101;
assign LUT_1[11387] = 32'b00000000000000000011100011011001;
assign LUT_1[11388] = 32'b00000000000000010110011100100011;
assign LUT_1[11389] = 32'b00000000000000001111101110011111;
assign LUT_1[11390] = 32'b00000000000000010010001010110100;
assign LUT_1[11391] = 32'b00000000000000001011011100110000;
assign LUT_1[11392] = 32'b00000000000000001101100001010001;
assign LUT_1[11393] = 32'b00000000000000000110110011001101;
assign LUT_1[11394] = 32'b00000000000000001001001111100010;
assign LUT_1[11395] = 32'b00000000000000000010100001011110;
assign LUT_1[11396] = 32'b00000000000000010101011010101000;
assign LUT_1[11397] = 32'b00000000000000001110101100100100;
assign LUT_1[11398] = 32'b00000000000000010001001000111001;
assign LUT_1[11399] = 32'b00000000000000001010011010110101;
assign LUT_1[11400] = 32'b00000000000000001100101111000110;
assign LUT_1[11401] = 32'b00000000000000000110000001000010;
assign LUT_1[11402] = 32'b00000000000000001000011101010111;
assign LUT_1[11403] = 32'b00000000000000000001101111010011;
assign LUT_1[11404] = 32'b00000000000000010100101000011101;
assign LUT_1[11405] = 32'b00000000000000001101111010011001;
assign LUT_1[11406] = 32'b00000000000000010000010110101110;
assign LUT_1[11407] = 32'b00000000000000001001101000101010;
assign LUT_1[11408] = 32'b00000000000000001111011100110011;
assign LUT_1[11409] = 32'b00000000000000001000101110101111;
assign LUT_1[11410] = 32'b00000000000000001011001011000100;
assign LUT_1[11411] = 32'b00000000000000000100011101000000;
assign LUT_1[11412] = 32'b00000000000000010111010110001010;
assign LUT_1[11413] = 32'b00000000000000010000101000000110;
assign LUT_1[11414] = 32'b00000000000000010011000100011011;
assign LUT_1[11415] = 32'b00000000000000001100010110010111;
assign LUT_1[11416] = 32'b00000000000000001110101010101000;
assign LUT_1[11417] = 32'b00000000000000000111111100100100;
assign LUT_1[11418] = 32'b00000000000000001010011000111001;
assign LUT_1[11419] = 32'b00000000000000000011101010110101;
assign LUT_1[11420] = 32'b00000000000000010110100011111111;
assign LUT_1[11421] = 32'b00000000000000001111110101111011;
assign LUT_1[11422] = 32'b00000000000000010010010010010000;
assign LUT_1[11423] = 32'b00000000000000001011100100001100;
assign LUT_1[11424] = 32'b00000000000000001110011100010000;
assign LUT_1[11425] = 32'b00000000000000000111101110001100;
assign LUT_1[11426] = 32'b00000000000000001010001010100001;
assign LUT_1[11427] = 32'b00000000000000000011011100011101;
assign LUT_1[11428] = 32'b00000000000000010110010101100111;
assign LUT_1[11429] = 32'b00000000000000001111100111100011;
assign LUT_1[11430] = 32'b00000000000000010010000011111000;
assign LUT_1[11431] = 32'b00000000000000001011010101110100;
assign LUT_1[11432] = 32'b00000000000000001101101010000101;
assign LUT_1[11433] = 32'b00000000000000000110111100000001;
assign LUT_1[11434] = 32'b00000000000000001001011000010110;
assign LUT_1[11435] = 32'b00000000000000000010101010010010;
assign LUT_1[11436] = 32'b00000000000000010101100011011100;
assign LUT_1[11437] = 32'b00000000000000001110110101011000;
assign LUT_1[11438] = 32'b00000000000000010001010001101101;
assign LUT_1[11439] = 32'b00000000000000001010100011101001;
assign LUT_1[11440] = 32'b00000000000000010000010111110010;
assign LUT_1[11441] = 32'b00000000000000001001101001101110;
assign LUT_1[11442] = 32'b00000000000000001100000110000011;
assign LUT_1[11443] = 32'b00000000000000000101010111111111;
assign LUT_1[11444] = 32'b00000000000000011000010001001001;
assign LUT_1[11445] = 32'b00000000000000010001100011000101;
assign LUT_1[11446] = 32'b00000000000000010011111111011010;
assign LUT_1[11447] = 32'b00000000000000001101010001010110;
assign LUT_1[11448] = 32'b00000000000000001111100101100111;
assign LUT_1[11449] = 32'b00000000000000001000110111100011;
assign LUT_1[11450] = 32'b00000000000000001011010011111000;
assign LUT_1[11451] = 32'b00000000000000000100100101110100;
assign LUT_1[11452] = 32'b00000000000000010111011110111110;
assign LUT_1[11453] = 32'b00000000000000010000110000111010;
assign LUT_1[11454] = 32'b00000000000000010011001101001111;
assign LUT_1[11455] = 32'b00000000000000001100011111001011;
assign LUT_1[11456] = 32'b00000000000000001111011110111001;
assign LUT_1[11457] = 32'b00000000000000001000110000110101;
assign LUT_1[11458] = 32'b00000000000000001011001101001010;
assign LUT_1[11459] = 32'b00000000000000000100011111000110;
assign LUT_1[11460] = 32'b00000000000000010111011000010000;
assign LUT_1[11461] = 32'b00000000000000010000101010001100;
assign LUT_1[11462] = 32'b00000000000000010011000110100001;
assign LUT_1[11463] = 32'b00000000000000001100011000011101;
assign LUT_1[11464] = 32'b00000000000000001110101100101110;
assign LUT_1[11465] = 32'b00000000000000000111111110101010;
assign LUT_1[11466] = 32'b00000000000000001010011010111111;
assign LUT_1[11467] = 32'b00000000000000000011101100111011;
assign LUT_1[11468] = 32'b00000000000000010110100110000101;
assign LUT_1[11469] = 32'b00000000000000001111111000000001;
assign LUT_1[11470] = 32'b00000000000000010010010100010110;
assign LUT_1[11471] = 32'b00000000000000001011100110010010;
assign LUT_1[11472] = 32'b00000000000000010001011010011011;
assign LUT_1[11473] = 32'b00000000000000001010101100010111;
assign LUT_1[11474] = 32'b00000000000000001101001000101100;
assign LUT_1[11475] = 32'b00000000000000000110011010101000;
assign LUT_1[11476] = 32'b00000000000000011001010011110010;
assign LUT_1[11477] = 32'b00000000000000010010100101101110;
assign LUT_1[11478] = 32'b00000000000000010101000010000011;
assign LUT_1[11479] = 32'b00000000000000001110010011111111;
assign LUT_1[11480] = 32'b00000000000000010000101000010000;
assign LUT_1[11481] = 32'b00000000000000001001111010001100;
assign LUT_1[11482] = 32'b00000000000000001100010110100001;
assign LUT_1[11483] = 32'b00000000000000000101101000011101;
assign LUT_1[11484] = 32'b00000000000000011000100001100111;
assign LUT_1[11485] = 32'b00000000000000010001110011100011;
assign LUT_1[11486] = 32'b00000000000000010100001111111000;
assign LUT_1[11487] = 32'b00000000000000001101100001110100;
assign LUT_1[11488] = 32'b00000000000000010000011001111000;
assign LUT_1[11489] = 32'b00000000000000001001101011110100;
assign LUT_1[11490] = 32'b00000000000000001100001000001001;
assign LUT_1[11491] = 32'b00000000000000000101011010000101;
assign LUT_1[11492] = 32'b00000000000000011000010011001111;
assign LUT_1[11493] = 32'b00000000000000010001100101001011;
assign LUT_1[11494] = 32'b00000000000000010100000001100000;
assign LUT_1[11495] = 32'b00000000000000001101010011011100;
assign LUT_1[11496] = 32'b00000000000000001111100111101101;
assign LUT_1[11497] = 32'b00000000000000001000111001101001;
assign LUT_1[11498] = 32'b00000000000000001011010101111110;
assign LUT_1[11499] = 32'b00000000000000000100100111111010;
assign LUT_1[11500] = 32'b00000000000000010111100001000100;
assign LUT_1[11501] = 32'b00000000000000010000110011000000;
assign LUT_1[11502] = 32'b00000000000000010011001111010101;
assign LUT_1[11503] = 32'b00000000000000001100100001010001;
assign LUT_1[11504] = 32'b00000000000000010010010101011010;
assign LUT_1[11505] = 32'b00000000000000001011100111010110;
assign LUT_1[11506] = 32'b00000000000000001110000011101011;
assign LUT_1[11507] = 32'b00000000000000000111010101100111;
assign LUT_1[11508] = 32'b00000000000000011010001110110001;
assign LUT_1[11509] = 32'b00000000000000010011100000101101;
assign LUT_1[11510] = 32'b00000000000000010101111101000010;
assign LUT_1[11511] = 32'b00000000000000001111001110111110;
assign LUT_1[11512] = 32'b00000000000000010001100011001111;
assign LUT_1[11513] = 32'b00000000000000001010110101001011;
assign LUT_1[11514] = 32'b00000000000000001101010001100000;
assign LUT_1[11515] = 32'b00000000000000000110100011011100;
assign LUT_1[11516] = 32'b00000000000000011001011100100110;
assign LUT_1[11517] = 32'b00000000000000010010101110100010;
assign LUT_1[11518] = 32'b00000000000000010101001010110111;
assign LUT_1[11519] = 32'b00000000000000001110011100110011;
assign LUT_1[11520] = 32'b00000000000000001000010101011010;
assign LUT_1[11521] = 32'b00000000000000000001100111010110;
assign LUT_1[11522] = 32'b00000000000000000100000011101011;
assign LUT_1[11523] = 32'b11111111111111111101010101100111;
assign LUT_1[11524] = 32'b00000000000000010000001110110001;
assign LUT_1[11525] = 32'b00000000000000001001100000101101;
assign LUT_1[11526] = 32'b00000000000000001011111101000010;
assign LUT_1[11527] = 32'b00000000000000000101001110111110;
assign LUT_1[11528] = 32'b00000000000000000111100011001111;
assign LUT_1[11529] = 32'b00000000000000000000110101001011;
assign LUT_1[11530] = 32'b00000000000000000011010001100000;
assign LUT_1[11531] = 32'b11111111111111111100100011011100;
assign LUT_1[11532] = 32'b00000000000000001111011100100110;
assign LUT_1[11533] = 32'b00000000000000001000101110100010;
assign LUT_1[11534] = 32'b00000000000000001011001010110111;
assign LUT_1[11535] = 32'b00000000000000000100011100110011;
assign LUT_1[11536] = 32'b00000000000000001010010000111100;
assign LUT_1[11537] = 32'b00000000000000000011100010111000;
assign LUT_1[11538] = 32'b00000000000000000101111111001101;
assign LUT_1[11539] = 32'b11111111111111111111010001001001;
assign LUT_1[11540] = 32'b00000000000000010010001010010011;
assign LUT_1[11541] = 32'b00000000000000001011011100001111;
assign LUT_1[11542] = 32'b00000000000000001101111000100100;
assign LUT_1[11543] = 32'b00000000000000000111001010100000;
assign LUT_1[11544] = 32'b00000000000000001001011110110001;
assign LUT_1[11545] = 32'b00000000000000000010110000101101;
assign LUT_1[11546] = 32'b00000000000000000101001101000010;
assign LUT_1[11547] = 32'b11111111111111111110011110111110;
assign LUT_1[11548] = 32'b00000000000000010001011000001000;
assign LUT_1[11549] = 32'b00000000000000001010101010000100;
assign LUT_1[11550] = 32'b00000000000000001101000110011001;
assign LUT_1[11551] = 32'b00000000000000000110011000010101;
assign LUT_1[11552] = 32'b00000000000000001001010000011001;
assign LUT_1[11553] = 32'b00000000000000000010100010010101;
assign LUT_1[11554] = 32'b00000000000000000100111110101010;
assign LUT_1[11555] = 32'b11111111111111111110010000100110;
assign LUT_1[11556] = 32'b00000000000000010001001001110000;
assign LUT_1[11557] = 32'b00000000000000001010011011101100;
assign LUT_1[11558] = 32'b00000000000000001100111000000001;
assign LUT_1[11559] = 32'b00000000000000000110001001111101;
assign LUT_1[11560] = 32'b00000000000000001000011110001110;
assign LUT_1[11561] = 32'b00000000000000000001110000001010;
assign LUT_1[11562] = 32'b00000000000000000100001100011111;
assign LUT_1[11563] = 32'b11111111111111111101011110011011;
assign LUT_1[11564] = 32'b00000000000000010000010111100101;
assign LUT_1[11565] = 32'b00000000000000001001101001100001;
assign LUT_1[11566] = 32'b00000000000000001100000101110110;
assign LUT_1[11567] = 32'b00000000000000000101010111110010;
assign LUT_1[11568] = 32'b00000000000000001011001011111011;
assign LUT_1[11569] = 32'b00000000000000000100011101110111;
assign LUT_1[11570] = 32'b00000000000000000110111010001100;
assign LUT_1[11571] = 32'b00000000000000000000001100001000;
assign LUT_1[11572] = 32'b00000000000000010011000101010010;
assign LUT_1[11573] = 32'b00000000000000001100010111001110;
assign LUT_1[11574] = 32'b00000000000000001110110011100011;
assign LUT_1[11575] = 32'b00000000000000001000000101011111;
assign LUT_1[11576] = 32'b00000000000000001010011001110000;
assign LUT_1[11577] = 32'b00000000000000000011101011101100;
assign LUT_1[11578] = 32'b00000000000000000110001000000001;
assign LUT_1[11579] = 32'b11111111111111111111011001111101;
assign LUT_1[11580] = 32'b00000000000000010010010011000111;
assign LUT_1[11581] = 32'b00000000000000001011100101000011;
assign LUT_1[11582] = 32'b00000000000000001110000001011000;
assign LUT_1[11583] = 32'b00000000000000000111010011010100;
assign LUT_1[11584] = 32'b00000000000000001010010011000010;
assign LUT_1[11585] = 32'b00000000000000000011100100111110;
assign LUT_1[11586] = 32'b00000000000000000110000001010011;
assign LUT_1[11587] = 32'b11111111111111111111010011001111;
assign LUT_1[11588] = 32'b00000000000000010010001100011001;
assign LUT_1[11589] = 32'b00000000000000001011011110010101;
assign LUT_1[11590] = 32'b00000000000000001101111010101010;
assign LUT_1[11591] = 32'b00000000000000000111001100100110;
assign LUT_1[11592] = 32'b00000000000000001001100000110111;
assign LUT_1[11593] = 32'b00000000000000000010110010110011;
assign LUT_1[11594] = 32'b00000000000000000101001111001000;
assign LUT_1[11595] = 32'b11111111111111111110100001000100;
assign LUT_1[11596] = 32'b00000000000000010001011010001110;
assign LUT_1[11597] = 32'b00000000000000001010101100001010;
assign LUT_1[11598] = 32'b00000000000000001101001000011111;
assign LUT_1[11599] = 32'b00000000000000000110011010011011;
assign LUT_1[11600] = 32'b00000000000000001100001110100100;
assign LUT_1[11601] = 32'b00000000000000000101100000100000;
assign LUT_1[11602] = 32'b00000000000000000111111100110101;
assign LUT_1[11603] = 32'b00000000000000000001001110110001;
assign LUT_1[11604] = 32'b00000000000000010100000111111011;
assign LUT_1[11605] = 32'b00000000000000001101011001110111;
assign LUT_1[11606] = 32'b00000000000000001111110110001100;
assign LUT_1[11607] = 32'b00000000000000001001001000001000;
assign LUT_1[11608] = 32'b00000000000000001011011100011001;
assign LUT_1[11609] = 32'b00000000000000000100101110010101;
assign LUT_1[11610] = 32'b00000000000000000111001010101010;
assign LUT_1[11611] = 32'b00000000000000000000011100100110;
assign LUT_1[11612] = 32'b00000000000000010011010101110000;
assign LUT_1[11613] = 32'b00000000000000001100100111101100;
assign LUT_1[11614] = 32'b00000000000000001111000100000001;
assign LUT_1[11615] = 32'b00000000000000001000010101111101;
assign LUT_1[11616] = 32'b00000000000000001011001110000001;
assign LUT_1[11617] = 32'b00000000000000000100011111111101;
assign LUT_1[11618] = 32'b00000000000000000110111100010010;
assign LUT_1[11619] = 32'b00000000000000000000001110001110;
assign LUT_1[11620] = 32'b00000000000000010011000111011000;
assign LUT_1[11621] = 32'b00000000000000001100011001010100;
assign LUT_1[11622] = 32'b00000000000000001110110101101001;
assign LUT_1[11623] = 32'b00000000000000001000000111100101;
assign LUT_1[11624] = 32'b00000000000000001010011011110110;
assign LUT_1[11625] = 32'b00000000000000000011101101110010;
assign LUT_1[11626] = 32'b00000000000000000110001010000111;
assign LUT_1[11627] = 32'b11111111111111111111011100000011;
assign LUT_1[11628] = 32'b00000000000000010010010101001101;
assign LUT_1[11629] = 32'b00000000000000001011100111001001;
assign LUT_1[11630] = 32'b00000000000000001110000011011110;
assign LUT_1[11631] = 32'b00000000000000000111010101011010;
assign LUT_1[11632] = 32'b00000000000000001101001001100011;
assign LUT_1[11633] = 32'b00000000000000000110011011011111;
assign LUT_1[11634] = 32'b00000000000000001000110111110100;
assign LUT_1[11635] = 32'b00000000000000000010001001110000;
assign LUT_1[11636] = 32'b00000000000000010101000010111010;
assign LUT_1[11637] = 32'b00000000000000001110010100110110;
assign LUT_1[11638] = 32'b00000000000000010000110001001011;
assign LUT_1[11639] = 32'b00000000000000001010000011000111;
assign LUT_1[11640] = 32'b00000000000000001100010111011000;
assign LUT_1[11641] = 32'b00000000000000000101101001010100;
assign LUT_1[11642] = 32'b00000000000000001000000101101001;
assign LUT_1[11643] = 32'b00000000000000000001010111100101;
assign LUT_1[11644] = 32'b00000000000000010100010000101111;
assign LUT_1[11645] = 32'b00000000000000001101100010101011;
assign LUT_1[11646] = 32'b00000000000000001111111111000000;
assign LUT_1[11647] = 32'b00000000000000001001010000111100;
assign LUT_1[11648] = 32'b00000000000000001011010101011101;
assign LUT_1[11649] = 32'b00000000000000000100100111011001;
assign LUT_1[11650] = 32'b00000000000000000111000011101110;
assign LUT_1[11651] = 32'b00000000000000000000010101101010;
assign LUT_1[11652] = 32'b00000000000000010011001110110100;
assign LUT_1[11653] = 32'b00000000000000001100100000110000;
assign LUT_1[11654] = 32'b00000000000000001110111101000101;
assign LUT_1[11655] = 32'b00000000000000001000001111000001;
assign LUT_1[11656] = 32'b00000000000000001010100011010010;
assign LUT_1[11657] = 32'b00000000000000000011110101001110;
assign LUT_1[11658] = 32'b00000000000000000110010001100011;
assign LUT_1[11659] = 32'b11111111111111111111100011011111;
assign LUT_1[11660] = 32'b00000000000000010010011100101001;
assign LUT_1[11661] = 32'b00000000000000001011101110100101;
assign LUT_1[11662] = 32'b00000000000000001110001010111010;
assign LUT_1[11663] = 32'b00000000000000000111011100110110;
assign LUT_1[11664] = 32'b00000000000000001101010000111111;
assign LUT_1[11665] = 32'b00000000000000000110100010111011;
assign LUT_1[11666] = 32'b00000000000000001000111111010000;
assign LUT_1[11667] = 32'b00000000000000000010010001001100;
assign LUT_1[11668] = 32'b00000000000000010101001010010110;
assign LUT_1[11669] = 32'b00000000000000001110011100010010;
assign LUT_1[11670] = 32'b00000000000000010000111000100111;
assign LUT_1[11671] = 32'b00000000000000001010001010100011;
assign LUT_1[11672] = 32'b00000000000000001100011110110100;
assign LUT_1[11673] = 32'b00000000000000000101110000110000;
assign LUT_1[11674] = 32'b00000000000000001000001101000101;
assign LUT_1[11675] = 32'b00000000000000000001011111000001;
assign LUT_1[11676] = 32'b00000000000000010100011000001011;
assign LUT_1[11677] = 32'b00000000000000001101101010000111;
assign LUT_1[11678] = 32'b00000000000000010000000110011100;
assign LUT_1[11679] = 32'b00000000000000001001011000011000;
assign LUT_1[11680] = 32'b00000000000000001100010000011100;
assign LUT_1[11681] = 32'b00000000000000000101100010011000;
assign LUT_1[11682] = 32'b00000000000000000111111110101101;
assign LUT_1[11683] = 32'b00000000000000000001010000101001;
assign LUT_1[11684] = 32'b00000000000000010100001001110011;
assign LUT_1[11685] = 32'b00000000000000001101011011101111;
assign LUT_1[11686] = 32'b00000000000000001111111000000100;
assign LUT_1[11687] = 32'b00000000000000001001001010000000;
assign LUT_1[11688] = 32'b00000000000000001011011110010001;
assign LUT_1[11689] = 32'b00000000000000000100110000001101;
assign LUT_1[11690] = 32'b00000000000000000111001100100010;
assign LUT_1[11691] = 32'b00000000000000000000011110011110;
assign LUT_1[11692] = 32'b00000000000000010011010111101000;
assign LUT_1[11693] = 32'b00000000000000001100101001100100;
assign LUT_1[11694] = 32'b00000000000000001111000101111001;
assign LUT_1[11695] = 32'b00000000000000001000010111110101;
assign LUT_1[11696] = 32'b00000000000000001110001011111110;
assign LUT_1[11697] = 32'b00000000000000000111011101111010;
assign LUT_1[11698] = 32'b00000000000000001001111010001111;
assign LUT_1[11699] = 32'b00000000000000000011001100001011;
assign LUT_1[11700] = 32'b00000000000000010110000101010101;
assign LUT_1[11701] = 32'b00000000000000001111010111010001;
assign LUT_1[11702] = 32'b00000000000000010001110011100110;
assign LUT_1[11703] = 32'b00000000000000001011000101100010;
assign LUT_1[11704] = 32'b00000000000000001101011001110011;
assign LUT_1[11705] = 32'b00000000000000000110101011101111;
assign LUT_1[11706] = 32'b00000000000000001001001000000100;
assign LUT_1[11707] = 32'b00000000000000000010011010000000;
assign LUT_1[11708] = 32'b00000000000000010101010011001010;
assign LUT_1[11709] = 32'b00000000000000001110100101000110;
assign LUT_1[11710] = 32'b00000000000000010001000001011011;
assign LUT_1[11711] = 32'b00000000000000001010010011010111;
assign LUT_1[11712] = 32'b00000000000000001101010011000101;
assign LUT_1[11713] = 32'b00000000000000000110100101000001;
assign LUT_1[11714] = 32'b00000000000000001001000001010110;
assign LUT_1[11715] = 32'b00000000000000000010010011010010;
assign LUT_1[11716] = 32'b00000000000000010101001100011100;
assign LUT_1[11717] = 32'b00000000000000001110011110011000;
assign LUT_1[11718] = 32'b00000000000000010000111010101101;
assign LUT_1[11719] = 32'b00000000000000001010001100101001;
assign LUT_1[11720] = 32'b00000000000000001100100000111010;
assign LUT_1[11721] = 32'b00000000000000000101110010110110;
assign LUT_1[11722] = 32'b00000000000000001000001111001011;
assign LUT_1[11723] = 32'b00000000000000000001100001000111;
assign LUT_1[11724] = 32'b00000000000000010100011010010001;
assign LUT_1[11725] = 32'b00000000000000001101101100001101;
assign LUT_1[11726] = 32'b00000000000000010000001000100010;
assign LUT_1[11727] = 32'b00000000000000001001011010011110;
assign LUT_1[11728] = 32'b00000000000000001111001110100111;
assign LUT_1[11729] = 32'b00000000000000001000100000100011;
assign LUT_1[11730] = 32'b00000000000000001010111100111000;
assign LUT_1[11731] = 32'b00000000000000000100001110110100;
assign LUT_1[11732] = 32'b00000000000000010111000111111110;
assign LUT_1[11733] = 32'b00000000000000010000011001111010;
assign LUT_1[11734] = 32'b00000000000000010010110110001111;
assign LUT_1[11735] = 32'b00000000000000001100001000001011;
assign LUT_1[11736] = 32'b00000000000000001110011100011100;
assign LUT_1[11737] = 32'b00000000000000000111101110011000;
assign LUT_1[11738] = 32'b00000000000000001010001010101101;
assign LUT_1[11739] = 32'b00000000000000000011011100101001;
assign LUT_1[11740] = 32'b00000000000000010110010101110011;
assign LUT_1[11741] = 32'b00000000000000001111100111101111;
assign LUT_1[11742] = 32'b00000000000000010010000100000100;
assign LUT_1[11743] = 32'b00000000000000001011010110000000;
assign LUT_1[11744] = 32'b00000000000000001110001110000100;
assign LUT_1[11745] = 32'b00000000000000000111100000000000;
assign LUT_1[11746] = 32'b00000000000000001001111100010101;
assign LUT_1[11747] = 32'b00000000000000000011001110010001;
assign LUT_1[11748] = 32'b00000000000000010110000111011011;
assign LUT_1[11749] = 32'b00000000000000001111011001010111;
assign LUT_1[11750] = 32'b00000000000000010001110101101100;
assign LUT_1[11751] = 32'b00000000000000001011000111101000;
assign LUT_1[11752] = 32'b00000000000000001101011011111001;
assign LUT_1[11753] = 32'b00000000000000000110101101110101;
assign LUT_1[11754] = 32'b00000000000000001001001010001010;
assign LUT_1[11755] = 32'b00000000000000000010011100000110;
assign LUT_1[11756] = 32'b00000000000000010101010101010000;
assign LUT_1[11757] = 32'b00000000000000001110100111001100;
assign LUT_1[11758] = 32'b00000000000000010001000011100001;
assign LUT_1[11759] = 32'b00000000000000001010010101011101;
assign LUT_1[11760] = 32'b00000000000000010000001001100110;
assign LUT_1[11761] = 32'b00000000000000001001011011100010;
assign LUT_1[11762] = 32'b00000000000000001011110111110111;
assign LUT_1[11763] = 32'b00000000000000000101001001110011;
assign LUT_1[11764] = 32'b00000000000000011000000010111101;
assign LUT_1[11765] = 32'b00000000000000010001010100111001;
assign LUT_1[11766] = 32'b00000000000000010011110001001110;
assign LUT_1[11767] = 32'b00000000000000001101000011001010;
assign LUT_1[11768] = 32'b00000000000000001111010111011011;
assign LUT_1[11769] = 32'b00000000000000001000101001010111;
assign LUT_1[11770] = 32'b00000000000000001011000101101100;
assign LUT_1[11771] = 32'b00000000000000000100010111101000;
assign LUT_1[11772] = 32'b00000000000000010111010000110010;
assign LUT_1[11773] = 32'b00000000000000010000100010101110;
assign LUT_1[11774] = 32'b00000000000000010010111111000011;
assign LUT_1[11775] = 32'b00000000000000001100010000111111;
assign LUT_1[11776] = 32'b00000000000000000100001111101011;
assign LUT_1[11777] = 32'b11111111111111111101100001100111;
assign LUT_1[11778] = 32'b11111111111111111111111101111100;
assign LUT_1[11779] = 32'b11111111111111111001001111111000;
assign LUT_1[11780] = 32'b00000000000000001100001001000010;
assign LUT_1[11781] = 32'b00000000000000000101011010111110;
assign LUT_1[11782] = 32'b00000000000000000111110111010011;
assign LUT_1[11783] = 32'b00000000000000000001001001001111;
assign LUT_1[11784] = 32'b00000000000000000011011101100000;
assign LUT_1[11785] = 32'b11111111111111111100101111011100;
assign LUT_1[11786] = 32'b11111111111111111111001011110001;
assign LUT_1[11787] = 32'b11111111111111111000011101101101;
assign LUT_1[11788] = 32'b00000000000000001011010110110111;
assign LUT_1[11789] = 32'b00000000000000000100101000110011;
assign LUT_1[11790] = 32'b00000000000000000111000101001000;
assign LUT_1[11791] = 32'b00000000000000000000010111000100;
assign LUT_1[11792] = 32'b00000000000000000110001011001101;
assign LUT_1[11793] = 32'b11111111111111111111011101001001;
assign LUT_1[11794] = 32'b00000000000000000001111001011110;
assign LUT_1[11795] = 32'b11111111111111111011001011011010;
assign LUT_1[11796] = 32'b00000000000000001110000100100100;
assign LUT_1[11797] = 32'b00000000000000000111010110100000;
assign LUT_1[11798] = 32'b00000000000000001001110010110101;
assign LUT_1[11799] = 32'b00000000000000000011000100110001;
assign LUT_1[11800] = 32'b00000000000000000101011001000010;
assign LUT_1[11801] = 32'b11111111111111111110101010111110;
assign LUT_1[11802] = 32'b00000000000000000001000111010011;
assign LUT_1[11803] = 32'b11111111111111111010011001001111;
assign LUT_1[11804] = 32'b00000000000000001101010010011001;
assign LUT_1[11805] = 32'b00000000000000000110100100010101;
assign LUT_1[11806] = 32'b00000000000000001001000000101010;
assign LUT_1[11807] = 32'b00000000000000000010010010100110;
assign LUT_1[11808] = 32'b00000000000000000101001010101010;
assign LUT_1[11809] = 32'b11111111111111111110011100100110;
assign LUT_1[11810] = 32'b00000000000000000000111000111011;
assign LUT_1[11811] = 32'b11111111111111111010001010110111;
assign LUT_1[11812] = 32'b00000000000000001101000100000001;
assign LUT_1[11813] = 32'b00000000000000000110010101111101;
assign LUT_1[11814] = 32'b00000000000000001000110010010010;
assign LUT_1[11815] = 32'b00000000000000000010000100001110;
assign LUT_1[11816] = 32'b00000000000000000100011000011111;
assign LUT_1[11817] = 32'b11111111111111111101101010011011;
assign LUT_1[11818] = 32'b00000000000000000000000110110000;
assign LUT_1[11819] = 32'b11111111111111111001011000101100;
assign LUT_1[11820] = 32'b00000000000000001100010001110110;
assign LUT_1[11821] = 32'b00000000000000000101100011110010;
assign LUT_1[11822] = 32'b00000000000000001000000000000111;
assign LUT_1[11823] = 32'b00000000000000000001010010000011;
assign LUT_1[11824] = 32'b00000000000000000111000110001100;
assign LUT_1[11825] = 32'b00000000000000000000011000001000;
assign LUT_1[11826] = 32'b00000000000000000010110100011101;
assign LUT_1[11827] = 32'b11111111111111111100000110011001;
assign LUT_1[11828] = 32'b00000000000000001110111111100011;
assign LUT_1[11829] = 32'b00000000000000001000010001011111;
assign LUT_1[11830] = 32'b00000000000000001010101101110100;
assign LUT_1[11831] = 32'b00000000000000000011111111110000;
assign LUT_1[11832] = 32'b00000000000000000110010100000001;
assign LUT_1[11833] = 32'b11111111111111111111100101111101;
assign LUT_1[11834] = 32'b00000000000000000010000010010010;
assign LUT_1[11835] = 32'b11111111111111111011010100001110;
assign LUT_1[11836] = 32'b00000000000000001110001101011000;
assign LUT_1[11837] = 32'b00000000000000000111011111010100;
assign LUT_1[11838] = 32'b00000000000000001001111011101001;
assign LUT_1[11839] = 32'b00000000000000000011001101100101;
assign LUT_1[11840] = 32'b00000000000000000110001101010011;
assign LUT_1[11841] = 32'b11111111111111111111011111001111;
assign LUT_1[11842] = 32'b00000000000000000001111011100100;
assign LUT_1[11843] = 32'b11111111111111111011001101100000;
assign LUT_1[11844] = 32'b00000000000000001110000110101010;
assign LUT_1[11845] = 32'b00000000000000000111011000100110;
assign LUT_1[11846] = 32'b00000000000000001001110100111011;
assign LUT_1[11847] = 32'b00000000000000000011000110110111;
assign LUT_1[11848] = 32'b00000000000000000101011011001000;
assign LUT_1[11849] = 32'b11111111111111111110101101000100;
assign LUT_1[11850] = 32'b00000000000000000001001001011001;
assign LUT_1[11851] = 32'b11111111111111111010011011010101;
assign LUT_1[11852] = 32'b00000000000000001101010100011111;
assign LUT_1[11853] = 32'b00000000000000000110100110011011;
assign LUT_1[11854] = 32'b00000000000000001001000010110000;
assign LUT_1[11855] = 32'b00000000000000000010010100101100;
assign LUT_1[11856] = 32'b00000000000000001000001000110101;
assign LUT_1[11857] = 32'b00000000000000000001011010110001;
assign LUT_1[11858] = 32'b00000000000000000011110111000110;
assign LUT_1[11859] = 32'b11111111111111111101001001000010;
assign LUT_1[11860] = 32'b00000000000000010000000010001100;
assign LUT_1[11861] = 32'b00000000000000001001010100001000;
assign LUT_1[11862] = 32'b00000000000000001011110000011101;
assign LUT_1[11863] = 32'b00000000000000000101000010011001;
assign LUT_1[11864] = 32'b00000000000000000111010110101010;
assign LUT_1[11865] = 32'b00000000000000000000101000100110;
assign LUT_1[11866] = 32'b00000000000000000011000100111011;
assign LUT_1[11867] = 32'b11111111111111111100010110110111;
assign LUT_1[11868] = 32'b00000000000000001111010000000001;
assign LUT_1[11869] = 32'b00000000000000001000100001111101;
assign LUT_1[11870] = 32'b00000000000000001010111110010010;
assign LUT_1[11871] = 32'b00000000000000000100010000001110;
assign LUT_1[11872] = 32'b00000000000000000111001000010010;
assign LUT_1[11873] = 32'b00000000000000000000011010001110;
assign LUT_1[11874] = 32'b00000000000000000010110110100011;
assign LUT_1[11875] = 32'b11111111111111111100001000011111;
assign LUT_1[11876] = 32'b00000000000000001111000001101001;
assign LUT_1[11877] = 32'b00000000000000001000010011100101;
assign LUT_1[11878] = 32'b00000000000000001010101111111010;
assign LUT_1[11879] = 32'b00000000000000000100000001110110;
assign LUT_1[11880] = 32'b00000000000000000110010110000111;
assign LUT_1[11881] = 32'b11111111111111111111101000000011;
assign LUT_1[11882] = 32'b00000000000000000010000100011000;
assign LUT_1[11883] = 32'b11111111111111111011010110010100;
assign LUT_1[11884] = 32'b00000000000000001110001111011110;
assign LUT_1[11885] = 32'b00000000000000000111100001011010;
assign LUT_1[11886] = 32'b00000000000000001001111101101111;
assign LUT_1[11887] = 32'b00000000000000000011001111101011;
assign LUT_1[11888] = 32'b00000000000000001001000011110100;
assign LUT_1[11889] = 32'b00000000000000000010010101110000;
assign LUT_1[11890] = 32'b00000000000000000100110010000101;
assign LUT_1[11891] = 32'b11111111111111111110000100000001;
assign LUT_1[11892] = 32'b00000000000000010000111101001011;
assign LUT_1[11893] = 32'b00000000000000001010001111000111;
assign LUT_1[11894] = 32'b00000000000000001100101011011100;
assign LUT_1[11895] = 32'b00000000000000000101111101011000;
assign LUT_1[11896] = 32'b00000000000000001000010001101001;
assign LUT_1[11897] = 32'b00000000000000000001100011100101;
assign LUT_1[11898] = 32'b00000000000000000011111111111010;
assign LUT_1[11899] = 32'b11111111111111111101010001110110;
assign LUT_1[11900] = 32'b00000000000000010000001011000000;
assign LUT_1[11901] = 32'b00000000000000001001011100111100;
assign LUT_1[11902] = 32'b00000000000000001011111001010001;
assign LUT_1[11903] = 32'b00000000000000000101001011001101;
assign LUT_1[11904] = 32'b00000000000000000111001111101110;
assign LUT_1[11905] = 32'b00000000000000000000100001101010;
assign LUT_1[11906] = 32'b00000000000000000010111101111111;
assign LUT_1[11907] = 32'b11111111111111111100001111111011;
assign LUT_1[11908] = 32'b00000000000000001111001001000101;
assign LUT_1[11909] = 32'b00000000000000001000011011000001;
assign LUT_1[11910] = 32'b00000000000000001010110111010110;
assign LUT_1[11911] = 32'b00000000000000000100001001010010;
assign LUT_1[11912] = 32'b00000000000000000110011101100011;
assign LUT_1[11913] = 32'b11111111111111111111101111011111;
assign LUT_1[11914] = 32'b00000000000000000010001011110100;
assign LUT_1[11915] = 32'b11111111111111111011011101110000;
assign LUT_1[11916] = 32'b00000000000000001110010110111010;
assign LUT_1[11917] = 32'b00000000000000000111101000110110;
assign LUT_1[11918] = 32'b00000000000000001010000101001011;
assign LUT_1[11919] = 32'b00000000000000000011010111000111;
assign LUT_1[11920] = 32'b00000000000000001001001011010000;
assign LUT_1[11921] = 32'b00000000000000000010011101001100;
assign LUT_1[11922] = 32'b00000000000000000100111001100001;
assign LUT_1[11923] = 32'b11111111111111111110001011011101;
assign LUT_1[11924] = 32'b00000000000000010001000100100111;
assign LUT_1[11925] = 32'b00000000000000001010010110100011;
assign LUT_1[11926] = 32'b00000000000000001100110010111000;
assign LUT_1[11927] = 32'b00000000000000000110000100110100;
assign LUT_1[11928] = 32'b00000000000000001000011001000101;
assign LUT_1[11929] = 32'b00000000000000000001101011000001;
assign LUT_1[11930] = 32'b00000000000000000100000111010110;
assign LUT_1[11931] = 32'b11111111111111111101011001010010;
assign LUT_1[11932] = 32'b00000000000000010000010010011100;
assign LUT_1[11933] = 32'b00000000000000001001100100011000;
assign LUT_1[11934] = 32'b00000000000000001100000000101101;
assign LUT_1[11935] = 32'b00000000000000000101010010101001;
assign LUT_1[11936] = 32'b00000000000000001000001010101101;
assign LUT_1[11937] = 32'b00000000000000000001011100101001;
assign LUT_1[11938] = 32'b00000000000000000011111000111110;
assign LUT_1[11939] = 32'b11111111111111111101001010111010;
assign LUT_1[11940] = 32'b00000000000000010000000100000100;
assign LUT_1[11941] = 32'b00000000000000001001010110000000;
assign LUT_1[11942] = 32'b00000000000000001011110010010101;
assign LUT_1[11943] = 32'b00000000000000000101000100010001;
assign LUT_1[11944] = 32'b00000000000000000111011000100010;
assign LUT_1[11945] = 32'b00000000000000000000101010011110;
assign LUT_1[11946] = 32'b00000000000000000011000110110011;
assign LUT_1[11947] = 32'b11111111111111111100011000101111;
assign LUT_1[11948] = 32'b00000000000000001111010001111001;
assign LUT_1[11949] = 32'b00000000000000001000100011110101;
assign LUT_1[11950] = 32'b00000000000000001011000000001010;
assign LUT_1[11951] = 32'b00000000000000000100010010000110;
assign LUT_1[11952] = 32'b00000000000000001010000110001111;
assign LUT_1[11953] = 32'b00000000000000000011011000001011;
assign LUT_1[11954] = 32'b00000000000000000101110100100000;
assign LUT_1[11955] = 32'b11111111111111111111000110011100;
assign LUT_1[11956] = 32'b00000000000000010001111111100110;
assign LUT_1[11957] = 32'b00000000000000001011010001100010;
assign LUT_1[11958] = 32'b00000000000000001101101101110111;
assign LUT_1[11959] = 32'b00000000000000000110111111110011;
assign LUT_1[11960] = 32'b00000000000000001001010100000100;
assign LUT_1[11961] = 32'b00000000000000000010100110000000;
assign LUT_1[11962] = 32'b00000000000000000101000010010101;
assign LUT_1[11963] = 32'b11111111111111111110010100010001;
assign LUT_1[11964] = 32'b00000000000000010001001101011011;
assign LUT_1[11965] = 32'b00000000000000001010011111010111;
assign LUT_1[11966] = 32'b00000000000000001100111011101100;
assign LUT_1[11967] = 32'b00000000000000000110001101101000;
assign LUT_1[11968] = 32'b00000000000000001001001101010110;
assign LUT_1[11969] = 32'b00000000000000000010011111010010;
assign LUT_1[11970] = 32'b00000000000000000100111011100111;
assign LUT_1[11971] = 32'b11111111111111111110001101100011;
assign LUT_1[11972] = 32'b00000000000000010001000110101101;
assign LUT_1[11973] = 32'b00000000000000001010011000101001;
assign LUT_1[11974] = 32'b00000000000000001100110100111110;
assign LUT_1[11975] = 32'b00000000000000000110000110111010;
assign LUT_1[11976] = 32'b00000000000000001000011011001011;
assign LUT_1[11977] = 32'b00000000000000000001101101000111;
assign LUT_1[11978] = 32'b00000000000000000100001001011100;
assign LUT_1[11979] = 32'b11111111111111111101011011011000;
assign LUT_1[11980] = 32'b00000000000000010000010100100010;
assign LUT_1[11981] = 32'b00000000000000001001100110011110;
assign LUT_1[11982] = 32'b00000000000000001100000010110011;
assign LUT_1[11983] = 32'b00000000000000000101010100101111;
assign LUT_1[11984] = 32'b00000000000000001011001000111000;
assign LUT_1[11985] = 32'b00000000000000000100011010110100;
assign LUT_1[11986] = 32'b00000000000000000110110111001001;
assign LUT_1[11987] = 32'b00000000000000000000001001000101;
assign LUT_1[11988] = 32'b00000000000000010011000010001111;
assign LUT_1[11989] = 32'b00000000000000001100010100001011;
assign LUT_1[11990] = 32'b00000000000000001110110000100000;
assign LUT_1[11991] = 32'b00000000000000001000000010011100;
assign LUT_1[11992] = 32'b00000000000000001010010110101101;
assign LUT_1[11993] = 32'b00000000000000000011101000101001;
assign LUT_1[11994] = 32'b00000000000000000110000100111110;
assign LUT_1[11995] = 32'b11111111111111111111010110111010;
assign LUT_1[11996] = 32'b00000000000000010010010000000100;
assign LUT_1[11997] = 32'b00000000000000001011100010000000;
assign LUT_1[11998] = 32'b00000000000000001101111110010101;
assign LUT_1[11999] = 32'b00000000000000000111010000010001;
assign LUT_1[12000] = 32'b00000000000000001010001000010101;
assign LUT_1[12001] = 32'b00000000000000000011011010010001;
assign LUT_1[12002] = 32'b00000000000000000101110110100110;
assign LUT_1[12003] = 32'b11111111111111111111001000100010;
assign LUT_1[12004] = 32'b00000000000000010010000001101100;
assign LUT_1[12005] = 32'b00000000000000001011010011101000;
assign LUT_1[12006] = 32'b00000000000000001101101111111101;
assign LUT_1[12007] = 32'b00000000000000000111000001111001;
assign LUT_1[12008] = 32'b00000000000000001001010110001010;
assign LUT_1[12009] = 32'b00000000000000000010101000000110;
assign LUT_1[12010] = 32'b00000000000000000101000100011011;
assign LUT_1[12011] = 32'b11111111111111111110010110010111;
assign LUT_1[12012] = 32'b00000000000000010001001111100001;
assign LUT_1[12013] = 32'b00000000000000001010100001011101;
assign LUT_1[12014] = 32'b00000000000000001100111101110010;
assign LUT_1[12015] = 32'b00000000000000000110001111101110;
assign LUT_1[12016] = 32'b00000000000000001100000011110111;
assign LUT_1[12017] = 32'b00000000000000000101010101110011;
assign LUT_1[12018] = 32'b00000000000000000111110010001000;
assign LUT_1[12019] = 32'b00000000000000000001000100000100;
assign LUT_1[12020] = 32'b00000000000000010011111101001110;
assign LUT_1[12021] = 32'b00000000000000001101001111001010;
assign LUT_1[12022] = 32'b00000000000000001111101011011111;
assign LUT_1[12023] = 32'b00000000000000001000111101011011;
assign LUT_1[12024] = 32'b00000000000000001011010001101100;
assign LUT_1[12025] = 32'b00000000000000000100100011101000;
assign LUT_1[12026] = 32'b00000000000000000110111111111101;
assign LUT_1[12027] = 32'b00000000000000000000010001111001;
assign LUT_1[12028] = 32'b00000000000000010011001011000011;
assign LUT_1[12029] = 32'b00000000000000001100011100111111;
assign LUT_1[12030] = 32'b00000000000000001110111001010100;
assign LUT_1[12031] = 32'b00000000000000001000001011010000;
assign LUT_1[12032] = 32'b00000000000000000010000011110111;
assign LUT_1[12033] = 32'b11111111111111111011010101110011;
assign LUT_1[12034] = 32'b11111111111111111101110010001000;
assign LUT_1[12035] = 32'b11111111111111110111000100000100;
assign LUT_1[12036] = 32'b00000000000000001001111101001110;
assign LUT_1[12037] = 32'b00000000000000000011001111001010;
assign LUT_1[12038] = 32'b00000000000000000101101011011111;
assign LUT_1[12039] = 32'b11111111111111111110111101011011;
assign LUT_1[12040] = 32'b00000000000000000001010001101100;
assign LUT_1[12041] = 32'b11111111111111111010100011101000;
assign LUT_1[12042] = 32'b11111111111111111100111111111101;
assign LUT_1[12043] = 32'b11111111111111110110010001111001;
assign LUT_1[12044] = 32'b00000000000000001001001011000011;
assign LUT_1[12045] = 32'b00000000000000000010011100111111;
assign LUT_1[12046] = 32'b00000000000000000100111001010100;
assign LUT_1[12047] = 32'b11111111111111111110001011010000;
assign LUT_1[12048] = 32'b00000000000000000011111111011001;
assign LUT_1[12049] = 32'b11111111111111111101010001010101;
assign LUT_1[12050] = 32'b11111111111111111111101101101010;
assign LUT_1[12051] = 32'b11111111111111111000111111100110;
assign LUT_1[12052] = 32'b00000000000000001011111000110000;
assign LUT_1[12053] = 32'b00000000000000000101001010101100;
assign LUT_1[12054] = 32'b00000000000000000111100111000001;
assign LUT_1[12055] = 32'b00000000000000000000111000111101;
assign LUT_1[12056] = 32'b00000000000000000011001101001110;
assign LUT_1[12057] = 32'b11111111111111111100011111001010;
assign LUT_1[12058] = 32'b11111111111111111110111011011111;
assign LUT_1[12059] = 32'b11111111111111111000001101011011;
assign LUT_1[12060] = 32'b00000000000000001011000110100101;
assign LUT_1[12061] = 32'b00000000000000000100011000100001;
assign LUT_1[12062] = 32'b00000000000000000110110100110110;
assign LUT_1[12063] = 32'b00000000000000000000000110110010;
assign LUT_1[12064] = 32'b00000000000000000010111110110110;
assign LUT_1[12065] = 32'b11111111111111111100010000110010;
assign LUT_1[12066] = 32'b11111111111111111110101101000111;
assign LUT_1[12067] = 32'b11111111111111110111111111000011;
assign LUT_1[12068] = 32'b00000000000000001010111000001101;
assign LUT_1[12069] = 32'b00000000000000000100001010001001;
assign LUT_1[12070] = 32'b00000000000000000110100110011110;
assign LUT_1[12071] = 32'b11111111111111111111111000011010;
assign LUT_1[12072] = 32'b00000000000000000010001100101011;
assign LUT_1[12073] = 32'b11111111111111111011011110100111;
assign LUT_1[12074] = 32'b11111111111111111101111010111100;
assign LUT_1[12075] = 32'b11111111111111110111001100111000;
assign LUT_1[12076] = 32'b00000000000000001010000110000010;
assign LUT_1[12077] = 32'b00000000000000000011010111111110;
assign LUT_1[12078] = 32'b00000000000000000101110100010011;
assign LUT_1[12079] = 32'b11111111111111111111000110001111;
assign LUT_1[12080] = 32'b00000000000000000100111010011000;
assign LUT_1[12081] = 32'b11111111111111111110001100010100;
assign LUT_1[12082] = 32'b00000000000000000000101000101001;
assign LUT_1[12083] = 32'b11111111111111111001111010100101;
assign LUT_1[12084] = 32'b00000000000000001100110011101111;
assign LUT_1[12085] = 32'b00000000000000000110000101101011;
assign LUT_1[12086] = 32'b00000000000000001000100010000000;
assign LUT_1[12087] = 32'b00000000000000000001110011111100;
assign LUT_1[12088] = 32'b00000000000000000100001000001101;
assign LUT_1[12089] = 32'b11111111111111111101011010001001;
assign LUT_1[12090] = 32'b11111111111111111111110110011110;
assign LUT_1[12091] = 32'b11111111111111111001001000011010;
assign LUT_1[12092] = 32'b00000000000000001100000001100100;
assign LUT_1[12093] = 32'b00000000000000000101010011100000;
assign LUT_1[12094] = 32'b00000000000000000111101111110101;
assign LUT_1[12095] = 32'b00000000000000000001000001110001;
assign LUT_1[12096] = 32'b00000000000000000100000001011111;
assign LUT_1[12097] = 32'b11111111111111111101010011011011;
assign LUT_1[12098] = 32'b11111111111111111111101111110000;
assign LUT_1[12099] = 32'b11111111111111111001000001101100;
assign LUT_1[12100] = 32'b00000000000000001011111010110110;
assign LUT_1[12101] = 32'b00000000000000000101001100110010;
assign LUT_1[12102] = 32'b00000000000000000111101001000111;
assign LUT_1[12103] = 32'b00000000000000000000111011000011;
assign LUT_1[12104] = 32'b00000000000000000011001111010100;
assign LUT_1[12105] = 32'b11111111111111111100100001010000;
assign LUT_1[12106] = 32'b11111111111111111110111101100101;
assign LUT_1[12107] = 32'b11111111111111111000001111100001;
assign LUT_1[12108] = 32'b00000000000000001011001000101011;
assign LUT_1[12109] = 32'b00000000000000000100011010100111;
assign LUT_1[12110] = 32'b00000000000000000110110110111100;
assign LUT_1[12111] = 32'b00000000000000000000001000111000;
assign LUT_1[12112] = 32'b00000000000000000101111101000001;
assign LUT_1[12113] = 32'b11111111111111111111001110111101;
assign LUT_1[12114] = 32'b00000000000000000001101011010010;
assign LUT_1[12115] = 32'b11111111111111111010111101001110;
assign LUT_1[12116] = 32'b00000000000000001101110110011000;
assign LUT_1[12117] = 32'b00000000000000000111001000010100;
assign LUT_1[12118] = 32'b00000000000000001001100100101001;
assign LUT_1[12119] = 32'b00000000000000000010110110100101;
assign LUT_1[12120] = 32'b00000000000000000101001010110110;
assign LUT_1[12121] = 32'b11111111111111111110011100110010;
assign LUT_1[12122] = 32'b00000000000000000000111001000111;
assign LUT_1[12123] = 32'b11111111111111111010001011000011;
assign LUT_1[12124] = 32'b00000000000000001101000100001101;
assign LUT_1[12125] = 32'b00000000000000000110010110001001;
assign LUT_1[12126] = 32'b00000000000000001000110010011110;
assign LUT_1[12127] = 32'b00000000000000000010000100011010;
assign LUT_1[12128] = 32'b00000000000000000100111100011110;
assign LUT_1[12129] = 32'b11111111111111111110001110011010;
assign LUT_1[12130] = 32'b00000000000000000000101010101111;
assign LUT_1[12131] = 32'b11111111111111111001111100101011;
assign LUT_1[12132] = 32'b00000000000000001100110101110101;
assign LUT_1[12133] = 32'b00000000000000000110000111110001;
assign LUT_1[12134] = 32'b00000000000000001000100100000110;
assign LUT_1[12135] = 32'b00000000000000000001110110000010;
assign LUT_1[12136] = 32'b00000000000000000100001010010011;
assign LUT_1[12137] = 32'b11111111111111111101011100001111;
assign LUT_1[12138] = 32'b11111111111111111111111000100100;
assign LUT_1[12139] = 32'b11111111111111111001001010100000;
assign LUT_1[12140] = 32'b00000000000000001100000011101010;
assign LUT_1[12141] = 32'b00000000000000000101010101100110;
assign LUT_1[12142] = 32'b00000000000000000111110001111011;
assign LUT_1[12143] = 32'b00000000000000000001000011110111;
assign LUT_1[12144] = 32'b00000000000000000110111000000000;
assign LUT_1[12145] = 32'b00000000000000000000001001111100;
assign LUT_1[12146] = 32'b00000000000000000010100110010001;
assign LUT_1[12147] = 32'b11111111111111111011111000001101;
assign LUT_1[12148] = 32'b00000000000000001110110001010111;
assign LUT_1[12149] = 32'b00000000000000001000000011010011;
assign LUT_1[12150] = 32'b00000000000000001010011111101000;
assign LUT_1[12151] = 32'b00000000000000000011110001100100;
assign LUT_1[12152] = 32'b00000000000000000110000101110101;
assign LUT_1[12153] = 32'b11111111111111111111010111110001;
assign LUT_1[12154] = 32'b00000000000000000001110100000110;
assign LUT_1[12155] = 32'b11111111111111111011000110000010;
assign LUT_1[12156] = 32'b00000000000000001101111111001100;
assign LUT_1[12157] = 32'b00000000000000000111010001001000;
assign LUT_1[12158] = 32'b00000000000000001001101101011101;
assign LUT_1[12159] = 32'b00000000000000000010111111011001;
assign LUT_1[12160] = 32'b00000000000000000101000011111010;
assign LUT_1[12161] = 32'b11111111111111111110010101110110;
assign LUT_1[12162] = 32'b00000000000000000000110010001011;
assign LUT_1[12163] = 32'b11111111111111111010000100000111;
assign LUT_1[12164] = 32'b00000000000000001100111101010001;
assign LUT_1[12165] = 32'b00000000000000000110001111001101;
assign LUT_1[12166] = 32'b00000000000000001000101011100010;
assign LUT_1[12167] = 32'b00000000000000000001111101011110;
assign LUT_1[12168] = 32'b00000000000000000100010001101111;
assign LUT_1[12169] = 32'b11111111111111111101100011101011;
assign LUT_1[12170] = 32'b00000000000000000000000000000000;
assign LUT_1[12171] = 32'b11111111111111111001010001111100;
assign LUT_1[12172] = 32'b00000000000000001100001011000110;
assign LUT_1[12173] = 32'b00000000000000000101011101000010;
assign LUT_1[12174] = 32'b00000000000000000111111001010111;
assign LUT_1[12175] = 32'b00000000000000000001001011010011;
assign LUT_1[12176] = 32'b00000000000000000110111111011100;
assign LUT_1[12177] = 32'b00000000000000000000010001011000;
assign LUT_1[12178] = 32'b00000000000000000010101101101101;
assign LUT_1[12179] = 32'b11111111111111111011111111101001;
assign LUT_1[12180] = 32'b00000000000000001110111000110011;
assign LUT_1[12181] = 32'b00000000000000001000001010101111;
assign LUT_1[12182] = 32'b00000000000000001010100111000100;
assign LUT_1[12183] = 32'b00000000000000000011111001000000;
assign LUT_1[12184] = 32'b00000000000000000110001101010001;
assign LUT_1[12185] = 32'b11111111111111111111011111001101;
assign LUT_1[12186] = 32'b00000000000000000001111011100010;
assign LUT_1[12187] = 32'b11111111111111111011001101011110;
assign LUT_1[12188] = 32'b00000000000000001110000110101000;
assign LUT_1[12189] = 32'b00000000000000000111011000100100;
assign LUT_1[12190] = 32'b00000000000000001001110100111001;
assign LUT_1[12191] = 32'b00000000000000000011000110110101;
assign LUT_1[12192] = 32'b00000000000000000101111110111001;
assign LUT_1[12193] = 32'b11111111111111111111010000110101;
assign LUT_1[12194] = 32'b00000000000000000001101101001010;
assign LUT_1[12195] = 32'b11111111111111111010111111000110;
assign LUT_1[12196] = 32'b00000000000000001101111000010000;
assign LUT_1[12197] = 32'b00000000000000000111001010001100;
assign LUT_1[12198] = 32'b00000000000000001001100110100001;
assign LUT_1[12199] = 32'b00000000000000000010111000011101;
assign LUT_1[12200] = 32'b00000000000000000101001100101110;
assign LUT_1[12201] = 32'b11111111111111111110011110101010;
assign LUT_1[12202] = 32'b00000000000000000000111010111111;
assign LUT_1[12203] = 32'b11111111111111111010001100111011;
assign LUT_1[12204] = 32'b00000000000000001101000110000101;
assign LUT_1[12205] = 32'b00000000000000000110011000000001;
assign LUT_1[12206] = 32'b00000000000000001000110100010110;
assign LUT_1[12207] = 32'b00000000000000000010000110010010;
assign LUT_1[12208] = 32'b00000000000000000111111010011011;
assign LUT_1[12209] = 32'b00000000000000000001001100010111;
assign LUT_1[12210] = 32'b00000000000000000011101000101100;
assign LUT_1[12211] = 32'b11111111111111111100111010101000;
assign LUT_1[12212] = 32'b00000000000000001111110011110010;
assign LUT_1[12213] = 32'b00000000000000001001000101101110;
assign LUT_1[12214] = 32'b00000000000000001011100010000011;
assign LUT_1[12215] = 32'b00000000000000000100110011111111;
assign LUT_1[12216] = 32'b00000000000000000111001000010000;
assign LUT_1[12217] = 32'b00000000000000000000011010001100;
assign LUT_1[12218] = 32'b00000000000000000010110110100001;
assign LUT_1[12219] = 32'b11111111111111111100001000011101;
assign LUT_1[12220] = 32'b00000000000000001111000001100111;
assign LUT_1[12221] = 32'b00000000000000001000010011100011;
assign LUT_1[12222] = 32'b00000000000000001010101111111000;
assign LUT_1[12223] = 32'b00000000000000000100000001110100;
assign LUT_1[12224] = 32'b00000000000000000111000001100010;
assign LUT_1[12225] = 32'b00000000000000000000010011011110;
assign LUT_1[12226] = 32'b00000000000000000010101111110011;
assign LUT_1[12227] = 32'b11111111111111111100000001101111;
assign LUT_1[12228] = 32'b00000000000000001110111010111001;
assign LUT_1[12229] = 32'b00000000000000001000001100110101;
assign LUT_1[12230] = 32'b00000000000000001010101001001010;
assign LUT_1[12231] = 32'b00000000000000000011111011000110;
assign LUT_1[12232] = 32'b00000000000000000110001111010111;
assign LUT_1[12233] = 32'b11111111111111111111100001010011;
assign LUT_1[12234] = 32'b00000000000000000001111101101000;
assign LUT_1[12235] = 32'b11111111111111111011001111100100;
assign LUT_1[12236] = 32'b00000000000000001110001000101110;
assign LUT_1[12237] = 32'b00000000000000000111011010101010;
assign LUT_1[12238] = 32'b00000000000000001001110110111111;
assign LUT_1[12239] = 32'b00000000000000000011001000111011;
assign LUT_1[12240] = 32'b00000000000000001000111101000100;
assign LUT_1[12241] = 32'b00000000000000000010001111000000;
assign LUT_1[12242] = 32'b00000000000000000100101011010101;
assign LUT_1[12243] = 32'b11111111111111111101111101010001;
assign LUT_1[12244] = 32'b00000000000000010000110110011011;
assign LUT_1[12245] = 32'b00000000000000001010001000010111;
assign LUT_1[12246] = 32'b00000000000000001100100100101100;
assign LUT_1[12247] = 32'b00000000000000000101110110101000;
assign LUT_1[12248] = 32'b00000000000000001000001010111001;
assign LUT_1[12249] = 32'b00000000000000000001011100110101;
assign LUT_1[12250] = 32'b00000000000000000011111001001010;
assign LUT_1[12251] = 32'b11111111111111111101001011000110;
assign LUT_1[12252] = 32'b00000000000000010000000100010000;
assign LUT_1[12253] = 32'b00000000000000001001010110001100;
assign LUT_1[12254] = 32'b00000000000000001011110010100001;
assign LUT_1[12255] = 32'b00000000000000000101000100011101;
assign LUT_1[12256] = 32'b00000000000000000111111100100001;
assign LUT_1[12257] = 32'b00000000000000000001001110011101;
assign LUT_1[12258] = 32'b00000000000000000011101010110010;
assign LUT_1[12259] = 32'b11111111111111111100111100101110;
assign LUT_1[12260] = 32'b00000000000000001111110101111000;
assign LUT_1[12261] = 32'b00000000000000001001000111110100;
assign LUT_1[12262] = 32'b00000000000000001011100100001001;
assign LUT_1[12263] = 32'b00000000000000000100110110000101;
assign LUT_1[12264] = 32'b00000000000000000111001010010110;
assign LUT_1[12265] = 32'b00000000000000000000011100010010;
assign LUT_1[12266] = 32'b00000000000000000010111000100111;
assign LUT_1[12267] = 32'b11111111111111111100001010100011;
assign LUT_1[12268] = 32'b00000000000000001111000011101101;
assign LUT_1[12269] = 32'b00000000000000001000010101101001;
assign LUT_1[12270] = 32'b00000000000000001010110001111110;
assign LUT_1[12271] = 32'b00000000000000000100000011111010;
assign LUT_1[12272] = 32'b00000000000000001001111000000011;
assign LUT_1[12273] = 32'b00000000000000000011001001111111;
assign LUT_1[12274] = 32'b00000000000000000101100110010100;
assign LUT_1[12275] = 32'b11111111111111111110111000010000;
assign LUT_1[12276] = 32'b00000000000000010001110001011010;
assign LUT_1[12277] = 32'b00000000000000001011000011010110;
assign LUT_1[12278] = 32'b00000000000000001101011111101011;
assign LUT_1[12279] = 32'b00000000000000000110110001100111;
assign LUT_1[12280] = 32'b00000000000000001001000101111000;
assign LUT_1[12281] = 32'b00000000000000000010010111110100;
assign LUT_1[12282] = 32'b00000000000000000100110100001001;
assign LUT_1[12283] = 32'b11111111111111111110000110000101;
assign LUT_1[12284] = 32'b00000000000000010000111111001111;
assign LUT_1[12285] = 32'b00000000000000001010010001001011;
assign LUT_1[12286] = 32'b00000000000000001100101101100000;
assign LUT_1[12287] = 32'b00000000000000000101111111011100;
assign LUT_1[12288] = 32'b00000000000000000010111101101001;
assign LUT_1[12289] = 32'b11111111111111111100001111100101;
assign LUT_1[12290] = 32'b11111111111111111110101011111010;
assign LUT_1[12291] = 32'b11111111111111110111111101110110;
assign LUT_1[12292] = 32'b00000000000000001010110111000000;
assign LUT_1[12293] = 32'b00000000000000000100001000111100;
assign LUT_1[12294] = 32'b00000000000000000110100101010001;
assign LUT_1[12295] = 32'b11111111111111111111110111001101;
assign LUT_1[12296] = 32'b00000000000000000010001011011110;
assign LUT_1[12297] = 32'b11111111111111111011011101011010;
assign LUT_1[12298] = 32'b11111111111111111101111001101111;
assign LUT_1[12299] = 32'b11111111111111110111001011101011;
assign LUT_1[12300] = 32'b00000000000000001010000100110101;
assign LUT_1[12301] = 32'b00000000000000000011010110110001;
assign LUT_1[12302] = 32'b00000000000000000101110011000110;
assign LUT_1[12303] = 32'b11111111111111111111000101000010;
assign LUT_1[12304] = 32'b00000000000000000100111001001011;
assign LUT_1[12305] = 32'b11111111111111111110001011000111;
assign LUT_1[12306] = 32'b00000000000000000000100111011100;
assign LUT_1[12307] = 32'b11111111111111111001111001011000;
assign LUT_1[12308] = 32'b00000000000000001100110010100010;
assign LUT_1[12309] = 32'b00000000000000000110000100011110;
assign LUT_1[12310] = 32'b00000000000000001000100000110011;
assign LUT_1[12311] = 32'b00000000000000000001110010101111;
assign LUT_1[12312] = 32'b00000000000000000100000111000000;
assign LUT_1[12313] = 32'b11111111111111111101011000111100;
assign LUT_1[12314] = 32'b11111111111111111111110101010001;
assign LUT_1[12315] = 32'b11111111111111111001000111001101;
assign LUT_1[12316] = 32'b00000000000000001100000000010111;
assign LUT_1[12317] = 32'b00000000000000000101010010010011;
assign LUT_1[12318] = 32'b00000000000000000111101110101000;
assign LUT_1[12319] = 32'b00000000000000000001000000100100;
assign LUT_1[12320] = 32'b00000000000000000011111000101000;
assign LUT_1[12321] = 32'b11111111111111111101001010100100;
assign LUT_1[12322] = 32'b11111111111111111111100110111001;
assign LUT_1[12323] = 32'b11111111111111111000111000110101;
assign LUT_1[12324] = 32'b00000000000000001011110001111111;
assign LUT_1[12325] = 32'b00000000000000000101000011111011;
assign LUT_1[12326] = 32'b00000000000000000111100000010000;
assign LUT_1[12327] = 32'b00000000000000000000110010001100;
assign LUT_1[12328] = 32'b00000000000000000011000110011101;
assign LUT_1[12329] = 32'b11111111111111111100011000011001;
assign LUT_1[12330] = 32'b11111111111111111110110100101110;
assign LUT_1[12331] = 32'b11111111111111111000000110101010;
assign LUT_1[12332] = 32'b00000000000000001010111111110100;
assign LUT_1[12333] = 32'b00000000000000000100010001110000;
assign LUT_1[12334] = 32'b00000000000000000110101110000101;
assign LUT_1[12335] = 32'b00000000000000000000000000000001;
assign LUT_1[12336] = 32'b00000000000000000101110100001010;
assign LUT_1[12337] = 32'b11111111111111111111000110000110;
assign LUT_1[12338] = 32'b00000000000000000001100010011011;
assign LUT_1[12339] = 32'b11111111111111111010110100010111;
assign LUT_1[12340] = 32'b00000000000000001101101101100001;
assign LUT_1[12341] = 32'b00000000000000000110111111011101;
assign LUT_1[12342] = 32'b00000000000000001001011011110010;
assign LUT_1[12343] = 32'b00000000000000000010101101101110;
assign LUT_1[12344] = 32'b00000000000000000101000001111111;
assign LUT_1[12345] = 32'b11111111111111111110010011111011;
assign LUT_1[12346] = 32'b00000000000000000000110000010000;
assign LUT_1[12347] = 32'b11111111111111111010000010001100;
assign LUT_1[12348] = 32'b00000000000000001100111011010110;
assign LUT_1[12349] = 32'b00000000000000000110001101010010;
assign LUT_1[12350] = 32'b00000000000000001000101001100111;
assign LUT_1[12351] = 32'b00000000000000000001111011100011;
assign LUT_1[12352] = 32'b00000000000000000100111011010001;
assign LUT_1[12353] = 32'b11111111111111111110001101001101;
assign LUT_1[12354] = 32'b00000000000000000000101001100010;
assign LUT_1[12355] = 32'b11111111111111111001111011011110;
assign LUT_1[12356] = 32'b00000000000000001100110100101000;
assign LUT_1[12357] = 32'b00000000000000000110000110100100;
assign LUT_1[12358] = 32'b00000000000000001000100010111001;
assign LUT_1[12359] = 32'b00000000000000000001110100110101;
assign LUT_1[12360] = 32'b00000000000000000100001001000110;
assign LUT_1[12361] = 32'b11111111111111111101011011000010;
assign LUT_1[12362] = 32'b11111111111111111111110111010111;
assign LUT_1[12363] = 32'b11111111111111111001001001010011;
assign LUT_1[12364] = 32'b00000000000000001100000010011101;
assign LUT_1[12365] = 32'b00000000000000000101010100011001;
assign LUT_1[12366] = 32'b00000000000000000111110000101110;
assign LUT_1[12367] = 32'b00000000000000000001000010101010;
assign LUT_1[12368] = 32'b00000000000000000110110110110011;
assign LUT_1[12369] = 32'b00000000000000000000001000101111;
assign LUT_1[12370] = 32'b00000000000000000010100101000100;
assign LUT_1[12371] = 32'b11111111111111111011110111000000;
assign LUT_1[12372] = 32'b00000000000000001110110000001010;
assign LUT_1[12373] = 32'b00000000000000001000000010000110;
assign LUT_1[12374] = 32'b00000000000000001010011110011011;
assign LUT_1[12375] = 32'b00000000000000000011110000010111;
assign LUT_1[12376] = 32'b00000000000000000110000100101000;
assign LUT_1[12377] = 32'b11111111111111111111010110100100;
assign LUT_1[12378] = 32'b00000000000000000001110010111001;
assign LUT_1[12379] = 32'b11111111111111111011000100110101;
assign LUT_1[12380] = 32'b00000000000000001101111101111111;
assign LUT_1[12381] = 32'b00000000000000000111001111111011;
assign LUT_1[12382] = 32'b00000000000000001001101100010000;
assign LUT_1[12383] = 32'b00000000000000000010111110001100;
assign LUT_1[12384] = 32'b00000000000000000101110110010000;
assign LUT_1[12385] = 32'b11111111111111111111001000001100;
assign LUT_1[12386] = 32'b00000000000000000001100100100001;
assign LUT_1[12387] = 32'b11111111111111111010110110011101;
assign LUT_1[12388] = 32'b00000000000000001101101111100111;
assign LUT_1[12389] = 32'b00000000000000000111000001100011;
assign LUT_1[12390] = 32'b00000000000000001001011101111000;
assign LUT_1[12391] = 32'b00000000000000000010101111110100;
assign LUT_1[12392] = 32'b00000000000000000101000100000101;
assign LUT_1[12393] = 32'b11111111111111111110010110000001;
assign LUT_1[12394] = 32'b00000000000000000000110010010110;
assign LUT_1[12395] = 32'b11111111111111111010000100010010;
assign LUT_1[12396] = 32'b00000000000000001100111101011100;
assign LUT_1[12397] = 32'b00000000000000000110001111011000;
assign LUT_1[12398] = 32'b00000000000000001000101011101101;
assign LUT_1[12399] = 32'b00000000000000000001111101101001;
assign LUT_1[12400] = 32'b00000000000000000111110001110010;
assign LUT_1[12401] = 32'b00000000000000000001000011101110;
assign LUT_1[12402] = 32'b00000000000000000011100000000011;
assign LUT_1[12403] = 32'b11111111111111111100110001111111;
assign LUT_1[12404] = 32'b00000000000000001111101011001001;
assign LUT_1[12405] = 32'b00000000000000001000111101000101;
assign LUT_1[12406] = 32'b00000000000000001011011001011010;
assign LUT_1[12407] = 32'b00000000000000000100101011010110;
assign LUT_1[12408] = 32'b00000000000000000110111111100111;
assign LUT_1[12409] = 32'b00000000000000000000010001100011;
assign LUT_1[12410] = 32'b00000000000000000010101101111000;
assign LUT_1[12411] = 32'b11111111111111111011111111110100;
assign LUT_1[12412] = 32'b00000000000000001110111000111110;
assign LUT_1[12413] = 32'b00000000000000001000001010111010;
assign LUT_1[12414] = 32'b00000000000000001010100111001111;
assign LUT_1[12415] = 32'b00000000000000000011111001001011;
assign LUT_1[12416] = 32'b00000000000000000101111101101100;
assign LUT_1[12417] = 32'b11111111111111111111001111101000;
assign LUT_1[12418] = 32'b00000000000000000001101011111101;
assign LUT_1[12419] = 32'b11111111111111111010111101111001;
assign LUT_1[12420] = 32'b00000000000000001101110111000011;
assign LUT_1[12421] = 32'b00000000000000000111001000111111;
assign LUT_1[12422] = 32'b00000000000000001001100101010100;
assign LUT_1[12423] = 32'b00000000000000000010110111010000;
assign LUT_1[12424] = 32'b00000000000000000101001011100001;
assign LUT_1[12425] = 32'b11111111111111111110011101011101;
assign LUT_1[12426] = 32'b00000000000000000000111001110010;
assign LUT_1[12427] = 32'b11111111111111111010001011101110;
assign LUT_1[12428] = 32'b00000000000000001101000100111000;
assign LUT_1[12429] = 32'b00000000000000000110010110110100;
assign LUT_1[12430] = 32'b00000000000000001000110011001001;
assign LUT_1[12431] = 32'b00000000000000000010000101000101;
assign LUT_1[12432] = 32'b00000000000000000111111001001110;
assign LUT_1[12433] = 32'b00000000000000000001001011001010;
assign LUT_1[12434] = 32'b00000000000000000011100111011111;
assign LUT_1[12435] = 32'b11111111111111111100111001011011;
assign LUT_1[12436] = 32'b00000000000000001111110010100101;
assign LUT_1[12437] = 32'b00000000000000001001000100100001;
assign LUT_1[12438] = 32'b00000000000000001011100000110110;
assign LUT_1[12439] = 32'b00000000000000000100110010110010;
assign LUT_1[12440] = 32'b00000000000000000111000111000011;
assign LUT_1[12441] = 32'b00000000000000000000011000111111;
assign LUT_1[12442] = 32'b00000000000000000010110101010100;
assign LUT_1[12443] = 32'b11111111111111111100000111010000;
assign LUT_1[12444] = 32'b00000000000000001111000000011010;
assign LUT_1[12445] = 32'b00000000000000001000010010010110;
assign LUT_1[12446] = 32'b00000000000000001010101110101011;
assign LUT_1[12447] = 32'b00000000000000000100000000100111;
assign LUT_1[12448] = 32'b00000000000000000110111000101011;
assign LUT_1[12449] = 32'b00000000000000000000001010100111;
assign LUT_1[12450] = 32'b00000000000000000010100110111100;
assign LUT_1[12451] = 32'b11111111111111111011111000111000;
assign LUT_1[12452] = 32'b00000000000000001110110010000010;
assign LUT_1[12453] = 32'b00000000000000001000000011111110;
assign LUT_1[12454] = 32'b00000000000000001010100000010011;
assign LUT_1[12455] = 32'b00000000000000000011110010001111;
assign LUT_1[12456] = 32'b00000000000000000110000110100000;
assign LUT_1[12457] = 32'b11111111111111111111011000011100;
assign LUT_1[12458] = 32'b00000000000000000001110100110001;
assign LUT_1[12459] = 32'b11111111111111111011000110101101;
assign LUT_1[12460] = 32'b00000000000000001101111111110111;
assign LUT_1[12461] = 32'b00000000000000000111010001110011;
assign LUT_1[12462] = 32'b00000000000000001001101110001000;
assign LUT_1[12463] = 32'b00000000000000000011000000000100;
assign LUT_1[12464] = 32'b00000000000000001000110100001101;
assign LUT_1[12465] = 32'b00000000000000000010000110001001;
assign LUT_1[12466] = 32'b00000000000000000100100010011110;
assign LUT_1[12467] = 32'b11111111111111111101110100011010;
assign LUT_1[12468] = 32'b00000000000000010000101101100100;
assign LUT_1[12469] = 32'b00000000000000001001111111100000;
assign LUT_1[12470] = 32'b00000000000000001100011011110101;
assign LUT_1[12471] = 32'b00000000000000000101101101110001;
assign LUT_1[12472] = 32'b00000000000000001000000010000010;
assign LUT_1[12473] = 32'b00000000000000000001010011111110;
assign LUT_1[12474] = 32'b00000000000000000011110000010011;
assign LUT_1[12475] = 32'b11111111111111111101000010001111;
assign LUT_1[12476] = 32'b00000000000000001111111011011001;
assign LUT_1[12477] = 32'b00000000000000001001001101010101;
assign LUT_1[12478] = 32'b00000000000000001011101001101010;
assign LUT_1[12479] = 32'b00000000000000000100111011100110;
assign LUT_1[12480] = 32'b00000000000000000111111011010100;
assign LUT_1[12481] = 32'b00000000000000000001001101010000;
assign LUT_1[12482] = 32'b00000000000000000011101001100101;
assign LUT_1[12483] = 32'b11111111111111111100111011100001;
assign LUT_1[12484] = 32'b00000000000000001111110100101011;
assign LUT_1[12485] = 32'b00000000000000001001000110100111;
assign LUT_1[12486] = 32'b00000000000000001011100010111100;
assign LUT_1[12487] = 32'b00000000000000000100110100111000;
assign LUT_1[12488] = 32'b00000000000000000111001001001001;
assign LUT_1[12489] = 32'b00000000000000000000011011000101;
assign LUT_1[12490] = 32'b00000000000000000010110111011010;
assign LUT_1[12491] = 32'b11111111111111111100001001010110;
assign LUT_1[12492] = 32'b00000000000000001111000010100000;
assign LUT_1[12493] = 32'b00000000000000001000010100011100;
assign LUT_1[12494] = 32'b00000000000000001010110000110001;
assign LUT_1[12495] = 32'b00000000000000000100000010101101;
assign LUT_1[12496] = 32'b00000000000000001001110110110110;
assign LUT_1[12497] = 32'b00000000000000000011001000110010;
assign LUT_1[12498] = 32'b00000000000000000101100101000111;
assign LUT_1[12499] = 32'b11111111111111111110110111000011;
assign LUT_1[12500] = 32'b00000000000000010001110000001101;
assign LUT_1[12501] = 32'b00000000000000001011000010001001;
assign LUT_1[12502] = 32'b00000000000000001101011110011110;
assign LUT_1[12503] = 32'b00000000000000000110110000011010;
assign LUT_1[12504] = 32'b00000000000000001001000100101011;
assign LUT_1[12505] = 32'b00000000000000000010010110100111;
assign LUT_1[12506] = 32'b00000000000000000100110010111100;
assign LUT_1[12507] = 32'b11111111111111111110000100111000;
assign LUT_1[12508] = 32'b00000000000000010000111110000010;
assign LUT_1[12509] = 32'b00000000000000001010001111111110;
assign LUT_1[12510] = 32'b00000000000000001100101100010011;
assign LUT_1[12511] = 32'b00000000000000000101111110001111;
assign LUT_1[12512] = 32'b00000000000000001000110110010011;
assign LUT_1[12513] = 32'b00000000000000000010001000001111;
assign LUT_1[12514] = 32'b00000000000000000100100100100100;
assign LUT_1[12515] = 32'b11111111111111111101110110100000;
assign LUT_1[12516] = 32'b00000000000000010000101111101010;
assign LUT_1[12517] = 32'b00000000000000001010000001100110;
assign LUT_1[12518] = 32'b00000000000000001100011101111011;
assign LUT_1[12519] = 32'b00000000000000000101101111110111;
assign LUT_1[12520] = 32'b00000000000000001000000100001000;
assign LUT_1[12521] = 32'b00000000000000000001010110000100;
assign LUT_1[12522] = 32'b00000000000000000011110010011001;
assign LUT_1[12523] = 32'b11111111111111111101000100010101;
assign LUT_1[12524] = 32'b00000000000000001111111101011111;
assign LUT_1[12525] = 32'b00000000000000001001001111011011;
assign LUT_1[12526] = 32'b00000000000000001011101011110000;
assign LUT_1[12527] = 32'b00000000000000000100111101101100;
assign LUT_1[12528] = 32'b00000000000000001010110001110101;
assign LUT_1[12529] = 32'b00000000000000000100000011110001;
assign LUT_1[12530] = 32'b00000000000000000110100000000110;
assign LUT_1[12531] = 32'b11111111111111111111110010000010;
assign LUT_1[12532] = 32'b00000000000000010010101011001100;
assign LUT_1[12533] = 32'b00000000000000001011111101001000;
assign LUT_1[12534] = 32'b00000000000000001110011001011101;
assign LUT_1[12535] = 32'b00000000000000000111101011011001;
assign LUT_1[12536] = 32'b00000000000000001001111111101010;
assign LUT_1[12537] = 32'b00000000000000000011010001100110;
assign LUT_1[12538] = 32'b00000000000000000101101101111011;
assign LUT_1[12539] = 32'b11111111111111111110111111110111;
assign LUT_1[12540] = 32'b00000000000000010001111001000001;
assign LUT_1[12541] = 32'b00000000000000001011001010111101;
assign LUT_1[12542] = 32'b00000000000000001101100111010010;
assign LUT_1[12543] = 32'b00000000000000000110111001001110;
assign LUT_1[12544] = 32'b00000000000000000000110001110101;
assign LUT_1[12545] = 32'b11111111111111111010000011110001;
assign LUT_1[12546] = 32'b11111111111111111100100000000110;
assign LUT_1[12547] = 32'b11111111111111110101110010000010;
assign LUT_1[12548] = 32'b00000000000000001000101011001100;
assign LUT_1[12549] = 32'b00000000000000000001111101001000;
assign LUT_1[12550] = 32'b00000000000000000100011001011101;
assign LUT_1[12551] = 32'b11111111111111111101101011011001;
assign LUT_1[12552] = 32'b11111111111111111111111111101010;
assign LUT_1[12553] = 32'b11111111111111111001010001100110;
assign LUT_1[12554] = 32'b11111111111111111011101101111011;
assign LUT_1[12555] = 32'b11111111111111110100111111110111;
assign LUT_1[12556] = 32'b00000000000000000111111001000001;
assign LUT_1[12557] = 32'b00000000000000000001001010111101;
assign LUT_1[12558] = 32'b00000000000000000011100111010010;
assign LUT_1[12559] = 32'b11111111111111111100111001001110;
assign LUT_1[12560] = 32'b00000000000000000010101101010111;
assign LUT_1[12561] = 32'b11111111111111111011111111010011;
assign LUT_1[12562] = 32'b11111111111111111110011011101000;
assign LUT_1[12563] = 32'b11111111111111110111101101100100;
assign LUT_1[12564] = 32'b00000000000000001010100110101110;
assign LUT_1[12565] = 32'b00000000000000000011111000101010;
assign LUT_1[12566] = 32'b00000000000000000110010100111111;
assign LUT_1[12567] = 32'b11111111111111111111100110111011;
assign LUT_1[12568] = 32'b00000000000000000001111011001100;
assign LUT_1[12569] = 32'b11111111111111111011001101001000;
assign LUT_1[12570] = 32'b11111111111111111101101001011101;
assign LUT_1[12571] = 32'b11111111111111110110111011011001;
assign LUT_1[12572] = 32'b00000000000000001001110100100011;
assign LUT_1[12573] = 32'b00000000000000000011000110011111;
assign LUT_1[12574] = 32'b00000000000000000101100010110100;
assign LUT_1[12575] = 32'b11111111111111111110110100110000;
assign LUT_1[12576] = 32'b00000000000000000001101100110100;
assign LUT_1[12577] = 32'b11111111111111111010111110110000;
assign LUT_1[12578] = 32'b11111111111111111101011011000101;
assign LUT_1[12579] = 32'b11111111111111110110101101000001;
assign LUT_1[12580] = 32'b00000000000000001001100110001011;
assign LUT_1[12581] = 32'b00000000000000000010111000000111;
assign LUT_1[12582] = 32'b00000000000000000101010100011100;
assign LUT_1[12583] = 32'b11111111111111111110100110011000;
assign LUT_1[12584] = 32'b00000000000000000000111010101001;
assign LUT_1[12585] = 32'b11111111111111111010001100100101;
assign LUT_1[12586] = 32'b11111111111111111100101000111010;
assign LUT_1[12587] = 32'b11111111111111110101111010110110;
assign LUT_1[12588] = 32'b00000000000000001000110100000000;
assign LUT_1[12589] = 32'b00000000000000000010000101111100;
assign LUT_1[12590] = 32'b00000000000000000100100010010001;
assign LUT_1[12591] = 32'b11111111111111111101110100001101;
assign LUT_1[12592] = 32'b00000000000000000011101000010110;
assign LUT_1[12593] = 32'b11111111111111111100111010010010;
assign LUT_1[12594] = 32'b11111111111111111111010110100111;
assign LUT_1[12595] = 32'b11111111111111111000101000100011;
assign LUT_1[12596] = 32'b00000000000000001011100001101101;
assign LUT_1[12597] = 32'b00000000000000000100110011101001;
assign LUT_1[12598] = 32'b00000000000000000111001111111110;
assign LUT_1[12599] = 32'b00000000000000000000100001111010;
assign LUT_1[12600] = 32'b00000000000000000010110110001011;
assign LUT_1[12601] = 32'b11111111111111111100001000000111;
assign LUT_1[12602] = 32'b11111111111111111110100100011100;
assign LUT_1[12603] = 32'b11111111111111110111110110011000;
assign LUT_1[12604] = 32'b00000000000000001010101111100010;
assign LUT_1[12605] = 32'b00000000000000000100000001011110;
assign LUT_1[12606] = 32'b00000000000000000110011101110011;
assign LUT_1[12607] = 32'b11111111111111111111101111101111;
assign LUT_1[12608] = 32'b00000000000000000010101111011101;
assign LUT_1[12609] = 32'b11111111111111111100000001011001;
assign LUT_1[12610] = 32'b11111111111111111110011101101110;
assign LUT_1[12611] = 32'b11111111111111110111101111101010;
assign LUT_1[12612] = 32'b00000000000000001010101000110100;
assign LUT_1[12613] = 32'b00000000000000000011111010110000;
assign LUT_1[12614] = 32'b00000000000000000110010111000101;
assign LUT_1[12615] = 32'b11111111111111111111101001000001;
assign LUT_1[12616] = 32'b00000000000000000001111101010010;
assign LUT_1[12617] = 32'b11111111111111111011001111001110;
assign LUT_1[12618] = 32'b11111111111111111101101011100011;
assign LUT_1[12619] = 32'b11111111111111110110111101011111;
assign LUT_1[12620] = 32'b00000000000000001001110110101001;
assign LUT_1[12621] = 32'b00000000000000000011001000100101;
assign LUT_1[12622] = 32'b00000000000000000101100100111010;
assign LUT_1[12623] = 32'b11111111111111111110110110110110;
assign LUT_1[12624] = 32'b00000000000000000100101010111111;
assign LUT_1[12625] = 32'b11111111111111111101111100111011;
assign LUT_1[12626] = 32'b00000000000000000000011001010000;
assign LUT_1[12627] = 32'b11111111111111111001101011001100;
assign LUT_1[12628] = 32'b00000000000000001100100100010110;
assign LUT_1[12629] = 32'b00000000000000000101110110010010;
assign LUT_1[12630] = 32'b00000000000000001000010010100111;
assign LUT_1[12631] = 32'b00000000000000000001100100100011;
assign LUT_1[12632] = 32'b00000000000000000011111000110100;
assign LUT_1[12633] = 32'b11111111111111111101001010110000;
assign LUT_1[12634] = 32'b11111111111111111111100111000101;
assign LUT_1[12635] = 32'b11111111111111111000111001000001;
assign LUT_1[12636] = 32'b00000000000000001011110010001011;
assign LUT_1[12637] = 32'b00000000000000000101000100000111;
assign LUT_1[12638] = 32'b00000000000000000111100000011100;
assign LUT_1[12639] = 32'b00000000000000000000110010011000;
assign LUT_1[12640] = 32'b00000000000000000011101010011100;
assign LUT_1[12641] = 32'b11111111111111111100111100011000;
assign LUT_1[12642] = 32'b11111111111111111111011000101101;
assign LUT_1[12643] = 32'b11111111111111111000101010101001;
assign LUT_1[12644] = 32'b00000000000000001011100011110011;
assign LUT_1[12645] = 32'b00000000000000000100110101101111;
assign LUT_1[12646] = 32'b00000000000000000111010010000100;
assign LUT_1[12647] = 32'b00000000000000000000100100000000;
assign LUT_1[12648] = 32'b00000000000000000010111000010001;
assign LUT_1[12649] = 32'b11111111111111111100001010001101;
assign LUT_1[12650] = 32'b11111111111111111110100110100010;
assign LUT_1[12651] = 32'b11111111111111110111111000011110;
assign LUT_1[12652] = 32'b00000000000000001010110001101000;
assign LUT_1[12653] = 32'b00000000000000000100000011100100;
assign LUT_1[12654] = 32'b00000000000000000110011111111001;
assign LUT_1[12655] = 32'b11111111111111111111110001110101;
assign LUT_1[12656] = 32'b00000000000000000101100101111110;
assign LUT_1[12657] = 32'b11111111111111111110110111111010;
assign LUT_1[12658] = 32'b00000000000000000001010100001111;
assign LUT_1[12659] = 32'b11111111111111111010100110001011;
assign LUT_1[12660] = 32'b00000000000000001101011111010101;
assign LUT_1[12661] = 32'b00000000000000000110110001010001;
assign LUT_1[12662] = 32'b00000000000000001001001101100110;
assign LUT_1[12663] = 32'b00000000000000000010011111100010;
assign LUT_1[12664] = 32'b00000000000000000100110011110011;
assign LUT_1[12665] = 32'b11111111111111111110000101101111;
assign LUT_1[12666] = 32'b00000000000000000000100010000100;
assign LUT_1[12667] = 32'b11111111111111111001110100000000;
assign LUT_1[12668] = 32'b00000000000000001100101101001010;
assign LUT_1[12669] = 32'b00000000000000000101111111000110;
assign LUT_1[12670] = 32'b00000000000000001000011011011011;
assign LUT_1[12671] = 32'b00000000000000000001101101010111;
assign LUT_1[12672] = 32'b00000000000000000011110001111000;
assign LUT_1[12673] = 32'b11111111111111111101000011110100;
assign LUT_1[12674] = 32'b11111111111111111111100000001001;
assign LUT_1[12675] = 32'b11111111111111111000110010000101;
assign LUT_1[12676] = 32'b00000000000000001011101011001111;
assign LUT_1[12677] = 32'b00000000000000000100111101001011;
assign LUT_1[12678] = 32'b00000000000000000111011001100000;
assign LUT_1[12679] = 32'b00000000000000000000101011011100;
assign LUT_1[12680] = 32'b00000000000000000010111111101101;
assign LUT_1[12681] = 32'b11111111111111111100010001101001;
assign LUT_1[12682] = 32'b11111111111111111110101101111110;
assign LUT_1[12683] = 32'b11111111111111110111111111111010;
assign LUT_1[12684] = 32'b00000000000000001010111001000100;
assign LUT_1[12685] = 32'b00000000000000000100001011000000;
assign LUT_1[12686] = 32'b00000000000000000110100111010101;
assign LUT_1[12687] = 32'b11111111111111111111111001010001;
assign LUT_1[12688] = 32'b00000000000000000101101101011010;
assign LUT_1[12689] = 32'b11111111111111111110111111010110;
assign LUT_1[12690] = 32'b00000000000000000001011011101011;
assign LUT_1[12691] = 32'b11111111111111111010101101100111;
assign LUT_1[12692] = 32'b00000000000000001101100110110001;
assign LUT_1[12693] = 32'b00000000000000000110111000101101;
assign LUT_1[12694] = 32'b00000000000000001001010101000010;
assign LUT_1[12695] = 32'b00000000000000000010100110111110;
assign LUT_1[12696] = 32'b00000000000000000100111011001111;
assign LUT_1[12697] = 32'b11111111111111111110001101001011;
assign LUT_1[12698] = 32'b00000000000000000000101001100000;
assign LUT_1[12699] = 32'b11111111111111111001111011011100;
assign LUT_1[12700] = 32'b00000000000000001100110100100110;
assign LUT_1[12701] = 32'b00000000000000000110000110100010;
assign LUT_1[12702] = 32'b00000000000000001000100010110111;
assign LUT_1[12703] = 32'b00000000000000000001110100110011;
assign LUT_1[12704] = 32'b00000000000000000100101100110111;
assign LUT_1[12705] = 32'b11111111111111111101111110110011;
assign LUT_1[12706] = 32'b00000000000000000000011011001000;
assign LUT_1[12707] = 32'b11111111111111111001101101000100;
assign LUT_1[12708] = 32'b00000000000000001100100110001110;
assign LUT_1[12709] = 32'b00000000000000000101111000001010;
assign LUT_1[12710] = 32'b00000000000000001000010100011111;
assign LUT_1[12711] = 32'b00000000000000000001100110011011;
assign LUT_1[12712] = 32'b00000000000000000011111010101100;
assign LUT_1[12713] = 32'b11111111111111111101001100101000;
assign LUT_1[12714] = 32'b11111111111111111111101000111101;
assign LUT_1[12715] = 32'b11111111111111111000111010111001;
assign LUT_1[12716] = 32'b00000000000000001011110100000011;
assign LUT_1[12717] = 32'b00000000000000000101000101111111;
assign LUT_1[12718] = 32'b00000000000000000111100010010100;
assign LUT_1[12719] = 32'b00000000000000000000110100010000;
assign LUT_1[12720] = 32'b00000000000000000110101000011001;
assign LUT_1[12721] = 32'b11111111111111111111111010010101;
assign LUT_1[12722] = 32'b00000000000000000010010110101010;
assign LUT_1[12723] = 32'b11111111111111111011101000100110;
assign LUT_1[12724] = 32'b00000000000000001110100001110000;
assign LUT_1[12725] = 32'b00000000000000000111110011101100;
assign LUT_1[12726] = 32'b00000000000000001010010000000001;
assign LUT_1[12727] = 32'b00000000000000000011100001111101;
assign LUT_1[12728] = 32'b00000000000000000101110110001110;
assign LUT_1[12729] = 32'b11111111111111111111001000001010;
assign LUT_1[12730] = 32'b00000000000000000001100100011111;
assign LUT_1[12731] = 32'b11111111111111111010110110011011;
assign LUT_1[12732] = 32'b00000000000000001101101111100101;
assign LUT_1[12733] = 32'b00000000000000000111000001100001;
assign LUT_1[12734] = 32'b00000000000000001001011101110110;
assign LUT_1[12735] = 32'b00000000000000000010101111110010;
assign LUT_1[12736] = 32'b00000000000000000101101111100000;
assign LUT_1[12737] = 32'b11111111111111111111000001011100;
assign LUT_1[12738] = 32'b00000000000000000001011101110001;
assign LUT_1[12739] = 32'b11111111111111111010101111101101;
assign LUT_1[12740] = 32'b00000000000000001101101000110111;
assign LUT_1[12741] = 32'b00000000000000000110111010110011;
assign LUT_1[12742] = 32'b00000000000000001001010111001000;
assign LUT_1[12743] = 32'b00000000000000000010101001000100;
assign LUT_1[12744] = 32'b00000000000000000100111101010101;
assign LUT_1[12745] = 32'b11111111111111111110001111010001;
assign LUT_1[12746] = 32'b00000000000000000000101011100110;
assign LUT_1[12747] = 32'b11111111111111111001111101100010;
assign LUT_1[12748] = 32'b00000000000000001100110110101100;
assign LUT_1[12749] = 32'b00000000000000000110001000101000;
assign LUT_1[12750] = 32'b00000000000000001000100100111101;
assign LUT_1[12751] = 32'b00000000000000000001110110111001;
assign LUT_1[12752] = 32'b00000000000000000111101011000010;
assign LUT_1[12753] = 32'b00000000000000000000111100111110;
assign LUT_1[12754] = 32'b00000000000000000011011001010011;
assign LUT_1[12755] = 32'b11111111111111111100101011001111;
assign LUT_1[12756] = 32'b00000000000000001111100100011001;
assign LUT_1[12757] = 32'b00000000000000001000110110010101;
assign LUT_1[12758] = 32'b00000000000000001011010010101010;
assign LUT_1[12759] = 32'b00000000000000000100100100100110;
assign LUT_1[12760] = 32'b00000000000000000110111000110111;
assign LUT_1[12761] = 32'b00000000000000000000001010110011;
assign LUT_1[12762] = 32'b00000000000000000010100111001000;
assign LUT_1[12763] = 32'b11111111111111111011111001000100;
assign LUT_1[12764] = 32'b00000000000000001110110010001110;
assign LUT_1[12765] = 32'b00000000000000001000000100001010;
assign LUT_1[12766] = 32'b00000000000000001010100000011111;
assign LUT_1[12767] = 32'b00000000000000000011110010011011;
assign LUT_1[12768] = 32'b00000000000000000110101010011111;
assign LUT_1[12769] = 32'b11111111111111111111111100011011;
assign LUT_1[12770] = 32'b00000000000000000010011000110000;
assign LUT_1[12771] = 32'b11111111111111111011101010101100;
assign LUT_1[12772] = 32'b00000000000000001110100011110110;
assign LUT_1[12773] = 32'b00000000000000000111110101110010;
assign LUT_1[12774] = 32'b00000000000000001010010010000111;
assign LUT_1[12775] = 32'b00000000000000000011100100000011;
assign LUT_1[12776] = 32'b00000000000000000101111000010100;
assign LUT_1[12777] = 32'b11111111111111111111001010010000;
assign LUT_1[12778] = 32'b00000000000000000001100110100101;
assign LUT_1[12779] = 32'b11111111111111111010111000100001;
assign LUT_1[12780] = 32'b00000000000000001101110001101011;
assign LUT_1[12781] = 32'b00000000000000000111000011100111;
assign LUT_1[12782] = 32'b00000000000000001001011111111100;
assign LUT_1[12783] = 32'b00000000000000000010110001111000;
assign LUT_1[12784] = 32'b00000000000000001000100110000001;
assign LUT_1[12785] = 32'b00000000000000000001110111111101;
assign LUT_1[12786] = 32'b00000000000000000100010100010010;
assign LUT_1[12787] = 32'b11111111111111111101100110001110;
assign LUT_1[12788] = 32'b00000000000000010000011111011000;
assign LUT_1[12789] = 32'b00000000000000001001110001010100;
assign LUT_1[12790] = 32'b00000000000000001100001101101001;
assign LUT_1[12791] = 32'b00000000000000000101011111100101;
assign LUT_1[12792] = 32'b00000000000000000111110011110110;
assign LUT_1[12793] = 32'b00000000000000000001000101110010;
assign LUT_1[12794] = 32'b00000000000000000011100010000111;
assign LUT_1[12795] = 32'b11111111111111111100110100000011;
assign LUT_1[12796] = 32'b00000000000000001111101101001101;
assign LUT_1[12797] = 32'b00000000000000001000111111001001;
assign LUT_1[12798] = 32'b00000000000000001011011011011110;
assign LUT_1[12799] = 32'b00000000000000000100101101011010;
assign LUT_1[12800] = 32'b11111111111111111100101100000110;
assign LUT_1[12801] = 32'b11111111111111110101111110000010;
assign LUT_1[12802] = 32'b11111111111111111000011010010111;
assign LUT_1[12803] = 32'b11111111111111110001101100010011;
assign LUT_1[12804] = 32'b00000000000000000100100101011101;
assign LUT_1[12805] = 32'b11111111111111111101110111011001;
assign LUT_1[12806] = 32'b00000000000000000000010011101110;
assign LUT_1[12807] = 32'b11111111111111111001100101101010;
assign LUT_1[12808] = 32'b11111111111111111011111001111011;
assign LUT_1[12809] = 32'b11111111111111110101001011110111;
assign LUT_1[12810] = 32'b11111111111111110111101000001100;
assign LUT_1[12811] = 32'b11111111111111110000111010001000;
assign LUT_1[12812] = 32'b00000000000000000011110011010010;
assign LUT_1[12813] = 32'b11111111111111111101000101001110;
assign LUT_1[12814] = 32'b11111111111111111111100001100011;
assign LUT_1[12815] = 32'b11111111111111111000110011011111;
assign LUT_1[12816] = 32'b11111111111111111110100111101000;
assign LUT_1[12817] = 32'b11111111111111110111111001100100;
assign LUT_1[12818] = 32'b11111111111111111010010101111001;
assign LUT_1[12819] = 32'b11111111111111110011100111110101;
assign LUT_1[12820] = 32'b00000000000000000110100000111111;
assign LUT_1[12821] = 32'b11111111111111111111110010111011;
assign LUT_1[12822] = 32'b00000000000000000010001111010000;
assign LUT_1[12823] = 32'b11111111111111111011100001001100;
assign LUT_1[12824] = 32'b11111111111111111101110101011101;
assign LUT_1[12825] = 32'b11111111111111110111000111011001;
assign LUT_1[12826] = 32'b11111111111111111001100011101110;
assign LUT_1[12827] = 32'b11111111111111110010110101101010;
assign LUT_1[12828] = 32'b00000000000000000101101110110100;
assign LUT_1[12829] = 32'b11111111111111111111000000110000;
assign LUT_1[12830] = 32'b00000000000000000001011101000101;
assign LUT_1[12831] = 32'b11111111111111111010101111000001;
assign LUT_1[12832] = 32'b11111111111111111101100111000101;
assign LUT_1[12833] = 32'b11111111111111110110111001000001;
assign LUT_1[12834] = 32'b11111111111111111001010101010110;
assign LUT_1[12835] = 32'b11111111111111110010100111010010;
assign LUT_1[12836] = 32'b00000000000000000101100000011100;
assign LUT_1[12837] = 32'b11111111111111111110110010011000;
assign LUT_1[12838] = 32'b00000000000000000001001110101101;
assign LUT_1[12839] = 32'b11111111111111111010100000101001;
assign LUT_1[12840] = 32'b11111111111111111100110100111010;
assign LUT_1[12841] = 32'b11111111111111110110000110110110;
assign LUT_1[12842] = 32'b11111111111111111000100011001011;
assign LUT_1[12843] = 32'b11111111111111110001110101000111;
assign LUT_1[12844] = 32'b00000000000000000100101110010001;
assign LUT_1[12845] = 32'b11111111111111111110000000001101;
assign LUT_1[12846] = 32'b00000000000000000000011100100010;
assign LUT_1[12847] = 32'b11111111111111111001101110011110;
assign LUT_1[12848] = 32'b11111111111111111111100010100111;
assign LUT_1[12849] = 32'b11111111111111111000110100100011;
assign LUT_1[12850] = 32'b11111111111111111011010000111000;
assign LUT_1[12851] = 32'b11111111111111110100100010110100;
assign LUT_1[12852] = 32'b00000000000000000111011011111110;
assign LUT_1[12853] = 32'b00000000000000000000101101111010;
assign LUT_1[12854] = 32'b00000000000000000011001010001111;
assign LUT_1[12855] = 32'b11111111111111111100011100001011;
assign LUT_1[12856] = 32'b11111111111111111110110000011100;
assign LUT_1[12857] = 32'b11111111111111111000000010011000;
assign LUT_1[12858] = 32'b11111111111111111010011110101101;
assign LUT_1[12859] = 32'b11111111111111110011110000101001;
assign LUT_1[12860] = 32'b00000000000000000110101001110011;
assign LUT_1[12861] = 32'b11111111111111111111111011101111;
assign LUT_1[12862] = 32'b00000000000000000010011000000100;
assign LUT_1[12863] = 32'b11111111111111111011101010000000;
assign LUT_1[12864] = 32'b11111111111111111110101001101110;
assign LUT_1[12865] = 32'b11111111111111110111111011101010;
assign LUT_1[12866] = 32'b11111111111111111010010111111111;
assign LUT_1[12867] = 32'b11111111111111110011101001111011;
assign LUT_1[12868] = 32'b00000000000000000110100011000101;
assign LUT_1[12869] = 32'b11111111111111111111110101000001;
assign LUT_1[12870] = 32'b00000000000000000010010001010110;
assign LUT_1[12871] = 32'b11111111111111111011100011010010;
assign LUT_1[12872] = 32'b11111111111111111101110111100011;
assign LUT_1[12873] = 32'b11111111111111110111001001011111;
assign LUT_1[12874] = 32'b11111111111111111001100101110100;
assign LUT_1[12875] = 32'b11111111111111110010110111110000;
assign LUT_1[12876] = 32'b00000000000000000101110000111010;
assign LUT_1[12877] = 32'b11111111111111111111000010110110;
assign LUT_1[12878] = 32'b00000000000000000001011111001011;
assign LUT_1[12879] = 32'b11111111111111111010110001000111;
assign LUT_1[12880] = 32'b00000000000000000000100101010000;
assign LUT_1[12881] = 32'b11111111111111111001110111001100;
assign LUT_1[12882] = 32'b11111111111111111100010011100001;
assign LUT_1[12883] = 32'b11111111111111110101100101011101;
assign LUT_1[12884] = 32'b00000000000000001000011110100111;
assign LUT_1[12885] = 32'b00000000000000000001110000100011;
assign LUT_1[12886] = 32'b00000000000000000100001100111000;
assign LUT_1[12887] = 32'b11111111111111111101011110110100;
assign LUT_1[12888] = 32'b11111111111111111111110011000101;
assign LUT_1[12889] = 32'b11111111111111111001000101000001;
assign LUT_1[12890] = 32'b11111111111111111011100001010110;
assign LUT_1[12891] = 32'b11111111111111110100110011010010;
assign LUT_1[12892] = 32'b00000000000000000111101100011100;
assign LUT_1[12893] = 32'b00000000000000000000111110011000;
assign LUT_1[12894] = 32'b00000000000000000011011010101101;
assign LUT_1[12895] = 32'b11111111111111111100101100101001;
assign LUT_1[12896] = 32'b11111111111111111111100100101101;
assign LUT_1[12897] = 32'b11111111111111111000110110101001;
assign LUT_1[12898] = 32'b11111111111111111011010010111110;
assign LUT_1[12899] = 32'b11111111111111110100100100111010;
assign LUT_1[12900] = 32'b00000000000000000111011110000100;
assign LUT_1[12901] = 32'b00000000000000000000110000000000;
assign LUT_1[12902] = 32'b00000000000000000011001100010101;
assign LUT_1[12903] = 32'b11111111111111111100011110010001;
assign LUT_1[12904] = 32'b11111111111111111110110010100010;
assign LUT_1[12905] = 32'b11111111111111111000000100011110;
assign LUT_1[12906] = 32'b11111111111111111010100000110011;
assign LUT_1[12907] = 32'b11111111111111110011110010101111;
assign LUT_1[12908] = 32'b00000000000000000110101011111001;
assign LUT_1[12909] = 32'b11111111111111111111111101110101;
assign LUT_1[12910] = 32'b00000000000000000010011010001010;
assign LUT_1[12911] = 32'b11111111111111111011101100000110;
assign LUT_1[12912] = 32'b00000000000000000001100000001111;
assign LUT_1[12913] = 32'b11111111111111111010110010001011;
assign LUT_1[12914] = 32'b11111111111111111101001110100000;
assign LUT_1[12915] = 32'b11111111111111110110100000011100;
assign LUT_1[12916] = 32'b00000000000000001001011001100110;
assign LUT_1[12917] = 32'b00000000000000000010101011100010;
assign LUT_1[12918] = 32'b00000000000000000101000111110111;
assign LUT_1[12919] = 32'b11111111111111111110011001110011;
assign LUT_1[12920] = 32'b00000000000000000000101110000100;
assign LUT_1[12921] = 32'b11111111111111111010000000000000;
assign LUT_1[12922] = 32'b11111111111111111100011100010101;
assign LUT_1[12923] = 32'b11111111111111110101101110010001;
assign LUT_1[12924] = 32'b00000000000000001000100111011011;
assign LUT_1[12925] = 32'b00000000000000000001111001010111;
assign LUT_1[12926] = 32'b00000000000000000100010101101100;
assign LUT_1[12927] = 32'b11111111111111111101100111101000;
assign LUT_1[12928] = 32'b11111111111111111111101100001001;
assign LUT_1[12929] = 32'b11111111111111111000111110000101;
assign LUT_1[12930] = 32'b11111111111111111011011010011010;
assign LUT_1[12931] = 32'b11111111111111110100101100010110;
assign LUT_1[12932] = 32'b00000000000000000111100101100000;
assign LUT_1[12933] = 32'b00000000000000000000110111011100;
assign LUT_1[12934] = 32'b00000000000000000011010011110001;
assign LUT_1[12935] = 32'b11111111111111111100100101101101;
assign LUT_1[12936] = 32'b11111111111111111110111001111110;
assign LUT_1[12937] = 32'b11111111111111111000001011111010;
assign LUT_1[12938] = 32'b11111111111111111010101000001111;
assign LUT_1[12939] = 32'b11111111111111110011111010001011;
assign LUT_1[12940] = 32'b00000000000000000110110011010101;
assign LUT_1[12941] = 32'b00000000000000000000000101010001;
assign LUT_1[12942] = 32'b00000000000000000010100001100110;
assign LUT_1[12943] = 32'b11111111111111111011110011100010;
assign LUT_1[12944] = 32'b00000000000000000001100111101011;
assign LUT_1[12945] = 32'b11111111111111111010111001100111;
assign LUT_1[12946] = 32'b11111111111111111101010101111100;
assign LUT_1[12947] = 32'b11111111111111110110100111111000;
assign LUT_1[12948] = 32'b00000000000000001001100001000010;
assign LUT_1[12949] = 32'b00000000000000000010110010111110;
assign LUT_1[12950] = 32'b00000000000000000101001111010011;
assign LUT_1[12951] = 32'b11111111111111111110100001001111;
assign LUT_1[12952] = 32'b00000000000000000000110101100000;
assign LUT_1[12953] = 32'b11111111111111111010000111011100;
assign LUT_1[12954] = 32'b11111111111111111100100011110001;
assign LUT_1[12955] = 32'b11111111111111110101110101101101;
assign LUT_1[12956] = 32'b00000000000000001000101110110111;
assign LUT_1[12957] = 32'b00000000000000000010000000110011;
assign LUT_1[12958] = 32'b00000000000000000100011101001000;
assign LUT_1[12959] = 32'b11111111111111111101101111000100;
assign LUT_1[12960] = 32'b00000000000000000000100111001000;
assign LUT_1[12961] = 32'b11111111111111111001111001000100;
assign LUT_1[12962] = 32'b11111111111111111100010101011001;
assign LUT_1[12963] = 32'b11111111111111110101100111010101;
assign LUT_1[12964] = 32'b00000000000000001000100000011111;
assign LUT_1[12965] = 32'b00000000000000000001110010011011;
assign LUT_1[12966] = 32'b00000000000000000100001110110000;
assign LUT_1[12967] = 32'b11111111111111111101100000101100;
assign LUT_1[12968] = 32'b11111111111111111111110100111101;
assign LUT_1[12969] = 32'b11111111111111111001000110111001;
assign LUT_1[12970] = 32'b11111111111111111011100011001110;
assign LUT_1[12971] = 32'b11111111111111110100110101001010;
assign LUT_1[12972] = 32'b00000000000000000111101110010100;
assign LUT_1[12973] = 32'b00000000000000000001000000010000;
assign LUT_1[12974] = 32'b00000000000000000011011100100101;
assign LUT_1[12975] = 32'b11111111111111111100101110100001;
assign LUT_1[12976] = 32'b00000000000000000010100010101010;
assign LUT_1[12977] = 32'b11111111111111111011110100100110;
assign LUT_1[12978] = 32'b11111111111111111110010000111011;
assign LUT_1[12979] = 32'b11111111111111110111100010110111;
assign LUT_1[12980] = 32'b00000000000000001010011100000001;
assign LUT_1[12981] = 32'b00000000000000000011101101111101;
assign LUT_1[12982] = 32'b00000000000000000110001010010010;
assign LUT_1[12983] = 32'b11111111111111111111011100001110;
assign LUT_1[12984] = 32'b00000000000000000001110000011111;
assign LUT_1[12985] = 32'b11111111111111111011000010011011;
assign LUT_1[12986] = 32'b11111111111111111101011110110000;
assign LUT_1[12987] = 32'b11111111111111110110110000101100;
assign LUT_1[12988] = 32'b00000000000000001001101001110110;
assign LUT_1[12989] = 32'b00000000000000000010111011110010;
assign LUT_1[12990] = 32'b00000000000000000101011000000111;
assign LUT_1[12991] = 32'b11111111111111111110101010000011;
assign LUT_1[12992] = 32'b00000000000000000001101001110001;
assign LUT_1[12993] = 32'b11111111111111111010111011101101;
assign LUT_1[12994] = 32'b11111111111111111101011000000010;
assign LUT_1[12995] = 32'b11111111111111110110101001111110;
assign LUT_1[12996] = 32'b00000000000000001001100011001000;
assign LUT_1[12997] = 32'b00000000000000000010110101000100;
assign LUT_1[12998] = 32'b00000000000000000101010001011001;
assign LUT_1[12999] = 32'b11111111111111111110100011010101;
assign LUT_1[13000] = 32'b00000000000000000000110111100110;
assign LUT_1[13001] = 32'b11111111111111111010001001100010;
assign LUT_1[13002] = 32'b11111111111111111100100101110111;
assign LUT_1[13003] = 32'b11111111111111110101110111110011;
assign LUT_1[13004] = 32'b00000000000000001000110000111101;
assign LUT_1[13005] = 32'b00000000000000000010000010111001;
assign LUT_1[13006] = 32'b00000000000000000100011111001110;
assign LUT_1[13007] = 32'b11111111111111111101110001001010;
assign LUT_1[13008] = 32'b00000000000000000011100101010011;
assign LUT_1[13009] = 32'b11111111111111111100110111001111;
assign LUT_1[13010] = 32'b11111111111111111111010011100100;
assign LUT_1[13011] = 32'b11111111111111111000100101100000;
assign LUT_1[13012] = 32'b00000000000000001011011110101010;
assign LUT_1[13013] = 32'b00000000000000000100110000100110;
assign LUT_1[13014] = 32'b00000000000000000111001100111011;
assign LUT_1[13015] = 32'b00000000000000000000011110110111;
assign LUT_1[13016] = 32'b00000000000000000010110011001000;
assign LUT_1[13017] = 32'b11111111111111111100000101000100;
assign LUT_1[13018] = 32'b11111111111111111110100001011001;
assign LUT_1[13019] = 32'b11111111111111110111110011010101;
assign LUT_1[13020] = 32'b00000000000000001010101100011111;
assign LUT_1[13021] = 32'b00000000000000000011111110011011;
assign LUT_1[13022] = 32'b00000000000000000110011010110000;
assign LUT_1[13023] = 32'b11111111111111111111101100101100;
assign LUT_1[13024] = 32'b00000000000000000010100100110000;
assign LUT_1[13025] = 32'b11111111111111111011110110101100;
assign LUT_1[13026] = 32'b11111111111111111110010011000001;
assign LUT_1[13027] = 32'b11111111111111110111100100111101;
assign LUT_1[13028] = 32'b00000000000000001010011110000111;
assign LUT_1[13029] = 32'b00000000000000000011110000000011;
assign LUT_1[13030] = 32'b00000000000000000110001100011000;
assign LUT_1[13031] = 32'b11111111111111111111011110010100;
assign LUT_1[13032] = 32'b00000000000000000001110010100101;
assign LUT_1[13033] = 32'b11111111111111111011000100100001;
assign LUT_1[13034] = 32'b11111111111111111101100000110110;
assign LUT_1[13035] = 32'b11111111111111110110110010110010;
assign LUT_1[13036] = 32'b00000000000000001001101011111100;
assign LUT_1[13037] = 32'b00000000000000000010111101111000;
assign LUT_1[13038] = 32'b00000000000000000101011010001101;
assign LUT_1[13039] = 32'b11111111111111111110101100001001;
assign LUT_1[13040] = 32'b00000000000000000100100000010010;
assign LUT_1[13041] = 32'b11111111111111111101110010001110;
assign LUT_1[13042] = 32'b00000000000000000000001110100011;
assign LUT_1[13043] = 32'b11111111111111111001100000011111;
assign LUT_1[13044] = 32'b00000000000000001100011001101001;
assign LUT_1[13045] = 32'b00000000000000000101101011100101;
assign LUT_1[13046] = 32'b00000000000000001000000111111010;
assign LUT_1[13047] = 32'b00000000000000000001011001110110;
assign LUT_1[13048] = 32'b00000000000000000011101110000111;
assign LUT_1[13049] = 32'b11111111111111111101000000000011;
assign LUT_1[13050] = 32'b11111111111111111111011100011000;
assign LUT_1[13051] = 32'b11111111111111111000101110010100;
assign LUT_1[13052] = 32'b00000000000000001011100111011110;
assign LUT_1[13053] = 32'b00000000000000000100111001011010;
assign LUT_1[13054] = 32'b00000000000000000111010101101111;
assign LUT_1[13055] = 32'b00000000000000000000100111101011;
assign LUT_1[13056] = 32'b11111111111111111010100000010010;
assign LUT_1[13057] = 32'b11111111111111110011110010001110;
assign LUT_1[13058] = 32'b11111111111111110110001110100011;
assign LUT_1[13059] = 32'b11111111111111101111100000011111;
assign LUT_1[13060] = 32'b00000000000000000010011001101001;
assign LUT_1[13061] = 32'b11111111111111111011101011100101;
assign LUT_1[13062] = 32'b11111111111111111110000111111010;
assign LUT_1[13063] = 32'b11111111111111110111011001110110;
assign LUT_1[13064] = 32'b11111111111111111001101110000111;
assign LUT_1[13065] = 32'b11111111111111110011000000000011;
assign LUT_1[13066] = 32'b11111111111111110101011100011000;
assign LUT_1[13067] = 32'b11111111111111101110101110010100;
assign LUT_1[13068] = 32'b00000000000000000001100111011110;
assign LUT_1[13069] = 32'b11111111111111111010111001011010;
assign LUT_1[13070] = 32'b11111111111111111101010101101111;
assign LUT_1[13071] = 32'b11111111111111110110100111101011;
assign LUT_1[13072] = 32'b11111111111111111100011011110100;
assign LUT_1[13073] = 32'b11111111111111110101101101110000;
assign LUT_1[13074] = 32'b11111111111111111000001010000101;
assign LUT_1[13075] = 32'b11111111111111110001011100000001;
assign LUT_1[13076] = 32'b00000000000000000100010101001011;
assign LUT_1[13077] = 32'b11111111111111111101100111000111;
assign LUT_1[13078] = 32'b00000000000000000000000011011100;
assign LUT_1[13079] = 32'b11111111111111111001010101011000;
assign LUT_1[13080] = 32'b11111111111111111011101001101001;
assign LUT_1[13081] = 32'b11111111111111110100111011100101;
assign LUT_1[13082] = 32'b11111111111111110111010111111010;
assign LUT_1[13083] = 32'b11111111111111110000101001110110;
assign LUT_1[13084] = 32'b00000000000000000011100011000000;
assign LUT_1[13085] = 32'b11111111111111111100110100111100;
assign LUT_1[13086] = 32'b11111111111111111111010001010001;
assign LUT_1[13087] = 32'b11111111111111111000100011001101;
assign LUT_1[13088] = 32'b11111111111111111011011011010001;
assign LUT_1[13089] = 32'b11111111111111110100101101001101;
assign LUT_1[13090] = 32'b11111111111111110111001001100010;
assign LUT_1[13091] = 32'b11111111111111110000011011011110;
assign LUT_1[13092] = 32'b00000000000000000011010100101000;
assign LUT_1[13093] = 32'b11111111111111111100100110100100;
assign LUT_1[13094] = 32'b11111111111111111111000010111001;
assign LUT_1[13095] = 32'b11111111111111111000010100110101;
assign LUT_1[13096] = 32'b11111111111111111010101001000110;
assign LUT_1[13097] = 32'b11111111111111110011111011000010;
assign LUT_1[13098] = 32'b11111111111111110110010111010111;
assign LUT_1[13099] = 32'b11111111111111101111101001010011;
assign LUT_1[13100] = 32'b00000000000000000010100010011101;
assign LUT_1[13101] = 32'b11111111111111111011110100011001;
assign LUT_1[13102] = 32'b11111111111111111110010000101110;
assign LUT_1[13103] = 32'b11111111111111110111100010101010;
assign LUT_1[13104] = 32'b11111111111111111101010110110011;
assign LUT_1[13105] = 32'b11111111111111110110101000101111;
assign LUT_1[13106] = 32'b11111111111111111001000101000100;
assign LUT_1[13107] = 32'b11111111111111110010010111000000;
assign LUT_1[13108] = 32'b00000000000000000101010000001010;
assign LUT_1[13109] = 32'b11111111111111111110100010000110;
assign LUT_1[13110] = 32'b00000000000000000000111110011011;
assign LUT_1[13111] = 32'b11111111111111111010010000010111;
assign LUT_1[13112] = 32'b11111111111111111100100100101000;
assign LUT_1[13113] = 32'b11111111111111110101110110100100;
assign LUT_1[13114] = 32'b11111111111111111000010010111001;
assign LUT_1[13115] = 32'b11111111111111110001100100110101;
assign LUT_1[13116] = 32'b00000000000000000100011101111111;
assign LUT_1[13117] = 32'b11111111111111111101101111111011;
assign LUT_1[13118] = 32'b00000000000000000000001100010000;
assign LUT_1[13119] = 32'b11111111111111111001011110001100;
assign LUT_1[13120] = 32'b11111111111111111100011101111010;
assign LUT_1[13121] = 32'b11111111111111110101101111110110;
assign LUT_1[13122] = 32'b11111111111111111000001100001011;
assign LUT_1[13123] = 32'b11111111111111110001011110000111;
assign LUT_1[13124] = 32'b00000000000000000100010111010001;
assign LUT_1[13125] = 32'b11111111111111111101101001001101;
assign LUT_1[13126] = 32'b00000000000000000000000101100010;
assign LUT_1[13127] = 32'b11111111111111111001010111011110;
assign LUT_1[13128] = 32'b11111111111111111011101011101111;
assign LUT_1[13129] = 32'b11111111111111110100111101101011;
assign LUT_1[13130] = 32'b11111111111111110111011010000000;
assign LUT_1[13131] = 32'b11111111111111110000101011111100;
assign LUT_1[13132] = 32'b00000000000000000011100101000110;
assign LUT_1[13133] = 32'b11111111111111111100110111000010;
assign LUT_1[13134] = 32'b11111111111111111111010011010111;
assign LUT_1[13135] = 32'b11111111111111111000100101010011;
assign LUT_1[13136] = 32'b11111111111111111110011001011100;
assign LUT_1[13137] = 32'b11111111111111110111101011011000;
assign LUT_1[13138] = 32'b11111111111111111010000111101101;
assign LUT_1[13139] = 32'b11111111111111110011011001101001;
assign LUT_1[13140] = 32'b00000000000000000110010010110011;
assign LUT_1[13141] = 32'b11111111111111111111100100101111;
assign LUT_1[13142] = 32'b00000000000000000010000001000100;
assign LUT_1[13143] = 32'b11111111111111111011010011000000;
assign LUT_1[13144] = 32'b11111111111111111101100111010001;
assign LUT_1[13145] = 32'b11111111111111110110111001001101;
assign LUT_1[13146] = 32'b11111111111111111001010101100010;
assign LUT_1[13147] = 32'b11111111111111110010100111011110;
assign LUT_1[13148] = 32'b00000000000000000101100000101000;
assign LUT_1[13149] = 32'b11111111111111111110110010100100;
assign LUT_1[13150] = 32'b00000000000000000001001110111001;
assign LUT_1[13151] = 32'b11111111111111111010100000110101;
assign LUT_1[13152] = 32'b11111111111111111101011000111001;
assign LUT_1[13153] = 32'b11111111111111110110101010110101;
assign LUT_1[13154] = 32'b11111111111111111001000111001010;
assign LUT_1[13155] = 32'b11111111111111110010011001000110;
assign LUT_1[13156] = 32'b00000000000000000101010010010000;
assign LUT_1[13157] = 32'b11111111111111111110100100001100;
assign LUT_1[13158] = 32'b00000000000000000001000000100001;
assign LUT_1[13159] = 32'b11111111111111111010010010011101;
assign LUT_1[13160] = 32'b11111111111111111100100110101110;
assign LUT_1[13161] = 32'b11111111111111110101111000101010;
assign LUT_1[13162] = 32'b11111111111111111000010100111111;
assign LUT_1[13163] = 32'b11111111111111110001100110111011;
assign LUT_1[13164] = 32'b00000000000000000100100000000101;
assign LUT_1[13165] = 32'b11111111111111111101110010000001;
assign LUT_1[13166] = 32'b00000000000000000000001110010110;
assign LUT_1[13167] = 32'b11111111111111111001100000010010;
assign LUT_1[13168] = 32'b11111111111111111111010100011011;
assign LUT_1[13169] = 32'b11111111111111111000100110010111;
assign LUT_1[13170] = 32'b11111111111111111011000010101100;
assign LUT_1[13171] = 32'b11111111111111110100010100101000;
assign LUT_1[13172] = 32'b00000000000000000111001101110010;
assign LUT_1[13173] = 32'b00000000000000000000011111101110;
assign LUT_1[13174] = 32'b00000000000000000010111100000011;
assign LUT_1[13175] = 32'b11111111111111111100001101111111;
assign LUT_1[13176] = 32'b11111111111111111110100010010000;
assign LUT_1[13177] = 32'b11111111111111110111110100001100;
assign LUT_1[13178] = 32'b11111111111111111010010000100001;
assign LUT_1[13179] = 32'b11111111111111110011100010011101;
assign LUT_1[13180] = 32'b00000000000000000110011011100111;
assign LUT_1[13181] = 32'b11111111111111111111101101100011;
assign LUT_1[13182] = 32'b00000000000000000010001001111000;
assign LUT_1[13183] = 32'b11111111111111111011011011110100;
assign LUT_1[13184] = 32'b11111111111111111101100000010101;
assign LUT_1[13185] = 32'b11111111111111110110110010010001;
assign LUT_1[13186] = 32'b11111111111111111001001110100110;
assign LUT_1[13187] = 32'b11111111111111110010100000100010;
assign LUT_1[13188] = 32'b00000000000000000101011001101100;
assign LUT_1[13189] = 32'b11111111111111111110101011101000;
assign LUT_1[13190] = 32'b00000000000000000001000111111101;
assign LUT_1[13191] = 32'b11111111111111111010011001111001;
assign LUT_1[13192] = 32'b11111111111111111100101110001010;
assign LUT_1[13193] = 32'b11111111111111110110000000000110;
assign LUT_1[13194] = 32'b11111111111111111000011100011011;
assign LUT_1[13195] = 32'b11111111111111110001101110010111;
assign LUT_1[13196] = 32'b00000000000000000100100111100001;
assign LUT_1[13197] = 32'b11111111111111111101111001011101;
assign LUT_1[13198] = 32'b00000000000000000000010101110010;
assign LUT_1[13199] = 32'b11111111111111111001100111101110;
assign LUT_1[13200] = 32'b11111111111111111111011011110111;
assign LUT_1[13201] = 32'b11111111111111111000101101110011;
assign LUT_1[13202] = 32'b11111111111111111011001010001000;
assign LUT_1[13203] = 32'b11111111111111110100011100000100;
assign LUT_1[13204] = 32'b00000000000000000111010101001110;
assign LUT_1[13205] = 32'b00000000000000000000100111001010;
assign LUT_1[13206] = 32'b00000000000000000011000011011111;
assign LUT_1[13207] = 32'b11111111111111111100010101011011;
assign LUT_1[13208] = 32'b11111111111111111110101001101100;
assign LUT_1[13209] = 32'b11111111111111110111111011101000;
assign LUT_1[13210] = 32'b11111111111111111010010111111101;
assign LUT_1[13211] = 32'b11111111111111110011101001111001;
assign LUT_1[13212] = 32'b00000000000000000110100011000011;
assign LUT_1[13213] = 32'b11111111111111111111110100111111;
assign LUT_1[13214] = 32'b00000000000000000010010001010100;
assign LUT_1[13215] = 32'b11111111111111111011100011010000;
assign LUT_1[13216] = 32'b11111111111111111110011011010100;
assign LUT_1[13217] = 32'b11111111111111110111101101010000;
assign LUT_1[13218] = 32'b11111111111111111010001001100101;
assign LUT_1[13219] = 32'b11111111111111110011011011100001;
assign LUT_1[13220] = 32'b00000000000000000110010100101011;
assign LUT_1[13221] = 32'b11111111111111111111100110100111;
assign LUT_1[13222] = 32'b00000000000000000010000010111100;
assign LUT_1[13223] = 32'b11111111111111111011010100111000;
assign LUT_1[13224] = 32'b11111111111111111101101001001001;
assign LUT_1[13225] = 32'b11111111111111110110111011000101;
assign LUT_1[13226] = 32'b11111111111111111001010111011010;
assign LUT_1[13227] = 32'b11111111111111110010101001010110;
assign LUT_1[13228] = 32'b00000000000000000101100010100000;
assign LUT_1[13229] = 32'b11111111111111111110110100011100;
assign LUT_1[13230] = 32'b00000000000000000001010000110001;
assign LUT_1[13231] = 32'b11111111111111111010100010101101;
assign LUT_1[13232] = 32'b00000000000000000000010110110110;
assign LUT_1[13233] = 32'b11111111111111111001101000110010;
assign LUT_1[13234] = 32'b11111111111111111100000101000111;
assign LUT_1[13235] = 32'b11111111111111110101010111000011;
assign LUT_1[13236] = 32'b00000000000000001000010000001101;
assign LUT_1[13237] = 32'b00000000000000000001100010001001;
assign LUT_1[13238] = 32'b00000000000000000011111110011110;
assign LUT_1[13239] = 32'b11111111111111111101010000011010;
assign LUT_1[13240] = 32'b11111111111111111111100100101011;
assign LUT_1[13241] = 32'b11111111111111111000110110100111;
assign LUT_1[13242] = 32'b11111111111111111011010010111100;
assign LUT_1[13243] = 32'b11111111111111110100100100111000;
assign LUT_1[13244] = 32'b00000000000000000111011110000010;
assign LUT_1[13245] = 32'b00000000000000000000101111111110;
assign LUT_1[13246] = 32'b00000000000000000011001100010011;
assign LUT_1[13247] = 32'b11111111111111111100011110001111;
assign LUT_1[13248] = 32'b11111111111111111111011101111101;
assign LUT_1[13249] = 32'b11111111111111111000101111111001;
assign LUT_1[13250] = 32'b11111111111111111011001100001110;
assign LUT_1[13251] = 32'b11111111111111110100011110001010;
assign LUT_1[13252] = 32'b00000000000000000111010111010100;
assign LUT_1[13253] = 32'b00000000000000000000101001010000;
assign LUT_1[13254] = 32'b00000000000000000011000101100101;
assign LUT_1[13255] = 32'b11111111111111111100010111100001;
assign LUT_1[13256] = 32'b11111111111111111110101011110010;
assign LUT_1[13257] = 32'b11111111111111110111111101101110;
assign LUT_1[13258] = 32'b11111111111111111010011010000011;
assign LUT_1[13259] = 32'b11111111111111110011101011111111;
assign LUT_1[13260] = 32'b00000000000000000110100101001001;
assign LUT_1[13261] = 32'b11111111111111111111110111000101;
assign LUT_1[13262] = 32'b00000000000000000010010011011010;
assign LUT_1[13263] = 32'b11111111111111111011100101010110;
assign LUT_1[13264] = 32'b00000000000000000001011001011111;
assign LUT_1[13265] = 32'b11111111111111111010101011011011;
assign LUT_1[13266] = 32'b11111111111111111101000111110000;
assign LUT_1[13267] = 32'b11111111111111110110011001101100;
assign LUT_1[13268] = 32'b00000000000000001001010010110110;
assign LUT_1[13269] = 32'b00000000000000000010100100110010;
assign LUT_1[13270] = 32'b00000000000000000101000001000111;
assign LUT_1[13271] = 32'b11111111111111111110010011000011;
assign LUT_1[13272] = 32'b00000000000000000000100111010100;
assign LUT_1[13273] = 32'b11111111111111111001111001010000;
assign LUT_1[13274] = 32'b11111111111111111100010101100101;
assign LUT_1[13275] = 32'b11111111111111110101100111100001;
assign LUT_1[13276] = 32'b00000000000000001000100000101011;
assign LUT_1[13277] = 32'b00000000000000000001110010100111;
assign LUT_1[13278] = 32'b00000000000000000100001110111100;
assign LUT_1[13279] = 32'b11111111111111111101100000111000;
assign LUT_1[13280] = 32'b00000000000000000000011000111100;
assign LUT_1[13281] = 32'b11111111111111111001101010111000;
assign LUT_1[13282] = 32'b11111111111111111100000111001101;
assign LUT_1[13283] = 32'b11111111111111110101011001001001;
assign LUT_1[13284] = 32'b00000000000000001000010010010011;
assign LUT_1[13285] = 32'b00000000000000000001100100001111;
assign LUT_1[13286] = 32'b00000000000000000100000000100100;
assign LUT_1[13287] = 32'b11111111111111111101010010100000;
assign LUT_1[13288] = 32'b11111111111111111111100110110001;
assign LUT_1[13289] = 32'b11111111111111111000111000101101;
assign LUT_1[13290] = 32'b11111111111111111011010101000010;
assign LUT_1[13291] = 32'b11111111111111110100100110111110;
assign LUT_1[13292] = 32'b00000000000000000111100000001000;
assign LUT_1[13293] = 32'b00000000000000000000110010000100;
assign LUT_1[13294] = 32'b00000000000000000011001110011001;
assign LUT_1[13295] = 32'b11111111111111111100100000010101;
assign LUT_1[13296] = 32'b00000000000000000010010100011110;
assign LUT_1[13297] = 32'b11111111111111111011100110011010;
assign LUT_1[13298] = 32'b11111111111111111110000010101111;
assign LUT_1[13299] = 32'b11111111111111110111010100101011;
assign LUT_1[13300] = 32'b00000000000000001010001101110101;
assign LUT_1[13301] = 32'b00000000000000000011011111110001;
assign LUT_1[13302] = 32'b00000000000000000101111100000110;
assign LUT_1[13303] = 32'b11111111111111111111001110000010;
assign LUT_1[13304] = 32'b00000000000000000001100010010011;
assign LUT_1[13305] = 32'b11111111111111111010110100001111;
assign LUT_1[13306] = 32'b11111111111111111101010000100100;
assign LUT_1[13307] = 32'b11111111111111110110100010100000;
assign LUT_1[13308] = 32'b00000000000000001001011011101010;
assign LUT_1[13309] = 32'b00000000000000000010101101100110;
assign LUT_1[13310] = 32'b00000000000000000101001001111011;
assign LUT_1[13311] = 32'b11111111111111111110011011110111;
assign LUT_1[13312] = 32'b00000000000000001001010100011001;
assign LUT_1[13313] = 32'b00000000000000000010100110010101;
assign LUT_1[13314] = 32'b00000000000000000101000010101010;
assign LUT_1[13315] = 32'b11111111111111111110010100100110;
assign LUT_1[13316] = 32'b00000000000000010001001101110000;
assign LUT_1[13317] = 32'b00000000000000001010011111101100;
assign LUT_1[13318] = 32'b00000000000000001100111100000001;
assign LUT_1[13319] = 32'b00000000000000000110001101111101;
assign LUT_1[13320] = 32'b00000000000000001000100010001110;
assign LUT_1[13321] = 32'b00000000000000000001110100001010;
assign LUT_1[13322] = 32'b00000000000000000100010000011111;
assign LUT_1[13323] = 32'b11111111111111111101100010011011;
assign LUT_1[13324] = 32'b00000000000000010000011011100101;
assign LUT_1[13325] = 32'b00000000000000001001101101100001;
assign LUT_1[13326] = 32'b00000000000000001100001001110110;
assign LUT_1[13327] = 32'b00000000000000000101011011110010;
assign LUT_1[13328] = 32'b00000000000000001011001111111011;
assign LUT_1[13329] = 32'b00000000000000000100100001110111;
assign LUT_1[13330] = 32'b00000000000000000110111110001100;
assign LUT_1[13331] = 32'b00000000000000000000010000001000;
assign LUT_1[13332] = 32'b00000000000000010011001001010010;
assign LUT_1[13333] = 32'b00000000000000001100011011001110;
assign LUT_1[13334] = 32'b00000000000000001110110111100011;
assign LUT_1[13335] = 32'b00000000000000001000001001011111;
assign LUT_1[13336] = 32'b00000000000000001010011101110000;
assign LUT_1[13337] = 32'b00000000000000000011101111101100;
assign LUT_1[13338] = 32'b00000000000000000110001100000001;
assign LUT_1[13339] = 32'b11111111111111111111011101111101;
assign LUT_1[13340] = 32'b00000000000000010010010111000111;
assign LUT_1[13341] = 32'b00000000000000001011101001000011;
assign LUT_1[13342] = 32'b00000000000000001110000101011000;
assign LUT_1[13343] = 32'b00000000000000000111010111010100;
assign LUT_1[13344] = 32'b00000000000000001010001111011000;
assign LUT_1[13345] = 32'b00000000000000000011100001010100;
assign LUT_1[13346] = 32'b00000000000000000101111101101001;
assign LUT_1[13347] = 32'b11111111111111111111001111100101;
assign LUT_1[13348] = 32'b00000000000000010010001000101111;
assign LUT_1[13349] = 32'b00000000000000001011011010101011;
assign LUT_1[13350] = 32'b00000000000000001101110111000000;
assign LUT_1[13351] = 32'b00000000000000000111001000111100;
assign LUT_1[13352] = 32'b00000000000000001001011101001101;
assign LUT_1[13353] = 32'b00000000000000000010101111001001;
assign LUT_1[13354] = 32'b00000000000000000101001011011110;
assign LUT_1[13355] = 32'b11111111111111111110011101011010;
assign LUT_1[13356] = 32'b00000000000000010001010110100100;
assign LUT_1[13357] = 32'b00000000000000001010101000100000;
assign LUT_1[13358] = 32'b00000000000000001101000100110101;
assign LUT_1[13359] = 32'b00000000000000000110010110110001;
assign LUT_1[13360] = 32'b00000000000000001100001010111010;
assign LUT_1[13361] = 32'b00000000000000000101011100110110;
assign LUT_1[13362] = 32'b00000000000000000111111001001011;
assign LUT_1[13363] = 32'b00000000000000000001001011000111;
assign LUT_1[13364] = 32'b00000000000000010100000100010001;
assign LUT_1[13365] = 32'b00000000000000001101010110001101;
assign LUT_1[13366] = 32'b00000000000000001111110010100010;
assign LUT_1[13367] = 32'b00000000000000001001000100011110;
assign LUT_1[13368] = 32'b00000000000000001011011000101111;
assign LUT_1[13369] = 32'b00000000000000000100101010101011;
assign LUT_1[13370] = 32'b00000000000000000111000111000000;
assign LUT_1[13371] = 32'b00000000000000000000011000111100;
assign LUT_1[13372] = 32'b00000000000000010011010010000110;
assign LUT_1[13373] = 32'b00000000000000001100100100000010;
assign LUT_1[13374] = 32'b00000000000000001111000000010111;
assign LUT_1[13375] = 32'b00000000000000001000010010010011;
assign LUT_1[13376] = 32'b00000000000000001011010010000001;
assign LUT_1[13377] = 32'b00000000000000000100100011111101;
assign LUT_1[13378] = 32'b00000000000000000111000000010010;
assign LUT_1[13379] = 32'b00000000000000000000010010001110;
assign LUT_1[13380] = 32'b00000000000000010011001011011000;
assign LUT_1[13381] = 32'b00000000000000001100011101010100;
assign LUT_1[13382] = 32'b00000000000000001110111001101001;
assign LUT_1[13383] = 32'b00000000000000001000001011100101;
assign LUT_1[13384] = 32'b00000000000000001010011111110110;
assign LUT_1[13385] = 32'b00000000000000000011110001110010;
assign LUT_1[13386] = 32'b00000000000000000110001110000111;
assign LUT_1[13387] = 32'b11111111111111111111100000000011;
assign LUT_1[13388] = 32'b00000000000000010010011001001101;
assign LUT_1[13389] = 32'b00000000000000001011101011001001;
assign LUT_1[13390] = 32'b00000000000000001110000111011110;
assign LUT_1[13391] = 32'b00000000000000000111011001011010;
assign LUT_1[13392] = 32'b00000000000000001101001101100011;
assign LUT_1[13393] = 32'b00000000000000000110011111011111;
assign LUT_1[13394] = 32'b00000000000000001000111011110100;
assign LUT_1[13395] = 32'b00000000000000000010001101110000;
assign LUT_1[13396] = 32'b00000000000000010101000110111010;
assign LUT_1[13397] = 32'b00000000000000001110011000110110;
assign LUT_1[13398] = 32'b00000000000000010000110101001011;
assign LUT_1[13399] = 32'b00000000000000001010000111000111;
assign LUT_1[13400] = 32'b00000000000000001100011011011000;
assign LUT_1[13401] = 32'b00000000000000000101101101010100;
assign LUT_1[13402] = 32'b00000000000000001000001001101001;
assign LUT_1[13403] = 32'b00000000000000000001011011100101;
assign LUT_1[13404] = 32'b00000000000000010100010100101111;
assign LUT_1[13405] = 32'b00000000000000001101100110101011;
assign LUT_1[13406] = 32'b00000000000000010000000011000000;
assign LUT_1[13407] = 32'b00000000000000001001010100111100;
assign LUT_1[13408] = 32'b00000000000000001100001101000000;
assign LUT_1[13409] = 32'b00000000000000000101011110111100;
assign LUT_1[13410] = 32'b00000000000000000111111011010001;
assign LUT_1[13411] = 32'b00000000000000000001001101001101;
assign LUT_1[13412] = 32'b00000000000000010100000110010111;
assign LUT_1[13413] = 32'b00000000000000001101011000010011;
assign LUT_1[13414] = 32'b00000000000000001111110100101000;
assign LUT_1[13415] = 32'b00000000000000001001000110100100;
assign LUT_1[13416] = 32'b00000000000000001011011010110101;
assign LUT_1[13417] = 32'b00000000000000000100101100110001;
assign LUT_1[13418] = 32'b00000000000000000111001001000110;
assign LUT_1[13419] = 32'b00000000000000000000011011000010;
assign LUT_1[13420] = 32'b00000000000000010011010100001100;
assign LUT_1[13421] = 32'b00000000000000001100100110001000;
assign LUT_1[13422] = 32'b00000000000000001111000010011101;
assign LUT_1[13423] = 32'b00000000000000001000010100011001;
assign LUT_1[13424] = 32'b00000000000000001110001000100010;
assign LUT_1[13425] = 32'b00000000000000000111011010011110;
assign LUT_1[13426] = 32'b00000000000000001001110110110011;
assign LUT_1[13427] = 32'b00000000000000000011001000101111;
assign LUT_1[13428] = 32'b00000000000000010110000001111001;
assign LUT_1[13429] = 32'b00000000000000001111010011110101;
assign LUT_1[13430] = 32'b00000000000000010001110000001010;
assign LUT_1[13431] = 32'b00000000000000001011000010000110;
assign LUT_1[13432] = 32'b00000000000000001101010110010111;
assign LUT_1[13433] = 32'b00000000000000000110101000010011;
assign LUT_1[13434] = 32'b00000000000000001001000100101000;
assign LUT_1[13435] = 32'b00000000000000000010010110100100;
assign LUT_1[13436] = 32'b00000000000000010101001111101110;
assign LUT_1[13437] = 32'b00000000000000001110100001101010;
assign LUT_1[13438] = 32'b00000000000000010000111101111111;
assign LUT_1[13439] = 32'b00000000000000001010001111111011;
assign LUT_1[13440] = 32'b00000000000000001100010100011100;
assign LUT_1[13441] = 32'b00000000000000000101100110011000;
assign LUT_1[13442] = 32'b00000000000000001000000010101101;
assign LUT_1[13443] = 32'b00000000000000000001010100101001;
assign LUT_1[13444] = 32'b00000000000000010100001101110011;
assign LUT_1[13445] = 32'b00000000000000001101011111101111;
assign LUT_1[13446] = 32'b00000000000000001111111100000100;
assign LUT_1[13447] = 32'b00000000000000001001001110000000;
assign LUT_1[13448] = 32'b00000000000000001011100010010001;
assign LUT_1[13449] = 32'b00000000000000000100110100001101;
assign LUT_1[13450] = 32'b00000000000000000111010000100010;
assign LUT_1[13451] = 32'b00000000000000000000100010011110;
assign LUT_1[13452] = 32'b00000000000000010011011011101000;
assign LUT_1[13453] = 32'b00000000000000001100101101100100;
assign LUT_1[13454] = 32'b00000000000000001111001001111001;
assign LUT_1[13455] = 32'b00000000000000001000011011110101;
assign LUT_1[13456] = 32'b00000000000000001110001111111110;
assign LUT_1[13457] = 32'b00000000000000000111100001111010;
assign LUT_1[13458] = 32'b00000000000000001001111110001111;
assign LUT_1[13459] = 32'b00000000000000000011010000001011;
assign LUT_1[13460] = 32'b00000000000000010110001001010101;
assign LUT_1[13461] = 32'b00000000000000001111011011010001;
assign LUT_1[13462] = 32'b00000000000000010001110111100110;
assign LUT_1[13463] = 32'b00000000000000001011001001100010;
assign LUT_1[13464] = 32'b00000000000000001101011101110011;
assign LUT_1[13465] = 32'b00000000000000000110101111101111;
assign LUT_1[13466] = 32'b00000000000000001001001100000100;
assign LUT_1[13467] = 32'b00000000000000000010011110000000;
assign LUT_1[13468] = 32'b00000000000000010101010111001010;
assign LUT_1[13469] = 32'b00000000000000001110101001000110;
assign LUT_1[13470] = 32'b00000000000000010001000101011011;
assign LUT_1[13471] = 32'b00000000000000001010010111010111;
assign LUT_1[13472] = 32'b00000000000000001101001111011011;
assign LUT_1[13473] = 32'b00000000000000000110100001010111;
assign LUT_1[13474] = 32'b00000000000000001000111101101100;
assign LUT_1[13475] = 32'b00000000000000000010001111101000;
assign LUT_1[13476] = 32'b00000000000000010101001000110010;
assign LUT_1[13477] = 32'b00000000000000001110011010101110;
assign LUT_1[13478] = 32'b00000000000000010000110111000011;
assign LUT_1[13479] = 32'b00000000000000001010001000111111;
assign LUT_1[13480] = 32'b00000000000000001100011101010000;
assign LUT_1[13481] = 32'b00000000000000000101101111001100;
assign LUT_1[13482] = 32'b00000000000000001000001011100001;
assign LUT_1[13483] = 32'b00000000000000000001011101011101;
assign LUT_1[13484] = 32'b00000000000000010100010110100111;
assign LUT_1[13485] = 32'b00000000000000001101101000100011;
assign LUT_1[13486] = 32'b00000000000000010000000100111000;
assign LUT_1[13487] = 32'b00000000000000001001010110110100;
assign LUT_1[13488] = 32'b00000000000000001111001010111101;
assign LUT_1[13489] = 32'b00000000000000001000011100111001;
assign LUT_1[13490] = 32'b00000000000000001010111001001110;
assign LUT_1[13491] = 32'b00000000000000000100001011001010;
assign LUT_1[13492] = 32'b00000000000000010111000100010100;
assign LUT_1[13493] = 32'b00000000000000010000010110010000;
assign LUT_1[13494] = 32'b00000000000000010010110010100101;
assign LUT_1[13495] = 32'b00000000000000001100000100100001;
assign LUT_1[13496] = 32'b00000000000000001110011000110010;
assign LUT_1[13497] = 32'b00000000000000000111101010101110;
assign LUT_1[13498] = 32'b00000000000000001010000111000011;
assign LUT_1[13499] = 32'b00000000000000000011011000111111;
assign LUT_1[13500] = 32'b00000000000000010110010010001001;
assign LUT_1[13501] = 32'b00000000000000001111100100000101;
assign LUT_1[13502] = 32'b00000000000000010010000000011010;
assign LUT_1[13503] = 32'b00000000000000001011010010010110;
assign LUT_1[13504] = 32'b00000000000000001110010010000100;
assign LUT_1[13505] = 32'b00000000000000000111100100000000;
assign LUT_1[13506] = 32'b00000000000000001010000000010101;
assign LUT_1[13507] = 32'b00000000000000000011010010010001;
assign LUT_1[13508] = 32'b00000000000000010110001011011011;
assign LUT_1[13509] = 32'b00000000000000001111011101010111;
assign LUT_1[13510] = 32'b00000000000000010001111001101100;
assign LUT_1[13511] = 32'b00000000000000001011001011101000;
assign LUT_1[13512] = 32'b00000000000000001101011111111001;
assign LUT_1[13513] = 32'b00000000000000000110110001110101;
assign LUT_1[13514] = 32'b00000000000000001001001110001010;
assign LUT_1[13515] = 32'b00000000000000000010100000000110;
assign LUT_1[13516] = 32'b00000000000000010101011001010000;
assign LUT_1[13517] = 32'b00000000000000001110101011001100;
assign LUT_1[13518] = 32'b00000000000000010001000111100001;
assign LUT_1[13519] = 32'b00000000000000001010011001011101;
assign LUT_1[13520] = 32'b00000000000000010000001101100110;
assign LUT_1[13521] = 32'b00000000000000001001011111100010;
assign LUT_1[13522] = 32'b00000000000000001011111011110111;
assign LUT_1[13523] = 32'b00000000000000000101001101110011;
assign LUT_1[13524] = 32'b00000000000000011000000110111101;
assign LUT_1[13525] = 32'b00000000000000010001011000111001;
assign LUT_1[13526] = 32'b00000000000000010011110101001110;
assign LUT_1[13527] = 32'b00000000000000001101000111001010;
assign LUT_1[13528] = 32'b00000000000000001111011011011011;
assign LUT_1[13529] = 32'b00000000000000001000101101010111;
assign LUT_1[13530] = 32'b00000000000000001011001001101100;
assign LUT_1[13531] = 32'b00000000000000000100011011101000;
assign LUT_1[13532] = 32'b00000000000000010111010100110010;
assign LUT_1[13533] = 32'b00000000000000010000100110101110;
assign LUT_1[13534] = 32'b00000000000000010011000011000011;
assign LUT_1[13535] = 32'b00000000000000001100010100111111;
assign LUT_1[13536] = 32'b00000000000000001111001101000011;
assign LUT_1[13537] = 32'b00000000000000001000011110111111;
assign LUT_1[13538] = 32'b00000000000000001010111011010100;
assign LUT_1[13539] = 32'b00000000000000000100001101010000;
assign LUT_1[13540] = 32'b00000000000000010111000110011010;
assign LUT_1[13541] = 32'b00000000000000010000011000010110;
assign LUT_1[13542] = 32'b00000000000000010010110100101011;
assign LUT_1[13543] = 32'b00000000000000001100000110100111;
assign LUT_1[13544] = 32'b00000000000000001110011010111000;
assign LUT_1[13545] = 32'b00000000000000000111101100110100;
assign LUT_1[13546] = 32'b00000000000000001010001001001001;
assign LUT_1[13547] = 32'b00000000000000000011011011000101;
assign LUT_1[13548] = 32'b00000000000000010110010100001111;
assign LUT_1[13549] = 32'b00000000000000001111100110001011;
assign LUT_1[13550] = 32'b00000000000000010010000010100000;
assign LUT_1[13551] = 32'b00000000000000001011010100011100;
assign LUT_1[13552] = 32'b00000000000000010001001000100101;
assign LUT_1[13553] = 32'b00000000000000001010011010100001;
assign LUT_1[13554] = 32'b00000000000000001100110110110110;
assign LUT_1[13555] = 32'b00000000000000000110001000110010;
assign LUT_1[13556] = 32'b00000000000000011001000001111100;
assign LUT_1[13557] = 32'b00000000000000010010010011111000;
assign LUT_1[13558] = 32'b00000000000000010100110000001101;
assign LUT_1[13559] = 32'b00000000000000001110000010001001;
assign LUT_1[13560] = 32'b00000000000000010000010110011010;
assign LUT_1[13561] = 32'b00000000000000001001101000010110;
assign LUT_1[13562] = 32'b00000000000000001100000100101011;
assign LUT_1[13563] = 32'b00000000000000000101010110100111;
assign LUT_1[13564] = 32'b00000000000000011000001111110001;
assign LUT_1[13565] = 32'b00000000000000010001100001101101;
assign LUT_1[13566] = 32'b00000000000000010011111110000010;
assign LUT_1[13567] = 32'b00000000000000001101001111111110;
assign LUT_1[13568] = 32'b00000000000000000111001000100101;
assign LUT_1[13569] = 32'b00000000000000000000011010100001;
assign LUT_1[13570] = 32'b00000000000000000010110110110110;
assign LUT_1[13571] = 32'b11111111111111111100001000110010;
assign LUT_1[13572] = 32'b00000000000000001111000001111100;
assign LUT_1[13573] = 32'b00000000000000001000010011111000;
assign LUT_1[13574] = 32'b00000000000000001010110000001101;
assign LUT_1[13575] = 32'b00000000000000000100000010001001;
assign LUT_1[13576] = 32'b00000000000000000110010110011010;
assign LUT_1[13577] = 32'b11111111111111111111101000010110;
assign LUT_1[13578] = 32'b00000000000000000010000100101011;
assign LUT_1[13579] = 32'b11111111111111111011010110100111;
assign LUT_1[13580] = 32'b00000000000000001110001111110001;
assign LUT_1[13581] = 32'b00000000000000000111100001101101;
assign LUT_1[13582] = 32'b00000000000000001001111110000010;
assign LUT_1[13583] = 32'b00000000000000000011001111111110;
assign LUT_1[13584] = 32'b00000000000000001001000100000111;
assign LUT_1[13585] = 32'b00000000000000000010010110000011;
assign LUT_1[13586] = 32'b00000000000000000100110010011000;
assign LUT_1[13587] = 32'b11111111111111111110000100010100;
assign LUT_1[13588] = 32'b00000000000000010000111101011110;
assign LUT_1[13589] = 32'b00000000000000001010001111011010;
assign LUT_1[13590] = 32'b00000000000000001100101011101111;
assign LUT_1[13591] = 32'b00000000000000000101111101101011;
assign LUT_1[13592] = 32'b00000000000000001000010001111100;
assign LUT_1[13593] = 32'b00000000000000000001100011111000;
assign LUT_1[13594] = 32'b00000000000000000100000000001101;
assign LUT_1[13595] = 32'b11111111111111111101010010001001;
assign LUT_1[13596] = 32'b00000000000000010000001011010011;
assign LUT_1[13597] = 32'b00000000000000001001011101001111;
assign LUT_1[13598] = 32'b00000000000000001011111001100100;
assign LUT_1[13599] = 32'b00000000000000000101001011100000;
assign LUT_1[13600] = 32'b00000000000000001000000011100100;
assign LUT_1[13601] = 32'b00000000000000000001010101100000;
assign LUT_1[13602] = 32'b00000000000000000011110001110101;
assign LUT_1[13603] = 32'b11111111111111111101000011110001;
assign LUT_1[13604] = 32'b00000000000000001111111100111011;
assign LUT_1[13605] = 32'b00000000000000001001001110110111;
assign LUT_1[13606] = 32'b00000000000000001011101011001100;
assign LUT_1[13607] = 32'b00000000000000000100111101001000;
assign LUT_1[13608] = 32'b00000000000000000111010001011001;
assign LUT_1[13609] = 32'b00000000000000000000100011010101;
assign LUT_1[13610] = 32'b00000000000000000010111111101010;
assign LUT_1[13611] = 32'b11111111111111111100010001100110;
assign LUT_1[13612] = 32'b00000000000000001111001010110000;
assign LUT_1[13613] = 32'b00000000000000001000011100101100;
assign LUT_1[13614] = 32'b00000000000000001010111001000001;
assign LUT_1[13615] = 32'b00000000000000000100001010111101;
assign LUT_1[13616] = 32'b00000000000000001001111111000110;
assign LUT_1[13617] = 32'b00000000000000000011010001000010;
assign LUT_1[13618] = 32'b00000000000000000101101101010111;
assign LUT_1[13619] = 32'b11111111111111111110111111010011;
assign LUT_1[13620] = 32'b00000000000000010001111000011101;
assign LUT_1[13621] = 32'b00000000000000001011001010011001;
assign LUT_1[13622] = 32'b00000000000000001101100110101110;
assign LUT_1[13623] = 32'b00000000000000000110111000101010;
assign LUT_1[13624] = 32'b00000000000000001001001100111011;
assign LUT_1[13625] = 32'b00000000000000000010011110110111;
assign LUT_1[13626] = 32'b00000000000000000100111011001100;
assign LUT_1[13627] = 32'b11111111111111111110001101001000;
assign LUT_1[13628] = 32'b00000000000000010001000110010010;
assign LUT_1[13629] = 32'b00000000000000001010011000001110;
assign LUT_1[13630] = 32'b00000000000000001100110100100011;
assign LUT_1[13631] = 32'b00000000000000000110000110011111;
assign LUT_1[13632] = 32'b00000000000000001001000110001101;
assign LUT_1[13633] = 32'b00000000000000000010011000001001;
assign LUT_1[13634] = 32'b00000000000000000100110100011110;
assign LUT_1[13635] = 32'b11111111111111111110000110011010;
assign LUT_1[13636] = 32'b00000000000000010000111111100100;
assign LUT_1[13637] = 32'b00000000000000001010010001100000;
assign LUT_1[13638] = 32'b00000000000000001100101101110101;
assign LUT_1[13639] = 32'b00000000000000000101111111110001;
assign LUT_1[13640] = 32'b00000000000000001000010100000010;
assign LUT_1[13641] = 32'b00000000000000000001100101111110;
assign LUT_1[13642] = 32'b00000000000000000100000010010011;
assign LUT_1[13643] = 32'b11111111111111111101010100001111;
assign LUT_1[13644] = 32'b00000000000000010000001101011001;
assign LUT_1[13645] = 32'b00000000000000001001011111010101;
assign LUT_1[13646] = 32'b00000000000000001011111011101010;
assign LUT_1[13647] = 32'b00000000000000000101001101100110;
assign LUT_1[13648] = 32'b00000000000000001011000001101111;
assign LUT_1[13649] = 32'b00000000000000000100010011101011;
assign LUT_1[13650] = 32'b00000000000000000110110000000000;
assign LUT_1[13651] = 32'b00000000000000000000000001111100;
assign LUT_1[13652] = 32'b00000000000000010010111011000110;
assign LUT_1[13653] = 32'b00000000000000001100001101000010;
assign LUT_1[13654] = 32'b00000000000000001110101001010111;
assign LUT_1[13655] = 32'b00000000000000000111111011010011;
assign LUT_1[13656] = 32'b00000000000000001010001111100100;
assign LUT_1[13657] = 32'b00000000000000000011100001100000;
assign LUT_1[13658] = 32'b00000000000000000101111101110101;
assign LUT_1[13659] = 32'b11111111111111111111001111110001;
assign LUT_1[13660] = 32'b00000000000000010010001000111011;
assign LUT_1[13661] = 32'b00000000000000001011011010110111;
assign LUT_1[13662] = 32'b00000000000000001101110111001100;
assign LUT_1[13663] = 32'b00000000000000000111001001001000;
assign LUT_1[13664] = 32'b00000000000000001010000001001100;
assign LUT_1[13665] = 32'b00000000000000000011010011001000;
assign LUT_1[13666] = 32'b00000000000000000101101111011101;
assign LUT_1[13667] = 32'b11111111111111111111000001011001;
assign LUT_1[13668] = 32'b00000000000000010001111010100011;
assign LUT_1[13669] = 32'b00000000000000001011001100011111;
assign LUT_1[13670] = 32'b00000000000000001101101000110100;
assign LUT_1[13671] = 32'b00000000000000000110111010110000;
assign LUT_1[13672] = 32'b00000000000000001001001111000001;
assign LUT_1[13673] = 32'b00000000000000000010100000111101;
assign LUT_1[13674] = 32'b00000000000000000100111101010010;
assign LUT_1[13675] = 32'b11111111111111111110001111001110;
assign LUT_1[13676] = 32'b00000000000000010001001000011000;
assign LUT_1[13677] = 32'b00000000000000001010011010010100;
assign LUT_1[13678] = 32'b00000000000000001100110110101001;
assign LUT_1[13679] = 32'b00000000000000000110001000100101;
assign LUT_1[13680] = 32'b00000000000000001011111100101110;
assign LUT_1[13681] = 32'b00000000000000000101001110101010;
assign LUT_1[13682] = 32'b00000000000000000111101010111111;
assign LUT_1[13683] = 32'b00000000000000000000111100111011;
assign LUT_1[13684] = 32'b00000000000000010011110110000101;
assign LUT_1[13685] = 32'b00000000000000001101001000000001;
assign LUT_1[13686] = 32'b00000000000000001111100100010110;
assign LUT_1[13687] = 32'b00000000000000001000110110010010;
assign LUT_1[13688] = 32'b00000000000000001011001010100011;
assign LUT_1[13689] = 32'b00000000000000000100011100011111;
assign LUT_1[13690] = 32'b00000000000000000110111000110100;
assign LUT_1[13691] = 32'b00000000000000000000001010110000;
assign LUT_1[13692] = 32'b00000000000000010011000011111010;
assign LUT_1[13693] = 32'b00000000000000001100010101110110;
assign LUT_1[13694] = 32'b00000000000000001110110010001011;
assign LUT_1[13695] = 32'b00000000000000001000000100000111;
assign LUT_1[13696] = 32'b00000000000000001010001000101000;
assign LUT_1[13697] = 32'b00000000000000000011011010100100;
assign LUT_1[13698] = 32'b00000000000000000101110110111001;
assign LUT_1[13699] = 32'b11111111111111111111001000110101;
assign LUT_1[13700] = 32'b00000000000000010010000001111111;
assign LUT_1[13701] = 32'b00000000000000001011010011111011;
assign LUT_1[13702] = 32'b00000000000000001101110000010000;
assign LUT_1[13703] = 32'b00000000000000000111000010001100;
assign LUT_1[13704] = 32'b00000000000000001001010110011101;
assign LUT_1[13705] = 32'b00000000000000000010101000011001;
assign LUT_1[13706] = 32'b00000000000000000101000100101110;
assign LUT_1[13707] = 32'b11111111111111111110010110101010;
assign LUT_1[13708] = 32'b00000000000000010001001111110100;
assign LUT_1[13709] = 32'b00000000000000001010100001110000;
assign LUT_1[13710] = 32'b00000000000000001100111110000101;
assign LUT_1[13711] = 32'b00000000000000000110010000000001;
assign LUT_1[13712] = 32'b00000000000000001100000100001010;
assign LUT_1[13713] = 32'b00000000000000000101010110000110;
assign LUT_1[13714] = 32'b00000000000000000111110010011011;
assign LUT_1[13715] = 32'b00000000000000000001000100010111;
assign LUT_1[13716] = 32'b00000000000000010011111101100001;
assign LUT_1[13717] = 32'b00000000000000001101001111011101;
assign LUT_1[13718] = 32'b00000000000000001111101011110010;
assign LUT_1[13719] = 32'b00000000000000001000111101101110;
assign LUT_1[13720] = 32'b00000000000000001011010001111111;
assign LUT_1[13721] = 32'b00000000000000000100100011111011;
assign LUT_1[13722] = 32'b00000000000000000111000000010000;
assign LUT_1[13723] = 32'b00000000000000000000010010001100;
assign LUT_1[13724] = 32'b00000000000000010011001011010110;
assign LUT_1[13725] = 32'b00000000000000001100011101010010;
assign LUT_1[13726] = 32'b00000000000000001110111001100111;
assign LUT_1[13727] = 32'b00000000000000001000001011100011;
assign LUT_1[13728] = 32'b00000000000000001011000011100111;
assign LUT_1[13729] = 32'b00000000000000000100010101100011;
assign LUT_1[13730] = 32'b00000000000000000110110001111000;
assign LUT_1[13731] = 32'b00000000000000000000000011110100;
assign LUT_1[13732] = 32'b00000000000000010010111100111110;
assign LUT_1[13733] = 32'b00000000000000001100001110111010;
assign LUT_1[13734] = 32'b00000000000000001110101011001111;
assign LUT_1[13735] = 32'b00000000000000000111111101001011;
assign LUT_1[13736] = 32'b00000000000000001010010001011100;
assign LUT_1[13737] = 32'b00000000000000000011100011011000;
assign LUT_1[13738] = 32'b00000000000000000101111111101101;
assign LUT_1[13739] = 32'b11111111111111111111010001101001;
assign LUT_1[13740] = 32'b00000000000000010010001010110011;
assign LUT_1[13741] = 32'b00000000000000001011011100101111;
assign LUT_1[13742] = 32'b00000000000000001101111001000100;
assign LUT_1[13743] = 32'b00000000000000000111001011000000;
assign LUT_1[13744] = 32'b00000000000000001100111111001001;
assign LUT_1[13745] = 32'b00000000000000000110010001000101;
assign LUT_1[13746] = 32'b00000000000000001000101101011010;
assign LUT_1[13747] = 32'b00000000000000000001111111010110;
assign LUT_1[13748] = 32'b00000000000000010100111000100000;
assign LUT_1[13749] = 32'b00000000000000001110001010011100;
assign LUT_1[13750] = 32'b00000000000000010000100110110001;
assign LUT_1[13751] = 32'b00000000000000001001111000101101;
assign LUT_1[13752] = 32'b00000000000000001100001100111110;
assign LUT_1[13753] = 32'b00000000000000000101011110111010;
assign LUT_1[13754] = 32'b00000000000000000111111011001111;
assign LUT_1[13755] = 32'b00000000000000000001001101001011;
assign LUT_1[13756] = 32'b00000000000000010100000110010101;
assign LUT_1[13757] = 32'b00000000000000001101011000010001;
assign LUT_1[13758] = 32'b00000000000000001111110100100110;
assign LUT_1[13759] = 32'b00000000000000001001000110100010;
assign LUT_1[13760] = 32'b00000000000000001100000110010000;
assign LUT_1[13761] = 32'b00000000000000000101011000001100;
assign LUT_1[13762] = 32'b00000000000000000111110100100001;
assign LUT_1[13763] = 32'b00000000000000000001000110011101;
assign LUT_1[13764] = 32'b00000000000000010011111111100111;
assign LUT_1[13765] = 32'b00000000000000001101010001100011;
assign LUT_1[13766] = 32'b00000000000000001111101101111000;
assign LUT_1[13767] = 32'b00000000000000001000111111110100;
assign LUT_1[13768] = 32'b00000000000000001011010100000101;
assign LUT_1[13769] = 32'b00000000000000000100100110000001;
assign LUT_1[13770] = 32'b00000000000000000111000010010110;
assign LUT_1[13771] = 32'b00000000000000000000010100010010;
assign LUT_1[13772] = 32'b00000000000000010011001101011100;
assign LUT_1[13773] = 32'b00000000000000001100011111011000;
assign LUT_1[13774] = 32'b00000000000000001110111011101101;
assign LUT_1[13775] = 32'b00000000000000001000001101101001;
assign LUT_1[13776] = 32'b00000000000000001110000001110010;
assign LUT_1[13777] = 32'b00000000000000000111010011101110;
assign LUT_1[13778] = 32'b00000000000000001001110000000011;
assign LUT_1[13779] = 32'b00000000000000000011000001111111;
assign LUT_1[13780] = 32'b00000000000000010101111011001001;
assign LUT_1[13781] = 32'b00000000000000001111001101000101;
assign LUT_1[13782] = 32'b00000000000000010001101001011010;
assign LUT_1[13783] = 32'b00000000000000001010111011010110;
assign LUT_1[13784] = 32'b00000000000000001101001111100111;
assign LUT_1[13785] = 32'b00000000000000000110100001100011;
assign LUT_1[13786] = 32'b00000000000000001000111101111000;
assign LUT_1[13787] = 32'b00000000000000000010001111110100;
assign LUT_1[13788] = 32'b00000000000000010101001000111110;
assign LUT_1[13789] = 32'b00000000000000001110011010111010;
assign LUT_1[13790] = 32'b00000000000000010000110111001111;
assign LUT_1[13791] = 32'b00000000000000001010001001001011;
assign LUT_1[13792] = 32'b00000000000000001101000001001111;
assign LUT_1[13793] = 32'b00000000000000000110010011001011;
assign LUT_1[13794] = 32'b00000000000000001000101111100000;
assign LUT_1[13795] = 32'b00000000000000000010000001011100;
assign LUT_1[13796] = 32'b00000000000000010100111010100110;
assign LUT_1[13797] = 32'b00000000000000001110001100100010;
assign LUT_1[13798] = 32'b00000000000000010000101000110111;
assign LUT_1[13799] = 32'b00000000000000001001111010110011;
assign LUT_1[13800] = 32'b00000000000000001100001111000100;
assign LUT_1[13801] = 32'b00000000000000000101100001000000;
assign LUT_1[13802] = 32'b00000000000000000111111101010101;
assign LUT_1[13803] = 32'b00000000000000000001001111010001;
assign LUT_1[13804] = 32'b00000000000000010100001000011011;
assign LUT_1[13805] = 32'b00000000000000001101011010010111;
assign LUT_1[13806] = 32'b00000000000000001111110110101100;
assign LUT_1[13807] = 32'b00000000000000001001001000101000;
assign LUT_1[13808] = 32'b00000000000000001110111100110001;
assign LUT_1[13809] = 32'b00000000000000001000001110101101;
assign LUT_1[13810] = 32'b00000000000000001010101011000010;
assign LUT_1[13811] = 32'b00000000000000000011111100111110;
assign LUT_1[13812] = 32'b00000000000000010110110110001000;
assign LUT_1[13813] = 32'b00000000000000010000001000000100;
assign LUT_1[13814] = 32'b00000000000000010010100100011001;
assign LUT_1[13815] = 32'b00000000000000001011110110010101;
assign LUT_1[13816] = 32'b00000000000000001110001010100110;
assign LUT_1[13817] = 32'b00000000000000000111011100100010;
assign LUT_1[13818] = 32'b00000000000000001001111000110111;
assign LUT_1[13819] = 32'b00000000000000000011001010110011;
assign LUT_1[13820] = 32'b00000000000000010110000011111101;
assign LUT_1[13821] = 32'b00000000000000001111010101111001;
assign LUT_1[13822] = 32'b00000000000000010001110010001110;
assign LUT_1[13823] = 32'b00000000000000001011000100001010;
assign LUT_1[13824] = 32'b00000000000000000011000010110110;
assign LUT_1[13825] = 32'b11111111111111111100010100110010;
assign LUT_1[13826] = 32'b11111111111111111110110001000111;
assign LUT_1[13827] = 32'b11111111111111111000000011000011;
assign LUT_1[13828] = 32'b00000000000000001010111100001101;
assign LUT_1[13829] = 32'b00000000000000000100001110001001;
assign LUT_1[13830] = 32'b00000000000000000110101010011110;
assign LUT_1[13831] = 32'b11111111111111111111111100011010;
assign LUT_1[13832] = 32'b00000000000000000010010000101011;
assign LUT_1[13833] = 32'b11111111111111111011100010100111;
assign LUT_1[13834] = 32'b11111111111111111101111110111100;
assign LUT_1[13835] = 32'b11111111111111110111010000111000;
assign LUT_1[13836] = 32'b00000000000000001010001010000010;
assign LUT_1[13837] = 32'b00000000000000000011011011111110;
assign LUT_1[13838] = 32'b00000000000000000101111000010011;
assign LUT_1[13839] = 32'b11111111111111111111001010001111;
assign LUT_1[13840] = 32'b00000000000000000100111110011000;
assign LUT_1[13841] = 32'b11111111111111111110010000010100;
assign LUT_1[13842] = 32'b00000000000000000000101100101001;
assign LUT_1[13843] = 32'b11111111111111111001111110100101;
assign LUT_1[13844] = 32'b00000000000000001100110111101111;
assign LUT_1[13845] = 32'b00000000000000000110001001101011;
assign LUT_1[13846] = 32'b00000000000000001000100110000000;
assign LUT_1[13847] = 32'b00000000000000000001110111111100;
assign LUT_1[13848] = 32'b00000000000000000100001100001101;
assign LUT_1[13849] = 32'b11111111111111111101011110001001;
assign LUT_1[13850] = 32'b11111111111111111111111010011110;
assign LUT_1[13851] = 32'b11111111111111111001001100011010;
assign LUT_1[13852] = 32'b00000000000000001100000101100100;
assign LUT_1[13853] = 32'b00000000000000000101010111100000;
assign LUT_1[13854] = 32'b00000000000000000111110011110101;
assign LUT_1[13855] = 32'b00000000000000000001000101110001;
assign LUT_1[13856] = 32'b00000000000000000011111101110101;
assign LUT_1[13857] = 32'b11111111111111111101001111110001;
assign LUT_1[13858] = 32'b11111111111111111111101100000110;
assign LUT_1[13859] = 32'b11111111111111111000111110000010;
assign LUT_1[13860] = 32'b00000000000000001011110111001100;
assign LUT_1[13861] = 32'b00000000000000000101001001001000;
assign LUT_1[13862] = 32'b00000000000000000111100101011101;
assign LUT_1[13863] = 32'b00000000000000000000110111011001;
assign LUT_1[13864] = 32'b00000000000000000011001011101010;
assign LUT_1[13865] = 32'b11111111111111111100011101100110;
assign LUT_1[13866] = 32'b11111111111111111110111001111011;
assign LUT_1[13867] = 32'b11111111111111111000001011110111;
assign LUT_1[13868] = 32'b00000000000000001011000101000001;
assign LUT_1[13869] = 32'b00000000000000000100010110111101;
assign LUT_1[13870] = 32'b00000000000000000110110011010010;
assign LUT_1[13871] = 32'b00000000000000000000000101001110;
assign LUT_1[13872] = 32'b00000000000000000101111001010111;
assign LUT_1[13873] = 32'b11111111111111111111001011010011;
assign LUT_1[13874] = 32'b00000000000000000001100111101000;
assign LUT_1[13875] = 32'b11111111111111111010111001100100;
assign LUT_1[13876] = 32'b00000000000000001101110010101110;
assign LUT_1[13877] = 32'b00000000000000000111000100101010;
assign LUT_1[13878] = 32'b00000000000000001001100000111111;
assign LUT_1[13879] = 32'b00000000000000000010110010111011;
assign LUT_1[13880] = 32'b00000000000000000101000111001100;
assign LUT_1[13881] = 32'b11111111111111111110011001001000;
assign LUT_1[13882] = 32'b00000000000000000000110101011101;
assign LUT_1[13883] = 32'b11111111111111111010000111011001;
assign LUT_1[13884] = 32'b00000000000000001101000000100011;
assign LUT_1[13885] = 32'b00000000000000000110010010011111;
assign LUT_1[13886] = 32'b00000000000000001000101110110100;
assign LUT_1[13887] = 32'b00000000000000000010000000110000;
assign LUT_1[13888] = 32'b00000000000000000101000000011110;
assign LUT_1[13889] = 32'b11111111111111111110010010011010;
assign LUT_1[13890] = 32'b00000000000000000000101110101111;
assign LUT_1[13891] = 32'b11111111111111111010000000101011;
assign LUT_1[13892] = 32'b00000000000000001100111001110101;
assign LUT_1[13893] = 32'b00000000000000000110001011110001;
assign LUT_1[13894] = 32'b00000000000000001000101000000110;
assign LUT_1[13895] = 32'b00000000000000000001111010000010;
assign LUT_1[13896] = 32'b00000000000000000100001110010011;
assign LUT_1[13897] = 32'b11111111111111111101100000001111;
assign LUT_1[13898] = 32'b11111111111111111111111100100100;
assign LUT_1[13899] = 32'b11111111111111111001001110100000;
assign LUT_1[13900] = 32'b00000000000000001100000111101010;
assign LUT_1[13901] = 32'b00000000000000000101011001100110;
assign LUT_1[13902] = 32'b00000000000000000111110101111011;
assign LUT_1[13903] = 32'b00000000000000000001000111110111;
assign LUT_1[13904] = 32'b00000000000000000110111100000000;
assign LUT_1[13905] = 32'b00000000000000000000001101111100;
assign LUT_1[13906] = 32'b00000000000000000010101010010001;
assign LUT_1[13907] = 32'b11111111111111111011111100001101;
assign LUT_1[13908] = 32'b00000000000000001110110101010111;
assign LUT_1[13909] = 32'b00000000000000001000000111010011;
assign LUT_1[13910] = 32'b00000000000000001010100011101000;
assign LUT_1[13911] = 32'b00000000000000000011110101100100;
assign LUT_1[13912] = 32'b00000000000000000110001001110101;
assign LUT_1[13913] = 32'b11111111111111111111011011110001;
assign LUT_1[13914] = 32'b00000000000000000001111000000110;
assign LUT_1[13915] = 32'b11111111111111111011001010000010;
assign LUT_1[13916] = 32'b00000000000000001110000011001100;
assign LUT_1[13917] = 32'b00000000000000000111010101001000;
assign LUT_1[13918] = 32'b00000000000000001001110001011101;
assign LUT_1[13919] = 32'b00000000000000000011000011011001;
assign LUT_1[13920] = 32'b00000000000000000101111011011101;
assign LUT_1[13921] = 32'b11111111111111111111001101011001;
assign LUT_1[13922] = 32'b00000000000000000001101001101110;
assign LUT_1[13923] = 32'b11111111111111111010111011101010;
assign LUT_1[13924] = 32'b00000000000000001101110100110100;
assign LUT_1[13925] = 32'b00000000000000000111000110110000;
assign LUT_1[13926] = 32'b00000000000000001001100011000101;
assign LUT_1[13927] = 32'b00000000000000000010110101000001;
assign LUT_1[13928] = 32'b00000000000000000101001001010010;
assign LUT_1[13929] = 32'b11111111111111111110011011001110;
assign LUT_1[13930] = 32'b00000000000000000000110111100011;
assign LUT_1[13931] = 32'b11111111111111111010001001011111;
assign LUT_1[13932] = 32'b00000000000000001101000010101001;
assign LUT_1[13933] = 32'b00000000000000000110010100100101;
assign LUT_1[13934] = 32'b00000000000000001000110000111010;
assign LUT_1[13935] = 32'b00000000000000000010000010110110;
assign LUT_1[13936] = 32'b00000000000000000111110110111111;
assign LUT_1[13937] = 32'b00000000000000000001001000111011;
assign LUT_1[13938] = 32'b00000000000000000011100101010000;
assign LUT_1[13939] = 32'b11111111111111111100110111001100;
assign LUT_1[13940] = 32'b00000000000000001111110000010110;
assign LUT_1[13941] = 32'b00000000000000001001000010010010;
assign LUT_1[13942] = 32'b00000000000000001011011110100111;
assign LUT_1[13943] = 32'b00000000000000000100110000100011;
assign LUT_1[13944] = 32'b00000000000000000111000100110100;
assign LUT_1[13945] = 32'b00000000000000000000010110110000;
assign LUT_1[13946] = 32'b00000000000000000010110011000101;
assign LUT_1[13947] = 32'b11111111111111111100000101000001;
assign LUT_1[13948] = 32'b00000000000000001110111110001011;
assign LUT_1[13949] = 32'b00000000000000001000010000000111;
assign LUT_1[13950] = 32'b00000000000000001010101100011100;
assign LUT_1[13951] = 32'b00000000000000000011111110011000;
assign LUT_1[13952] = 32'b00000000000000000110000010111001;
assign LUT_1[13953] = 32'b11111111111111111111010100110101;
assign LUT_1[13954] = 32'b00000000000000000001110001001010;
assign LUT_1[13955] = 32'b11111111111111111011000011000110;
assign LUT_1[13956] = 32'b00000000000000001101111100010000;
assign LUT_1[13957] = 32'b00000000000000000111001110001100;
assign LUT_1[13958] = 32'b00000000000000001001101010100001;
assign LUT_1[13959] = 32'b00000000000000000010111100011101;
assign LUT_1[13960] = 32'b00000000000000000101010000101110;
assign LUT_1[13961] = 32'b11111111111111111110100010101010;
assign LUT_1[13962] = 32'b00000000000000000000111110111111;
assign LUT_1[13963] = 32'b11111111111111111010010000111011;
assign LUT_1[13964] = 32'b00000000000000001101001010000101;
assign LUT_1[13965] = 32'b00000000000000000110011100000001;
assign LUT_1[13966] = 32'b00000000000000001000111000010110;
assign LUT_1[13967] = 32'b00000000000000000010001010010010;
assign LUT_1[13968] = 32'b00000000000000000111111110011011;
assign LUT_1[13969] = 32'b00000000000000000001010000010111;
assign LUT_1[13970] = 32'b00000000000000000011101100101100;
assign LUT_1[13971] = 32'b11111111111111111100111110101000;
assign LUT_1[13972] = 32'b00000000000000001111110111110010;
assign LUT_1[13973] = 32'b00000000000000001001001001101110;
assign LUT_1[13974] = 32'b00000000000000001011100110000011;
assign LUT_1[13975] = 32'b00000000000000000100110111111111;
assign LUT_1[13976] = 32'b00000000000000000111001100010000;
assign LUT_1[13977] = 32'b00000000000000000000011110001100;
assign LUT_1[13978] = 32'b00000000000000000010111010100001;
assign LUT_1[13979] = 32'b11111111111111111100001100011101;
assign LUT_1[13980] = 32'b00000000000000001111000101100111;
assign LUT_1[13981] = 32'b00000000000000001000010111100011;
assign LUT_1[13982] = 32'b00000000000000001010110011111000;
assign LUT_1[13983] = 32'b00000000000000000100000101110100;
assign LUT_1[13984] = 32'b00000000000000000110111101111000;
assign LUT_1[13985] = 32'b00000000000000000000001111110100;
assign LUT_1[13986] = 32'b00000000000000000010101100001001;
assign LUT_1[13987] = 32'b11111111111111111011111110000101;
assign LUT_1[13988] = 32'b00000000000000001110110111001111;
assign LUT_1[13989] = 32'b00000000000000001000001001001011;
assign LUT_1[13990] = 32'b00000000000000001010100101100000;
assign LUT_1[13991] = 32'b00000000000000000011110111011100;
assign LUT_1[13992] = 32'b00000000000000000110001011101101;
assign LUT_1[13993] = 32'b11111111111111111111011101101001;
assign LUT_1[13994] = 32'b00000000000000000001111001111110;
assign LUT_1[13995] = 32'b11111111111111111011001011111010;
assign LUT_1[13996] = 32'b00000000000000001110000101000100;
assign LUT_1[13997] = 32'b00000000000000000111010111000000;
assign LUT_1[13998] = 32'b00000000000000001001110011010101;
assign LUT_1[13999] = 32'b00000000000000000011000101010001;
assign LUT_1[14000] = 32'b00000000000000001000111001011010;
assign LUT_1[14001] = 32'b00000000000000000010001011010110;
assign LUT_1[14002] = 32'b00000000000000000100100111101011;
assign LUT_1[14003] = 32'b11111111111111111101111001100111;
assign LUT_1[14004] = 32'b00000000000000010000110010110001;
assign LUT_1[14005] = 32'b00000000000000001010000100101101;
assign LUT_1[14006] = 32'b00000000000000001100100001000010;
assign LUT_1[14007] = 32'b00000000000000000101110010111110;
assign LUT_1[14008] = 32'b00000000000000001000000111001111;
assign LUT_1[14009] = 32'b00000000000000000001011001001011;
assign LUT_1[14010] = 32'b00000000000000000011110101100000;
assign LUT_1[14011] = 32'b11111111111111111101000111011100;
assign LUT_1[14012] = 32'b00000000000000010000000000100110;
assign LUT_1[14013] = 32'b00000000000000001001010010100010;
assign LUT_1[14014] = 32'b00000000000000001011101110110111;
assign LUT_1[14015] = 32'b00000000000000000101000000110011;
assign LUT_1[14016] = 32'b00000000000000001000000000100001;
assign LUT_1[14017] = 32'b00000000000000000001010010011101;
assign LUT_1[14018] = 32'b00000000000000000011101110110010;
assign LUT_1[14019] = 32'b11111111111111111101000000101110;
assign LUT_1[14020] = 32'b00000000000000001111111001111000;
assign LUT_1[14021] = 32'b00000000000000001001001011110100;
assign LUT_1[14022] = 32'b00000000000000001011101000001001;
assign LUT_1[14023] = 32'b00000000000000000100111010000101;
assign LUT_1[14024] = 32'b00000000000000000111001110010110;
assign LUT_1[14025] = 32'b00000000000000000000100000010010;
assign LUT_1[14026] = 32'b00000000000000000010111100100111;
assign LUT_1[14027] = 32'b11111111111111111100001110100011;
assign LUT_1[14028] = 32'b00000000000000001111000111101101;
assign LUT_1[14029] = 32'b00000000000000001000011001101001;
assign LUT_1[14030] = 32'b00000000000000001010110101111110;
assign LUT_1[14031] = 32'b00000000000000000100000111111010;
assign LUT_1[14032] = 32'b00000000000000001001111100000011;
assign LUT_1[14033] = 32'b00000000000000000011001101111111;
assign LUT_1[14034] = 32'b00000000000000000101101010010100;
assign LUT_1[14035] = 32'b11111111111111111110111100010000;
assign LUT_1[14036] = 32'b00000000000000010001110101011010;
assign LUT_1[14037] = 32'b00000000000000001011000111010110;
assign LUT_1[14038] = 32'b00000000000000001101100011101011;
assign LUT_1[14039] = 32'b00000000000000000110110101100111;
assign LUT_1[14040] = 32'b00000000000000001001001001111000;
assign LUT_1[14041] = 32'b00000000000000000010011011110100;
assign LUT_1[14042] = 32'b00000000000000000100111000001001;
assign LUT_1[14043] = 32'b11111111111111111110001010000101;
assign LUT_1[14044] = 32'b00000000000000010001000011001111;
assign LUT_1[14045] = 32'b00000000000000001010010101001011;
assign LUT_1[14046] = 32'b00000000000000001100110001100000;
assign LUT_1[14047] = 32'b00000000000000000110000011011100;
assign LUT_1[14048] = 32'b00000000000000001000111011100000;
assign LUT_1[14049] = 32'b00000000000000000010001101011100;
assign LUT_1[14050] = 32'b00000000000000000100101001110001;
assign LUT_1[14051] = 32'b11111111111111111101111011101101;
assign LUT_1[14052] = 32'b00000000000000010000110100110111;
assign LUT_1[14053] = 32'b00000000000000001010000110110011;
assign LUT_1[14054] = 32'b00000000000000001100100011001000;
assign LUT_1[14055] = 32'b00000000000000000101110101000100;
assign LUT_1[14056] = 32'b00000000000000001000001001010101;
assign LUT_1[14057] = 32'b00000000000000000001011011010001;
assign LUT_1[14058] = 32'b00000000000000000011110111100110;
assign LUT_1[14059] = 32'b11111111111111111101001001100010;
assign LUT_1[14060] = 32'b00000000000000010000000010101100;
assign LUT_1[14061] = 32'b00000000000000001001010100101000;
assign LUT_1[14062] = 32'b00000000000000001011110000111101;
assign LUT_1[14063] = 32'b00000000000000000101000010111001;
assign LUT_1[14064] = 32'b00000000000000001010110111000010;
assign LUT_1[14065] = 32'b00000000000000000100001000111110;
assign LUT_1[14066] = 32'b00000000000000000110100101010011;
assign LUT_1[14067] = 32'b11111111111111111111110111001111;
assign LUT_1[14068] = 32'b00000000000000010010110000011001;
assign LUT_1[14069] = 32'b00000000000000001100000010010101;
assign LUT_1[14070] = 32'b00000000000000001110011110101010;
assign LUT_1[14071] = 32'b00000000000000000111110000100110;
assign LUT_1[14072] = 32'b00000000000000001010000100110111;
assign LUT_1[14073] = 32'b00000000000000000011010110110011;
assign LUT_1[14074] = 32'b00000000000000000101110011001000;
assign LUT_1[14075] = 32'b11111111111111111111000101000100;
assign LUT_1[14076] = 32'b00000000000000010001111110001110;
assign LUT_1[14077] = 32'b00000000000000001011010000001010;
assign LUT_1[14078] = 32'b00000000000000001101101100011111;
assign LUT_1[14079] = 32'b00000000000000000110111110011011;
assign LUT_1[14080] = 32'b00000000000000000000110111000010;
assign LUT_1[14081] = 32'b11111111111111111010001000111110;
assign LUT_1[14082] = 32'b11111111111111111100100101010011;
assign LUT_1[14083] = 32'b11111111111111110101110111001111;
assign LUT_1[14084] = 32'b00000000000000001000110000011001;
assign LUT_1[14085] = 32'b00000000000000000010000010010101;
assign LUT_1[14086] = 32'b00000000000000000100011110101010;
assign LUT_1[14087] = 32'b11111111111111111101110000100110;
assign LUT_1[14088] = 32'b00000000000000000000000100110111;
assign LUT_1[14089] = 32'b11111111111111111001010110110011;
assign LUT_1[14090] = 32'b11111111111111111011110011001000;
assign LUT_1[14091] = 32'b11111111111111110101000101000100;
assign LUT_1[14092] = 32'b00000000000000000111111110001110;
assign LUT_1[14093] = 32'b00000000000000000001010000001010;
assign LUT_1[14094] = 32'b00000000000000000011101100011111;
assign LUT_1[14095] = 32'b11111111111111111100111110011011;
assign LUT_1[14096] = 32'b00000000000000000010110010100100;
assign LUT_1[14097] = 32'b11111111111111111100000100100000;
assign LUT_1[14098] = 32'b11111111111111111110100000110101;
assign LUT_1[14099] = 32'b11111111111111110111110010110001;
assign LUT_1[14100] = 32'b00000000000000001010101011111011;
assign LUT_1[14101] = 32'b00000000000000000011111101110111;
assign LUT_1[14102] = 32'b00000000000000000110011010001100;
assign LUT_1[14103] = 32'b11111111111111111111101100001000;
assign LUT_1[14104] = 32'b00000000000000000010000000011001;
assign LUT_1[14105] = 32'b11111111111111111011010010010101;
assign LUT_1[14106] = 32'b11111111111111111101101110101010;
assign LUT_1[14107] = 32'b11111111111111110111000000100110;
assign LUT_1[14108] = 32'b00000000000000001001111001110000;
assign LUT_1[14109] = 32'b00000000000000000011001011101100;
assign LUT_1[14110] = 32'b00000000000000000101101000000001;
assign LUT_1[14111] = 32'b11111111111111111110111001111101;
assign LUT_1[14112] = 32'b00000000000000000001110010000001;
assign LUT_1[14113] = 32'b11111111111111111011000011111101;
assign LUT_1[14114] = 32'b11111111111111111101100000010010;
assign LUT_1[14115] = 32'b11111111111111110110110010001110;
assign LUT_1[14116] = 32'b00000000000000001001101011011000;
assign LUT_1[14117] = 32'b00000000000000000010111101010100;
assign LUT_1[14118] = 32'b00000000000000000101011001101001;
assign LUT_1[14119] = 32'b11111111111111111110101011100101;
assign LUT_1[14120] = 32'b00000000000000000000111111110110;
assign LUT_1[14121] = 32'b11111111111111111010010001110010;
assign LUT_1[14122] = 32'b11111111111111111100101110000111;
assign LUT_1[14123] = 32'b11111111111111110110000000000011;
assign LUT_1[14124] = 32'b00000000000000001000111001001101;
assign LUT_1[14125] = 32'b00000000000000000010001011001001;
assign LUT_1[14126] = 32'b00000000000000000100100111011110;
assign LUT_1[14127] = 32'b11111111111111111101111001011010;
assign LUT_1[14128] = 32'b00000000000000000011101101100011;
assign LUT_1[14129] = 32'b11111111111111111100111111011111;
assign LUT_1[14130] = 32'b11111111111111111111011011110100;
assign LUT_1[14131] = 32'b11111111111111111000101101110000;
assign LUT_1[14132] = 32'b00000000000000001011100110111010;
assign LUT_1[14133] = 32'b00000000000000000100111000110110;
assign LUT_1[14134] = 32'b00000000000000000111010101001011;
assign LUT_1[14135] = 32'b00000000000000000000100111000111;
assign LUT_1[14136] = 32'b00000000000000000010111011011000;
assign LUT_1[14137] = 32'b11111111111111111100001101010100;
assign LUT_1[14138] = 32'b11111111111111111110101001101001;
assign LUT_1[14139] = 32'b11111111111111110111111011100101;
assign LUT_1[14140] = 32'b00000000000000001010110100101111;
assign LUT_1[14141] = 32'b00000000000000000100000110101011;
assign LUT_1[14142] = 32'b00000000000000000110100011000000;
assign LUT_1[14143] = 32'b11111111111111111111110100111100;
assign LUT_1[14144] = 32'b00000000000000000010110100101010;
assign LUT_1[14145] = 32'b11111111111111111100000110100110;
assign LUT_1[14146] = 32'b11111111111111111110100010111011;
assign LUT_1[14147] = 32'b11111111111111110111110100110111;
assign LUT_1[14148] = 32'b00000000000000001010101110000001;
assign LUT_1[14149] = 32'b00000000000000000011111111111101;
assign LUT_1[14150] = 32'b00000000000000000110011100010010;
assign LUT_1[14151] = 32'b11111111111111111111101110001110;
assign LUT_1[14152] = 32'b00000000000000000010000010011111;
assign LUT_1[14153] = 32'b11111111111111111011010100011011;
assign LUT_1[14154] = 32'b11111111111111111101110000110000;
assign LUT_1[14155] = 32'b11111111111111110111000010101100;
assign LUT_1[14156] = 32'b00000000000000001001111011110110;
assign LUT_1[14157] = 32'b00000000000000000011001101110010;
assign LUT_1[14158] = 32'b00000000000000000101101010000111;
assign LUT_1[14159] = 32'b11111111111111111110111100000011;
assign LUT_1[14160] = 32'b00000000000000000100110000001100;
assign LUT_1[14161] = 32'b11111111111111111110000010001000;
assign LUT_1[14162] = 32'b00000000000000000000011110011101;
assign LUT_1[14163] = 32'b11111111111111111001110000011001;
assign LUT_1[14164] = 32'b00000000000000001100101001100011;
assign LUT_1[14165] = 32'b00000000000000000101111011011111;
assign LUT_1[14166] = 32'b00000000000000001000010111110100;
assign LUT_1[14167] = 32'b00000000000000000001101001110000;
assign LUT_1[14168] = 32'b00000000000000000011111110000001;
assign LUT_1[14169] = 32'b11111111111111111101001111111101;
assign LUT_1[14170] = 32'b11111111111111111111101100010010;
assign LUT_1[14171] = 32'b11111111111111111000111110001110;
assign LUT_1[14172] = 32'b00000000000000001011110111011000;
assign LUT_1[14173] = 32'b00000000000000000101001001010100;
assign LUT_1[14174] = 32'b00000000000000000111100101101001;
assign LUT_1[14175] = 32'b00000000000000000000110111100101;
assign LUT_1[14176] = 32'b00000000000000000011101111101001;
assign LUT_1[14177] = 32'b11111111111111111101000001100101;
assign LUT_1[14178] = 32'b11111111111111111111011101111010;
assign LUT_1[14179] = 32'b11111111111111111000101111110110;
assign LUT_1[14180] = 32'b00000000000000001011101001000000;
assign LUT_1[14181] = 32'b00000000000000000100111010111100;
assign LUT_1[14182] = 32'b00000000000000000111010111010001;
assign LUT_1[14183] = 32'b00000000000000000000101001001101;
assign LUT_1[14184] = 32'b00000000000000000010111101011110;
assign LUT_1[14185] = 32'b11111111111111111100001111011010;
assign LUT_1[14186] = 32'b11111111111111111110101011101111;
assign LUT_1[14187] = 32'b11111111111111110111111101101011;
assign LUT_1[14188] = 32'b00000000000000001010110110110101;
assign LUT_1[14189] = 32'b00000000000000000100001000110001;
assign LUT_1[14190] = 32'b00000000000000000110100101000110;
assign LUT_1[14191] = 32'b11111111111111111111110111000010;
assign LUT_1[14192] = 32'b00000000000000000101101011001011;
assign LUT_1[14193] = 32'b11111111111111111110111101000111;
assign LUT_1[14194] = 32'b00000000000000000001011001011100;
assign LUT_1[14195] = 32'b11111111111111111010101011011000;
assign LUT_1[14196] = 32'b00000000000000001101100100100010;
assign LUT_1[14197] = 32'b00000000000000000110110110011110;
assign LUT_1[14198] = 32'b00000000000000001001010010110011;
assign LUT_1[14199] = 32'b00000000000000000010100100101111;
assign LUT_1[14200] = 32'b00000000000000000100111001000000;
assign LUT_1[14201] = 32'b11111111111111111110001010111100;
assign LUT_1[14202] = 32'b00000000000000000000100111010001;
assign LUT_1[14203] = 32'b11111111111111111001111001001101;
assign LUT_1[14204] = 32'b00000000000000001100110010010111;
assign LUT_1[14205] = 32'b00000000000000000110000100010011;
assign LUT_1[14206] = 32'b00000000000000001000100000101000;
assign LUT_1[14207] = 32'b00000000000000000001110010100100;
assign LUT_1[14208] = 32'b00000000000000000011110111000101;
assign LUT_1[14209] = 32'b11111111111111111101001001000001;
assign LUT_1[14210] = 32'b11111111111111111111100101010110;
assign LUT_1[14211] = 32'b11111111111111111000110111010010;
assign LUT_1[14212] = 32'b00000000000000001011110000011100;
assign LUT_1[14213] = 32'b00000000000000000101000010011000;
assign LUT_1[14214] = 32'b00000000000000000111011110101101;
assign LUT_1[14215] = 32'b00000000000000000000110000101001;
assign LUT_1[14216] = 32'b00000000000000000011000100111010;
assign LUT_1[14217] = 32'b11111111111111111100010110110110;
assign LUT_1[14218] = 32'b11111111111111111110110011001011;
assign LUT_1[14219] = 32'b11111111111111111000000101000111;
assign LUT_1[14220] = 32'b00000000000000001010111110010001;
assign LUT_1[14221] = 32'b00000000000000000100010000001101;
assign LUT_1[14222] = 32'b00000000000000000110101100100010;
assign LUT_1[14223] = 32'b11111111111111111111111110011110;
assign LUT_1[14224] = 32'b00000000000000000101110010100111;
assign LUT_1[14225] = 32'b11111111111111111111000100100011;
assign LUT_1[14226] = 32'b00000000000000000001100000111000;
assign LUT_1[14227] = 32'b11111111111111111010110010110100;
assign LUT_1[14228] = 32'b00000000000000001101101011111110;
assign LUT_1[14229] = 32'b00000000000000000110111101111010;
assign LUT_1[14230] = 32'b00000000000000001001011010001111;
assign LUT_1[14231] = 32'b00000000000000000010101100001011;
assign LUT_1[14232] = 32'b00000000000000000101000000011100;
assign LUT_1[14233] = 32'b11111111111111111110010010011000;
assign LUT_1[14234] = 32'b00000000000000000000101110101101;
assign LUT_1[14235] = 32'b11111111111111111010000000101001;
assign LUT_1[14236] = 32'b00000000000000001100111001110011;
assign LUT_1[14237] = 32'b00000000000000000110001011101111;
assign LUT_1[14238] = 32'b00000000000000001000101000000100;
assign LUT_1[14239] = 32'b00000000000000000001111010000000;
assign LUT_1[14240] = 32'b00000000000000000100110010000100;
assign LUT_1[14241] = 32'b11111111111111111110000100000000;
assign LUT_1[14242] = 32'b00000000000000000000100000010101;
assign LUT_1[14243] = 32'b11111111111111111001110010010001;
assign LUT_1[14244] = 32'b00000000000000001100101011011011;
assign LUT_1[14245] = 32'b00000000000000000101111101010111;
assign LUT_1[14246] = 32'b00000000000000001000011001101100;
assign LUT_1[14247] = 32'b00000000000000000001101011101000;
assign LUT_1[14248] = 32'b00000000000000000011111111111001;
assign LUT_1[14249] = 32'b11111111111111111101010001110101;
assign LUT_1[14250] = 32'b11111111111111111111101110001010;
assign LUT_1[14251] = 32'b11111111111111111001000000000110;
assign LUT_1[14252] = 32'b00000000000000001011111001010000;
assign LUT_1[14253] = 32'b00000000000000000101001011001100;
assign LUT_1[14254] = 32'b00000000000000000111100111100001;
assign LUT_1[14255] = 32'b00000000000000000000111001011101;
assign LUT_1[14256] = 32'b00000000000000000110101101100110;
assign LUT_1[14257] = 32'b11111111111111111111111111100010;
assign LUT_1[14258] = 32'b00000000000000000010011011110111;
assign LUT_1[14259] = 32'b11111111111111111011101101110011;
assign LUT_1[14260] = 32'b00000000000000001110100110111101;
assign LUT_1[14261] = 32'b00000000000000000111111000111001;
assign LUT_1[14262] = 32'b00000000000000001010010101001110;
assign LUT_1[14263] = 32'b00000000000000000011100111001010;
assign LUT_1[14264] = 32'b00000000000000000101111011011011;
assign LUT_1[14265] = 32'b11111111111111111111001101010111;
assign LUT_1[14266] = 32'b00000000000000000001101001101100;
assign LUT_1[14267] = 32'b11111111111111111010111011101000;
assign LUT_1[14268] = 32'b00000000000000001101110100110010;
assign LUT_1[14269] = 32'b00000000000000000111000110101110;
assign LUT_1[14270] = 32'b00000000000000001001100011000011;
assign LUT_1[14271] = 32'b00000000000000000010110100111111;
assign LUT_1[14272] = 32'b00000000000000000101110100101101;
assign LUT_1[14273] = 32'b11111111111111111111000110101001;
assign LUT_1[14274] = 32'b00000000000000000001100010111110;
assign LUT_1[14275] = 32'b11111111111111111010110100111010;
assign LUT_1[14276] = 32'b00000000000000001101101110000100;
assign LUT_1[14277] = 32'b00000000000000000111000000000000;
assign LUT_1[14278] = 32'b00000000000000001001011100010101;
assign LUT_1[14279] = 32'b00000000000000000010101110010001;
assign LUT_1[14280] = 32'b00000000000000000101000010100010;
assign LUT_1[14281] = 32'b11111111111111111110010100011110;
assign LUT_1[14282] = 32'b00000000000000000000110000110011;
assign LUT_1[14283] = 32'b11111111111111111010000010101111;
assign LUT_1[14284] = 32'b00000000000000001100111011111001;
assign LUT_1[14285] = 32'b00000000000000000110001101110101;
assign LUT_1[14286] = 32'b00000000000000001000101010001010;
assign LUT_1[14287] = 32'b00000000000000000001111100000110;
assign LUT_1[14288] = 32'b00000000000000000111110000001111;
assign LUT_1[14289] = 32'b00000000000000000001000010001011;
assign LUT_1[14290] = 32'b00000000000000000011011110100000;
assign LUT_1[14291] = 32'b11111111111111111100110000011100;
assign LUT_1[14292] = 32'b00000000000000001111101001100110;
assign LUT_1[14293] = 32'b00000000000000001000111011100010;
assign LUT_1[14294] = 32'b00000000000000001011010111110111;
assign LUT_1[14295] = 32'b00000000000000000100101001110011;
assign LUT_1[14296] = 32'b00000000000000000110111110000100;
assign LUT_1[14297] = 32'b00000000000000000000010000000000;
assign LUT_1[14298] = 32'b00000000000000000010101100010101;
assign LUT_1[14299] = 32'b11111111111111111011111110010001;
assign LUT_1[14300] = 32'b00000000000000001110110111011011;
assign LUT_1[14301] = 32'b00000000000000001000001001010111;
assign LUT_1[14302] = 32'b00000000000000001010100101101100;
assign LUT_1[14303] = 32'b00000000000000000011110111101000;
assign LUT_1[14304] = 32'b00000000000000000110101111101100;
assign LUT_1[14305] = 32'b00000000000000000000000001101000;
assign LUT_1[14306] = 32'b00000000000000000010011101111101;
assign LUT_1[14307] = 32'b11111111111111111011101111111001;
assign LUT_1[14308] = 32'b00000000000000001110101001000011;
assign LUT_1[14309] = 32'b00000000000000000111111010111111;
assign LUT_1[14310] = 32'b00000000000000001010010111010100;
assign LUT_1[14311] = 32'b00000000000000000011101001010000;
assign LUT_1[14312] = 32'b00000000000000000101111101100001;
assign LUT_1[14313] = 32'b11111111111111111111001111011101;
assign LUT_1[14314] = 32'b00000000000000000001101011110010;
assign LUT_1[14315] = 32'b11111111111111111010111101101110;
assign LUT_1[14316] = 32'b00000000000000001101110110111000;
assign LUT_1[14317] = 32'b00000000000000000111001000110100;
assign LUT_1[14318] = 32'b00000000000000001001100101001001;
assign LUT_1[14319] = 32'b00000000000000000010110111000101;
assign LUT_1[14320] = 32'b00000000000000001000101011001110;
assign LUT_1[14321] = 32'b00000000000000000001111101001010;
assign LUT_1[14322] = 32'b00000000000000000100011001011111;
assign LUT_1[14323] = 32'b11111111111111111101101011011011;
assign LUT_1[14324] = 32'b00000000000000010000100100100101;
assign LUT_1[14325] = 32'b00000000000000001001110110100001;
assign LUT_1[14326] = 32'b00000000000000001100010010110110;
assign LUT_1[14327] = 32'b00000000000000000101100100110010;
assign LUT_1[14328] = 32'b00000000000000000111111001000011;
assign LUT_1[14329] = 32'b00000000000000000001001010111111;
assign LUT_1[14330] = 32'b00000000000000000011100111010100;
assign LUT_1[14331] = 32'b11111111111111111100111001010000;
assign LUT_1[14332] = 32'b00000000000000001111110010011010;
assign LUT_1[14333] = 32'b00000000000000001001000100010110;
assign LUT_1[14334] = 32'b00000000000000001011100000101011;
assign LUT_1[14335] = 32'b00000000000000000100110010100111;
assign LUT_1[14336] = 32'b00000000000000000011111111100100;
assign LUT_1[14337] = 32'b11111111111111111101010001100000;
assign LUT_1[14338] = 32'b11111111111111111111101101110101;
assign LUT_1[14339] = 32'b11111111111111111000111111110001;
assign LUT_1[14340] = 32'b00000000000000001011111000111011;
assign LUT_1[14341] = 32'b00000000000000000101001010110111;
assign LUT_1[14342] = 32'b00000000000000000111100111001100;
assign LUT_1[14343] = 32'b00000000000000000000111001001000;
assign LUT_1[14344] = 32'b00000000000000000011001101011001;
assign LUT_1[14345] = 32'b11111111111111111100011111010101;
assign LUT_1[14346] = 32'b11111111111111111110111011101010;
assign LUT_1[14347] = 32'b11111111111111111000001101100110;
assign LUT_1[14348] = 32'b00000000000000001011000110110000;
assign LUT_1[14349] = 32'b00000000000000000100011000101100;
assign LUT_1[14350] = 32'b00000000000000000110110101000001;
assign LUT_1[14351] = 32'b00000000000000000000000110111101;
assign LUT_1[14352] = 32'b00000000000000000101111011000110;
assign LUT_1[14353] = 32'b11111111111111111111001101000010;
assign LUT_1[14354] = 32'b00000000000000000001101001010111;
assign LUT_1[14355] = 32'b11111111111111111010111011010011;
assign LUT_1[14356] = 32'b00000000000000001101110100011101;
assign LUT_1[14357] = 32'b00000000000000000111000110011001;
assign LUT_1[14358] = 32'b00000000000000001001100010101110;
assign LUT_1[14359] = 32'b00000000000000000010110100101010;
assign LUT_1[14360] = 32'b00000000000000000101001000111011;
assign LUT_1[14361] = 32'b11111111111111111110011010110111;
assign LUT_1[14362] = 32'b00000000000000000000110111001100;
assign LUT_1[14363] = 32'b11111111111111111010001001001000;
assign LUT_1[14364] = 32'b00000000000000001101000010010010;
assign LUT_1[14365] = 32'b00000000000000000110010100001110;
assign LUT_1[14366] = 32'b00000000000000001000110000100011;
assign LUT_1[14367] = 32'b00000000000000000010000010011111;
assign LUT_1[14368] = 32'b00000000000000000100111010100011;
assign LUT_1[14369] = 32'b11111111111111111110001100011111;
assign LUT_1[14370] = 32'b00000000000000000000101000110100;
assign LUT_1[14371] = 32'b11111111111111111001111010110000;
assign LUT_1[14372] = 32'b00000000000000001100110011111010;
assign LUT_1[14373] = 32'b00000000000000000110000101110110;
assign LUT_1[14374] = 32'b00000000000000001000100010001011;
assign LUT_1[14375] = 32'b00000000000000000001110100000111;
assign LUT_1[14376] = 32'b00000000000000000100001000011000;
assign LUT_1[14377] = 32'b11111111111111111101011010010100;
assign LUT_1[14378] = 32'b11111111111111111111110110101001;
assign LUT_1[14379] = 32'b11111111111111111001001000100101;
assign LUT_1[14380] = 32'b00000000000000001100000001101111;
assign LUT_1[14381] = 32'b00000000000000000101010011101011;
assign LUT_1[14382] = 32'b00000000000000000111110000000000;
assign LUT_1[14383] = 32'b00000000000000000001000001111100;
assign LUT_1[14384] = 32'b00000000000000000110110110000101;
assign LUT_1[14385] = 32'b00000000000000000000001000000001;
assign LUT_1[14386] = 32'b00000000000000000010100100010110;
assign LUT_1[14387] = 32'b11111111111111111011110110010010;
assign LUT_1[14388] = 32'b00000000000000001110101111011100;
assign LUT_1[14389] = 32'b00000000000000001000000001011000;
assign LUT_1[14390] = 32'b00000000000000001010011101101101;
assign LUT_1[14391] = 32'b00000000000000000011101111101001;
assign LUT_1[14392] = 32'b00000000000000000110000011111010;
assign LUT_1[14393] = 32'b11111111111111111111010101110110;
assign LUT_1[14394] = 32'b00000000000000000001110010001011;
assign LUT_1[14395] = 32'b11111111111111111011000100000111;
assign LUT_1[14396] = 32'b00000000000000001101111101010001;
assign LUT_1[14397] = 32'b00000000000000000111001111001101;
assign LUT_1[14398] = 32'b00000000000000001001101011100010;
assign LUT_1[14399] = 32'b00000000000000000010111101011110;
assign LUT_1[14400] = 32'b00000000000000000101111101001100;
assign LUT_1[14401] = 32'b11111111111111111111001111001000;
assign LUT_1[14402] = 32'b00000000000000000001101011011101;
assign LUT_1[14403] = 32'b11111111111111111010111101011001;
assign LUT_1[14404] = 32'b00000000000000001101110110100011;
assign LUT_1[14405] = 32'b00000000000000000111001000011111;
assign LUT_1[14406] = 32'b00000000000000001001100100110100;
assign LUT_1[14407] = 32'b00000000000000000010110110110000;
assign LUT_1[14408] = 32'b00000000000000000101001011000001;
assign LUT_1[14409] = 32'b11111111111111111110011100111101;
assign LUT_1[14410] = 32'b00000000000000000000111001010010;
assign LUT_1[14411] = 32'b11111111111111111010001011001110;
assign LUT_1[14412] = 32'b00000000000000001101000100011000;
assign LUT_1[14413] = 32'b00000000000000000110010110010100;
assign LUT_1[14414] = 32'b00000000000000001000110010101001;
assign LUT_1[14415] = 32'b00000000000000000010000100100101;
assign LUT_1[14416] = 32'b00000000000000000111111000101110;
assign LUT_1[14417] = 32'b00000000000000000001001010101010;
assign LUT_1[14418] = 32'b00000000000000000011100110111111;
assign LUT_1[14419] = 32'b11111111111111111100111000111011;
assign LUT_1[14420] = 32'b00000000000000001111110010000101;
assign LUT_1[14421] = 32'b00000000000000001001000100000001;
assign LUT_1[14422] = 32'b00000000000000001011100000010110;
assign LUT_1[14423] = 32'b00000000000000000100110010010010;
assign LUT_1[14424] = 32'b00000000000000000111000110100011;
assign LUT_1[14425] = 32'b00000000000000000000011000011111;
assign LUT_1[14426] = 32'b00000000000000000010110100110100;
assign LUT_1[14427] = 32'b11111111111111111100000110110000;
assign LUT_1[14428] = 32'b00000000000000001110111111111010;
assign LUT_1[14429] = 32'b00000000000000001000010001110110;
assign LUT_1[14430] = 32'b00000000000000001010101110001011;
assign LUT_1[14431] = 32'b00000000000000000100000000000111;
assign LUT_1[14432] = 32'b00000000000000000110111000001011;
assign LUT_1[14433] = 32'b00000000000000000000001010000111;
assign LUT_1[14434] = 32'b00000000000000000010100110011100;
assign LUT_1[14435] = 32'b11111111111111111011111000011000;
assign LUT_1[14436] = 32'b00000000000000001110110001100010;
assign LUT_1[14437] = 32'b00000000000000001000000011011110;
assign LUT_1[14438] = 32'b00000000000000001010011111110011;
assign LUT_1[14439] = 32'b00000000000000000011110001101111;
assign LUT_1[14440] = 32'b00000000000000000110000110000000;
assign LUT_1[14441] = 32'b11111111111111111111010111111100;
assign LUT_1[14442] = 32'b00000000000000000001110100010001;
assign LUT_1[14443] = 32'b11111111111111111011000110001101;
assign LUT_1[14444] = 32'b00000000000000001101111111010111;
assign LUT_1[14445] = 32'b00000000000000000111010001010011;
assign LUT_1[14446] = 32'b00000000000000001001101101101000;
assign LUT_1[14447] = 32'b00000000000000000010111111100100;
assign LUT_1[14448] = 32'b00000000000000001000110011101101;
assign LUT_1[14449] = 32'b00000000000000000010000101101001;
assign LUT_1[14450] = 32'b00000000000000000100100001111110;
assign LUT_1[14451] = 32'b11111111111111111101110011111010;
assign LUT_1[14452] = 32'b00000000000000010000101101000100;
assign LUT_1[14453] = 32'b00000000000000001001111111000000;
assign LUT_1[14454] = 32'b00000000000000001100011011010101;
assign LUT_1[14455] = 32'b00000000000000000101101101010001;
assign LUT_1[14456] = 32'b00000000000000001000000001100010;
assign LUT_1[14457] = 32'b00000000000000000001010011011110;
assign LUT_1[14458] = 32'b00000000000000000011101111110011;
assign LUT_1[14459] = 32'b11111111111111111101000001101111;
assign LUT_1[14460] = 32'b00000000000000001111111010111001;
assign LUT_1[14461] = 32'b00000000000000001001001100110101;
assign LUT_1[14462] = 32'b00000000000000001011101001001010;
assign LUT_1[14463] = 32'b00000000000000000100111011000110;
assign LUT_1[14464] = 32'b00000000000000000110111111100111;
assign LUT_1[14465] = 32'b00000000000000000000010001100011;
assign LUT_1[14466] = 32'b00000000000000000010101101111000;
assign LUT_1[14467] = 32'b11111111111111111011111111110100;
assign LUT_1[14468] = 32'b00000000000000001110111000111110;
assign LUT_1[14469] = 32'b00000000000000001000001010111010;
assign LUT_1[14470] = 32'b00000000000000001010100111001111;
assign LUT_1[14471] = 32'b00000000000000000011111001001011;
assign LUT_1[14472] = 32'b00000000000000000110001101011100;
assign LUT_1[14473] = 32'b11111111111111111111011111011000;
assign LUT_1[14474] = 32'b00000000000000000001111011101101;
assign LUT_1[14475] = 32'b11111111111111111011001101101001;
assign LUT_1[14476] = 32'b00000000000000001110000110110011;
assign LUT_1[14477] = 32'b00000000000000000111011000101111;
assign LUT_1[14478] = 32'b00000000000000001001110101000100;
assign LUT_1[14479] = 32'b00000000000000000011000111000000;
assign LUT_1[14480] = 32'b00000000000000001000111011001001;
assign LUT_1[14481] = 32'b00000000000000000010001101000101;
assign LUT_1[14482] = 32'b00000000000000000100101001011010;
assign LUT_1[14483] = 32'b11111111111111111101111011010110;
assign LUT_1[14484] = 32'b00000000000000010000110100100000;
assign LUT_1[14485] = 32'b00000000000000001010000110011100;
assign LUT_1[14486] = 32'b00000000000000001100100010110001;
assign LUT_1[14487] = 32'b00000000000000000101110100101101;
assign LUT_1[14488] = 32'b00000000000000001000001000111110;
assign LUT_1[14489] = 32'b00000000000000000001011010111010;
assign LUT_1[14490] = 32'b00000000000000000011110111001111;
assign LUT_1[14491] = 32'b11111111111111111101001001001011;
assign LUT_1[14492] = 32'b00000000000000010000000010010101;
assign LUT_1[14493] = 32'b00000000000000001001010100010001;
assign LUT_1[14494] = 32'b00000000000000001011110000100110;
assign LUT_1[14495] = 32'b00000000000000000101000010100010;
assign LUT_1[14496] = 32'b00000000000000000111111010100110;
assign LUT_1[14497] = 32'b00000000000000000001001100100010;
assign LUT_1[14498] = 32'b00000000000000000011101000110111;
assign LUT_1[14499] = 32'b11111111111111111100111010110011;
assign LUT_1[14500] = 32'b00000000000000001111110011111101;
assign LUT_1[14501] = 32'b00000000000000001001000101111001;
assign LUT_1[14502] = 32'b00000000000000001011100010001110;
assign LUT_1[14503] = 32'b00000000000000000100110100001010;
assign LUT_1[14504] = 32'b00000000000000000111001000011011;
assign LUT_1[14505] = 32'b00000000000000000000011010010111;
assign LUT_1[14506] = 32'b00000000000000000010110110101100;
assign LUT_1[14507] = 32'b11111111111111111100001000101000;
assign LUT_1[14508] = 32'b00000000000000001111000001110010;
assign LUT_1[14509] = 32'b00000000000000001000010011101110;
assign LUT_1[14510] = 32'b00000000000000001010110000000011;
assign LUT_1[14511] = 32'b00000000000000000100000001111111;
assign LUT_1[14512] = 32'b00000000000000001001110110001000;
assign LUT_1[14513] = 32'b00000000000000000011001000000100;
assign LUT_1[14514] = 32'b00000000000000000101100100011001;
assign LUT_1[14515] = 32'b11111111111111111110110110010101;
assign LUT_1[14516] = 32'b00000000000000010001101111011111;
assign LUT_1[14517] = 32'b00000000000000001011000001011011;
assign LUT_1[14518] = 32'b00000000000000001101011101110000;
assign LUT_1[14519] = 32'b00000000000000000110101111101100;
assign LUT_1[14520] = 32'b00000000000000001001000011111101;
assign LUT_1[14521] = 32'b00000000000000000010010101111001;
assign LUT_1[14522] = 32'b00000000000000000100110010001110;
assign LUT_1[14523] = 32'b11111111111111111110000100001010;
assign LUT_1[14524] = 32'b00000000000000010000111101010100;
assign LUT_1[14525] = 32'b00000000000000001010001111010000;
assign LUT_1[14526] = 32'b00000000000000001100101011100101;
assign LUT_1[14527] = 32'b00000000000000000101111101100001;
assign LUT_1[14528] = 32'b00000000000000001000111101001111;
assign LUT_1[14529] = 32'b00000000000000000010001111001011;
assign LUT_1[14530] = 32'b00000000000000000100101011100000;
assign LUT_1[14531] = 32'b11111111111111111101111101011100;
assign LUT_1[14532] = 32'b00000000000000010000110110100110;
assign LUT_1[14533] = 32'b00000000000000001010001000100010;
assign LUT_1[14534] = 32'b00000000000000001100100100110111;
assign LUT_1[14535] = 32'b00000000000000000101110110110011;
assign LUT_1[14536] = 32'b00000000000000001000001011000100;
assign LUT_1[14537] = 32'b00000000000000000001011101000000;
assign LUT_1[14538] = 32'b00000000000000000011111001010101;
assign LUT_1[14539] = 32'b11111111111111111101001011010001;
assign LUT_1[14540] = 32'b00000000000000010000000100011011;
assign LUT_1[14541] = 32'b00000000000000001001010110010111;
assign LUT_1[14542] = 32'b00000000000000001011110010101100;
assign LUT_1[14543] = 32'b00000000000000000101000100101000;
assign LUT_1[14544] = 32'b00000000000000001010111000110001;
assign LUT_1[14545] = 32'b00000000000000000100001010101101;
assign LUT_1[14546] = 32'b00000000000000000110100111000010;
assign LUT_1[14547] = 32'b11111111111111111111111000111110;
assign LUT_1[14548] = 32'b00000000000000010010110010001000;
assign LUT_1[14549] = 32'b00000000000000001100000100000100;
assign LUT_1[14550] = 32'b00000000000000001110100000011001;
assign LUT_1[14551] = 32'b00000000000000000111110010010101;
assign LUT_1[14552] = 32'b00000000000000001010000110100110;
assign LUT_1[14553] = 32'b00000000000000000011011000100010;
assign LUT_1[14554] = 32'b00000000000000000101110100110111;
assign LUT_1[14555] = 32'b11111111111111111111000110110011;
assign LUT_1[14556] = 32'b00000000000000010001111111111101;
assign LUT_1[14557] = 32'b00000000000000001011010001111001;
assign LUT_1[14558] = 32'b00000000000000001101101110001110;
assign LUT_1[14559] = 32'b00000000000000000111000000001010;
assign LUT_1[14560] = 32'b00000000000000001001111000001110;
assign LUT_1[14561] = 32'b00000000000000000011001010001010;
assign LUT_1[14562] = 32'b00000000000000000101100110011111;
assign LUT_1[14563] = 32'b11111111111111111110111000011011;
assign LUT_1[14564] = 32'b00000000000000010001110001100101;
assign LUT_1[14565] = 32'b00000000000000001011000011100001;
assign LUT_1[14566] = 32'b00000000000000001101011111110110;
assign LUT_1[14567] = 32'b00000000000000000110110001110010;
assign LUT_1[14568] = 32'b00000000000000001001000110000011;
assign LUT_1[14569] = 32'b00000000000000000010010111111111;
assign LUT_1[14570] = 32'b00000000000000000100110100010100;
assign LUT_1[14571] = 32'b11111111111111111110000110010000;
assign LUT_1[14572] = 32'b00000000000000010000111111011010;
assign LUT_1[14573] = 32'b00000000000000001010010001010110;
assign LUT_1[14574] = 32'b00000000000000001100101101101011;
assign LUT_1[14575] = 32'b00000000000000000101111111100111;
assign LUT_1[14576] = 32'b00000000000000001011110011110000;
assign LUT_1[14577] = 32'b00000000000000000101000101101100;
assign LUT_1[14578] = 32'b00000000000000000111100010000001;
assign LUT_1[14579] = 32'b00000000000000000000110011111101;
assign LUT_1[14580] = 32'b00000000000000010011101101000111;
assign LUT_1[14581] = 32'b00000000000000001100111111000011;
assign LUT_1[14582] = 32'b00000000000000001111011011011000;
assign LUT_1[14583] = 32'b00000000000000001000101101010100;
assign LUT_1[14584] = 32'b00000000000000001011000001100101;
assign LUT_1[14585] = 32'b00000000000000000100010011100001;
assign LUT_1[14586] = 32'b00000000000000000110101111110110;
assign LUT_1[14587] = 32'b00000000000000000000000001110010;
assign LUT_1[14588] = 32'b00000000000000010010111010111100;
assign LUT_1[14589] = 32'b00000000000000001100001100111000;
assign LUT_1[14590] = 32'b00000000000000001110101001001101;
assign LUT_1[14591] = 32'b00000000000000000111111011001001;
assign LUT_1[14592] = 32'b00000000000000000001110011110000;
assign LUT_1[14593] = 32'b11111111111111111011000101101100;
assign LUT_1[14594] = 32'b11111111111111111101100010000001;
assign LUT_1[14595] = 32'b11111111111111110110110011111101;
assign LUT_1[14596] = 32'b00000000000000001001101101000111;
assign LUT_1[14597] = 32'b00000000000000000010111111000011;
assign LUT_1[14598] = 32'b00000000000000000101011011011000;
assign LUT_1[14599] = 32'b11111111111111111110101101010100;
assign LUT_1[14600] = 32'b00000000000000000001000001100101;
assign LUT_1[14601] = 32'b11111111111111111010010011100001;
assign LUT_1[14602] = 32'b11111111111111111100101111110110;
assign LUT_1[14603] = 32'b11111111111111110110000001110010;
assign LUT_1[14604] = 32'b00000000000000001000111010111100;
assign LUT_1[14605] = 32'b00000000000000000010001100111000;
assign LUT_1[14606] = 32'b00000000000000000100101001001101;
assign LUT_1[14607] = 32'b11111111111111111101111011001001;
assign LUT_1[14608] = 32'b00000000000000000011101111010010;
assign LUT_1[14609] = 32'b11111111111111111101000001001110;
assign LUT_1[14610] = 32'b11111111111111111111011101100011;
assign LUT_1[14611] = 32'b11111111111111111000101111011111;
assign LUT_1[14612] = 32'b00000000000000001011101000101001;
assign LUT_1[14613] = 32'b00000000000000000100111010100101;
assign LUT_1[14614] = 32'b00000000000000000111010110111010;
assign LUT_1[14615] = 32'b00000000000000000000101000110110;
assign LUT_1[14616] = 32'b00000000000000000010111101000111;
assign LUT_1[14617] = 32'b11111111111111111100001111000011;
assign LUT_1[14618] = 32'b11111111111111111110101011011000;
assign LUT_1[14619] = 32'b11111111111111110111111101010100;
assign LUT_1[14620] = 32'b00000000000000001010110110011110;
assign LUT_1[14621] = 32'b00000000000000000100001000011010;
assign LUT_1[14622] = 32'b00000000000000000110100100101111;
assign LUT_1[14623] = 32'b11111111111111111111110110101011;
assign LUT_1[14624] = 32'b00000000000000000010101110101111;
assign LUT_1[14625] = 32'b11111111111111111100000000101011;
assign LUT_1[14626] = 32'b11111111111111111110011101000000;
assign LUT_1[14627] = 32'b11111111111111110111101110111100;
assign LUT_1[14628] = 32'b00000000000000001010101000000110;
assign LUT_1[14629] = 32'b00000000000000000011111010000010;
assign LUT_1[14630] = 32'b00000000000000000110010110010111;
assign LUT_1[14631] = 32'b11111111111111111111101000010011;
assign LUT_1[14632] = 32'b00000000000000000001111100100100;
assign LUT_1[14633] = 32'b11111111111111111011001110100000;
assign LUT_1[14634] = 32'b11111111111111111101101010110101;
assign LUT_1[14635] = 32'b11111111111111110110111100110001;
assign LUT_1[14636] = 32'b00000000000000001001110101111011;
assign LUT_1[14637] = 32'b00000000000000000011000111110111;
assign LUT_1[14638] = 32'b00000000000000000101100100001100;
assign LUT_1[14639] = 32'b11111111111111111110110110001000;
assign LUT_1[14640] = 32'b00000000000000000100101010010001;
assign LUT_1[14641] = 32'b11111111111111111101111100001101;
assign LUT_1[14642] = 32'b00000000000000000000011000100010;
assign LUT_1[14643] = 32'b11111111111111111001101010011110;
assign LUT_1[14644] = 32'b00000000000000001100100011101000;
assign LUT_1[14645] = 32'b00000000000000000101110101100100;
assign LUT_1[14646] = 32'b00000000000000001000010001111001;
assign LUT_1[14647] = 32'b00000000000000000001100011110101;
assign LUT_1[14648] = 32'b00000000000000000011111000000110;
assign LUT_1[14649] = 32'b11111111111111111101001010000010;
assign LUT_1[14650] = 32'b11111111111111111111100110010111;
assign LUT_1[14651] = 32'b11111111111111111000111000010011;
assign LUT_1[14652] = 32'b00000000000000001011110001011101;
assign LUT_1[14653] = 32'b00000000000000000101000011011001;
assign LUT_1[14654] = 32'b00000000000000000111011111101110;
assign LUT_1[14655] = 32'b00000000000000000000110001101010;
assign LUT_1[14656] = 32'b00000000000000000011110001011000;
assign LUT_1[14657] = 32'b11111111111111111101000011010100;
assign LUT_1[14658] = 32'b11111111111111111111011111101001;
assign LUT_1[14659] = 32'b11111111111111111000110001100101;
assign LUT_1[14660] = 32'b00000000000000001011101010101111;
assign LUT_1[14661] = 32'b00000000000000000100111100101011;
assign LUT_1[14662] = 32'b00000000000000000111011001000000;
assign LUT_1[14663] = 32'b00000000000000000000101010111100;
assign LUT_1[14664] = 32'b00000000000000000010111111001101;
assign LUT_1[14665] = 32'b11111111111111111100010001001001;
assign LUT_1[14666] = 32'b11111111111111111110101101011110;
assign LUT_1[14667] = 32'b11111111111111110111111111011010;
assign LUT_1[14668] = 32'b00000000000000001010111000100100;
assign LUT_1[14669] = 32'b00000000000000000100001010100000;
assign LUT_1[14670] = 32'b00000000000000000110100110110101;
assign LUT_1[14671] = 32'b11111111111111111111111000110001;
assign LUT_1[14672] = 32'b00000000000000000101101100111010;
assign LUT_1[14673] = 32'b11111111111111111110111110110110;
assign LUT_1[14674] = 32'b00000000000000000001011011001011;
assign LUT_1[14675] = 32'b11111111111111111010101101000111;
assign LUT_1[14676] = 32'b00000000000000001101100110010001;
assign LUT_1[14677] = 32'b00000000000000000110111000001101;
assign LUT_1[14678] = 32'b00000000000000001001010100100010;
assign LUT_1[14679] = 32'b00000000000000000010100110011110;
assign LUT_1[14680] = 32'b00000000000000000100111010101111;
assign LUT_1[14681] = 32'b11111111111111111110001100101011;
assign LUT_1[14682] = 32'b00000000000000000000101001000000;
assign LUT_1[14683] = 32'b11111111111111111001111010111100;
assign LUT_1[14684] = 32'b00000000000000001100110100000110;
assign LUT_1[14685] = 32'b00000000000000000110000110000010;
assign LUT_1[14686] = 32'b00000000000000001000100010010111;
assign LUT_1[14687] = 32'b00000000000000000001110100010011;
assign LUT_1[14688] = 32'b00000000000000000100101100010111;
assign LUT_1[14689] = 32'b11111111111111111101111110010011;
assign LUT_1[14690] = 32'b00000000000000000000011010101000;
assign LUT_1[14691] = 32'b11111111111111111001101100100100;
assign LUT_1[14692] = 32'b00000000000000001100100101101110;
assign LUT_1[14693] = 32'b00000000000000000101110111101010;
assign LUT_1[14694] = 32'b00000000000000001000010011111111;
assign LUT_1[14695] = 32'b00000000000000000001100101111011;
assign LUT_1[14696] = 32'b00000000000000000011111010001100;
assign LUT_1[14697] = 32'b11111111111111111101001100001000;
assign LUT_1[14698] = 32'b11111111111111111111101000011101;
assign LUT_1[14699] = 32'b11111111111111111000111010011001;
assign LUT_1[14700] = 32'b00000000000000001011110011100011;
assign LUT_1[14701] = 32'b00000000000000000101000101011111;
assign LUT_1[14702] = 32'b00000000000000000111100001110100;
assign LUT_1[14703] = 32'b00000000000000000000110011110000;
assign LUT_1[14704] = 32'b00000000000000000110100111111001;
assign LUT_1[14705] = 32'b11111111111111111111111001110101;
assign LUT_1[14706] = 32'b00000000000000000010010110001010;
assign LUT_1[14707] = 32'b11111111111111111011101000000110;
assign LUT_1[14708] = 32'b00000000000000001110100001010000;
assign LUT_1[14709] = 32'b00000000000000000111110011001100;
assign LUT_1[14710] = 32'b00000000000000001010001111100001;
assign LUT_1[14711] = 32'b00000000000000000011100001011101;
assign LUT_1[14712] = 32'b00000000000000000101110101101110;
assign LUT_1[14713] = 32'b11111111111111111111000111101010;
assign LUT_1[14714] = 32'b00000000000000000001100011111111;
assign LUT_1[14715] = 32'b11111111111111111010110101111011;
assign LUT_1[14716] = 32'b00000000000000001101101111000101;
assign LUT_1[14717] = 32'b00000000000000000111000001000001;
assign LUT_1[14718] = 32'b00000000000000001001011101010110;
assign LUT_1[14719] = 32'b00000000000000000010101111010010;
assign LUT_1[14720] = 32'b00000000000000000100110011110011;
assign LUT_1[14721] = 32'b11111111111111111110000101101111;
assign LUT_1[14722] = 32'b00000000000000000000100010000100;
assign LUT_1[14723] = 32'b11111111111111111001110100000000;
assign LUT_1[14724] = 32'b00000000000000001100101101001010;
assign LUT_1[14725] = 32'b00000000000000000101111111000110;
assign LUT_1[14726] = 32'b00000000000000001000011011011011;
assign LUT_1[14727] = 32'b00000000000000000001101101010111;
assign LUT_1[14728] = 32'b00000000000000000100000001101000;
assign LUT_1[14729] = 32'b11111111111111111101010011100100;
assign LUT_1[14730] = 32'b11111111111111111111101111111001;
assign LUT_1[14731] = 32'b11111111111111111001000001110101;
assign LUT_1[14732] = 32'b00000000000000001011111010111111;
assign LUT_1[14733] = 32'b00000000000000000101001100111011;
assign LUT_1[14734] = 32'b00000000000000000111101001010000;
assign LUT_1[14735] = 32'b00000000000000000000111011001100;
assign LUT_1[14736] = 32'b00000000000000000110101111010101;
assign LUT_1[14737] = 32'b00000000000000000000000001010001;
assign LUT_1[14738] = 32'b00000000000000000010011101100110;
assign LUT_1[14739] = 32'b11111111111111111011101111100010;
assign LUT_1[14740] = 32'b00000000000000001110101000101100;
assign LUT_1[14741] = 32'b00000000000000000111111010101000;
assign LUT_1[14742] = 32'b00000000000000001010010110111101;
assign LUT_1[14743] = 32'b00000000000000000011101000111001;
assign LUT_1[14744] = 32'b00000000000000000101111101001010;
assign LUT_1[14745] = 32'b11111111111111111111001111000110;
assign LUT_1[14746] = 32'b00000000000000000001101011011011;
assign LUT_1[14747] = 32'b11111111111111111010111101010111;
assign LUT_1[14748] = 32'b00000000000000001101110110100001;
assign LUT_1[14749] = 32'b00000000000000000111001000011101;
assign LUT_1[14750] = 32'b00000000000000001001100100110010;
assign LUT_1[14751] = 32'b00000000000000000010110110101110;
assign LUT_1[14752] = 32'b00000000000000000101101110110010;
assign LUT_1[14753] = 32'b11111111111111111111000000101110;
assign LUT_1[14754] = 32'b00000000000000000001011101000011;
assign LUT_1[14755] = 32'b11111111111111111010101110111111;
assign LUT_1[14756] = 32'b00000000000000001101101000001001;
assign LUT_1[14757] = 32'b00000000000000000110111010000101;
assign LUT_1[14758] = 32'b00000000000000001001010110011010;
assign LUT_1[14759] = 32'b00000000000000000010101000010110;
assign LUT_1[14760] = 32'b00000000000000000100111100100111;
assign LUT_1[14761] = 32'b11111111111111111110001110100011;
assign LUT_1[14762] = 32'b00000000000000000000101010111000;
assign LUT_1[14763] = 32'b11111111111111111001111100110100;
assign LUT_1[14764] = 32'b00000000000000001100110101111110;
assign LUT_1[14765] = 32'b00000000000000000110000111111010;
assign LUT_1[14766] = 32'b00000000000000001000100100001111;
assign LUT_1[14767] = 32'b00000000000000000001110110001011;
assign LUT_1[14768] = 32'b00000000000000000111101010010100;
assign LUT_1[14769] = 32'b00000000000000000000111100010000;
assign LUT_1[14770] = 32'b00000000000000000011011000100101;
assign LUT_1[14771] = 32'b11111111111111111100101010100001;
assign LUT_1[14772] = 32'b00000000000000001111100011101011;
assign LUT_1[14773] = 32'b00000000000000001000110101100111;
assign LUT_1[14774] = 32'b00000000000000001011010001111100;
assign LUT_1[14775] = 32'b00000000000000000100100011111000;
assign LUT_1[14776] = 32'b00000000000000000110111000001001;
assign LUT_1[14777] = 32'b00000000000000000000001010000101;
assign LUT_1[14778] = 32'b00000000000000000010100110011010;
assign LUT_1[14779] = 32'b11111111111111111011111000010110;
assign LUT_1[14780] = 32'b00000000000000001110110001100000;
assign LUT_1[14781] = 32'b00000000000000001000000011011100;
assign LUT_1[14782] = 32'b00000000000000001010011111110001;
assign LUT_1[14783] = 32'b00000000000000000011110001101101;
assign LUT_1[14784] = 32'b00000000000000000110110001011011;
assign LUT_1[14785] = 32'b00000000000000000000000011010111;
assign LUT_1[14786] = 32'b00000000000000000010011111101100;
assign LUT_1[14787] = 32'b11111111111111111011110001101000;
assign LUT_1[14788] = 32'b00000000000000001110101010110010;
assign LUT_1[14789] = 32'b00000000000000000111111100101110;
assign LUT_1[14790] = 32'b00000000000000001010011001000011;
assign LUT_1[14791] = 32'b00000000000000000011101010111111;
assign LUT_1[14792] = 32'b00000000000000000101111111010000;
assign LUT_1[14793] = 32'b11111111111111111111010001001100;
assign LUT_1[14794] = 32'b00000000000000000001101101100001;
assign LUT_1[14795] = 32'b11111111111111111010111111011101;
assign LUT_1[14796] = 32'b00000000000000001101111000100111;
assign LUT_1[14797] = 32'b00000000000000000111001010100011;
assign LUT_1[14798] = 32'b00000000000000001001100110111000;
assign LUT_1[14799] = 32'b00000000000000000010111000110100;
assign LUT_1[14800] = 32'b00000000000000001000101100111101;
assign LUT_1[14801] = 32'b00000000000000000001111110111001;
assign LUT_1[14802] = 32'b00000000000000000100011011001110;
assign LUT_1[14803] = 32'b11111111111111111101101101001010;
assign LUT_1[14804] = 32'b00000000000000010000100110010100;
assign LUT_1[14805] = 32'b00000000000000001001111000010000;
assign LUT_1[14806] = 32'b00000000000000001100010100100101;
assign LUT_1[14807] = 32'b00000000000000000101100110100001;
assign LUT_1[14808] = 32'b00000000000000000111111010110010;
assign LUT_1[14809] = 32'b00000000000000000001001100101110;
assign LUT_1[14810] = 32'b00000000000000000011101001000011;
assign LUT_1[14811] = 32'b11111111111111111100111010111111;
assign LUT_1[14812] = 32'b00000000000000001111110100001001;
assign LUT_1[14813] = 32'b00000000000000001001000110000101;
assign LUT_1[14814] = 32'b00000000000000001011100010011010;
assign LUT_1[14815] = 32'b00000000000000000100110100010110;
assign LUT_1[14816] = 32'b00000000000000000111101100011010;
assign LUT_1[14817] = 32'b00000000000000000000111110010110;
assign LUT_1[14818] = 32'b00000000000000000011011010101011;
assign LUT_1[14819] = 32'b11111111111111111100101100100111;
assign LUT_1[14820] = 32'b00000000000000001111100101110001;
assign LUT_1[14821] = 32'b00000000000000001000110111101101;
assign LUT_1[14822] = 32'b00000000000000001011010100000010;
assign LUT_1[14823] = 32'b00000000000000000100100101111110;
assign LUT_1[14824] = 32'b00000000000000000110111010001111;
assign LUT_1[14825] = 32'b00000000000000000000001100001011;
assign LUT_1[14826] = 32'b00000000000000000010101000100000;
assign LUT_1[14827] = 32'b11111111111111111011111010011100;
assign LUT_1[14828] = 32'b00000000000000001110110011100110;
assign LUT_1[14829] = 32'b00000000000000001000000101100010;
assign LUT_1[14830] = 32'b00000000000000001010100001110111;
assign LUT_1[14831] = 32'b00000000000000000011110011110011;
assign LUT_1[14832] = 32'b00000000000000001001100111111100;
assign LUT_1[14833] = 32'b00000000000000000010111001111000;
assign LUT_1[14834] = 32'b00000000000000000101010110001101;
assign LUT_1[14835] = 32'b11111111111111111110101000001001;
assign LUT_1[14836] = 32'b00000000000000010001100001010011;
assign LUT_1[14837] = 32'b00000000000000001010110011001111;
assign LUT_1[14838] = 32'b00000000000000001101001111100100;
assign LUT_1[14839] = 32'b00000000000000000110100001100000;
assign LUT_1[14840] = 32'b00000000000000001000110101110001;
assign LUT_1[14841] = 32'b00000000000000000010000111101101;
assign LUT_1[14842] = 32'b00000000000000000100100100000010;
assign LUT_1[14843] = 32'b11111111111111111101110101111110;
assign LUT_1[14844] = 32'b00000000000000010000101111001000;
assign LUT_1[14845] = 32'b00000000000000001010000001000100;
assign LUT_1[14846] = 32'b00000000000000001100011101011001;
assign LUT_1[14847] = 32'b00000000000000000101101111010101;
assign LUT_1[14848] = 32'b11111111111111111101101110000001;
assign LUT_1[14849] = 32'b11111111111111110110111111111101;
assign LUT_1[14850] = 32'b11111111111111111001011100010010;
assign LUT_1[14851] = 32'b11111111111111110010101110001110;
assign LUT_1[14852] = 32'b00000000000000000101100111011000;
assign LUT_1[14853] = 32'b11111111111111111110111001010100;
assign LUT_1[14854] = 32'b00000000000000000001010101101001;
assign LUT_1[14855] = 32'b11111111111111111010100111100101;
assign LUT_1[14856] = 32'b11111111111111111100111011110110;
assign LUT_1[14857] = 32'b11111111111111110110001101110010;
assign LUT_1[14858] = 32'b11111111111111111000101010000111;
assign LUT_1[14859] = 32'b11111111111111110001111100000011;
assign LUT_1[14860] = 32'b00000000000000000100110101001101;
assign LUT_1[14861] = 32'b11111111111111111110000111001001;
assign LUT_1[14862] = 32'b00000000000000000000100011011110;
assign LUT_1[14863] = 32'b11111111111111111001110101011010;
assign LUT_1[14864] = 32'b11111111111111111111101001100011;
assign LUT_1[14865] = 32'b11111111111111111000111011011111;
assign LUT_1[14866] = 32'b11111111111111111011010111110100;
assign LUT_1[14867] = 32'b11111111111111110100101001110000;
assign LUT_1[14868] = 32'b00000000000000000111100010111010;
assign LUT_1[14869] = 32'b00000000000000000000110100110110;
assign LUT_1[14870] = 32'b00000000000000000011010001001011;
assign LUT_1[14871] = 32'b11111111111111111100100011000111;
assign LUT_1[14872] = 32'b11111111111111111110110111011000;
assign LUT_1[14873] = 32'b11111111111111111000001001010100;
assign LUT_1[14874] = 32'b11111111111111111010100101101001;
assign LUT_1[14875] = 32'b11111111111111110011110111100101;
assign LUT_1[14876] = 32'b00000000000000000110110000101111;
assign LUT_1[14877] = 32'b00000000000000000000000010101011;
assign LUT_1[14878] = 32'b00000000000000000010011111000000;
assign LUT_1[14879] = 32'b11111111111111111011110000111100;
assign LUT_1[14880] = 32'b11111111111111111110101001000000;
assign LUT_1[14881] = 32'b11111111111111110111111010111100;
assign LUT_1[14882] = 32'b11111111111111111010010111010001;
assign LUT_1[14883] = 32'b11111111111111110011101001001101;
assign LUT_1[14884] = 32'b00000000000000000110100010010111;
assign LUT_1[14885] = 32'b11111111111111111111110100010011;
assign LUT_1[14886] = 32'b00000000000000000010010000101000;
assign LUT_1[14887] = 32'b11111111111111111011100010100100;
assign LUT_1[14888] = 32'b11111111111111111101110110110101;
assign LUT_1[14889] = 32'b11111111111111110111001000110001;
assign LUT_1[14890] = 32'b11111111111111111001100101000110;
assign LUT_1[14891] = 32'b11111111111111110010110111000010;
assign LUT_1[14892] = 32'b00000000000000000101110000001100;
assign LUT_1[14893] = 32'b11111111111111111111000010001000;
assign LUT_1[14894] = 32'b00000000000000000001011110011101;
assign LUT_1[14895] = 32'b11111111111111111010110000011001;
assign LUT_1[14896] = 32'b00000000000000000000100100100010;
assign LUT_1[14897] = 32'b11111111111111111001110110011110;
assign LUT_1[14898] = 32'b11111111111111111100010010110011;
assign LUT_1[14899] = 32'b11111111111111110101100100101111;
assign LUT_1[14900] = 32'b00000000000000001000011101111001;
assign LUT_1[14901] = 32'b00000000000000000001101111110101;
assign LUT_1[14902] = 32'b00000000000000000100001100001010;
assign LUT_1[14903] = 32'b11111111111111111101011110000110;
assign LUT_1[14904] = 32'b11111111111111111111110010010111;
assign LUT_1[14905] = 32'b11111111111111111001000100010011;
assign LUT_1[14906] = 32'b11111111111111111011100000101000;
assign LUT_1[14907] = 32'b11111111111111110100110010100100;
assign LUT_1[14908] = 32'b00000000000000000111101011101110;
assign LUT_1[14909] = 32'b00000000000000000000111101101010;
assign LUT_1[14910] = 32'b00000000000000000011011001111111;
assign LUT_1[14911] = 32'b11111111111111111100101011111011;
assign LUT_1[14912] = 32'b11111111111111111111101011101001;
assign LUT_1[14913] = 32'b11111111111111111000111101100101;
assign LUT_1[14914] = 32'b11111111111111111011011001111010;
assign LUT_1[14915] = 32'b11111111111111110100101011110110;
assign LUT_1[14916] = 32'b00000000000000000111100101000000;
assign LUT_1[14917] = 32'b00000000000000000000110110111100;
assign LUT_1[14918] = 32'b00000000000000000011010011010001;
assign LUT_1[14919] = 32'b11111111111111111100100101001101;
assign LUT_1[14920] = 32'b11111111111111111110111001011110;
assign LUT_1[14921] = 32'b11111111111111111000001011011010;
assign LUT_1[14922] = 32'b11111111111111111010100111101111;
assign LUT_1[14923] = 32'b11111111111111110011111001101011;
assign LUT_1[14924] = 32'b00000000000000000110110010110101;
assign LUT_1[14925] = 32'b00000000000000000000000100110001;
assign LUT_1[14926] = 32'b00000000000000000010100001000110;
assign LUT_1[14927] = 32'b11111111111111111011110011000010;
assign LUT_1[14928] = 32'b00000000000000000001100111001011;
assign LUT_1[14929] = 32'b11111111111111111010111001000111;
assign LUT_1[14930] = 32'b11111111111111111101010101011100;
assign LUT_1[14931] = 32'b11111111111111110110100111011000;
assign LUT_1[14932] = 32'b00000000000000001001100000100010;
assign LUT_1[14933] = 32'b00000000000000000010110010011110;
assign LUT_1[14934] = 32'b00000000000000000101001110110011;
assign LUT_1[14935] = 32'b11111111111111111110100000101111;
assign LUT_1[14936] = 32'b00000000000000000000110101000000;
assign LUT_1[14937] = 32'b11111111111111111010000110111100;
assign LUT_1[14938] = 32'b11111111111111111100100011010001;
assign LUT_1[14939] = 32'b11111111111111110101110101001101;
assign LUT_1[14940] = 32'b00000000000000001000101110010111;
assign LUT_1[14941] = 32'b00000000000000000010000000010011;
assign LUT_1[14942] = 32'b00000000000000000100011100101000;
assign LUT_1[14943] = 32'b11111111111111111101101110100100;
assign LUT_1[14944] = 32'b00000000000000000000100110101000;
assign LUT_1[14945] = 32'b11111111111111111001111000100100;
assign LUT_1[14946] = 32'b11111111111111111100010100111001;
assign LUT_1[14947] = 32'b11111111111111110101100110110101;
assign LUT_1[14948] = 32'b00000000000000001000011111111111;
assign LUT_1[14949] = 32'b00000000000000000001110001111011;
assign LUT_1[14950] = 32'b00000000000000000100001110010000;
assign LUT_1[14951] = 32'b11111111111111111101100000001100;
assign LUT_1[14952] = 32'b11111111111111111111110100011101;
assign LUT_1[14953] = 32'b11111111111111111001000110011001;
assign LUT_1[14954] = 32'b11111111111111111011100010101110;
assign LUT_1[14955] = 32'b11111111111111110100110100101010;
assign LUT_1[14956] = 32'b00000000000000000111101101110100;
assign LUT_1[14957] = 32'b00000000000000000000111111110000;
assign LUT_1[14958] = 32'b00000000000000000011011100000101;
assign LUT_1[14959] = 32'b11111111111111111100101110000001;
assign LUT_1[14960] = 32'b00000000000000000010100010001010;
assign LUT_1[14961] = 32'b11111111111111111011110100000110;
assign LUT_1[14962] = 32'b11111111111111111110010000011011;
assign LUT_1[14963] = 32'b11111111111111110111100010010111;
assign LUT_1[14964] = 32'b00000000000000001010011011100001;
assign LUT_1[14965] = 32'b00000000000000000011101101011101;
assign LUT_1[14966] = 32'b00000000000000000110001001110010;
assign LUT_1[14967] = 32'b11111111111111111111011011101110;
assign LUT_1[14968] = 32'b00000000000000000001101111111111;
assign LUT_1[14969] = 32'b11111111111111111011000001111011;
assign LUT_1[14970] = 32'b11111111111111111101011110010000;
assign LUT_1[14971] = 32'b11111111111111110110110000001100;
assign LUT_1[14972] = 32'b00000000000000001001101001010110;
assign LUT_1[14973] = 32'b00000000000000000010111011010010;
assign LUT_1[14974] = 32'b00000000000000000101010111100111;
assign LUT_1[14975] = 32'b11111111111111111110101001100011;
assign LUT_1[14976] = 32'b00000000000000000000101110000100;
assign LUT_1[14977] = 32'b11111111111111111010000000000000;
assign LUT_1[14978] = 32'b11111111111111111100011100010101;
assign LUT_1[14979] = 32'b11111111111111110101101110010001;
assign LUT_1[14980] = 32'b00000000000000001000100111011011;
assign LUT_1[14981] = 32'b00000000000000000001111001010111;
assign LUT_1[14982] = 32'b00000000000000000100010101101100;
assign LUT_1[14983] = 32'b11111111111111111101100111101000;
assign LUT_1[14984] = 32'b11111111111111111111111011111001;
assign LUT_1[14985] = 32'b11111111111111111001001101110101;
assign LUT_1[14986] = 32'b11111111111111111011101010001010;
assign LUT_1[14987] = 32'b11111111111111110100111100000110;
assign LUT_1[14988] = 32'b00000000000000000111110101010000;
assign LUT_1[14989] = 32'b00000000000000000001000111001100;
assign LUT_1[14990] = 32'b00000000000000000011100011100001;
assign LUT_1[14991] = 32'b11111111111111111100110101011101;
assign LUT_1[14992] = 32'b00000000000000000010101001100110;
assign LUT_1[14993] = 32'b11111111111111111011111011100010;
assign LUT_1[14994] = 32'b11111111111111111110010111110111;
assign LUT_1[14995] = 32'b11111111111111110111101001110011;
assign LUT_1[14996] = 32'b00000000000000001010100010111101;
assign LUT_1[14997] = 32'b00000000000000000011110100111001;
assign LUT_1[14998] = 32'b00000000000000000110010001001110;
assign LUT_1[14999] = 32'b11111111111111111111100011001010;
assign LUT_1[15000] = 32'b00000000000000000001110111011011;
assign LUT_1[15001] = 32'b11111111111111111011001001010111;
assign LUT_1[15002] = 32'b11111111111111111101100101101100;
assign LUT_1[15003] = 32'b11111111111111110110110111101000;
assign LUT_1[15004] = 32'b00000000000000001001110000110010;
assign LUT_1[15005] = 32'b00000000000000000011000010101110;
assign LUT_1[15006] = 32'b00000000000000000101011111000011;
assign LUT_1[15007] = 32'b11111111111111111110110000111111;
assign LUT_1[15008] = 32'b00000000000000000001101001000011;
assign LUT_1[15009] = 32'b11111111111111111010111010111111;
assign LUT_1[15010] = 32'b11111111111111111101010111010100;
assign LUT_1[15011] = 32'b11111111111111110110101001010000;
assign LUT_1[15012] = 32'b00000000000000001001100010011010;
assign LUT_1[15013] = 32'b00000000000000000010110100010110;
assign LUT_1[15014] = 32'b00000000000000000101010000101011;
assign LUT_1[15015] = 32'b11111111111111111110100010100111;
assign LUT_1[15016] = 32'b00000000000000000000110110111000;
assign LUT_1[15017] = 32'b11111111111111111010001000110100;
assign LUT_1[15018] = 32'b11111111111111111100100101001001;
assign LUT_1[15019] = 32'b11111111111111110101110111000101;
assign LUT_1[15020] = 32'b00000000000000001000110000001111;
assign LUT_1[15021] = 32'b00000000000000000010000010001011;
assign LUT_1[15022] = 32'b00000000000000000100011110100000;
assign LUT_1[15023] = 32'b11111111111111111101110000011100;
assign LUT_1[15024] = 32'b00000000000000000011100100100101;
assign LUT_1[15025] = 32'b11111111111111111100110110100001;
assign LUT_1[15026] = 32'b11111111111111111111010010110110;
assign LUT_1[15027] = 32'b11111111111111111000100100110010;
assign LUT_1[15028] = 32'b00000000000000001011011101111100;
assign LUT_1[15029] = 32'b00000000000000000100101111111000;
assign LUT_1[15030] = 32'b00000000000000000111001100001101;
assign LUT_1[15031] = 32'b00000000000000000000011110001001;
assign LUT_1[15032] = 32'b00000000000000000010110010011010;
assign LUT_1[15033] = 32'b11111111111111111100000100010110;
assign LUT_1[15034] = 32'b11111111111111111110100000101011;
assign LUT_1[15035] = 32'b11111111111111110111110010100111;
assign LUT_1[15036] = 32'b00000000000000001010101011110001;
assign LUT_1[15037] = 32'b00000000000000000011111101101101;
assign LUT_1[15038] = 32'b00000000000000000110011010000010;
assign LUT_1[15039] = 32'b11111111111111111111101011111110;
assign LUT_1[15040] = 32'b00000000000000000010101011101100;
assign LUT_1[15041] = 32'b11111111111111111011111101101000;
assign LUT_1[15042] = 32'b11111111111111111110011001111101;
assign LUT_1[15043] = 32'b11111111111111110111101011111001;
assign LUT_1[15044] = 32'b00000000000000001010100101000011;
assign LUT_1[15045] = 32'b00000000000000000011110110111111;
assign LUT_1[15046] = 32'b00000000000000000110010011010100;
assign LUT_1[15047] = 32'b11111111111111111111100101010000;
assign LUT_1[15048] = 32'b00000000000000000001111001100001;
assign LUT_1[15049] = 32'b11111111111111111011001011011101;
assign LUT_1[15050] = 32'b11111111111111111101100111110010;
assign LUT_1[15051] = 32'b11111111111111110110111001101110;
assign LUT_1[15052] = 32'b00000000000000001001110010111000;
assign LUT_1[15053] = 32'b00000000000000000011000100110100;
assign LUT_1[15054] = 32'b00000000000000000101100001001001;
assign LUT_1[15055] = 32'b11111111111111111110110011000101;
assign LUT_1[15056] = 32'b00000000000000000100100111001110;
assign LUT_1[15057] = 32'b11111111111111111101111001001010;
assign LUT_1[15058] = 32'b00000000000000000000010101011111;
assign LUT_1[15059] = 32'b11111111111111111001100111011011;
assign LUT_1[15060] = 32'b00000000000000001100100000100101;
assign LUT_1[15061] = 32'b00000000000000000101110010100001;
assign LUT_1[15062] = 32'b00000000000000001000001110110110;
assign LUT_1[15063] = 32'b00000000000000000001100000110010;
assign LUT_1[15064] = 32'b00000000000000000011110101000011;
assign LUT_1[15065] = 32'b11111111111111111101000110111111;
assign LUT_1[15066] = 32'b11111111111111111111100011010100;
assign LUT_1[15067] = 32'b11111111111111111000110101010000;
assign LUT_1[15068] = 32'b00000000000000001011101110011010;
assign LUT_1[15069] = 32'b00000000000000000101000000010110;
assign LUT_1[15070] = 32'b00000000000000000111011100101011;
assign LUT_1[15071] = 32'b00000000000000000000101110100111;
assign LUT_1[15072] = 32'b00000000000000000011100110101011;
assign LUT_1[15073] = 32'b11111111111111111100111000100111;
assign LUT_1[15074] = 32'b11111111111111111111010100111100;
assign LUT_1[15075] = 32'b11111111111111111000100110111000;
assign LUT_1[15076] = 32'b00000000000000001011100000000010;
assign LUT_1[15077] = 32'b00000000000000000100110001111110;
assign LUT_1[15078] = 32'b00000000000000000111001110010011;
assign LUT_1[15079] = 32'b00000000000000000000100000001111;
assign LUT_1[15080] = 32'b00000000000000000010110100100000;
assign LUT_1[15081] = 32'b11111111111111111100000110011100;
assign LUT_1[15082] = 32'b11111111111111111110100010110001;
assign LUT_1[15083] = 32'b11111111111111110111110100101101;
assign LUT_1[15084] = 32'b00000000000000001010101101110111;
assign LUT_1[15085] = 32'b00000000000000000011111111110011;
assign LUT_1[15086] = 32'b00000000000000000110011100001000;
assign LUT_1[15087] = 32'b11111111111111111111101110000100;
assign LUT_1[15088] = 32'b00000000000000000101100010001101;
assign LUT_1[15089] = 32'b11111111111111111110110100001001;
assign LUT_1[15090] = 32'b00000000000000000001010000011110;
assign LUT_1[15091] = 32'b11111111111111111010100010011010;
assign LUT_1[15092] = 32'b00000000000000001101011011100100;
assign LUT_1[15093] = 32'b00000000000000000110101101100000;
assign LUT_1[15094] = 32'b00000000000000001001001001110101;
assign LUT_1[15095] = 32'b00000000000000000010011011110001;
assign LUT_1[15096] = 32'b00000000000000000100110000000010;
assign LUT_1[15097] = 32'b11111111111111111110000001111110;
assign LUT_1[15098] = 32'b00000000000000000000011110010011;
assign LUT_1[15099] = 32'b11111111111111111001110000001111;
assign LUT_1[15100] = 32'b00000000000000001100101001011001;
assign LUT_1[15101] = 32'b00000000000000000101111011010101;
assign LUT_1[15102] = 32'b00000000000000001000010111101010;
assign LUT_1[15103] = 32'b00000000000000000001101001100110;
assign LUT_1[15104] = 32'b11111111111111111011100010001101;
assign LUT_1[15105] = 32'b11111111111111110100110100001001;
assign LUT_1[15106] = 32'b11111111111111110111010000011110;
assign LUT_1[15107] = 32'b11111111111111110000100010011010;
assign LUT_1[15108] = 32'b00000000000000000011011011100100;
assign LUT_1[15109] = 32'b11111111111111111100101101100000;
assign LUT_1[15110] = 32'b11111111111111111111001001110101;
assign LUT_1[15111] = 32'b11111111111111111000011011110001;
assign LUT_1[15112] = 32'b11111111111111111010110000000010;
assign LUT_1[15113] = 32'b11111111111111110100000001111110;
assign LUT_1[15114] = 32'b11111111111111110110011110010011;
assign LUT_1[15115] = 32'b11111111111111101111110000001111;
assign LUT_1[15116] = 32'b00000000000000000010101001011001;
assign LUT_1[15117] = 32'b11111111111111111011111011010101;
assign LUT_1[15118] = 32'b11111111111111111110010111101010;
assign LUT_1[15119] = 32'b11111111111111110111101001100110;
assign LUT_1[15120] = 32'b11111111111111111101011101101111;
assign LUT_1[15121] = 32'b11111111111111110110101111101011;
assign LUT_1[15122] = 32'b11111111111111111001001100000000;
assign LUT_1[15123] = 32'b11111111111111110010011101111100;
assign LUT_1[15124] = 32'b00000000000000000101010111000110;
assign LUT_1[15125] = 32'b11111111111111111110101001000010;
assign LUT_1[15126] = 32'b00000000000000000001000101010111;
assign LUT_1[15127] = 32'b11111111111111111010010111010011;
assign LUT_1[15128] = 32'b11111111111111111100101011100100;
assign LUT_1[15129] = 32'b11111111111111110101111101100000;
assign LUT_1[15130] = 32'b11111111111111111000011001110101;
assign LUT_1[15131] = 32'b11111111111111110001101011110001;
assign LUT_1[15132] = 32'b00000000000000000100100100111011;
assign LUT_1[15133] = 32'b11111111111111111101110110110111;
assign LUT_1[15134] = 32'b00000000000000000000010011001100;
assign LUT_1[15135] = 32'b11111111111111111001100101001000;
assign LUT_1[15136] = 32'b11111111111111111100011101001100;
assign LUT_1[15137] = 32'b11111111111111110101101111001000;
assign LUT_1[15138] = 32'b11111111111111111000001011011101;
assign LUT_1[15139] = 32'b11111111111111110001011101011001;
assign LUT_1[15140] = 32'b00000000000000000100010110100011;
assign LUT_1[15141] = 32'b11111111111111111101101000011111;
assign LUT_1[15142] = 32'b00000000000000000000000100110100;
assign LUT_1[15143] = 32'b11111111111111111001010110110000;
assign LUT_1[15144] = 32'b11111111111111111011101011000001;
assign LUT_1[15145] = 32'b11111111111111110100111100111101;
assign LUT_1[15146] = 32'b11111111111111110111011001010010;
assign LUT_1[15147] = 32'b11111111111111110000101011001110;
assign LUT_1[15148] = 32'b00000000000000000011100100011000;
assign LUT_1[15149] = 32'b11111111111111111100110110010100;
assign LUT_1[15150] = 32'b11111111111111111111010010101001;
assign LUT_1[15151] = 32'b11111111111111111000100100100101;
assign LUT_1[15152] = 32'b11111111111111111110011000101110;
assign LUT_1[15153] = 32'b11111111111111110111101010101010;
assign LUT_1[15154] = 32'b11111111111111111010000110111111;
assign LUT_1[15155] = 32'b11111111111111110011011000111011;
assign LUT_1[15156] = 32'b00000000000000000110010010000101;
assign LUT_1[15157] = 32'b11111111111111111111100100000001;
assign LUT_1[15158] = 32'b00000000000000000010000000010110;
assign LUT_1[15159] = 32'b11111111111111111011010010010010;
assign LUT_1[15160] = 32'b11111111111111111101100110100011;
assign LUT_1[15161] = 32'b11111111111111110110111000011111;
assign LUT_1[15162] = 32'b11111111111111111001010100110100;
assign LUT_1[15163] = 32'b11111111111111110010100110110000;
assign LUT_1[15164] = 32'b00000000000000000101011111111010;
assign LUT_1[15165] = 32'b11111111111111111110110001110110;
assign LUT_1[15166] = 32'b00000000000000000001001110001011;
assign LUT_1[15167] = 32'b11111111111111111010100000000111;
assign LUT_1[15168] = 32'b11111111111111111101011111110101;
assign LUT_1[15169] = 32'b11111111111111110110110001110001;
assign LUT_1[15170] = 32'b11111111111111111001001110000110;
assign LUT_1[15171] = 32'b11111111111111110010100000000010;
assign LUT_1[15172] = 32'b00000000000000000101011001001100;
assign LUT_1[15173] = 32'b11111111111111111110101011001000;
assign LUT_1[15174] = 32'b00000000000000000001000111011101;
assign LUT_1[15175] = 32'b11111111111111111010011001011001;
assign LUT_1[15176] = 32'b11111111111111111100101101101010;
assign LUT_1[15177] = 32'b11111111111111110101111111100110;
assign LUT_1[15178] = 32'b11111111111111111000011011111011;
assign LUT_1[15179] = 32'b11111111111111110001101101110111;
assign LUT_1[15180] = 32'b00000000000000000100100111000001;
assign LUT_1[15181] = 32'b11111111111111111101111000111101;
assign LUT_1[15182] = 32'b00000000000000000000010101010010;
assign LUT_1[15183] = 32'b11111111111111111001100111001110;
assign LUT_1[15184] = 32'b11111111111111111111011011010111;
assign LUT_1[15185] = 32'b11111111111111111000101101010011;
assign LUT_1[15186] = 32'b11111111111111111011001001101000;
assign LUT_1[15187] = 32'b11111111111111110100011011100100;
assign LUT_1[15188] = 32'b00000000000000000111010100101110;
assign LUT_1[15189] = 32'b00000000000000000000100110101010;
assign LUT_1[15190] = 32'b00000000000000000011000010111111;
assign LUT_1[15191] = 32'b11111111111111111100010100111011;
assign LUT_1[15192] = 32'b11111111111111111110101001001100;
assign LUT_1[15193] = 32'b11111111111111110111111011001000;
assign LUT_1[15194] = 32'b11111111111111111010010111011101;
assign LUT_1[15195] = 32'b11111111111111110011101001011001;
assign LUT_1[15196] = 32'b00000000000000000110100010100011;
assign LUT_1[15197] = 32'b11111111111111111111110100011111;
assign LUT_1[15198] = 32'b00000000000000000010010000110100;
assign LUT_1[15199] = 32'b11111111111111111011100010110000;
assign LUT_1[15200] = 32'b11111111111111111110011010110100;
assign LUT_1[15201] = 32'b11111111111111110111101100110000;
assign LUT_1[15202] = 32'b11111111111111111010001001000101;
assign LUT_1[15203] = 32'b11111111111111110011011011000001;
assign LUT_1[15204] = 32'b00000000000000000110010100001011;
assign LUT_1[15205] = 32'b11111111111111111111100110000111;
assign LUT_1[15206] = 32'b00000000000000000010000010011100;
assign LUT_1[15207] = 32'b11111111111111111011010100011000;
assign LUT_1[15208] = 32'b11111111111111111101101000101001;
assign LUT_1[15209] = 32'b11111111111111110110111010100101;
assign LUT_1[15210] = 32'b11111111111111111001010110111010;
assign LUT_1[15211] = 32'b11111111111111110010101000110110;
assign LUT_1[15212] = 32'b00000000000000000101100010000000;
assign LUT_1[15213] = 32'b11111111111111111110110011111100;
assign LUT_1[15214] = 32'b00000000000000000001010000010001;
assign LUT_1[15215] = 32'b11111111111111111010100010001101;
assign LUT_1[15216] = 32'b00000000000000000000010110010110;
assign LUT_1[15217] = 32'b11111111111111111001101000010010;
assign LUT_1[15218] = 32'b11111111111111111100000100100111;
assign LUT_1[15219] = 32'b11111111111111110101010110100011;
assign LUT_1[15220] = 32'b00000000000000001000001111101101;
assign LUT_1[15221] = 32'b00000000000000000001100001101001;
assign LUT_1[15222] = 32'b00000000000000000011111101111110;
assign LUT_1[15223] = 32'b11111111111111111101001111111010;
assign LUT_1[15224] = 32'b11111111111111111111100100001011;
assign LUT_1[15225] = 32'b11111111111111111000110110000111;
assign LUT_1[15226] = 32'b11111111111111111011010010011100;
assign LUT_1[15227] = 32'b11111111111111110100100100011000;
assign LUT_1[15228] = 32'b00000000000000000111011101100010;
assign LUT_1[15229] = 32'b00000000000000000000101111011110;
assign LUT_1[15230] = 32'b00000000000000000011001011110011;
assign LUT_1[15231] = 32'b11111111111111111100011101101111;
assign LUT_1[15232] = 32'b11111111111111111110100010010000;
assign LUT_1[15233] = 32'b11111111111111110111110100001100;
assign LUT_1[15234] = 32'b11111111111111111010010000100001;
assign LUT_1[15235] = 32'b11111111111111110011100010011101;
assign LUT_1[15236] = 32'b00000000000000000110011011100111;
assign LUT_1[15237] = 32'b11111111111111111111101101100011;
assign LUT_1[15238] = 32'b00000000000000000010001001111000;
assign LUT_1[15239] = 32'b11111111111111111011011011110100;
assign LUT_1[15240] = 32'b11111111111111111101110000000101;
assign LUT_1[15241] = 32'b11111111111111110111000010000001;
assign LUT_1[15242] = 32'b11111111111111111001011110010110;
assign LUT_1[15243] = 32'b11111111111111110010110000010010;
assign LUT_1[15244] = 32'b00000000000000000101101001011100;
assign LUT_1[15245] = 32'b11111111111111111110111011011000;
assign LUT_1[15246] = 32'b00000000000000000001010111101101;
assign LUT_1[15247] = 32'b11111111111111111010101001101001;
assign LUT_1[15248] = 32'b00000000000000000000011101110010;
assign LUT_1[15249] = 32'b11111111111111111001101111101110;
assign LUT_1[15250] = 32'b11111111111111111100001100000011;
assign LUT_1[15251] = 32'b11111111111111110101011101111111;
assign LUT_1[15252] = 32'b00000000000000001000010111001001;
assign LUT_1[15253] = 32'b00000000000000000001101001000101;
assign LUT_1[15254] = 32'b00000000000000000100000101011010;
assign LUT_1[15255] = 32'b11111111111111111101010111010110;
assign LUT_1[15256] = 32'b11111111111111111111101011100111;
assign LUT_1[15257] = 32'b11111111111111111000111101100011;
assign LUT_1[15258] = 32'b11111111111111111011011001111000;
assign LUT_1[15259] = 32'b11111111111111110100101011110100;
assign LUT_1[15260] = 32'b00000000000000000111100100111110;
assign LUT_1[15261] = 32'b00000000000000000000110110111010;
assign LUT_1[15262] = 32'b00000000000000000011010011001111;
assign LUT_1[15263] = 32'b11111111111111111100100101001011;
assign LUT_1[15264] = 32'b11111111111111111111011101001111;
assign LUT_1[15265] = 32'b11111111111111111000101111001011;
assign LUT_1[15266] = 32'b11111111111111111011001011100000;
assign LUT_1[15267] = 32'b11111111111111110100011101011100;
assign LUT_1[15268] = 32'b00000000000000000111010110100110;
assign LUT_1[15269] = 32'b00000000000000000000101000100010;
assign LUT_1[15270] = 32'b00000000000000000011000100110111;
assign LUT_1[15271] = 32'b11111111111111111100010110110011;
assign LUT_1[15272] = 32'b11111111111111111110101011000100;
assign LUT_1[15273] = 32'b11111111111111110111111101000000;
assign LUT_1[15274] = 32'b11111111111111111010011001010101;
assign LUT_1[15275] = 32'b11111111111111110011101011010001;
assign LUT_1[15276] = 32'b00000000000000000110100100011011;
assign LUT_1[15277] = 32'b11111111111111111111110110010111;
assign LUT_1[15278] = 32'b00000000000000000010010010101100;
assign LUT_1[15279] = 32'b11111111111111111011100100101000;
assign LUT_1[15280] = 32'b00000000000000000001011000110001;
assign LUT_1[15281] = 32'b11111111111111111010101010101101;
assign LUT_1[15282] = 32'b11111111111111111101000111000010;
assign LUT_1[15283] = 32'b11111111111111110110011000111110;
assign LUT_1[15284] = 32'b00000000000000001001010010001000;
assign LUT_1[15285] = 32'b00000000000000000010100100000100;
assign LUT_1[15286] = 32'b00000000000000000101000000011001;
assign LUT_1[15287] = 32'b11111111111111111110010010010101;
assign LUT_1[15288] = 32'b00000000000000000000100110100110;
assign LUT_1[15289] = 32'b11111111111111111001111000100010;
assign LUT_1[15290] = 32'b11111111111111111100010100110111;
assign LUT_1[15291] = 32'b11111111111111110101100110110011;
assign LUT_1[15292] = 32'b00000000000000001000011111111101;
assign LUT_1[15293] = 32'b00000000000000000001110001111001;
assign LUT_1[15294] = 32'b00000000000000000100001110001110;
assign LUT_1[15295] = 32'b11111111111111111101100000001010;
assign LUT_1[15296] = 32'b00000000000000000000011111111000;
assign LUT_1[15297] = 32'b11111111111111111001110001110100;
assign LUT_1[15298] = 32'b11111111111111111100001110001001;
assign LUT_1[15299] = 32'b11111111111111110101100000000101;
assign LUT_1[15300] = 32'b00000000000000001000011001001111;
assign LUT_1[15301] = 32'b00000000000000000001101011001011;
assign LUT_1[15302] = 32'b00000000000000000100000111100000;
assign LUT_1[15303] = 32'b11111111111111111101011001011100;
assign LUT_1[15304] = 32'b11111111111111111111101101101101;
assign LUT_1[15305] = 32'b11111111111111111000111111101001;
assign LUT_1[15306] = 32'b11111111111111111011011011111110;
assign LUT_1[15307] = 32'b11111111111111110100101101111010;
assign LUT_1[15308] = 32'b00000000000000000111100111000100;
assign LUT_1[15309] = 32'b00000000000000000000111001000000;
assign LUT_1[15310] = 32'b00000000000000000011010101010101;
assign LUT_1[15311] = 32'b11111111111111111100100111010001;
assign LUT_1[15312] = 32'b00000000000000000010011011011010;
assign LUT_1[15313] = 32'b11111111111111111011101101010110;
assign LUT_1[15314] = 32'b11111111111111111110001001101011;
assign LUT_1[15315] = 32'b11111111111111110111011011100111;
assign LUT_1[15316] = 32'b00000000000000001010010100110001;
assign LUT_1[15317] = 32'b00000000000000000011100110101101;
assign LUT_1[15318] = 32'b00000000000000000110000011000010;
assign LUT_1[15319] = 32'b11111111111111111111010100111110;
assign LUT_1[15320] = 32'b00000000000000000001101001001111;
assign LUT_1[15321] = 32'b11111111111111111010111011001011;
assign LUT_1[15322] = 32'b11111111111111111101010111100000;
assign LUT_1[15323] = 32'b11111111111111110110101001011100;
assign LUT_1[15324] = 32'b00000000000000001001100010100110;
assign LUT_1[15325] = 32'b00000000000000000010110100100010;
assign LUT_1[15326] = 32'b00000000000000000101010000110111;
assign LUT_1[15327] = 32'b11111111111111111110100010110011;
assign LUT_1[15328] = 32'b00000000000000000001011010110111;
assign LUT_1[15329] = 32'b11111111111111111010101100110011;
assign LUT_1[15330] = 32'b11111111111111111101001001001000;
assign LUT_1[15331] = 32'b11111111111111110110011011000100;
assign LUT_1[15332] = 32'b00000000000000001001010100001110;
assign LUT_1[15333] = 32'b00000000000000000010100110001010;
assign LUT_1[15334] = 32'b00000000000000000101000010011111;
assign LUT_1[15335] = 32'b11111111111111111110010100011011;
assign LUT_1[15336] = 32'b00000000000000000000101000101100;
assign LUT_1[15337] = 32'b11111111111111111001111010101000;
assign LUT_1[15338] = 32'b11111111111111111100010110111101;
assign LUT_1[15339] = 32'b11111111111111110101101000111001;
assign LUT_1[15340] = 32'b00000000000000001000100010000011;
assign LUT_1[15341] = 32'b00000000000000000001110011111111;
assign LUT_1[15342] = 32'b00000000000000000100010000010100;
assign LUT_1[15343] = 32'b11111111111111111101100010010000;
assign LUT_1[15344] = 32'b00000000000000000011010110011001;
assign LUT_1[15345] = 32'b11111111111111111100101000010101;
assign LUT_1[15346] = 32'b11111111111111111111000100101010;
assign LUT_1[15347] = 32'b11111111111111111000010110100110;
assign LUT_1[15348] = 32'b00000000000000001011001111110000;
assign LUT_1[15349] = 32'b00000000000000000100100001101100;
assign LUT_1[15350] = 32'b00000000000000000110111110000001;
assign LUT_1[15351] = 32'b00000000000000000000001111111101;
assign LUT_1[15352] = 32'b00000000000000000010100100001110;
assign LUT_1[15353] = 32'b11111111111111111011110110001010;
assign LUT_1[15354] = 32'b11111111111111111110010010011111;
assign LUT_1[15355] = 32'b11111111111111110111100100011011;
assign LUT_1[15356] = 32'b00000000000000001010011101100101;
assign LUT_1[15357] = 32'b00000000000000000011101111100001;
assign LUT_1[15358] = 32'b00000000000000000110001011110110;
assign LUT_1[15359] = 32'b11111111111111111111011101110010;
assign LUT_1[15360] = 32'b00000000000000001010010110010100;
assign LUT_1[15361] = 32'b00000000000000000011101000010000;
assign LUT_1[15362] = 32'b00000000000000000110000100100101;
assign LUT_1[15363] = 32'b11111111111111111111010110100001;
assign LUT_1[15364] = 32'b00000000000000010010001111101011;
assign LUT_1[15365] = 32'b00000000000000001011100001100111;
assign LUT_1[15366] = 32'b00000000000000001101111101111100;
assign LUT_1[15367] = 32'b00000000000000000111001111111000;
assign LUT_1[15368] = 32'b00000000000000001001100100001001;
assign LUT_1[15369] = 32'b00000000000000000010110110000101;
assign LUT_1[15370] = 32'b00000000000000000101010010011010;
assign LUT_1[15371] = 32'b11111111111111111110100100010110;
assign LUT_1[15372] = 32'b00000000000000010001011101100000;
assign LUT_1[15373] = 32'b00000000000000001010101111011100;
assign LUT_1[15374] = 32'b00000000000000001101001011110001;
assign LUT_1[15375] = 32'b00000000000000000110011101101101;
assign LUT_1[15376] = 32'b00000000000000001100010001110110;
assign LUT_1[15377] = 32'b00000000000000000101100011110010;
assign LUT_1[15378] = 32'b00000000000000001000000000000111;
assign LUT_1[15379] = 32'b00000000000000000001010010000011;
assign LUT_1[15380] = 32'b00000000000000010100001011001101;
assign LUT_1[15381] = 32'b00000000000000001101011101001001;
assign LUT_1[15382] = 32'b00000000000000001111111001011110;
assign LUT_1[15383] = 32'b00000000000000001001001011011010;
assign LUT_1[15384] = 32'b00000000000000001011011111101011;
assign LUT_1[15385] = 32'b00000000000000000100110001100111;
assign LUT_1[15386] = 32'b00000000000000000111001101111100;
assign LUT_1[15387] = 32'b00000000000000000000011111111000;
assign LUT_1[15388] = 32'b00000000000000010011011001000010;
assign LUT_1[15389] = 32'b00000000000000001100101010111110;
assign LUT_1[15390] = 32'b00000000000000001111000111010011;
assign LUT_1[15391] = 32'b00000000000000001000011001001111;
assign LUT_1[15392] = 32'b00000000000000001011010001010011;
assign LUT_1[15393] = 32'b00000000000000000100100011001111;
assign LUT_1[15394] = 32'b00000000000000000110111111100100;
assign LUT_1[15395] = 32'b00000000000000000000010001100000;
assign LUT_1[15396] = 32'b00000000000000010011001010101010;
assign LUT_1[15397] = 32'b00000000000000001100011100100110;
assign LUT_1[15398] = 32'b00000000000000001110111000111011;
assign LUT_1[15399] = 32'b00000000000000001000001010110111;
assign LUT_1[15400] = 32'b00000000000000001010011111001000;
assign LUT_1[15401] = 32'b00000000000000000011110001000100;
assign LUT_1[15402] = 32'b00000000000000000110001101011001;
assign LUT_1[15403] = 32'b11111111111111111111011111010101;
assign LUT_1[15404] = 32'b00000000000000010010011000011111;
assign LUT_1[15405] = 32'b00000000000000001011101010011011;
assign LUT_1[15406] = 32'b00000000000000001110000110110000;
assign LUT_1[15407] = 32'b00000000000000000111011000101100;
assign LUT_1[15408] = 32'b00000000000000001101001100110101;
assign LUT_1[15409] = 32'b00000000000000000110011110110001;
assign LUT_1[15410] = 32'b00000000000000001000111011000110;
assign LUT_1[15411] = 32'b00000000000000000010001101000010;
assign LUT_1[15412] = 32'b00000000000000010101000110001100;
assign LUT_1[15413] = 32'b00000000000000001110011000001000;
assign LUT_1[15414] = 32'b00000000000000010000110100011101;
assign LUT_1[15415] = 32'b00000000000000001010000110011001;
assign LUT_1[15416] = 32'b00000000000000001100011010101010;
assign LUT_1[15417] = 32'b00000000000000000101101100100110;
assign LUT_1[15418] = 32'b00000000000000001000001000111011;
assign LUT_1[15419] = 32'b00000000000000000001011010110111;
assign LUT_1[15420] = 32'b00000000000000010100010100000001;
assign LUT_1[15421] = 32'b00000000000000001101100101111101;
assign LUT_1[15422] = 32'b00000000000000010000000010010010;
assign LUT_1[15423] = 32'b00000000000000001001010100001110;
assign LUT_1[15424] = 32'b00000000000000001100010011111100;
assign LUT_1[15425] = 32'b00000000000000000101100101111000;
assign LUT_1[15426] = 32'b00000000000000001000000010001101;
assign LUT_1[15427] = 32'b00000000000000000001010100001001;
assign LUT_1[15428] = 32'b00000000000000010100001101010011;
assign LUT_1[15429] = 32'b00000000000000001101011111001111;
assign LUT_1[15430] = 32'b00000000000000001111111011100100;
assign LUT_1[15431] = 32'b00000000000000001001001101100000;
assign LUT_1[15432] = 32'b00000000000000001011100001110001;
assign LUT_1[15433] = 32'b00000000000000000100110011101101;
assign LUT_1[15434] = 32'b00000000000000000111010000000010;
assign LUT_1[15435] = 32'b00000000000000000000100001111110;
assign LUT_1[15436] = 32'b00000000000000010011011011001000;
assign LUT_1[15437] = 32'b00000000000000001100101101000100;
assign LUT_1[15438] = 32'b00000000000000001111001001011001;
assign LUT_1[15439] = 32'b00000000000000001000011011010101;
assign LUT_1[15440] = 32'b00000000000000001110001111011110;
assign LUT_1[15441] = 32'b00000000000000000111100001011010;
assign LUT_1[15442] = 32'b00000000000000001001111101101111;
assign LUT_1[15443] = 32'b00000000000000000011001111101011;
assign LUT_1[15444] = 32'b00000000000000010110001000110101;
assign LUT_1[15445] = 32'b00000000000000001111011010110001;
assign LUT_1[15446] = 32'b00000000000000010001110111000110;
assign LUT_1[15447] = 32'b00000000000000001011001001000010;
assign LUT_1[15448] = 32'b00000000000000001101011101010011;
assign LUT_1[15449] = 32'b00000000000000000110101111001111;
assign LUT_1[15450] = 32'b00000000000000001001001011100100;
assign LUT_1[15451] = 32'b00000000000000000010011101100000;
assign LUT_1[15452] = 32'b00000000000000010101010110101010;
assign LUT_1[15453] = 32'b00000000000000001110101000100110;
assign LUT_1[15454] = 32'b00000000000000010001000100111011;
assign LUT_1[15455] = 32'b00000000000000001010010110110111;
assign LUT_1[15456] = 32'b00000000000000001101001110111011;
assign LUT_1[15457] = 32'b00000000000000000110100000110111;
assign LUT_1[15458] = 32'b00000000000000001000111101001100;
assign LUT_1[15459] = 32'b00000000000000000010001111001000;
assign LUT_1[15460] = 32'b00000000000000010101001000010010;
assign LUT_1[15461] = 32'b00000000000000001110011010001110;
assign LUT_1[15462] = 32'b00000000000000010000110110100011;
assign LUT_1[15463] = 32'b00000000000000001010001000011111;
assign LUT_1[15464] = 32'b00000000000000001100011100110000;
assign LUT_1[15465] = 32'b00000000000000000101101110101100;
assign LUT_1[15466] = 32'b00000000000000001000001011000001;
assign LUT_1[15467] = 32'b00000000000000000001011100111101;
assign LUT_1[15468] = 32'b00000000000000010100010110000111;
assign LUT_1[15469] = 32'b00000000000000001101101000000011;
assign LUT_1[15470] = 32'b00000000000000010000000100011000;
assign LUT_1[15471] = 32'b00000000000000001001010110010100;
assign LUT_1[15472] = 32'b00000000000000001111001010011101;
assign LUT_1[15473] = 32'b00000000000000001000011100011001;
assign LUT_1[15474] = 32'b00000000000000001010111000101110;
assign LUT_1[15475] = 32'b00000000000000000100001010101010;
assign LUT_1[15476] = 32'b00000000000000010111000011110100;
assign LUT_1[15477] = 32'b00000000000000010000010101110000;
assign LUT_1[15478] = 32'b00000000000000010010110010000101;
assign LUT_1[15479] = 32'b00000000000000001100000100000001;
assign LUT_1[15480] = 32'b00000000000000001110011000010010;
assign LUT_1[15481] = 32'b00000000000000000111101010001110;
assign LUT_1[15482] = 32'b00000000000000001010000110100011;
assign LUT_1[15483] = 32'b00000000000000000011011000011111;
assign LUT_1[15484] = 32'b00000000000000010110010001101001;
assign LUT_1[15485] = 32'b00000000000000001111100011100101;
assign LUT_1[15486] = 32'b00000000000000010001111111111010;
assign LUT_1[15487] = 32'b00000000000000001011010001110110;
assign LUT_1[15488] = 32'b00000000000000001101010110010111;
assign LUT_1[15489] = 32'b00000000000000000110101000010011;
assign LUT_1[15490] = 32'b00000000000000001001000100101000;
assign LUT_1[15491] = 32'b00000000000000000010010110100100;
assign LUT_1[15492] = 32'b00000000000000010101001111101110;
assign LUT_1[15493] = 32'b00000000000000001110100001101010;
assign LUT_1[15494] = 32'b00000000000000010000111101111111;
assign LUT_1[15495] = 32'b00000000000000001010001111111011;
assign LUT_1[15496] = 32'b00000000000000001100100100001100;
assign LUT_1[15497] = 32'b00000000000000000101110110001000;
assign LUT_1[15498] = 32'b00000000000000001000010010011101;
assign LUT_1[15499] = 32'b00000000000000000001100100011001;
assign LUT_1[15500] = 32'b00000000000000010100011101100011;
assign LUT_1[15501] = 32'b00000000000000001101101111011111;
assign LUT_1[15502] = 32'b00000000000000010000001011110100;
assign LUT_1[15503] = 32'b00000000000000001001011101110000;
assign LUT_1[15504] = 32'b00000000000000001111010001111001;
assign LUT_1[15505] = 32'b00000000000000001000100011110101;
assign LUT_1[15506] = 32'b00000000000000001011000000001010;
assign LUT_1[15507] = 32'b00000000000000000100010010000110;
assign LUT_1[15508] = 32'b00000000000000010111001011010000;
assign LUT_1[15509] = 32'b00000000000000010000011101001100;
assign LUT_1[15510] = 32'b00000000000000010010111001100001;
assign LUT_1[15511] = 32'b00000000000000001100001011011101;
assign LUT_1[15512] = 32'b00000000000000001110011111101110;
assign LUT_1[15513] = 32'b00000000000000000111110001101010;
assign LUT_1[15514] = 32'b00000000000000001010001101111111;
assign LUT_1[15515] = 32'b00000000000000000011011111111011;
assign LUT_1[15516] = 32'b00000000000000010110011001000101;
assign LUT_1[15517] = 32'b00000000000000001111101011000001;
assign LUT_1[15518] = 32'b00000000000000010010000111010110;
assign LUT_1[15519] = 32'b00000000000000001011011001010010;
assign LUT_1[15520] = 32'b00000000000000001110010001010110;
assign LUT_1[15521] = 32'b00000000000000000111100011010010;
assign LUT_1[15522] = 32'b00000000000000001001111111100111;
assign LUT_1[15523] = 32'b00000000000000000011010001100011;
assign LUT_1[15524] = 32'b00000000000000010110001010101101;
assign LUT_1[15525] = 32'b00000000000000001111011100101001;
assign LUT_1[15526] = 32'b00000000000000010001111000111110;
assign LUT_1[15527] = 32'b00000000000000001011001010111010;
assign LUT_1[15528] = 32'b00000000000000001101011111001011;
assign LUT_1[15529] = 32'b00000000000000000110110001000111;
assign LUT_1[15530] = 32'b00000000000000001001001101011100;
assign LUT_1[15531] = 32'b00000000000000000010011111011000;
assign LUT_1[15532] = 32'b00000000000000010101011000100010;
assign LUT_1[15533] = 32'b00000000000000001110101010011110;
assign LUT_1[15534] = 32'b00000000000000010001000110110011;
assign LUT_1[15535] = 32'b00000000000000001010011000101111;
assign LUT_1[15536] = 32'b00000000000000010000001100111000;
assign LUT_1[15537] = 32'b00000000000000001001011110110100;
assign LUT_1[15538] = 32'b00000000000000001011111011001001;
assign LUT_1[15539] = 32'b00000000000000000101001101000101;
assign LUT_1[15540] = 32'b00000000000000011000000110001111;
assign LUT_1[15541] = 32'b00000000000000010001011000001011;
assign LUT_1[15542] = 32'b00000000000000010011110100100000;
assign LUT_1[15543] = 32'b00000000000000001101000110011100;
assign LUT_1[15544] = 32'b00000000000000001111011010101101;
assign LUT_1[15545] = 32'b00000000000000001000101100101001;
assign LUT_1[15546] = 32'b00000000000000001011001000111110;
assign LUT_1[15547] = 32'b00000000000000000100011010111010;
assign LUT_1[15548] = 32'b00000000000000010111010100000100;
assign LUT_1[15549] = 32'b00000000000000010000100110000000;
assign LUT_1[15550] = 32'b00000000000000010011000010010101;
assign LUT_1[15551] = 32'b00000000000000001100010100010001;
assign LUT_1[15552] = 32'b00000000000000001111010011111111;
assign LUT_1[15553] = 32'b00000000000000001000100101111011;
assign LUT_1[15554] = 32'b00000000000000001011000010010000;
assign LUT_1[15555] = 32'b00000000000000000100010100001100;
assign LUT_1[15556] = 32'b00000000000000010111001101010110;
assign LUT_1[15557] = 32'b00000000000000010000011111010010;
assign LUT_1[15558] = 32'b00000000000000010010111011100111;
assign LUT_1[15559] = 32'b00000000000000001100001101100011;
assign LUT_1[15560] = 32'b00000000000000001110100001110100;
assign LUT_1[15561] = 32'b00000000000000000111110011110000;
assign LUT_1[15562] = 32'b00000000000000001010010000000101;
assign LUT_1[15563] = 32'b00000000000000000011100010000001;
assign LUT_1[15564] = 32'b00000000000000010110011011001011;
assign LUT_1[15565] = 32'b00000000000000001111101101000111;
assign LUT_1[15566] = 32'b00000000000000010010001001011100;
assign LUT_1[15567] = 32'b00000000000000001011011011011000;
assign LUT_1[15568] = 32'b00000000000000010001001111100001;
assign LUT_1[15569] = 32'b00000000000000001010100001011101;
assign LUT_1[15570] = 32'b00000000000000001100111101110010;
assign LUT_1[15571] = 32'b00000000000000000110001111101110;
assign LUT_1[15572] = 32'b00000000000000011001001000111000;
assign LUT_1[15573] = 32'b00000000000000010010011010110100;
assign LUT_1[15574] = 32'b00000000000000010100110111001001;
assign LUT_1[15575] = 32'b00000000000000001110001001000101;
assign LUT_1[15576] = 32'b00000000000000010000011101010110;
assign LUT_1[15577] = 32'b00000000000000001001101111010010;
assign LUT_1[15578] = 32'b00000000000000001100001011100111;
assign LUT_1[15579] = 32'b00000000000000000101011101100011;
assign LUT_1[15580] = 32'b00000000000000011000010110101101;
assign LUT_1[15581] = 32'b00000000000000010001101000101001;
assign LUT_1[15582] = 32'b00000000000000010100000100111110;
assign LUT_1[15583] = 32'b00000000000000001101010110111010;
assign LUT_1[15584] = 32'b00000000000000010000001110111110;
assign LUT_1[15585] = 32'b00000000000000001001100000111010;
assign LUT_1[15586] = 32'b00000000000000001011111101001111;
assign LUT_1[15587] = 32'b00000000000000000101001111001011;
assign LUT_1[15588] = 32'b00000000000000011000001000010101;
assign LUT_1[15589] = 32'b00000000000000010001011010010001;
assign LUT_1[15590] = 32'b00000000000000010011110110100110;
assign LUT_1[15591] = 32'b00000000000000001101001000100010;
assign LUT_1[15592] = 32'b00000000000000001111011100110011;
assign LUT_1[15593] = 32'b00000000000000001000101110101111;
assign LUT_1[15594] = 32'b00000000000000001011001011000100;
assign LUT_1[15595] = 32'b00000000000000000100011101000000;
assign LUT_1[15596] = 32'b00000000000000010111010110001010;
assign LUT_1[15597] = 32'b00000000000000010000101000000110;
assign LUT_1[15598] = 32'b00000000000000010011000100011011;
assign LUT_1[15599] = 32'b00000000000000001100010110010111;
assign LUT_1[15600] = 32'b00000000000000010010001010100000;
assign LUT_1[15601] = 32'b00000000000000001011011100011100;
assign LUT_1[15602] = 32'b00000000000000001101111000110001;
assign LUT_1[15603] = 32'b00000000000000000111001010101101;
assign LUT_1[15604] = 32'b00000000000000011010000011110111;
assign LUT_1[15605] = 32'b00000000000000010011010101110011;
assign LUT_1[15606] = 32'b00000000000000010101110010001000;
assign LUT_1[15607] = 32'b00000000000000001111000100000100;
assign LUT_1[15608] = 32'b00000000000000010001011000010101;
assign LUT_1[15609] = 32'b00000000000000001010101010010001;
assign LUT_1[15610] = 32'b00000000000000001101000110100110;
assign LUT_1[15611] = 32'b00000000000000000110011000100010;
assign LUT_1[15612] = 32'b00000000000000011001010001101100;
assign LUT_1[15613] = 32'b00000000000000010010100011101000;
assign LUT_1[15614] = 32'b00000000000000010100111111111101;
assign LUT_1[15615] = 32'b00000000000000001110010001111001;
assign LUT_1[15616] = 32'b00000000000000001000001010100000;
assign LUT_1[15617] = 32'b00000000000000000001011100011100;
assign LUT_1[15618] = 32'b00000000000000000011111000110001;
assign LUT_1[15619] = 32'b11111111111111111101001010101101;
assign LUT_1[15620] = 32'b00000000000000010000000011110111;
assign LUT_1[15621] = 32'b00000000000000001001010101110011;
assign LUT_1[15622] = 32'b00000000000000001011110010001000;
assign LUT_1[15623] = 32'b00000000000000000101000100000100;
assign LUT_1[15624] = 32'b00000000000000000111011000010101;
assign LUT_1[15625] = 32'b00000000000000000000101010010001;
assign LUT_1[15626] = 32'b00000000000000000011000110100110;
assign LUT_1[15627] = 32'b11111111111111111100011000100010;
assign LUT_1[15628] = 32'b00000000000000001111010001101100;
assign LUT_1[15629] = 32'b00000000000000001000100011101000;
assign LUT_1[15630] = 32'b00000000000000001010111111111101;
assign LUT_1[15631] = 32'b00000000000000000100010001111001;
assign LUT_1[15632] = 32'b00000000000000001010000110000010;
assign LUT_1[15633] = 32'b00000000000000000011010111111110;
assign LUT_1[15634] = 32'b00000000000000000101110100010011;
assign LUT_1[15635] = 32'b11111111111111111111000110001111;
assign LUT_1[15636] = 32'b00000000000000010001111111011001;
assign LUT_1[15637] = 32'b00000000000000001011010001010101;
assign LUT_1[15638] = 32'b00000000000000001101101101101010;
assign LUT_1[15639] = 32'b00000000000000000110111111100110;
assign LUT_1[15640] = 32'b00000000000000001001010011110111;
assign LUT_1[15641] = 32'b00000000000000000010100101110011;
assign LUT_1[15642] = 32'b00000000000000000101000010001000;
assign LUT_1[15643] = 32'b11111111111111111110010100000100;
assign LUT_1[15644] = 32'b00000000000000010001001101001110;
assign LUT_1[15645] = 32'b00000000000000001010011111001010;
assign LUT_1[15646] = 32'b00000000000000001100111011011111;
assign LUT_1[15647] = 32'b00000000000000000110001101011011;
assign LUT_1[15648] = 32'b00000000000000001001000101011111;
assign LUT_1[15649] = 32'b00000000000000000010010111011011;
assign LUT_1[15650] = 32'b00000000000000000100110011110000;
assign LUT_1[15651] = 32'b11111111111111111110000101101100;
assign LUT_1[15652] = 32'b00000000000000010000111110110110;
assign LUT_1[15653] = 32'b00000000000000001010010000110010;
assign LUT_1[15654] = 32'b00000000000000001100101101000111;
assign LUT_1[15655] = 32'b00000000000000000101111111000011;
assign LUT_1[15656] = 32'b00000000000000001000010011010100;
assign LUT_1[15657] = 32'b00000000000000000001100101010000;
assign LUT_1[15658] = 32'b00000000000000000100000001100101;
assign LUT_1[15659] = 32'b11111111111111111101010011100001;
assign LUT_1[15660] = 32'b00000000000000010000001100101011;
assign LUT_1[15661] = 32'b00000000000000001001011110100111;
assign LUT_1[15662] = 32'b00000000000000001011111010111100;
assign LUT_1[15663] = 32'b00000000000000000101001100111000;
assign LUT_1[15664] = 32'b00000000000000001011000001000001;
assign LUT_1[15665] = 32'b00000000000000000100010010111101;
assign LUT_1[15666] = 32'b00000000000000000110101111010010;
assign LUT_1[15667] = 32'b00000000000000000000000001001110;
assign LUT_1[15668] = 32'b00000000000000010010111010011000;
assign LUT_1[15669] = 32'b00000000000000001100001100010100;
assign LUT_1[15670] = 32'b00000000000000001110101000101001;
assign LUT_1[15671] = 32'b00000000000000000111111010100101;
assign LUT_1[15672] = 32'b00000000000000001010001110110110;
assign LUT_1[15673] = 32'b00000000000000000011100000110010;
assign LUT_1[15674] = 32'b00000000000000000101111101000111;
assign LUT_1[15675] = 32'b11111111111111111111001111000011;
assign LUT_1[15676] = 32'b00000000000000010010001000001101;
assign LUT_1[15677] = 32'b00000000000000001011011010001001;
assign LUT_1[15678] = 32'b00000000000000001101110110011110;
assign LUT_1[15679] = 32'b00000000000000000111001000011010;
assign LUT_1[15680] = 32'b00000000000000001010001000001000;
assign LUT_1[15681] = 32'b00000000000000000011011010000100;
assign LUT_1[15682] = 32'b00000000000000000101110110011001;
assign LUT_1[15683] = 32'b11111111111111111111001000010101;
assign LUT_1[15684] = 32'b00000000000000010010000001011111;
assign LUT_1[15685] = 32'b00000000000000001011010011011011;
assign LUT_1[15686] = 32'b00000000000000001101101111110000;
assign LUT_1[15687] = 32'b00000000000000000111000001101100;
assign LUT_1[15688] = 32'b00000000000000001001010101111101;
assign LUT_1[15689] = 32'b00000000000000000010100111111001;
assign LUT_1[15690] = 32'b00000000000000000101000100001110;
assign LUT_1[15691] = 32'b11111111111111111110010110001010;
assign LUT_1[15692] = 32'b00000000000000010001001111010100;
assign LUT_1[15693] = 32'b00000000000000001010100001010000;
assign LUT_1[15694] = 32'b00000000000000001100111101100101;
assign LUT_1[15695] = 32'b00000000000000000110001111100001;
assign LUT_1[15696] = 32'b00000000000000001100000011101010;
assign LUT_1[15697] = 32'b00000000000000000101010101100110;
assign LUT_1[15698] = 32'b00000000000000000111110001111011;
assign LUT_1[15699] = 32'b00000000000000000001000011110111;
assign LUT_1[15700] = 32'b00000000000000010011111101000001;
assign LUT_1[15701] = 32'b00000000000000001101001110111101;
assign LUT_1[15702] = 32'b00000000000000001111101011010010;
assign LUT_1[15703] = 32'b00000000000000001000111101001110;
assign LUT_1[15704] = 32'b00000000000000001011010001011111;
assign LUT_1[15705] = 32'b00000000000000000100100011011011;
assign LUT_1[15706] = 32'b00000000000000000110111111110000;
assign LUT_1[15707] = 32'b00000000000000000000010001101100;
assign LUT_1[15708] = 32'b00000000000000010011001010110110;
assign LUT_1[15709] = 32'b00000000000000001100011100110010;
assign LUT_1[15710] = 32'b00000000000000001110111001000111;
assign LUT_1[15711] = 32'b00000000000000001000001011000011;
assign LUT_1[15712] = 32'b00000000000000001011000011000111;
assign LUT_1[15713] = 32'b00000000000000000100010101000011;
assign LUT_1[15714] = 32'b00000000000000000110110001011000;
assign LUT_1[15715] = 32'b00000000000000000000000011010100;
assign LUT_1[15716] = 32'b00000000000000010010111100011110;
assign LUT_1[15717] = 32'b00000000000000001100001110011010;
assign LUT_1[15718] = 32'b00000000000000001110101010101111;
assign LUT_1[15719] = 32'b00000000000000000111111100101011;
assign LUT_1[15720] = 32'b00000000000000001010010000111100;
assign LUT_1[15721] = 32'b00000000000000000011100010111000;
assign LUT_1[15722] = 32'b00000000000000000101111111001101;
assign LUT_1[15723] = 32'b11111111111111111111010001001001;
assign LUT_1[15724] = 32'b00000000000000010010001010010011;
assign LUT_1[15725] = 32'b00000000000000001011011100001111;
assign LUT_1[15726] = 32'b00000000000000001101111000100100;
assign LUT_1[15727] = 32'b00000000000000000111001010100000;
assign LUT_1[15728] = 32'b00000000000000001100111110101001;
assign LUT_1[15729] = 32'b00000000000000000110010000100101;
assign LUT_1[15730] = 32'b00000000000000001000101100111010;
assign LUT_1[15731] = 32'b00000000000000000001111110110110;
assign LUT_1[15732] = 32'b00000000000000010100111000000000;
assign LUT_1[15733] = 32'b00000000000000001110001001111100;
assign LUT_1[15734] = 32'b00000000000000010000100110010001;
assign LUT_1[15735] = 32'b00000000000000001001111000001101;
assign LUT_1[15736] = 32'b00000000000000001100001100011110;
assign LUT_1[15737] = 32'b00000000000000000101011110011010;
assign LUT_1[15738] = 32'b00000000000000000111111010101111;
assign LUT_1[15739] = 32'b00000000000000000001001100101011;
assign LUT_1[15740] = 32'b00000000000000010100000101110101;
assign LUT_1[15741] = 32'b00000000000000001101010111110001;
assign LUT_1[15742] = 32'b00000000000000001111110100000110;
assign LUT_1[15743] = 32'b00000000000000001001000110000010;
assign LUT_1[15744] = 32'b00000000000000001011001010100011;
assign LUT_1[15745] = 32'b00000000000000000100011100011111;
assign LUT_1[15746] = 32'b00000000000000000110111000110100;
assign LUT_1[15747] = 32'b00000000000000000000001010110000;
assign LUT_1[15748] = 32'b00000000000000010011000011111010;
assign LUT_1[15749] = 32'b00000000000000001100010101110110;
assign LUT_1[15750] = 32'b00000000000000001110110010001011;
assign LUT_1[15751] = 32'b00000000000000001000000100000111;
assign LUT_1[15752] = 32'b00000000000000001010011000011000;
assign LUT_1[15753] = 32'b00000000000000000011101010010100;
assign LUT_1[15754] = 32'b00000000000000000110000110101001;
assign LUT_1[15755] = 32'b11111111111111111111011000100101;
assign LUT_1[15756] = 32'b00000000000000010010010001101111;
assign LUT_1[15757] = 32'b00000000000000001011100011101011;
assign LUT_1[15758] = 32'b00000000000000001110000000000000;
assign LUT_1[15759] = 32'b00000000000000000111010001111100;
assign LUT_1[15760] = 32'b00000000000000001101000110000101;
assign LUT_1[15761] = 32'b00000000000000000110011000000001;
assign LUT_1[15762] = 32'b00000000000000001000110100010110;
assign LUT_1[15763] = 32'b00000000000000000010000110010010;
assign LUT_1[15764] = 32'b00000000000000010100111111011100;
assign LUT_1[15765] = 32'b00000000000000001110010001011000;
assign LUT_1[15766] = 32'b00000000000000010000101101101101;
assign LUT_1[15767] = 32'b00000000000000001001111111101001;
assign LUT_1[15768] = 32'b00000000000000001100010011111010;
assign LUT_1[15769] = 32'b00000000000000000101100101110110;
assign LUT_1[15770] = 32'b00000000000000001000000010001011;
assign LUT_1[15771] = 32'b00000000000000000001010100000111;
assign LUT_1[15772] = 32'b00000000000000010100001101010001;
assign LUT_1[15773] = 32'b00000000000000001101011111001101;
assign LUT_1[15774] = 32'b00000000000000001111111011100010;
assign LUT_1[15775] = 32'b00000000000000001001001101011110;
assign LUT_1[15776] = 32'b00000000000000001100000101100010;
assign LUT_1[15777] = 32'b00000000000000000101010111011110;
assign LUT_1[15778] = 32'b00000000000000000111110011110011;
assign LUT_1[15779] = 32'b00000000000000000001000101101111;
assign LUT_1[15780] = 32'b00000000000000010011111110111001;
assign LUT_1[15781] = 32'b00000000000000001101010000110101;
assign LUT_1[15782] = 32'b00000000000000001111101101001010;
assign LUT_1[15783] = 32'b00000000000000001000111111000110;
assign LUT_1[15784] = 32'b00000000000000001011010011010111;
assign LUT_1[15785] = 32'b00000000000000000100100101010011;
assign LUT_1[15786] = 32'b00000000000000000111000001101000;
assign LUT_1[15787] = 32'b00000000000000000000010011100100;
assign LUT_1[15788] = 32'b00000000000000010011001100101110;
assign LUT_1[15789] = 32'b00000000000000001100011110101010;
assign LUT_1[15790] = 32'b00000000000000001110111010111111;
assign LUT_1[15791] = 32'b00000000000000001000001100111011;
assign LUT_1[15792] = 32'b00000000000000001110000001000100;
assign LUT_1[15793] = 32'b00000000000000000111010011000000;
assign LUT_1[15794] = 32'b00000000000000001001101111010101;
assign LUT_1[15795] = 32'b00000000000000000011000001010001;
assign LUT_1[15796] = 32'b00000000000000010101111010011011;
assign LUT_1[15797] = 32'b00000000000000001111001100010111;
assign LUT_1[15798] = 32'b00000000000000010001101000101100;
assign LUT_1[15799] = 32'b00000000000000001010111010101000;
assign LUT_1[15800] = 32'b00000000000000001101001110111001;
assign LUT_1[15801] = 32'b00000000000000000110100000110101;
assign LUT_1[15802] = 32'b00000000000000001000111101001010;
assign LUT_1[15803] = 32'b00000000000000000010001111000110;
assign LUT_1[15804] = 32'b00000000000000010101001000010000;
assign LUT_1[15805] = 32'b00000000000000001110011010001100;
assign LUT_1[15806] = 32'b00000000000000010000110110100001;
assign LUT_1[15807] = 32'b00000000000000001010001000011101;
assign LUT_1[15808] = 32'b00000000000000001101001000001011;
assign LUT_1[15809] = 32'b00000000000000000110011010000111;
assign LUT_1[15810] = 32'b00000000000000001000110110011100;
assign LUT_1[15811] = 32'b00000000000000000010001000011000;
assign LUT_1[15812] = 32'b00000000000000010101000001100010;
assign LUT_1[15813] = 32'b00000000000000001110010011011110;
assign LUT_1[15814] = 32'b00000000000000010000101111110011;
assign LUT_1[15815] = 32'b00000000000000001010000001101111;
assign LUT_1[15816] = 32'b00000000000000001100010110000000;
assign LUT_1[15817] = 32'b00000000000000000101100111111100;
assign LUT_1[15818] = 32'b00000000000000001000000100010001;
assign LUT_1[15819] = 32'b00000000000000000001010110001101;
assign LUT_1[15820] = 32'b00000000000000010100001111010111;
assign LUT_1[15821] = 32'b00000000000000001101100001010011;
assign LUT_1[15822] = 32'b00000000000000001111111101101000;
assign LUT_1[15823] = 32'b00000000000000001001001111100100;
assign LUT_1[15824] = 32'b00000000000000001111000011101101;
assign LUT_1[15825] = 32'b00000000000000001000010101101001;
assign LUT_1[15826] = 32'b00000000000000001010110001111110;
assign LUT_1[15827] = 32'b00000000000000000100000011111010;
assign LUT_1[15828] = 32'b00000000000000010110111101000100;
assign LUT_1[15829] = 32'b00000000000000010000001111000000;
assign LUT_1[15830] = 32'b00000000000000010010101011010101;
assign LUT_1[15831] = 32'b00000000000000001011111101010001;
assign LUT_1[15832] = 32'b00000000000000001110010001100010;
assign LUT_1[15833] = 32'b00000000000000000111100011011110;
assign LUT_1[15834] = 32'b00000000000000001001111111110011;
assign LUT_1[15835] = 32'b00000000000000000011010001101111;
assign LUT_1[15836] = 32'b00000000000000010110001010111001;
assign LUT_1[15837] = 32'b00000000000000001111011100110101;
assign LUT_1[15838] = 32'b00000000000000010001111001001010;
assign LUT_1[15839] = 32'b00000000000000001011001011000110;
assign LUT_1[15840] = 32'b00000000000000001110000011001010;
assign LUT_1[15841] = 32'b00000000000000000111010101000110;
assign LUT_1[15842] = 32'b00000000000000001001110001011011;
assign LUT_1[15843] = 32'b00000000000000000011000011010111;
assign LUT_1[15844] = 32'b00000000000000010101111100100001;
assign LUT_1[15845] = 32'b00000000000000001111001110011101;
assign LUT_1[15846] = 32'b00000000000000010001101010110010;
assign LUT_1[15847] = 32'b00000000000000001010111100101110;
assign LUT_1[15848] = 32'b00000000000000001101010000111111;
assign LUT_1[15849] = 32'b00000000000000000110100010111011;
assign LUT_1[15850] = 32'b00000000000000001000111111010000;
assign LUT_1[15851] = 32'b00000000000000000010010001001100;
assign LUT_1[15852] = 32'b00000000000000010101001010010110;
assign LUT_1[15853] = 32'b00000000000000001110011100010010;
assign LUT_1[15854] = 32'b00000000000000010000111000100111;
assign LUT_1[15855] = 32'b00000000000000001010001010100011;
assign LUT_1[15856] = 32'b00000000000000001111111110101100;
assign LUT_1[15857] = 32'b00000000000000001001010000101000;
assign LUT_1[15858] = 32'b00000000000000001011101100111101;
assign LUT_1[15859] = 32'b00000000000000000100111110111001;
assign LUT_1[15860] = 32'b00000000000000010111111000000011;
assign LUT_1[15861] = 32'b00000000000000010001001001111111;
assign LUT_1[15862] = 32'b00000000000000010011100110010100;
assign LUT_1[15863] = 32'b00000000000000001100111000010000;
assign LUT_1[15864] = 32'b00000000000000001111001100100001;
assign LUT_1[15865] = 32'b00000000000000001000011110011101;
assign LUT_1[15866] = 32'b00000000000000001010111010110010;
assign LUT_1[15867] = 32'b00000000000000000100001100101110;
assign LUT_1[15868] = 32'b00000000000000010111000101111000;
assign LUT_1[15869] = 32'b00000000000000010000010111110100;
assign LUT_1[15870] = 32'b00000000000000010010110100001001;
assign LUT_1[15871] = 32'b00000000000000001100000110000101;
assign LUT_1[15872] = 32'b00000000000000000100000100110001;
assign LUT_1[15873] = 32'b11111111111111111101010110101101;
assign LUT_1[15874] = 32'b11111111111111111111110011000010;
assign LUT_1[15875] = 32'b11111111111111111001000100111110;
assign LUT_1[15876] = 32'b00000000000000001011111110001000;
assign LUT_1[15877] = 32'b00000000000000000101010000000100;
assign LUT_1[15878] = 32'b00000000000000000111101100011001;
assign LUT_1[15879] = 32'b00000000000000000000111110010101;
assign LUT_1[15880] = 32'b00000000000000000011010010100110;
assign LUT_1[15881] = 32'b11111111111111111100100100100010;
assign LUT_1[15882] = 32'b11111111111111111111000000110111;
assign LUT_1[15883] = 32'b11111111111111111000010010110011;
assign LUT_1[15884] = 32'b00000000000000001011001011111101;
assign LUT_1[15885] = 32'b00000000000000000100011101111001;
assign LUT_1[15886] = 32'b00000000000000000110111010001110;
assign LUT_1[15887] = 32'b00000000000000000000001100001010;
assign LUT_1[15888] = 32'b00000000000000000110000000010011;
assign LUT_1[15889] = 32'b11111111111111111111010010001111;
assign LUT_1[15890] = 32'b00000000000000000001101110100100;
assign LUT_1[15891] = 32'b11111111111111111011000000100000;
assign LUT_1[15892] = 32'b00000000000000001101111001101010;
assign LUT_1[15893] = 32'b00000000000000000111001011100110;
assign LUT_1[15894] = 32'b00000000000000001001100111111011;
assign LUT_1[15895] = 32'b00000000000000000010111001110111;
assign LUT_1[15896] = 32'b00000000000000000101001110001000;
assign LUT_1[15897] = 32'b11111111111111111110100000000100;
assign LUT_1[15898] = 32'b00000000000000000000111100011001;
assign LUT_1[15899] = 32'b11111111111111111010001110010101;
assign LUT_1[15900] = 32'b00000000000000001101000111011111;
assign LUT_1[15901] = 32'b00000000000000000110011001011011;
assign LUT_1[15902] = 32'b00000000000000001000110101110000;
assign LUT_1[15903] = 32'b00000000000000000010000111101100;
assign LUT_1[15904] = 32'b00000000000000000100111111110000;
assign LUT_1[15905] = 32'b11111111111111111110010001101100;
assign LUT_1[15906] = 32'b00000000000000000000101110000001;
assign LUT_1[15907] = 32'b11111111111111111001111111111101;
assign LUT_1[15908] = 32'b00000000000000001100111001000111;
assign LUT_1[15909] = 32'b00000000000000000110001011000011;
assign LUT_1[15910] = 32'b00000000000000001000100111011000;
assign LUT_1[15911] = 32'b00000000000000000001111001010100;
assign LUT_1[15912] = 32'b00000000000000000100001101100101;
assign LUT_1[15913] = 32'b11111111111111111101011111100001;
assign LUT_1[15914] = 32'b11111111111111111111111011110110;
assign LUT_1[15915] = 32'b11111111111111111001001101110010;
assign LUT_1[15916] = 32'b00000000000000001100000110111100;
assign LUT_1[15917] = 32'b00000000000000000101011000111000;
assign LUT_1[15918] = 32'b00000000000000000111110101001101;
assign LUT_1[15919] = 32'b00000000000000000001000111001001;
assign LUT_1[15920] = 32'b00000000000000000110111011010010;
assign LUT_1[15921] = 32'b00000000000000000000001101001110;
assign LUT_1[15922] = 32'b00000000000000000010101001100011;
assign LUT_1[15923] = 32'b11111111111111111011111011011111;
assign LUT_1[15924] = 32'b00000000000000001110110100101001;
assign LUT_1[15925] = 32'b00000000000000001000000110100101;
assign LUT_1[15926] = 32'b00000000000000001010100010111010;
assign LUT_1[15927] = 32'b00000000000000000011110100110110;
assign LUT_1[15928] = 32'b00000000000000000110001001000111;
assign LUT_1[15929] = 32'b11111111111111111111011011000011;
assign LUT_1[15930] = 32'b00000000000000000001110111011000;
assign LUT_1[15931] = 32'b11111111111111111011001001010100;
assign LUT_1[15932] = 32'b00000000000000001110000010011110;
assign LUT_1[15933] = 32'b00000000000000000111010100011010;
assign LUT_1[15934] = 32'b00000000000000001001110000101111;
assign LUT_1[15935] = 32'b00000000000000000011000010101011;
assign LUT_1[15936] = 32'b00000000000000000110000010011001;
assign LUT_1[15937] = 32'b11111111111111111111010100010101;
assign LUT_1[15938] = 32'b00000000000000000001110000101010;
assign LUT_1[15939] = 32'b11111111111111111011000010100110;
assign LUT_1[15940] = 32'b00000000000000001101111011110000;
assign LUT_1[15941] = 32'b00000000000000000111001101101100;
assign LUT_1[15942] = 32'b00000000000000001001101010000001;
assign LUT_1[15943] = 32'b00000000000000000010111011111101;
assign LUT_1[15944] = 32'b00000000000000000101010000001110;
assign LUT_1[15945] = 32'b11111111111111111110100010001010;
assign LUT_1[15946] = 32'b00000000000000000000111110011111;
assign LUT_1[15947] = 32'b11111111111111111010010000011011;
assign LUT_1[15948] = 32'b00000000000000001101001001100101;
assign LUT_1[15949] = 32'b00000000000000000110011011100001;
assign LUT_1[15950] = 32'b00000000000000001000110111110110;
assign LUT_1[15951] = 32'b00000000000000000010001001110010;
assign LUT_1[15952] = 32'b00000000000000000111111101111011;
assign LUT_1[15953] = 32'b00000000000000000001001111110111;
assign LUT_1[15954] = 32'b00000000000000000011101100001100;
assign LUT_1[15955] = 32'b11111111111111111100111110001000;
assign LUT_1[15956] = 32'b00000000000000001111110111010010;
assign LUT_1[15957] = 32'b00000000000000001001001001001110;
assign LUT_1[15958] = 32'b00000000000000001011100101100011;
assign LUT_1[15959] = 32'b00000000000000000100110111011111;
assign LUT_1[15960] = 32'b00000000000000000111001011110000;
assign LUT_1[15961] = 32'b00000000000000000000011101101100;
assign LUT_1[15962] = 32'b00000000000000000010111010000001;
assign LUT_1[15963] = 32'b11111111111111111100001011111101;
assign LUT_1[15964] = 32'b00000000000000001111000101000111;
assign LUT_1[15965] = 32'b00000000000000001000010111000011;
assign LUT_1[15966] = 32'b00000000000000001010110011011000;
assign LUT_1[15967] = 32'b00000000000000000100000101010100;
assign LUT_1[15968] = 32'b00000000000000000110111101011000;
assign LUT_1[15969] = 32'b00000000000000000000001111010100;
assign LUT_1[15970] = 32'b00000000000000000010101011101001;
assign LUT_1[15971] = 32'b11111111111111111011111101100101;
assign LUT_1[15972] = 32'b00000000000000001110110110101111;
assign LUT_1[15973] = 32'b00000000000000001000001000101011;
assign LUT_1[15974] = 32'b00000000000000001010100101000000;
assign LUT_1[15975] = 32'b00000000000000000011110110111100;
assign LUT_1[15976] = 32'b00000000000000000110001011001101;
assign LUT_1[15977] = 32'b11111111111111111111011101001001;
assign LUT_1[15978] = 32'b00000000000000000001111001011110;
assign LUT_1[15979] = 32'b11111111111111111011001011011010;
assign LUT_1[15980] = 32'b00000000000000001110000100100100;
assign LUT_1[15981] = 32'b00000000000000000111010110100000;
assign LUT_1[15982] = 32'b00000000000000001001110010110101;
assign LUT_1[15983] = 32'b00000000000000000011000100110001;
assign LUT_1[15984] = 32'b00000000000000001000111000111010;
assign LUT_1[15985] = 32'b00000000000000000010001010110110;
assign LUT_1[15986] = 32'b00000000000000000100100111001011;
assign LUT_1[15987] = 32'b11111111111111111101111001000111;
assign LUT_1[15988] = 32'b00000000000000010000110010010001;
assign LUT_1[15989] = 32'b00000000000000001010000100001101;
assign LUT_1[15990] = 32'b00000000000000001100100000100010;
assign LUT_1[15991] = 32'b00000000000000000101110010011110;
assign LUT_1[15992] = 32'b00000000000000001000000110101111;
assign LUT_1[15993] = 32'b00000000000000000001011000101011;
assign LUT_1[15994] = 32'b00000000000000000011110101000000;
assign LUT_1[15995] = 32'b11111111111111111101000110111100;
assign LUT_1[15996] = 32'b00000000000000010000000000000110;
assign LUT_1[15997] = 32'b00000000000000001001010010000010;
assign LUT_1[15998] = 32'b00000000000000001011101110010111;
assign LUT_1[15999] = 32'b00000000000000000101000000010011;
assign LUT_1[16000] = 32'b00000000000000000111000100110100;
assign LUT_1[16001] = 32'b00000000000000000000010110110000;
assign LUT_1[16002] = 32'b00000000000000000010110011000101;
assign LUT_1[16003] = 32'b11111111111111111100000101000001;
assign LUT_1[16004] = 32'b00000000000000001110111110001011;
assign LUT_1[16005] = 32'b00000000000000001000010000000111;
assign LUT_1[16006] = 32'b00000000000000001010101100011100;
assign LUT_1[16007] = 32'b00000000000000000011111110011000;
assign LUT_1[16008] = 32'b00000000000000000110010010101001;
assign LUT_1[16009] = 32'b11111111111111111111100100100101;
assign LUT_1[16010] = 32'b00000000000000000010000000111010;
assign LUT_1[16011] = 32'b11111111111111111011010010110110;
assign LUT_1[16012] = 32'b00000000000000001110001100000000;
assign LUT_1[16013] = 32'b00000000000000000111011101111100;
assign LUT_1[16014] = 32'b00000000000000001001111010010001;
assign LUT_1[16015] = 32'b00000000000000000011001100001101;
assign LUT_1[16016] = 32'b00000000000000001001000000010110;
assign LUT_1[16017] = 32'b00000000000000000010010010010010;
assign LUT_1[16018] = 32'b00000000000000000100101110100111;
assign LUT_1[16019] = 32'b11111111111111111110000000100011;
assign LUT_1[16020] = 32'b00000000000000010000111001101101;
assign LUT_1[16021] = 32'b00000000000000001010001011101001;
assign LUT_1[16022] = 32'b00000000000000001100100111111110;
assign LUT_1[16023] = 32'b00000000000000000101111001111010;
assign LUT_1[16024] = 32'b00000000000000001000001110001011;
assign LUT_1[16025] = 32'b00000000000000000001100000000111;
assign LUT_1[16026] = 32'b00000000000000000011111100011100;
assign LUT_1[16027] = 32'b11111111111111111101001110011000;
assign LUT_1[16028] = 32'b00000000000000010000000111100010;
assign LUT_1[16029] = 32'b00000000000000001001011001011110;
assign LUT_1[16030] = 32'b00000000000000001011110101110011;
assign LUT_1[16031] = 32'b00000000000000000101000111101111;
assign LUT_1[16032] = 32'b00000000000000000111111111110011;
assign LUT_1[16033] = 32'b00000000000000000001010001101111;
assign LUT_1[16034] = 32'b00000000000000000011101110000100;
assign LUT_1[16035] = 32'b11111111111111111101000000000000;
assign LUT_1[16036] = 32'b00000000000000001111111001001010;
assign LUT_1[16037] = 32'b00000000000000001001001011000110;
assign LUT_1[16038] = 32'b00000000000000001011100111011011;
assign LUT_1[16039] = 32'b00000000000000000100111001010111;
assign LUT_1[16040] = 32'b00000000000000000111001101101000;
assign LUT_1[16041] = 32'b00000000000000000000011111100100;
assign LUT_1[16042] = 32'b00000000000000000010111011111001;
assign LUT_1[16043] = 32'b11111111111111111100001101110101;
assign LUT_1[16044] = 32'b00000000000000001111000110111111;
assign LUT_1[16045] = 32'b00000000000000001000011000111011;
assign LUT_1[16046] = 32'b00000000000000001010110101010000;
assign LUT_1[16047] = 32'b00000000000000000100000111001100;
assign LUT_1[16048] = 32'b00000000000000001001111011010101;
assign LUT_1[16049] = 32'b00000000000000000011001101010001;
assign LUT_1[16050] = 32'b00000000000000000101101001100110;
assign LUT_1[16051] = 32'b11111111111111111110111011100010;
assign LUT_1[16052] = 32'b00000000000000010001110100101100;
assign LUT_1[16053] = 32'b00000000000000001011000110101000;
assign LUT_1[16054] = 32'b00000000000000001101100010111101;
assign LUT_1[16055] = 32'b00000000000000000110110100111001;
assign LUT_1[16056] = 32'b00000000000000001001001001001010;
assign LUT_1[16057] = 32'b00000000000000000010011011000110;
assign LUT_1[16058] = 32'b00000000000000000100110111011011;
assign LUT_1[16059] = 32'b11111111111111111110001001010111;
assign LUT_1[16060] = 32'b00000000000000010001000010100001;
assign LUT_1[16061] = 32'b00000000000000001010010100011101;
assign LUT_1[16062] = 32'b00000000000000001100110000110010;
assign LUT_1[16063] = 32'b00000000000000000110000010101110;
assign LUT_1[16064] = 32'b00000000000000001001000010011100;
assign LUT_1[16065] = 32'b00000000000000000010010100011000;
assign LUT_1[16066] = 32'b00000000000000000100110000101101;
assign LUT_1[16067] = 32'b11111111111111111110000010101001;
assign LUT_1[16068] = 32'b00000000000000010000111011110011;
assign LUT_1[16069] = 32'b00000000000000001010001101101111;
assign LUT_1[16070] = 32'b00000000000000001100101010000100;
assign LUT_1[16071] = 32'b00000000000000000101111100000000;
assign LUT_1[16072] = 32'b00000000000000001000010000010001;
assign LUT_1[16073] = 32'b00000000000000000001100010001101;
assign LUT_1[16074] = 32'b00000000000000000011111110100010;
assign LUT_1[16075] = 32'b11111111111111111101010000011110;
assign LUT_1[16076] = 32'b00000000000000010000001001101000;
assign LUT_1[16077] = 32'b00000000000000001001011011100100;
assign LUT_1[16078] = 32'b00000000000000001011110111111001;
assign LUT_1[16079] = 32'b00000000000000000101001001110101;
assign LUT_1[16080] = 32'b00000000000000001010111101111110;
assign LUT_1[16081] = 32'b00000000000000000100001111111010;
assign LUT_1[16082] = 32'b00000000000000000110101100001111;
assign LUT_1[16083] = 32'b11111111111111111111111110001011;
assign LUT_1[16084] = 32'b00000000000000010010110111010101;
assign LUT_1[16085] = 32'b00000000000000001100001001010001;
assign LUT_1[16086] = 32'b00000000000000001110100101100110;
assign LUT_1[16087] = 32'b00000000000000000111110111100010;
assign LUT_1[16088] = 32'b00000000000000001010001011110011;
assign LUT_1[16089] = 32'b00000000000000000011011101101111;
assign LUT_1[16090] = 32'b00000000000000000101111010000100;
assign LUT_1[16091] = 32'b11111111111111111111001100000000;
assign LUT_1[16092] = 32'b00000000000000010010000101001010;
assign LUT_1[16093] = 32'b00000000000000001011010111000110;
assign LUT_1[16094] = 32'b00000000000000001101110011011011;
assign LUT_1[16095] = 32'b00000000000000000111000101010111;
assign LUT_1[16096] = 32'b00000000000000001001111101011011;
assign LUT_1[16097] = 32'b00000000000000000011001111010111;
assign LUT_1[16098] = 32'b00000000000000000101101011101100;
assign LUT_1[16099] = 32'b11111111111111111110111101101000;
assign LUT_1[16100] = 32'b00000000000000010001110110110010;
assign LUT_1[16101] = 32'b00000000000000001011001000101110;
assign LUT_1[16102] = 32'b00000000000000001101100101000011;
assign LUT_1[16103] = 32'b00000000000000000110110110111111;
assign LUT_1[16104] = 32'b00000000000000001001001011010000;
assign LUT_1[16105] = 32'b00000000000000000010011101001100;
assign LUT_1[16106] = 32'b00000000000000000100111001100001;
assign LUT_1[16107] = 32'b11111111111111111110001011011101;
assign LUT_1[16108] = 32'b00000000000000010001000100100111;
assign LUT_1[16109] = 32'b00000000000000001010010110100011;
assign LUT_1[16110] = 32'b00000000000000001100110010111000;
assign LUT_1[16111] = 32'b00000000000000000110000100110100;
assign LUT_1[16112] = 32'b00000000000000001011111000111101;
assign LUT_1[16113] = 32'b00000000000000000101001010111001;
assign LUT_1[16114] = 32'b00000000000000000111100111001110;
assign LUT_1[16115] = 32'b00000000000000000000111001001010;
assign LUT_1[16116] = 32'b00000000000000010011110010010100;
assign LUT_1[16117] = 32'b00000000000000001101000100010000;
assign LUT_1[16118] = 32'b00000000000000001111100000100101;
assign LUT_1[16119] = 32'b00000000000000001000110010100001;
assign LUT_1[16120] = 32'b00000000000000001011000110110010;
assign LUT_1[16121] = 32'b00000000000000000100011000101110;
assign LUT_1[16122] = 32'b00000000000000000110110101000011;
assign LUT_1[16123] = 32'b00000000000000000000000110111111;
assign LUT_1[16124] = 32'b00000000000000010011000000001001;
assign LUT_1[16125] = 32'b00000000000000001100010010000101;
assign LUT_1[16126] = 32'b00000000000000001110101110011010;
assign LUT_1[16127] = 32'b00000000000000001000000000010110;
assign LUT_1[16128] = 32'b00000000000000000001111000111101;
assign LUT_1[16129] = 32'b11111111111111111011001010111001;
assign LUT_1[16130] = 32'b11111111111111111101100111001110;
assign LUT_1[16131] = 32'b11111111111111110110111001001010;
assign LUT_1[16132] = 32'b00000000000000001001110010010100;
assign LUT_1[16133] = 32'b00000000000000000011000100010000;
assign LUT_1[16134] = 32'b00000000000000000101100000100101;
assign LUT_1[16135] = 32'b11111111111111111110110010100001;
assign LUT_1[16136] = 32'b00000000000000000001000110110010;
assign LUT_1[16137] = 32'b11111111111111111010011000101110;
assign LUT_1[16138] = 32'b11111111111111111100110101000011;
assign LUT_1[16139] = 32'b11111111111111110110000110111111;
assign LUT_1[16140] = 32'b00000000000000001001000000001001;
assign LUT_1[16141] = 32'b00000000000000000010010010000101;
assign LUT_1[16142] = 32'b00000000000000000100101110011010;
assign LUT_1[16143] = 32'b11111111111111111110000000010110;
assign LUT_1[16144] = 32'b00000000000000000011110100011111;
assign LUT_1[16145] = 32'b11111111111111111101000110011011;
assign LUT_1[16146] = 32'b11111111111111111111100010110000;
assign LUT_1[16147] = 32'b11111111111111111000110100101100;
assign LUT_1[16148] = 32'b00000000000000001011101101110110;
assign LUT_1[16149] = 32'b00000000000000000100111111110010;
assign LUT_1[16150] = 32'b00000000000000000111011100000111;
assign LUT_1[16151] = 32'b00000000000000000000101110000011;
assign LUT_1[16152] = 32'b00000000000000000011000010010100;
assign LUT_1[16153] = 32'b11111111111111111100010100010000;
assign LUT_1[16154] = 32'b11111111111111111110110000100101;
assign LUT_1[16155] = 32'b11111111111111111000000010100001;
assign LUT_1[16156] = 32'b00000000000000001010111011101011;
assign LUT_1[16157] = 32'b00000000000000000100001101100111;
assign LUT_1[16158] = 32'b00000000000000000110101001111100;
assign LUT_1[16159] = 32'b11111111111111111111111011111000;
assign LUT_1[16160] = 32'b00000000000000000010110011111100;
assign LUT_1[16161] = 32'b11111111111111111100000101111000;
assign LUT_1[16162] = 32'b11111111111111111110100010001101;
assign LUT_1[16163] = 32'b11111111111111110111110100001001;
assign LUT_1[16164] = 32'b00000000000000001010101101010011;
assign LUT_1[16165] = 32'b00000000000000000011111111001111;
assign LUT_1[16166] = 32'b00000000000000000110011011100100;
assign LUT_1[16167] = 32'b11111111111111111111101101100000;
assign LUT_1[16168] = 32'b00000000000000000010000001110001;
assign LUT_1[16169] = 32'b11111111111111111011010011101101;
assign LUT_1[16170] = 32'b11111111111111111101110000000010;
assign LUT_1[16171] = 32'b11111111111111110111000001111110;
assign LUT_1[16172] = 32'b00000000000000001001111011001000;
assign LUT_1[16173] = 32'b00000000000000000011001101000100;
assign LUT_1[16174] = 32'b00000000000000000101101001011001;
assign LUT_1[16175] = 32'b11111111111111111110111011010101;
assign LUT_1[16176] = 32'b00000000000000000100101111011110;
assign LUT_1[16177] = 32'b11111111111111111110000001011010;
assign LUT_1[16178] = 32'b00000000000000000000011101101111;
assign LUT_1[16179] = 32'b11111111111111111001101111101011;
assign LUT_1[16180] = 32'b00000000000000001100101000110101;
assign LUT_1[16181] = 32'b00000000000000000101111010110001;
assign LUT_1[16182] = 32'b00000000000000001000010111000110;
assign LUT_1[16183] = 32'b00000000000000000001101001000010;
assign LUT_1[16184] = 32'b00000000000000000011111101010011;
assign LUT_1[16185] = 32'b11111111111111111101001111001111;
assign LUT_1[16186] = 32'b11111111111111111111101011100100;
assign LUT_1[16187] = 32'b11111111111111111000111101100000;
assign LUT_1[16188] = 32'b00000000000000001011110110101010;
assign LUT_1[16189] = 32'b00000000000000000101001000100110;
assign LUT_1[16190] = 32'b00000000000000000111100100111011;
assign LUT_1[16191] = 32'b00000000000000000000110110110111;
assign LUT_1[16192] = 32'b00000000000000000011110110100101;
assign LUT_1[16193] = 32'b11111111111111111101001000100001;
assign LUT_1[16194] = 32'b11111111111111111111100100110110;
assign LUT_1[16195] = 32'b11111111111111111000110110110010;
assign LUT_1[16196] = 32'b00000000000000001011101111111100;
assign LUT_1[16197] = 32'b00000000000000000101000001111000;
assign LUT_1[16198] = 32'b00000000000000000111011110001101;
assign LUT_1[16199] = 32'b00000000000000000000110000001001;
assign LUT_1[16200] = 32'b00000000000000000011000100011010;
assign LUT_1[16201] = 32'b11111111111111111100010110010110;
assign LUT_1[16202] = 32'b11111111111111111110110010101011;
assign LUT_1[16203] = 32'b11111111111111111000000100100111;
assign LUT_1[16204] = 32'b00000000000000001010111101110001;
assign LUT_1[16205] = 32'b00000000000000000100001111101101;
assign LUT_1[16206] = 32'b00000000000000000110101100000010;
assign LUT_1[16207] = 32'b11111111111111111111111101111110;
assign LUT_1[16208] = 32'b00000000000000000101110010000111;
assign LUT_1[16209] = 32'b11111111111111111111000100000011;
assign LUT_1[16210] = 32'b00000000000000000001100000011000;
assign LUT_1[16211] = 32'b11111111111111111010110010010100;
assign LUT_1[16212] = 32'b00000000000000001101101011011110;
assign LUT_1[16213] = 32'b00000000000000000110111101011010;
assign LUT_1[16214] = 32'b00000000000000001001011001101111;
assign LUT_1[16215] = 32'b00000000000000000010101011101011;
assign LUT_1[16216] = 32'b00000000000000000100111111111100;
assign LUT_1[16217] = 32'b11111111111111111110010001111000;
assign LUT_1[16218] = 32'b00000000000000000000101110001101;
assign LUT_1[16219] = 32'b11111111111111111010000000001001;
assign LUT_1[16220] = 32'b00000000000000001100111001010011;
assign LUT_1[16221] = 32'b00000000000000000110001011001111;
assign LUT_1[16222] = 32'b00000000000000001000100111100100;
assign LUT_1[16223] = 32'b00000000000000000001111001100000;
assign LUT_1[16224] = 32'b00000000000000000100110001100100;
assign LUT_1[16225] = 32'b11111111111111111110000011100000;
assign LUT_1[16226] = 32'b00000000000000000000011111110101;
assign LUT_1[16227] = 32'b11111111111111111001110001110001;
assign LUT_1[16228] = 32'b00000000000000001100101010111011;
assign LUT_1[16229] = 32'b00000000000000000101111100110111;
assign LUT_1[16230] = 32'b00000000000000001000011001001100;
assign LUT_1[16231] = 32'b00000000000000000001101011001000;
assign LUT_1[16232] = 32'b00000000000000000011111111011001;
assign LUT_1[16233] = 32'b11111111111111111101010001010101;
assign LUT_1[16234] = 32'b11111111111111111111101101101010;
assign LUT_1[16235] = 32'b11111111111111111000111111100110;
assign LUT_1[16236] = 32'b00000000000000001011111000110000;
assign LUT_1[16237] = 32'b00000000000000000101001010101100;
assign LUT_1[16238] = 32'b00000000000000000111100111000001;
assign LUT_1[16239] = 32'b00000000000000000000111000111101;
assign LUT_1[16240] = 32'b00000000000000000110101101000110;
assign LUT_1[16241] = 32'b11111111111111111111111111000010;
assign LUT_1[16242] = 32'b00000000000000000010011011010111;
assign LUT_1[16243] = 32'b11111111111111111011101101010011;
assign LUT_1[16244] = 32'b00000000000000001110100110011101;
assign LUT_1[16245] = 32'b00000000000000000111111000011001;
assign LUT_1[16246] = 32'b00000000000000001010010100101110;
assign LUT_1[16247] = 32'b00000000000000000011100110101010;
assign LUT_1[16248] = 32'b00000000000000000101111010111011;
assign LUT_1[16249] = 32'b11111111111111111111001100110111;
assign LUT_1[16250] = 32'b00000000000000000001101001001100;
assign LUT_1[16251] = 32'b11111111111111111010111011001000;
assign LUT_1[16252] = 32'b00000000000000001101110100010010;
assign LUT_1[16253] = 32'b00000000000000000111000110001110;
assign LUT_1[16254] = 32'b00000000000000001001100010100011;
assign LUT_1[16255] = 32'b00000000000000000010110100011111;
assign LUT_1[16256] = 32'b00000000000000000100111001000000;
assign LUT_1[16257] = 32'b11111111111111111110001010111100;
assign LUT_1[16258] = 32'b00000000000000000000100111010001;
assign LUT_1[16259] = 32'b11111111111111111001111001001101;
assign LUT_1[16260] = 32'b00000000000000001100110010010111;
assign LUT_1[16261] = 32'b00000000000000000110000100010011;
assign LUT_1[16262] = 32'b00000000000000001000100000101000;
assign LUT_1[16263] = 32'b00000000000000000001110010100100;
assign LUT_1[16264] = 32'b00000000000000000100000110110101;
assign LUT_1[16265] = 32'b11111111111111111101011000110001;
assign LUT_1[16266] = 32'b11111111111111111111110101000110;
assign LUT_1[16267] = 32'b11111111111111111001000111000010;
assign LUT_1[16268] = 32'b00000000000000001100000000001100;
assign LUT_1[16269] = 32'b00000000000000000101010010001000;
assign LUT_1[16270] = 32'b00000000000000000111101110011101;
assign LUT_1[16271] = 32'b00000000000000000001000000011001;
assign LUT_1[16272] = 32'b00000000000000000110110100100010;
assign LUT_1[16273] = 32'b00000000000000000000000110011110;
assign LUT_1[16274] = 32'b00000000000000000010100010110011;
assign LUT_1[16275] = 32'b11111111111111111011110100101111;
assign LUT_1[16276] = 32'b00000000000000001110101101111001;
assign LUT_1[16277] = 32'b00000000000000000111111111110101;
assign LUT_1[16278] = 32'b00000000000000001010011100001010;
assign LUT_1[16279] = 32'b00000000000000000011101110000110;
assign LUT_1[16280] = 32'b00000000000000000110000010010111;
assign LUT_1[16281] = 32'b11111111111111111111010100010011;
assign LUT_1[16282] = 32'b00000000000000000001110000101000;
assign LUT_1[16283] = 32'b11111111111111111011000010100100;
assign LUT_1[16284] = 32'b00000000000000001101111011101110;
assign LUT_1[16285] = 32'b00000000000000000111001101101010;
assign LUT_1[16286] = 32'b00000000000000001001101001111111;
assign LUT_1[16287] = 32'b00000000000000000010111011111011;
assign LUT_1[16288] = 32'b00000000000000000101110011111111;
assign LUT_1[16289] = 32'b11111111111111111111000101111011;
assign LUT_1[16290] = 32'b00000000000000000001100010010000;
assign LUT_1[16291] = 32'b11111111111111111010110100001100;
assign LUT_1[16292] = 32'b00000000000000001101101101010110;
assign LUT_1[16293] = 32'b00000000000000000110111111010010;
assign LUT_1[16294] = 32'b00000000000000001001011011100111;
assign LUT_1[16295] = 32'b00000000000000000010101101100011;
assign LUT_1[16296] = 32'b00000000000000000101000001110100;
assign LUT_1[16297] = 32'b11111111111111111110010011110000;
assign LUT_1[16298] = 32'b00000000000000000000110000000101;
assign LUT_1[16299] = 32'b11111111111111111010000010000001;
assign LUT_1[16300] = 32'b00000000000000001100111011001011;
assign LUT_1[16301] = 32'b00000000000000000110001101000111;
assign LUT_1[16302] = 32'b00000000000000001000101001011100;
assign LUT_1[16303] = 32'b00000000000000000001111011011000;
assign LUT_1[16304] = 32'b00000000000000000111101111100001;
assign LUT_1[16305] = 32'b00000000000000000001000001011101;
assign LUT_1[16306] = 32'b00000000000000000011011101110010;
assign LUT_1[16307] = 32'b11111111111111111100101111101110;
assign LUT_1[16308] = 32'b00000000000000001111101000111000;
assign LUT_1[16309] = 32'b00000000000000001000111010110100;
assign LUT_1[16310] = 32'b00000000000000001011010111001001;
assign LUT_1[16311] = 32'b00000000000000000100101001000101;
assign LUT_1[16312] = 32'b00000000000000000110111101010110;
assign LUT_1[16313] = 32'b00000000000000000000001111010010;
assign LUT_1[16314] = 32'b00000000000000000010101011100111;
assign LUT_1[16315] = 32'b11111111111111111011111101100011;
assign LUT_1[16316] = 32'b00000000000000001110110110101101;
assign LUT_1[16317] = 32'b00000000000000001000001000101001;
assign LUT_1[16318] = 32'b00000000000000001010100100111110;
assign LUT_1[16319] = 32'b00000000000000000011110110111010;
assign LUT_1[16320] = 32'b00000000000000000110110110101000;
assign LUT_1[16321] = 32'b00000000000000000000001000100100;
assign LUT_1[16322] = 32'b00000000000000000010100100111001;
assign LUT_1[16323] = 32'b11111111111111111011110110110101;
assign LUT_1[16324] = 32'b00000000000000001110101111111111;
assign LUT_1[16325] = 32'b00000000000000001000000001111011;
assign LUT_1[16326] = 32'b00000000000000001010011110010000;
assign LUT_1[16327] = 32'b00000000000000000011110000001100;
assign LUT_1[16328] = 32'b00000000000000000110000100011101;
assign LUT_1[16329] = 32'b11111111111111111111010110011001;
assign LUT_1[16330] = 32'b00000000000000000001110010101110;
assign LUT_1[16331] = 32'b11111111111111111011000100101010;
assign LUT_1[16332] = 32'b00000000000000001101111101110100;
assign LUT_1[16333] = 32'b00000000000000000111001111110000;
assign LUT_1[16334] = 32'b00000000000000001001101100000101;
assign LUT_1[16335] = 32'b00000000000000000010111110000001;
assign LUT_1[16336] = 32'b00000000000000001000110010001010;
assign LUT_1[16337] = 32'b00000000000000000010000100000110;
assign LUT_1[16338] = 32'b00000000000000000100100000011011;
assign LUT_1[16339] = 32'b11111111111111111101110010010111;
assign LUT_1[16340] = 32'b00000000000000010000101011100001;
assign LUT_1[16341] = 32'b00000000000000001001111101011101;
assign LUT_1[16342] = 32'b00000000000000001100011001110010;
assign LUT_1[16343] = 32'b00000000000000000101101011101110;
assign LUT_1[16344] = 32'b00000000000000000111111111111111;
assign LUT_1[16345] = 32'b00000000000000000001010001111011;
assign LUT_1[16346] = 32'b00000000000000000011101110010000;
assign LUT_1[16347] = 32'b11111111111111111101000000001100;
assign LUT_1[16348] = 32'b00000000000000001111111001010110;
assign LUT_1[16349] = 32'b00000000000000001001001011010010;
assign LUT_1[16350] = 32'b00000000000000001011100111100111;
assign LUT_1[16351] = 32'b00000000000000000100111001100011;
assign LUT_1[16352] = 32'b00000000000000000111110001100111;
assign LUT_1[16353] = 32'b00000000000000000001000011100011;
assign LUT_1[16354] = 32'b00000000000000000011011111111000;
assign LUT_1[16355] = 32'b11111111111111111100110001110100;
assign LUT_1[16356] = 32'b00000000000000001111101010111110;
assign LUT_1[16357] = 32'b00000000000000001000111100111010;
assign LUT_1[16358] = 32'b00000000000000001011011001001111;
assign LUT_1[16359] = 32'b00000000000000000100101011001011;
assign LUT_1[16360] = 32'b00000000000000000110111111011100;
assign LUT_1[16361] = 32'b00000000000000000000010001011000;
assign LUT_1[16362] = 32'b00000000000000000010101101101101;
assign LUT_1[16363] = 32'b11111111111111111011111111101001;
assign LUT_1[16364] = 32'b00000000000000001110111000110011;
assign LUT_1[16365] = 32'b00000000000000001000001010101111;
assign LUT_1[16366] = 32'b00000000000000001010100111000100;
assign LUT_1[16367] = 32'b00000000000000000011111001000000;
assign LUT_1[16368] = 32'b00000000000000001001101101001001;
assign LUT_1[16369] = 32'b00000000000000000010111111000101;
assign LUT_1[16370] = 32'b00000000000000000101011011011010;
assign LUT_1[16371] = 32'b11111111111111111110101101010110;
assign LUT_1[16372] = 32'b00000000000000010001100110100000;
assign LUT_1[16373] = 32'b00000000000000001010111000011100;
assign LUT_1[16374] = 32'b00000000000000001101010100110001;
assign LUT_1[16375] = 32'b00000000000000000110100110101101;
assign LUT_1[16376] = 32'b00000000000000001000111010111110;
assign LUT_1[16377] = 32'b00000000000000000010001100111010;
assign LUT_1[16378] = 32'b00000000000000000100101001001111;
assign LUT_1[16379] = 32'b11111111111111111101111011001011;
assign LUT_1[16380] = 32'b00000000000000010000110100010101;
assign LUT_1[16381] = 32'b00000000000000001010000110010001;
assign LUT_1[16382] = 32'b00000000000000001100100010100110;
assign LUT_1[16383] = 32'b00000000000000000101110100100010;
assign LUT_1[16384] = 32'b11111111111111111110010011111101;
assign LUT_1[16385] = 32'b11111111111111110111100101111001;
assign LUT_1[16386] = 32'b11111111111111111010000010001110;
assign LUT_1[16387] = 32'b11111111111111110011010100001010;
assign LUT_1[16388] = 32'b00000000000000000110001101010100;
assign LUT_1[16389] = 32'b11111111111111111111011111010000;
assign LUT_1[16390] = 32'b00000000000000000001111011100101;
assign LUT_1[16391] = 32'b11111111111111111011001101100001;
assign LUT_1[16392] = 32'b11111111111111111101100001110010;
assign LUT_1[16393] = 32'b11111111111111110110110011101110;
assign LUT_1[16394] = 32'b11111111111111111001010000000011;
assign LUT_1[16395] = 32'b11111111111111110010100001111111;
assign LUT_1[16396] = 32'b00000000000000000101011011001001;
assign LUT_1[16397] = 32'b11111111111111111110101101000101;
assign LUT_1[16398] = 32'b00000000000000000001001001011010;
assign LUT_1[16399] = 32'b11111111111111111010011011010110;
assign LUT_1[16400] = 32'b00000000000000000000001111011111;
assign LUT_1[16401] = 32'b11111111111111111001100001011011;
assign LUT_1[16402] = 32'b11111111111111111011111101110000;
assign LUT_1[16403] = 32'b11111111111111110101001111101100;
assign LUT_1[16404] = 32'b00000000000000001000001000110110;
assign LUT_1[16405] = 32'b00000000000000000001011010110010;
assign LUT_1[16406] = 32'b00000000000000000011110111000111;
assign LUT_1[16407] = 32'b11111111111111111101001001000011;
assign LUT_1[16408] = 32'b11111111111111111111011101010100;
assign LUT_1[16409] = 32'b11111111111111111000101111010000;
assign LUT_1[16410] = 32'b11111111111111111011001011100101;
assign LUT_1[16411] = 32'b11111111111111110100011101100001;
assign LUT_1[16412] = 32'b00000000000000000111010110101011;
assign LUT_1[16413] = 32'b00000000000000000000101000100111;
assign LUT_1[16414] = 32'b00000000000000000011000100111100;
assign LUT_1[16415] = 32'b11111111111111111100010110111000;
assign LUT_1[16416] = 32'b11111111111111111111001110111100;
assign LUT_1[16417] = 32'b11111111111111111000100000111000;
assign LUT_1[16418] = 32'b11111111111111111010111101001101;
assign LUT_1[16419] = 32'b11111111111111110100001111001001;
assign LUT_1[16420] = 32'b00000000000000000111001000010011;
assign LUT_1[16421] = 32'b00000000000000000000011010001111;
assign LUT_1[16422] = 32'b00000000000000000010110110100100;
assign LUT_1[16423] = 32'b11111111111111111100001000100000;
assign LUT_1[16424] = 32'b11111111111111111110011100110001;
assign LUT_1[16425] = 32'b11111111111111110111101110101101;
assign LUT_1[16426] = 32'b11111111111111111010001011000010;
assign LUT_1[16427] = 32'b11111111111111110011011100111110;
assign LUT_1[16428] = 32'b00000000000000000110010110001000;
assign LUT_1[16429] = 32'b11111111111111111111101000000100;
assign LUT_1[16430] = 32'b00000000000000000010000100011001;
assign LUT_1[16431] = 32'b11111111111111111011010110010101;
assign LUT_1[16432] = 32'b00000000000000000001001010011110;
assign LUT_1[16433] = 32'b11111111111111111010011100011010;
assign LUT_1[16434] = 32'b11111111111111111100111000101111;
assign LUT_1[16435] = 32'b11111111111111110110001010101011;
assign LUT_1[16436] = 32'b00000000000000001001000011110101;
assign LUT_1[16437] = 32'b00000000000000000010010101110001;
assign LUT_1[16438] = 32'b00000000000000000100110010000110;
assign LUT_1[16439] = 32'b11111111111111111110000100000010;
assign LUT_1[16440] = 32'b00000000000000000000011000010011;
assign LUT_1[16441] = 32'b11111111111111111001101010001111;
assign LUT_1[16442] = 32'b11111111111111111100000110100100;
assign LUT_1[16443] = 32'b11111111111111110101011000100000;
assign LUT_1[16444] = 32'b00000000000000001000010001101010;
assign LUT_1[16445] = 32'b00000000000000000001100011100110;
assign LUT_1[16446] = 32'b00000000000000000011111111111011;
assign LUT_1[16447] = 32'b11111111111111111101010001110111;
assign LUT_1[16448] = 32'b00000000000000000000010001100101;
assign LUT_1[16449] = 32'b11111111111111111001100011100001;
assign LUT_1[16450] = 32'b11111111111111111011111111110110;
assign LUT_1[16451] = 32'b11111111111111110101010001110010;
assign LUT_1[16452] = 32'b00000000000000001000001010111100;
assign LUT_1[16453] = 32'b00000000000000000001011100111000;
assign LUT_1[16454] = 32'b00000000000000000011111001001101;
assign LUT_1[16455] = 32'b11111111111111111101001011001001;
assign LUT_1[16456] = 32'b11111111111111111111011111011010;
assign LUT_1[16457] = 32'b11111111111111111000110001010110;
assign LUT_1[16458] = 32'b11111111111111111011001101101011;
assign LUT_1[16459] = 32'b11111111111111110100011111100111;
assign LUT_1[16460] = 32'b00000000000000000111011000110001;
assign LUT_1[16461] = 32'b00000000000000000000101010101101;
assign LUT_1[16462] = 32'b00000000000000000011000111000010;
assign LUT_1[16463] = 32'b11111111111111111100011000111110;
assign LUT_1[16464] = 32'b00000000000000000010001101000111;
assign LUT_1[16465] = 32'b11111111111111111011011111000011;
assign LUT_1[16466] = 32'b11111111111111111101111011011000;
assign LUT_1[16467] = 32'b11111111111111110111001101010100;
assign LUT_1[16468] = 32'b00000000000000001010000110011110;
assign LUT_1[16469] = 32'b00000000000000000011011000011010;
assign LUT_1[16470] = 32'b00000000000000000101110100101111;
assign LUT_1[16471] = 32'b11111111111111111111000110101011;
assign LUT_1[16472] = 32'b00000000000000000001011010111100;
assign LUT_1[16473] = 32'b11111111111111111010101100111000;
assign LUT_1[16474] = 32'b11111111111111111101001001001101;
assign LUT_1[16475] = 32'b11111111111111110110011011001001;
assign LUT_1[16476] = 32'b00000000000000001001010100010011;
assign LUT_1[16477] = 32'b00000000000000000010100110001111;
assign LUT_1[16478] = 32'b00000000000000000101000010100100;
assign LUT_1[16479] = 32'b11111111111111111110010100100000;
assign LUT_1[16480] = 32'b00000000000000000001001100100100;
assign LUT_1[16481] = 32'b11111111111111111010011110100000;
assign LUT_1[16482] = 32'b11111111111111111100111010110101;
assign LUT_1[16483] = 32'b11111111111111110110001100110001;
assign LUT_1[16484] = 32'b00000000000000001001000101111011;
assign LUT_1[16485] = 32'b00000000000000000010010111110111;
assign LUT_1[16486] = 32'b00000000000000000100110100001100;
assign LUT_1[16487] = 32'b11111111111111111110000110001000;
assign LUT_1[16488] = 32'b00000000000000000000011010011001;
assign LUT_1[16489] = 32'b11111111111111111001101100010101;
assign LUT_1[16490] = 32'b11111111111111111100001000101010;
assign LUT_1[16491] = 32'b11111111111111110101011010100110;
assign LUT_1[16492] = 32'b00000000000000001000010011110000;
assign LUT_1[16493] = 32'b00000000000000000001100101101100;
assign LUT_1[16494] = 32'b00000000000000000100000010000001;
assign LUT_1[16495] = 32'b11111111111111111101010011111101;
assign LUT_1[16496] = 32'b00000000000000000011001000000110;
assign LUT_1[16497] = 32'b11111111111111111100011010000010;
assign LUT_1[16498] = 32'b11111111111111111110110110010111;
assign LUT_1[16499] = 32'b11111111111111111000001000010011;
assign LUT_1[16500] = 32'b00000000000000001011000001011101;
assign LUT_1[16501] = 32'b00000000000000000100010011011001;
assign LUT_1[16502] = 32'b00000000000000000110101111101110;
assign LUT_1[16503] = 32'b00000000000000000000000001101010;
assign LUT_1[16504] = 32'b00000000000000000010010101111011;
assign LUT_1[16505] = 32'b11111111111111111011100111110111;
assign LUT_1[16506] = 32'b11111111111111111110000100001100;
assign LUT_1[16507] = 32'b11111111111111110111010110001000;
assign LUT_1[16508] = 32'b00000000000000001010001111010010;
assign LUT_1[16509] = 32'b00000000000000000011100001001110;
assign LUT_1[16510] = 32'b00000000000000000101111101100011;
assign LUT_1[16511] = 32'b11111111111111111111001111011111;
assign LUT_1[16512] = 32'b00000000000000000001010100000000;
assign LUT_1[16513] = 32'b11111111111111111010100101111100;
assign LUT_1[16514] = 32'b11111111111111111101000010010001;
assign LUT_1[16515] = 32'b11111111111111110110010100001101;
assign LUT_1[16516] = 32'b00000000000000001001001101010111;
assign LUT_1[16517] = 32'b00000000000000000010011111010011;
assign LUT_1[16518] = 32'b00000000000000000100111011101000;
assign LUT_1[16519] = 32'b11111111111111111110001101100100;
assign LUT_1[16520] = 32'b00000000000000000000100001110101;
assign LUT_1[16521] = 32'b11111111111111111001110011110001;
assign LUT_1[16522] = 32'b11111111111111111100010000000110;
assign LUT_1[16523] = 32'b11111111111111110101100010000010;
assign LUT_1[16524] = 32'b00000000000000001000011011001100;
assign LUT_1[16525] = 32'b00000000000000000001101101001000;
assign LUT_1[16526] = 32'b00000000000000000100001001011101;
assign LUT_1[16527] = 32'b11111111111111111101011011011001;
assign LUT_1[16528] = 32'b00000000000000000011001111100010;
assign LUT_1[16529] = 32'b11111111111111111100100001011110;
assign LUT_1[16530] = 32'b11111111111111111110111101110011;
assign LUT_1[16531] = 32'b11111111111111111000001111101111;
assign LUT_1[16532] = 32'b00000000000000001011001000111001;
assign LUT_1[16533] = 32'b00000000000000000100011010110101;
assign LUT_1[16534] = 32'b00000000000000000110110111001010;
assign LUT_1[16535] = 32'b00000000000000000000001001000110;
assign LUT_1[16536] = 32'b00000000000000000010011101010111;
assign LUT_1[16537] = 32'b11111111111111111011101111010011;
assign LUT_1[16538] = 32'b11111111111111111110001011101000;
assign LUT_1[16539] = 32'b11111111111111110111011101100100;
assign LUT_1[16540] = 32'b00000000000000001010010110101110;
assign LUT_1[16541] = 32'b00000000000000000011101000101010;
assign LUT_1[16542] = 32'b00000000000000000110000100111111;
assign LUT_1[16543] = 32'b11111111111111111111010110111011;
assign LUT_1[16544] = 32'b00000000000000000010001110111111;
assign LUT_1[16545] = 32'b11111111111111111011100000111011;
assign LUT_1[16546] = 32'b11111111111111111101111101010000;
assign LUT_1[16547] = 32'b11111111111111110111001111001100;
assign LUT_1[16548] = 32'b00000000000000001010001000010110;
assign LUT_1[16549] = 32'b00000000000000000011011010010010;
assign LUT_1[16550] = 32'b00000000000000000101110110100111;
assign LUT_1[16551] = 32'b11111111111111111111001000100011;
assign LUT_1[16552] = 32'b00000000000000000001011100110100;
assign LUT_1[16553] = 32'b11111111111111111010101110110000;
assign LUT_1[16554] = 32'b11111111111111111101001011000101;
assign LUT_1[16555] = 32'b11111111111111110110011101000001;
assign LUT_1[16556] = 32'b00000000000000001001010110001011;
assign LUT_1[16557] = 32'b00000000000000000010101000000111;
assign LUT_1[16558] = 32'b00000000000000000101000100011100;
assign LUT_1[16559] = 32'b11111111111111111110010110011000;
assign LUT_1[16560] = 32'b00000000000000000100001010100001;
assign LUT_1[16561] = 32'b11111111111111111101011100011101;
assign LUT_1[16562] = 32'b11111111111111111111111000110010;
assign LUT_1[16563] = 32'b11111111111111111001001010101110;
assign LUT_1[16564] = 32'b00000000000000001100000011111000;
assign LUT_1[16565] = 32'b00000000000000000101010101110100;
assign LUT_1[16566] = 32'b00000000000000000111110010001001;
assign LUT_1[16567] = 32'b00000000000000000001000100000101;
assign LUT_1[16568] = 32'b00000000000000000011011000010110;
assign LUT_1[16569] = 32'b11111111111111111100101010010010;
assign LUT_1[16570] = 32'b11111111111111111111000110100111;
assign LUT_1[16571] = 32'b11111111111111111000011000100011;
assign LUT_1[16572] = 32'b00000000000000001011010001101101;
assign LUT_1[16573] = 32'b00000000000000000100100011101001;
assign LUT_1[16574] = 32'b00000000000000000110111111111110;
assign LUT_1[16575] = 32'b00000000000000000000010001111010;
assign LUT_1[16576] = 32'b00000000000000000011010001101000;
assign LUT_1[16577] = 32'b11111111111111111100100011100100;
assign LUT_1[16578] = 32'b11111111111111111110111111111001;
assign LUT_1[16579] = 32'b11111111111111111000010001110101;
assign LUT_1[16580] = 32'b00000000000000001011001010111111;
assign LUT_1[16581] = 32'b00000000000000000100011100111011;
assign LUT_1[16582] = 32'b00000000000000000110111001010000;
assign LUT_1[16583] = 32'b00000000000000000000001011001100;
assign LUT_1[16584] = 32'b00000000000000000010011111011101;
assign LUT_1[16585] = 32'b11111111111111111011110001011001;
assign LUT_1[16586] = 32'b11111111111111111110001101101110;
assign LUT_1[16587] = 32'b11111111111111110111011111101010;
assign LUT_1[16588] = 32'b00000000000000001010011000110100;
assign LUT_1[16589] = 32'b00000000000000000011101010110000;
assign LUT_1[16590] = 32'b00000000000000000110000111000101;
assign LUT_1[16591] = 32'b11111111111111111111011001000001;
assign LUT_1[16592] = 32'b00000000000000000101001101001010;
assign LUT_1[16593] = 32'b11111111111111111110011111000110;
assign LUT_1[16594] = 32'b00000000000000000000111011011011;
assign LUT_1[16595] = 32'b11111111111111111010001101010111;
assign LUT_1[16596] = 32'b00000000000000001101000110100001;
assign LUT_1[16597] = 32'b00000000000000000110011000011101;
assign LUT_1[16598] = 32'b00000000000000001000110100110010;
assign LUT_1[16599] = 32'b00000000000000000010000110101110;
assign LUT_1[16600] = 32'b00000000000000000100011010111111;
assign LUT_1[16601] = 32'b11111111111111111101101100111011;
assign LUT_1[16602] = 32'b00000000000000000000001001010000;
assign LUT_1[16603] = 32'b11111111111111111001011011001100;
assign LUT_1[16604] = 32'b00000000000000001100010100010110;
assign LUT_1[16605] = 32'b00000000000000000101100110010010;
assign LUT_1[16606] = 32'b00000000000000001000000010100111;
assign LUT_1[16607] = 32'b00000000000000000001010100100011;
assign LUT_1[16608] = 32'b00000000000000000100001100100111;
assign LUT_1[16609] = 32'b11111111111111111101011110100011;
assign LUT_1[16610] = 32'b11111111111111111111111010111000;
assign LUT_1[16611] = 32'b11111111111111111001001100110100;
assign LUT_1[16612] = 32'b00000000000000001100000101111110;
assign LUT_1[16613] = 32'b00000000000000000101010111111010;
assign LUT_1[16614] = 32'b00000000000000000111110100001111;
assign LUT_1[16615] = 32'b00000000000000000001000110001011;
assign LUT_1[16616] = 32'b00000000000000000011011010011100;
assign LUT_1[16617] = 32'b11111111111111111100101100011000;
assign LUT_1[16618] = 32'b11111111111111111111001000101101;
assign LUT_1[16619] = 32'b11111111111111111000011010101001;
assign LUT_1[16620] = 32'b00000000000000001011010011110011;
assign LUT_1[16621] = 32'b00000000000000000100100101101111;
assign LUT_1[16622] = 32'b00000000000000000111000010000100;
assign LUT_1[16623] = 32'b00000000000000000000010100000000;
assign LUT_1[16624] = 32'b00000000000000000110001000001001;
assign LUT_1[16625] = 32'b11111111111111111111011010000101;
assign LUT_1[16626] = 32'b00000000000000000001110110011010;
assign LUT_1[16627] = 32'b11111111111111111011001000010110;
assign LUT_1[16628] = 32'b00000000000000001110000001100000;
assign LUT_1[16629] = 32'b00000000000000000111010011011100;
assign LUT_1[16630] = 32'b00000000000000001001101111110001;
assign LUT_1[16631] = 32'b00000000000000000011000001101101;
assign LUT_1[16632] = 32'b00000000000000000101010101111110;
assign LUT_1[16633] = 32'b11111111111111111110100111111010;
assign LUT_1[16634] = 32'b00000000000000000001000100001111;
assign LUT_1[16635] = 32'b11111111111111111010010110001011;
assign LUT_1[16636] = 32'b00000000000000001101001111010101;
assign LUT_1[16637] = 32'b00000000000000000110100001010001;
assign LUT_1[16638] = 32'b00000000000000001000111101100110;
assign LUT_1[16639] = 32'b00000000000000000010001111100010;
assign LUT_1[16640] = 32'b11111111111111111100001000001001;
assign LUT_1[16641] = 32'b11111111111111110101011010000101;
assign LUT_1[16642] = 32'b11111111111111110111110110011010;
assign LUT_1[16643] = 32'b11111111111111110001001000010110;
assign LUT_1[16644] = 32'b00000000000000000100000001100000;
assign LUT_1[16645] = 32'b11111111111111111101010011011100;
assign LUT_1[16646] = 32'b11111111111111111111101111110001;
assign LUT_1[16647] = 32'b11111111111111111001000001101101;
assign LUT_1[16648] = 32'b11111111111111111011010101111110;
assign LUT_1[16649] = 32'b11111111111111110100100111111010;
assign LUT_1[16650] = 32'b11111111111111110111000100001111;
assign LUT_1[16651] = 32'b11111111111111110000010110001011;
assign LUT_1[16652] = 32'b00000000000000000011001111010101;
assign LUT_1[16653] = 32'b11111111111111111100100001010001;
assign LUT_1[16654] = 32'b11111111111111111110111101100110;
assign LUT_1[16655] = 32'b11111111111111111000001111100010;
assign LUT_1[16656] = 32'b11111111111111111110000011101011;
assign LUT_1[16657] = 32'b11111111111111110111010101100111;
assign LUT_1[16658] = 32'b11111111111111111001110001111100;
assign LUT_1[16659] = 32'b11111111111111110011000011111000;
assign LUT_1[16660] = 32'b00000000000000000101111101000010;
assign LUT_1[16661] = 32'b11111111111111111111001110111110;
assign LUT_1[16662] = 32'b00000000000000000001101011010011;
assign LUT_1[16663] = 32'b11111111111111111010111101001111;
assign LUT_1[16664] = 32'b11111111111111111101010001100000;
assign LUT_1[16665] = 32'b11111111111111110110100011011100;
assign LUT_1[16666] = 32'b11111111111111111000111111110001;
assign LUT_1[16667] = 32'b11111111111111110010010001101101;
assign LUT_1[16668] = 32'b00000000000000000101001010110111;
assign LUT_1[16669] = 32'b11111111111111111110011100110011;
assign LUT_1[16670] = 32'b00000000000000000000111001001000;
assign LUT_1[16671] = 32'b11111111111111111010001011000100;
assign LUT_1[16672] = 32'b11111111111111111101000011001000;
assign LUT_1[16673] = 32'b11111111111111110110010101000100;
assign LUT_1[16674] = 32'b11111111111111111000110001011001;
assign LUT_1[16675] = 32'b11111111111111110010000011010101;
assign LUT_1[16676] = 32'b00000000000000000100111100011111;
assign LUT_1[16677] = 32'b11111111111111111110001110011011;
assign LUT_1[16678] = 32'b00000000000000000000101010110000;
assign LUT_1[16679] = 32'b11111111111111111001111100101100;
assign LUT_1[16680] = 32'b11111111111111111100010000111101;
assign LUT_1[16681] = 32'b11111111111111110101100010111001;
assign LUT_1[16682] = 32'b11111111111111110111111111001110;
assign LUT_1[16683] = 32'b11111111111111110001010001001010;
assign LUT_1[16684] = 32'b00000000000000000100001010010100;
assign LUT_1[16685] = 32'b11111111111111111101011100010000;
assign LUT_1[16686] = 32'b11111111111111111111111000100101;
assign LUT_1[16687] = 32'b11111111111111111001001010100001;
assign LUT_1[16688] = 32'b11111111111111111110111110101010;
assign LUT_1[16689] = 32'b11111111111111111000010000100110;
assign LUT_1[16690] = 32'b11111111111111111010101100111011;
assign LUT_1[16691] = 32'b11111111111111110011111110110111;
assign LUT_1[16692] = 32'b00000000000000000110111000000001;
assign LUT_1[16693] = 32'b00000000000000000000001001111101;
assign LUT_1[16694] = 32'b00000000000000000010100110010010;
assign LUT_1[16695] = 32'b11111111111111111011111000001110;
assign LUT_1[16696] = 32'b11111111111111111110001100011111;
assign LUT_1[16697] = 32'b11111111111111110111011110011011;
assign LUT_1[16698] = 32'b11111111111111111001111010110000;
assign LUT_1[16699] = 32'b11111111111111110011001100101100;
assign LUT_1[16700] = 32'b00000000000000000110000101110110;
assign LUT_1[16701] = 32'b11111111111111111111010111110010;
assign LUT_1[16702] = 32'b00000000000000000001110100000111;
assign LUT_1[16703] = 32'b11111111111111111011000110000011;
assign LUT_1[16704] = 32'b11111111111111111110000101110001;
assign LUT_1[16705] = 32'b11111111111111110111010111101101;
assign LUT_1[16706] = 32'b11111111111111111001110100000010;
assign LUT_1[16707] = 32'b11111111111111110011000101111110;
assign LUT_1[16708] = 32'b00000000000000000101111111001000;
assign LUT_1[16709] = 32'b11111111111111111111010001000100;
assign LUT_1[16710] = 32'b00000000000000000001101101011001;
assign LUT_1[16711] = 32'b11111111111111111010111111010101;
assign LUT_1[16712] = 32'b11111111111111111101010011100110;
assign LUT_1[16713] = 32'b11111111111111110110100101100010;
assign LUT_1[16714] = 32'b11111111111111111001000001110111;
assign LUT_1[16715] = 32'b11111111111111110010010011110011;
assign LUT_1[16716] = 32'b00000000000000000101001100111101;
assign LUT_1[16717] = 32'b11111111111111111110011110111001;
assign LUT_1[16718] = 32'b00000000000000000000111011001110;
assign LUT_1[16719] = 32'b11111111111111111010001101001010;
assign LUT_1[16720] = 32'b00000000000000000000000001010011;
assign LUT_1[16721] = 32'b11111111111111111001010011001111;
assign LUT_1[16722] = 32'b11111111111111111011101111100100;
assign LUT_1[16723] = 32'b11111111111111110101000001100000;
assign LUT_1[16724] = 32'b00000000000000000111111010101010;
assign LUT_1[16725] = 32'b00000000000000000001001100100110;
assign LUT_1[16726] = 32'b00000000000000000011101000111011;
assign LUT_1[16727] = 32'b11111111111111111100111010110111;
assign LUT_1[16728] = 32'b11111111111111111111001111001000;
assign LUT_1[16729] = 32'b11111111111111111000100001000100;
assign LUT_1[16730] = 32'b11111111111111111010111101011001;
assign LUT_1[16731] = 32'b11111111111111110100001111010101;
assign LUT_1[16732] = 32'b00000000000000000111001000011111;
assign LUT_1[16733] = 32'b00000000000000000000011010011011;
assign LUT_1[16734] = 32'b00000000000000000010110110110000;
assign LUT_1[16735] = 32'b11111111111111111100001000101100;
assign LUT_1[16736] = 32'b11111111111111111111000000110000;
assign LUT_1[16737] = 32'b11111111111111111000010010101100;
assign LUT_1[16738] = 32'b11111111111111111010101111000001;
assign LUT_1[16739] = 32'b11111111111111110100000000111101;
assign LUT_1[16740] = 32'b00000000000000000110111010000111;
assign LUT_1[16741] = 32'b00000000000000000000001100000011;
assign LUT_1[16742] = 32'b00000000000000000010101000011000;
assign LUT_1[16743] = 32'b11111111111111111011111010010100;
assign LUT_1[16744] = 32'b11111111111111111110001110100101;
assign LUT_1[16745] = 32'b11111111111111110111100000100001;
assign LUT_1[16746] = 32'b11111111111111111001111100110110;
assign LUT_1[16747] = 32'b11111111111111110011001110110010;
assign LUT_1[16748] = 32'b00000000000000000110000111111100;
assign LUT_1[16749] = 32'b11111111111111111111011001111000;
assign LUT_1[16750] = 32'b00000000000000000001110110001101;
assign LUT_1[16751] = 32'b11111111111111111011001000001001;
assign LUT_1[16752] = 32'b00000000000000000000111100010010;
assign LUT_1[16753] = 32'b11111111111111111010001110001110;
assign LUT_1[16754] = 32'b11111111111111111100101010100011;
assign LUT_1[16755] = 32'b11111111111111110101111100011111;
assign LUT_1[16756] = 32'b00000000000000001000110101101001;
assign LUT_1[16757] = 32'b00000000000000000010000111100101;
assign LUT_1[16758] = 32'b00000000000000000100100011111010;
assign LUT_1[16759] = 32'b11111111111111111101110101110110;
assign LUT_1[16760] = 32'b00000000000000000000001010000111;
assign LUT_1[16761] = 32'b11111111111111111001011100000011;
assign LUT_1[16762] = 32'b11111111111111111011111000011000;
assign LUT_1[16763] = 32'b11111111111111110101001010010100;
assign LUT_1[16764] = 32'b00000000000000001000000011011110;
assign LUT_1[16765] = 32'b00000000000000000001010101011010;
assign LUT_1[16766] = 32'b00000000000000000011110001101111;
assign LUT_1[16767] = 32'b11111111111111111101000011101011;
assign LUT_1[16768] = 32'b11111111111111111111001000001100;
assign LUT_1[16769] = 32'b11111111111111111000011010001000;
assign LUT_1[16770] = 32'b11111111111111111010110110011101;
assign LUT_1[16771] = 32'b11111111111111110100001000011001;
assign LUT_1[16772] = 32'b00000000000000000111000001100011;
assign LUT_1[16773] = 32'b00000000000000000000010011011111;
assign LUT_1[16774] = 32'b00000000000000000010101111110100;
assign LUT_1[16775] = 32'b11111111111111111100000001110000;
assign LUT_1[16776] = 32'b11111111111111111110010110000001;
assign LUT_1[16777] = 32'b11111111111111110111100111111101;
assign LUT_1[16778] = 32'b11111111111111111010000100010010;
assign LUT_1[16779] = 32'b11111111111111110011010110001110;
assign LUT_1[16780] = 32'b00000000000000000110001111011000;
assign LUT_1[16781] = 32'b11111111111111111111100001010100;
assign LUT_1[16782] = 32'b00000000000000000001111101101001;
assign LUT_1[16783] = 32'b11111111111111111011001111100101;
assign LUT_1[16784] = 32'b00000000000000000001000011101110;
assign LUT_1[16785] = 32'b11111111111111111010010101101010;
assign LUT_1[16786] = 32'b11111111111111111100110001111111;
assign LUT_1[16787] = 32'b11111111111111110110000011111011;
assign LUT_1[16788] = 32'b00000000000000001000111101000101;
assign LUT_1[16789] = 32'b00000000000000000010001111000001;
assign LUT_1[16790] = 32'b00000000000000000100101011010110;
assign LUT_1[16791] = 32'b11111111111111111101111101010010;
assign LUT_1[16792] = 32'b00000000000000000000010001100011;
assign LUT_1[16793] = 32'b11111111111111111001100011011111;
assign LUT_1[16794] = 32'b11111111111111111011111111110100;
assign LUT_1[16795] = 32'b11111111111111110101010001110000;
assign LUT_1[16796] = 32'b00000000000000001000001010111010;
assign LUT_1[16797] = 32'b00000000000000000001011100110110;
assign LUT_1[16798] = 32'b00000000000000000011111001001011;
assign LUT_1[16799] = 32'b11111111111111111101001011000111;
assign LUT_1[16800] = 32'b00000000000000000000000011001011;
assign LUT_1[16801] = 32'b11111111111111111001010101000111;
assign LUT_1[16802] = 32'b11111111111111111011110001011100;
assign LUT_1[16803] = 32'b11111111111111110101000011011000;
assign LUT_1[16804] = 32'b00000000000000000111111100100010;
assign LUT_1[16805] = 32'b00000000000000000001001110011110;
assign LUT_1[16806] = 32'b00000000000000000011101010110011;
assign LUT_1[16807] = 32'b11111111111111111100111100101111;
assign LUT_1[16808] = 32'b11111111111111111111010001000000;
assign LUT_1[16809] = 32'b11111111111111111000100010111100;
assign LUT_1[16810] = 32'b11111111111111111010111111010001;
assign LUT_1[16811] = 32'b11111111111111110100010001001101;
assign LUT_1[16812] = 32'b00000000000000000111001010010111;
assign LUT_1[16813] = 32'b00000000000000000000011100010011;
assign LUT_1[16814] = 32'b00000000000000000010111000101000;
assign LUT_1[16815] = 32'b11111111111111111100001010100100;
assign LUT_1[16816] = 32'b00000000000000000001111110101101;
assign LUT_1[16817] = 32'b11111111111111111011010000101001;
assign LUT_1[16818] = 32'b11111111111111111101101100111110;
assign LUT_1[16819] = 32'b11111111111111110110111110111010;
assign LUT_1[16820] = 32'b00000000000000001001111000000100;
assign LUT_1[16821] = 32'b00000000000000000011001010000000;
assign LUT_1[16822] = 32'b00000000000000000101100110010101;
assign LUT_1[16823] = 32'b11111111111111111110111000010001;
assign LUT_1[16824] = 32'b00000000000000000001001100100010;
assign LUT_1[16825] = 32'b11111111111111111010011110011110;
assign LUT_1[16826] = 32'b11111111111111111100111010110011;
assign LUT_1[16827] = 32'b11111111111111110110001100101111;
assign LUT_1[16828] = 32'b00000000000000001001000101111001;
assign LUT_1[16829] = 32'b00000000000000000010010111110101;
assign LUT_1[16830] = 32'b00000000000000000100110100001010;
assign LUT_1[16831] = 32'b11111111111111111110000110000110;
assign LUT_1[16832] = 32'b00000000000000000001000101110100;
assign LUT_1[16833] = 32'b11111111111111111010010111110000;
assign LUT_1[16834] = 32'b11111111111111111100110100000101;
assign LUT_1[16835] = 32'b11111111111111110110000110000001;
assign LUT_1[16836] = 32'b00000000000000001000111111001011;
assign LUT_1[16837] = 32'b00000000000000000010010001000111;
assign LUT_1[16838] = 32'b00000000000000000100101101011100;
assign LUT_1[16839] = 32'b11111111111111111101111111011000;
assign LUT_1[16840] = 32'b00000000000000000000010011101001;
assign LUT_1[16841] = 32'b11111111111111111001100101100101;
assign LUT_1[16842] = 32'b11111111111111111100000001111010;
assign LUT_1[16843] = 32'b11111111111111110101010011110110;
assign LUT_1[16844] = 32'b00000000000000001000001101000000;
assign LUT_1[16845] = 32'b00000000000000000001011110111100;
assign LUT_1[16846] = 32'b00000000000000000011111011010001;
assign LUT_1[16847] = 32'b11111111111111111101001101001101;
assign LUT_1[16848] = 32'b00000000000000000011000001010110;
assign LUT_1[16849] = 32'b11111111111111111100010011010010;
assign LUT_1[16850] = 32'b11111111111111111110101111100111;
assign LUT_1[16851] = 32'b11111111111111111000000001100011;
assign LUT_1[16852] = 32'b00000000000000001010111010101101;
assign LUT_1[16853] = 32'b00000000000000000100001100101001;
assign LUT_1[16854] = 32'b00000000000000000110101000111110;
assign LUT_1[16855] = 32'b11111111111111111111111010111010;
assign LUT_1[16856] = 32'b00000000000000000010001111001011;
assign LUT_1[16857] = 32'b11111111111111111011100001000111;
assign LUT_1[16858] = 32'b11111111111111111101111101011100;
assign LUT_1[16859] = 32'b11111111111111110111001111011000;
assign LUT_1[16860] = 32'b00000000000000001010001000100010;
assign LUT_1[16861] = 32'b00000000000000000011011010011110;
assign LUT_1[16862] = 32'b00000000000000000101110110110011;
assign LUT_1[16863] = 32'b11111111111111111111001000101111;
assign LUT_1[16864] = 32'b00000000000000000010000000110011;
assign LUT_1[16865] = 32'b11111111111111111011010010101111;
assign LUT_1[16866] = 32'b11111111111111111101101111000100;
assign LUT_1[16867] = 32'b11111111111111110111000001000000;
assign LUT_1[16868] = 32'b00000000000000001001111010001010;
assign LUT_1[16869] = 32'b00000000000000000011001100000110;
assign LUT_1[16870] = 32'b00000000000000000101101000011011;
assign LUT_1[16871] = 32'b11111111111111111110111010010111;
assign LUT_1[16872] = 32'b00000000000000000001001110101000;
assign LUT_1[16873] = 32'b11111111111111111010100000100100;
assign LUT_1[16874] = 32'b11111111111111111100111100111001;
assign LUT_1[16875] = 32'b11111111111111110110001110110101;
assign LUT_1[16876] = 32'b00000000000000001001000111111111;
assign LUT_1[16877] = 32'b00000000000000000010011001111011;
assign LUT_1[16878] = 32'b00000000000000000100110110010000;
assign LUT_1[16879] = 32'b11111111111111111110001000001100;
assign LUT_1[16880] = 32'b00000000000000000011111100010101;
assign LUT_1[16881] = 32'b11111111111111111101001110010001;
assign LUT_1[16882] = 32'b11111111111111111111101010100110;
assign LUT_1[16883] = 32'b11111111111111111000111100100010;
assign LUT_1[16884] = 32'b00000000000000001011110101101100;
assign LUT_1[16885] = 32'b00000000000000000101000111101000;
assign LUT_1[16886] = 32'b00000000000000000111100011111101;
assign LUT_1[16887] = 32'b00000000000000000000110101111001;
assign LUT_1[16888] = 32'b00000000000000000011001010001010;
assign LUT_1[16889] = 32'b11111111111111111100011100000110;
assign LUT_1[16890] = 32'b11111111111111111110111000011011;
assign LUT_1[16891] = 32'b11111111111111111000001010010111;
assign LUT_1[16892] = 32'b00000000000000001011000011100001;
assign LUT_1[16893] = 32'b00000000000000000100010101011101;
assign LUT_1[16894] = 32'b00000000000000000110110001110010;
assign LUT_1[16895] = 32'b00000000000000000000000011101110;
assign LUT_1[16896] = 32'b11111111111111111000000010011010;
assign LUT_1[16897] = 32'b11111111111111110001010100010110;
assign LUT_1[16898] = 32'b11111111111111110011110000101011;
assign LUT_1[16899] = 32'b11111111111111101101000010100111;
assign LUT_1[16900] = 32'b11111111111111111111111011110001;
assign LUT_1[16901] = 32'b11111111111111111001001101101101;
assign LUT_1[16902] = 32'b11111111111111111011101010000010;
assign LUT_1[16903] = 32'b11111111111111110100111011111110;
assign LUT_1[16904] = 32'b11111111111111110111010000001111;
assign LUT_1[16905] = 32'b11111111111111110000100010001011;
assign LUT_1[16906] = 32'b11111111111111110010111110100000;
assign LUT_1[16907] = 32'b11111111111111101100010000011100;
assign LUT_1[16908] = 32'b11111111111111111111001001100110;
assign LUT_1[16909] = 32'b11111111111111111000011011100010;
assign LUT_1[16910] = 32'b11111111111111111010110111110111;
assign LUT_1[16911] = 32'b11111111111111110100001001110011;
assign LUT_1[16912] = 32'b11111111111111111001111101111100;
assign LUT_1[16913] = 32'b11111111111111110011001111111000;
assign LUT_1[16914] = 32'b11111111111111110101101100001101;
assign LUT_1[16915] = 32'b11111111111111101110111110001001;
assign LUT_1[16916] = 32'b00000000000000000001110111010011;
assign LUT_1[16917] = 32'b11111111111111111011001001001111;
assign LUT_1[16918] = 32'b11111111111111111101100101100100;
assign LUT_1[16919] = 32'b11111111111111110110110111100000;
assign LUT_1[16920] = 32'b11111111111111111001001011110001;
assign LUT_1[16921] = 32'b11111111111111110010011101101101;
assign LUT_1[16922] = 32'b11111111111111110100111010000010;
assign LUT_1[16923] = 32'b11111111111111101110001011111110;
assign LUT_1[16924] = 32'b00000000000000000001000101001000;
assign LUT_1[16925] = 32'b11111111111111111010010111000100;
assign LUT_1[16926] = 32'b11111111111111111100110011011001;
assign LUT_1[16927] = 32'b11111111111111110110000101010101;
assign LUT_1[16928] = 32'b11111111111111111000111101011001;
assign LUT_1[16929] = 32'b11111111111111110010001111010101;
assign LUT_1[16930] = 32'b11111111111111110100101011101010;
assign LUT_1[16931] = 32'b11111111111111101101111101100110;
assign LUT_1[16932] = 32'b00000000000000000000110110110000;
assign LUT_1[16933] = 32'b11111111111111111010001000101100;
assign LUT_1[16934] = 32'b11111111111111111100100101000001;
assign LUT_1[16935] = 32'b11111111111111110101110110111101;
assign LUT_1[16936] = 32'b11111111111111111000001011001110;
assign LUT_1[16937] = 32'b11111111111111110001011101001010;
assign LUT_1[16938] = 32'b11111111111111110011111001011111;
assign LUT_1[16939] = 32'b11111111111111101101001011011011;
assign LUT_1[16940] = 32'b00000000000000000000000100100101;
assign LUT_1[16941] = 32'b11111111111111111001010110100001;
assign LUT_1[16942] = 32'b11111111111111111011110010110110;
assign LUT_1[16943] = 32'b11111111111111110101000100110010;
assign LUT_1[16944] = 32'b11111111111111111010111000111011;
assign LUT_1[16945] = 32'b11111111111111110100001010110111;
assign LUT_1[16946] = 32'b11111111111111110110100111001100;
assign LUT_1[16947] = 32'b11111111111111101111111001001000;
assign LUT_1[16948] = 32'b00000000000000000010110010010010;
assign LUT_1[16949] = 32'b11111111111111111100000100001110;
assign LUT_1[16950] = 32'b11111111111111111110100000100011;
assign LUT_1[16951] = 32'b11111111111111110111110010011111;
assign LUT_1[16952] = 32'b11111111111111111010000110110000;
assign LUT_1[16953] = 32'b11111111111111110011011000101100;
assign LUT_1[16954] = 32'b11111111111111110101110101000001;
assign LUT_1[16955] = 32'b11111111111111101111000110111101;
assign LUT_1[16956] = 32'b00000000000000000010000000000111;
assign LUT_1[16957] = 32'b11111111111111111011010010000011;
assign LUT_1[16958] = 32'b11111111111111111101101110011000;
assign LUT_1[16959] = 32'b11111111111111110111000000010100;
assign LUT_1[16960] = 32'b11111111111111111010000000000010;
assign LUT_1[16961] = 32'b11111111111111110011010001111110;
assign LUT_1[16962] = 32'b11111111111111110101101110010011;
assign LUT_1[16963] = 32'b11111111111111101111000000001111;
assign LUT_1[16964] = 32'b00000000000000000001111001011001;
assign LUT_1[16965] = 32'b11111111111111111011001011010101;
assign LUT_1[16966] = 32'b11111111111111111101100111101010;
assign LUT_1[16967] = 32'b11111111111111110110111001100110;
assign LUT_1[16968] = 32'b11111111111111111001001101110111;
assign LUT_1[16969] = 32'b11111111111111110010011111110011;
assign LUT_1[16970] = 32'b11111111111111110100111100001000;
assign LUT_1[16971] = 32'b11111111111111101110001110000100;
assign LUT_1[16972] = 32'b00000000000000000001000111001110;
assign LUT_1[16973] = 32'b11111111111111111010011001001010;
assign LUT_1[16974] = 32'b11111111111111111100110101011111;
assign LUT_1[16975] = 32'b11111111111111110110000111011011;
assign LUT_1[16976] = 32'b11111111111111111011111011100100;
assign LUT_1[16977] = 32'b11111111111111110101001101100000;
assign LUT_1[16978] = 32'b11111111111111110111101001110101;
assign LUT_1[16979] = 32'b11111111111111110000111011110001;
assign LUT_1[16980] = 32'b00000000000000000011110100111011;
assign LUT_1[16981] = 32'b11111111111111111101000110110111;
assign LUT_1[16982] = 32'b11111111111111111111100011001100;
assign LUT_1[16983] = 32'b11111111111111111000110101001000;
assign LUT_1[16984] = 32'b11111111111111111011001001011001;
assign LUT_1[16985] = 32'b11111111111111110100011011010101;
assign LUT_1[16986] = 32'b11111111111111110110110111101010;
assign LUT_1[16987] = 32'b11111111111111110000001001100110;
assign LUT_1[16988] = 32'b00000000000000000011000010110000;
assign LUT_1[16989] = 32'b11111111111111111100010100101100;
assign LUT_1[16990] = 32'b11111111111111111110110001000001;
assign LUT_1[16991] = 32'b11111111111111111000000010111101;
assign LUT_1[16992] = 32'b11111111111111111010111011000001;
assign LUT_1[16993] = 32'b11111111111111110100001100111101;
assign LUT_1[16994] = 32'b11111111111111110110101001010010;
assign LUT_1[16995] = 32'b11111111111111101111111011001110;
assign LUT_1[16996] = 32'b00000000000000000010110100011000;
assign LUT_1[16997] = 32'b11111111111111111100000110010100;
assign LUT_1[16998] = 32'b11111111111111111110100010101001;
assign LUT_1[16999] = 32'b11111111111111110111110100100101;
assign LUT_1[17000] = 32'b11111111111111111010001000110110;
assign LUT_1[17001] = 32'b11111111111111110011011010110010;
assign LUT_1[17002] = 32'b11111111111111110101110111000111;
assign LUT_1[17003] = 32'b11111111111111101111001001000011;
assign LUT_1[17004] = 32'b00000000000000000010000010001101;
assign LUT_1[17005] = 32'b11111111111111111011010100001001;
assign LUT_1[17006] = 32'b11111111111111111101110000011110;
assign LUT_1[17007] = 32'b11111111111111110111000010011010;
assign LUT_1[17008] = 32'b11111111111111111100110110100011;
assign LUT_1[17009] = 32'b11111111111111110110001000011111;
assign LUT_1[17010] = 32'b11111111111111111000100100110100;
assign LUT_1[17011] = 32'b11111111111111110001110110110000;
assign LUT_1[17012] = 32'b00000000000000000100101111111010;
assign LUT_1[17013] = 32'b11111111111111111110000001110110;
assign LUT_1[17014] = 32'b00000000000000000000011110001011;
assign LUT_1[17015] = 32'b11111111111111111001110000000111;
assign LUT_1[17016] = 32'b11111111111111111100000100011000;
assign LUT_1[17017] = 32'b11111111111111110101010110010100;
assign LUT_1[17018] = 32'b11111111111111110111110010101001;
assign LUT_1[17019] = 32'b11111111111111110001000100100101;
assign LUT_1[17020] = 32'b00000000000000000011111101101111;
assign LUT_1[17021] = 32'b11111111111111111101001111101011;
assign LUT_1[17022] = 32'b11111111111111111111101100000000;
assign LUT_1[17023] = 32'b11111111111111111000111101111100;
assign LUT_1[17024] = 32'b11111111111111111011000010011101;
assign LUT_1[17025] = 32'b11111111111111110100010100011001;
assign LUT_1[17026] = 32'b11111111111111110110110000101110;
assign LUT_1[17027] = 32'b11111111111111110000000010101010;
assign LUT_1[17028] = 32'b00000000000000000010111011110100;
assign LUT_1[17029] = 32'b11111111111111111100001101110000;
assign LUT_1[17030] = 32'b11111111111111111110101010000101;
assign LUT_1[17031] = 32'b11111111111111110111111100000001;
assign LUT_1[17032] = 32'b11111111111111111010010000010010;
assign LUT_1[17033] = 32'b11111111111111110011100010001110;
assign LUT_1[17034] = 32'b11111111111111110101111110100011;
assign LUT_1[17035] = 32'b11111111111111101111010000011111;
assign LUT_1[17036] = 32'b00000000000000000010001001101001;
assign LUT_1[17037] = 32'b11111111111111111011011011100101;
assign LUT_1[17038] = 32'b11111111111111111101110111111010;
assign LUT_1[17039] = 32'b11111111111111110111001001110110;
assign LUT_1[17040] = 32'b11111111111111111100111101111111;
assign LUT_1[17041] = 32'b11111111111111110110001111111011;
assign LUT_1[17042] = 32'b11111111111111111000101100010000;
assign LUT_1[17043] = 32'b11111111111111110001111110001100;
assign LUT_1[17044] = 32'b00000000000000000100110111010110;
assign LUT_1[17045] = 32'b11111111111111111110001001010010;
assign LUT_1[17046] = 32'b00000000000000000000100101100111;
assign LUT_1[17047] = 32'b11111111111111111001110111100011;
assign LUT_1[17048] = 32'b11111111111111111100001011110100;
assign LUT_1[17049] = 32'b11111111111111110101011101110000;
assign LUT_1[17050] = 32'b11111111111111110111111010000101;
assign LUT_1[17051] = 32'b11111111111111110001001100000001;
assign LUT_1[17052] = 32'b00000000000000000100000101001011;
assign LUT_1[17053] = 32'b11111111111111111101010111000111;
assign LUT_1[17054] = 32'b11111111111111111111110011011100;
assign LUT_1[17055] = 32'b11111111111111111001000101011000;
assign LUT_1[17056] = 32'b11111111111111111011111101011100;
assign LUT_1[17057] = 32'b11111111111111110101001111011000;
assign LUT_1[17058] = 32'b11111111111111110111101011101101;
assign LUT_1[17059] = 32'b11111111111111110000111101101001;
assign LUT_1[17060] = 32'b00000000000000000011110110110011;
assign LUT_1[17061] = 32'b11111111111111111101001000101111;
assign LUT_1[17062] = 32'b11111111111111111111100101000100;
assign LUT_1[17063] = 32'b11111111111111111000110111000000;
assign LUT_1[17064] = 32'b11111111111111111011001011010001;
assign LUT_1[17065] = 32'b11111111111111110100011101001101;
assign LUT_1[17066] = 32'b11111111111111110110111001100010;
assign LUT_1[17067] = 32'b11111111111111110000001011011110;
assign LUT_1[17068] = 32'b00000000000000000011000100101000;
assign LUT_1[17069] = 32'b11111111111111111100010110100100;
assign LUT_1[17070] = 32'b11111111111111111110110010111001;
assign LUT_1[17071] = 32'b11111111111111111000000100110101;
assign LUT_1[17072] = 32'b11111111111111111101111000111110;
assign LUT_1[17073] = 32'b11111111111111110111001010111010;
assign LUT_1[17074] = 32'b11111111111111111001100111001111;
assign LUT_1[17075] = 32'b11111111111111110010111001001011;
assign LUT_1[17076] = 32'b00000000000000000101110010010101;
assign LUT_1[17077] = 32'b11111111111111111111000100010001;
assign LUT_1[17078] = 32'b00000000000000000001100000100110;
assign LUT_1[17079] = 32'b11111111111111111010110010100010;
assign LUT_1[17080] = 32'b11111111111111111101000110110011;
assign LUT_1[17081] = 32'b11111111111111110110011000101111;
assign LUT_1[17082] = 32'b11111111111111111000110101000100;
assign LUT_1[17083] = 32'b11111111111111110010000111000000;
assign LUT_1[17084] = 32'b00000000000000000101000000001010;
assign LUT_1[17085] = 32'b11111111111111111110010010000110;
assign LUT_1[17086] = 32'b00000000000000000000101110011011;
assign LUT_1[17087] = 32'b11111111111111111010000000010111;
assign LUT_1[17088] = 32'b11111111111111111101000000000101;
assign LUT_1[17089] = 32'b11111111111111110110010010000001;
assign LUT_1[17090] = 32'b11111111111111111000101110010110;
assign LUT_1[17091] = 32'b11111111111111110010000000010010;
assign LUT_1[17092] = 32'b00000000000000000100111001011100;
assign LUT_1[17093] = 32'b11111111111111111110001011011000;
assign LUT_1[17094] = 32'b00000000000000000000100111101101;
assign LUT_1[17095] = 32'b11111111111111111001111001101001;
assign LUT_1[17096] = 32'b11111111111111111100001101111010;
assign LUT_1[17097] = 32'b11111111111111110101011111110110;
assign LUT_1[17098] = 32'b11111111111111110111111100001011;
assign LUT_1[17099] = 32'b11111111111111110001001110000111;
assign LUT_1[17100] = 32'b00000000000000000100000111010001;
assign LUT_1[17101] = 32'b11111111111111111101011001001101;
assign LUT_1[17102] = 32'b11111111111111111111110101100010;
assign LUT_1[17103] = 32'b11111111111111111001000111011110;
assign LUT_1[17104] = 32'b11111111111111111110111011100111;
assign LUT_1[17105] = 32'b11111111111111111000001101100011;
assign LUT_1[17106] = 32'b11111111111111111010101001111000;
assign LUT_1[17107] = 32'b11111111111111110011111011110100;
assign LUT_1[17108] = 32'b00000000000000000110110100111110;
assign LUT_1[17109] = 32'b00000000000000000000000110111010;
assign LUT_1[17110] = 32'b00000000000000000010100011001111;
assign LUT_1[17111] = 32'b11111111111111111011110101001011;
assign LUT_1[17112] = 32'b11111111111111111110001001011100;
assign LUT_1[17113] = 32'b11111111111111110111011011011000;
assign LUT_1[17114] = 32'b11111111111111111001110111101101;
assign LUT_1[17115] = 32'b11111111111111110011001001101001;
assign LUT_1[17116] = 32'b00000000000000000110000010110011;
assign LUT_1[17117] = 32'b11111111111111111111010100101111;
assign LUT_1[17118] = 32'b00000000000000000001110001000100;
assign LUT_1[17119] = 32'b11111111111111111011000011000000;
assign LUT_1[17120] = 32'b11111111111111111101111011000100;
assign LUT_1[17121] = 32'b11111111111111110111001101000000;
assign LUT_1[17122] = 32'b11111111111111111001101001010101;
assign LUT_1[17123] = 32'b11111111111111110010111011010001;
assign LUT_1[17124] = 32'b00000000000000000101110100011011;
assign LUT_1[17125] = 32'b11111111111111111111000110010111;
assign LUT_1[17126] = 32'b00000000000000000001100010101100;
assign LUT_1[17127] = 32'b11111111111111111010110100101000;
assign LUT_1[17128] = 32'b11111111111111111101001000111001;
assign LUT_1[17129] = 32'b11111111111111110110011010110101;
assign LUT_1[17130] = 32'b11111111111111111000110111001010;
assign LUT_1[17131] = 32'b11111111111111110010001001000110;
assign LUT_1[17132] = 32'b00000000000000000101000010010000;
assign LUT_1[17133] = 32'b11111111111111111110010100001100;
assign LUT_1[17134] = 32'b00000000000000000000110000100001;
assign LUT_1[17135] = 32'b11111111111111111010000010011101;
assign LUT_1[17136] = 32'b11111111111111111111110110100110;
assign LUT_1[17137] = 32'b11111111111111111001001000100010;
assign LUT_1[17138] = 32'b11111111111111111011100100110111;
assign LUT_1[17139] = 32'b11111111111111110100110110110011;
assign LUT_1[17140] = 32'b00000000000000000111101111111101;
assign LUT_1[17141] = 32'b00000000000000000001000001111001;
assign LUT_1[17142] = 32'b00000000000000000011011110001110;
assign LUT_1[17143] = 32'b11111111111111111100110000001010;
assign LUT_1[17144] = 32'b11111111111111111111000100011011;
assign LUT_1[17145] = 32'b11111111111111111000010110010111;
assign LUT_1[17146] = 32'b11111111111111111010110010101100;
assign LUT_1[17147] = 32'b11111111111111110100000100101000;
assign LUT_1[17148] = 32'b00000000000000000110111101110010;
assign LUT_1[17149] = 32'b00000000000000000000001111101110;
assign LUT_1[17150] = 32'b00000000000000000010101100000011;
assign LUT_1[17151] = 32'b11111111111111111011111101111111;
assign LUT_1[17152] = 32'b11111111111111110101110110100110;
assign LUT_1[17153] = 32'b11111111111111101111001000100010;
assign LUT_1[17154] = 32'b11111111111111110001100100110111;
assign LUT_1[17155] = 32'b11111111111111101010110110110011;
assign LUT_1[17156] = 32'b11111111111111111101101111111101;
assign LUT_1[17157] = 32'b11111111111111110111000001111001;
assign LUT_1[17158] = 32'b11111111111111111001011110001110;
assign LUT_1[17159] = 32'b11111111111111110010110000001010;
assign LUT_1[17160] = 32'b11111111111111110101000100011011;
assign LUT_1[17161] = 32'b11111111111111101110010110010111;
assign LUT_1[17162] = 32'b11111111111111110000110010101100;
assign LUT_1[17163] = 32'b11111111111111101010000100101000;
assign LUT_1[17164] = 32'b11111111111111111100111101110010;
assign LUT_1[17165] = 32'b11111111111111110110001111101110;
assign LUT_1[17166] = 32'b11111111111111111000101100000011;
assign LUT_1[17167] = 32'b11111111111111110001111101111111;
assign LUT_1[17168] = 32'b11111111111111110111110010001000;
assign LUT_1[17169] = 32'b11111111111111110001000100000100;
assign LUT_1[17170] = 32'b11111111111111110011100000011001;
assign LUT_1[17171] = 32'b11111111111111101100110010010101;
assign LUT_1[17172] = 32'b11111111111111111111101011011111;
assign LUT_1[17173] = 32'b11111111111111111000111101011011;
assign LUT_1[17174] = 32'b11111111111111111011011001110000;
assign LUT_1[17175] = 32'b11111111111111110100101011101100;
assign LUT_1[17176] = 32'b11111111111111110110111111111101;
assign LUT_1[17177] = 32'b11111111111111110000010001111001;
assign LUT_1[17178] = 32'b11111111111111110010101110001110;
assign LUT_1[17179] = 32'b11111111111111101100000000001010;
assign LUT_1[17180] = 32'b11111111111111111110111001010100;
assign LUT_1[17181] = 32'b11111111111111111000001011010000;
assign LUT_1[17182] = 32'b11111111111111111010100111100101;
assign LUT_1[17183] = 32'b11111111111111110011111001100001;
assign LUT_1[17184] = 32'b11111111111111110110110001100101;
assign LUT_1[17185] = 32'b11111111111111110000000011100001;
assign LUT_1[17186] = 32'b11111111111111110010011111110110;
assign LUT_1[17187] = 32'b11111111111111101011110001110010;
assign LUT_1[17188] = 32'b11111111111111111110101010111100;
assign LUT_1[17189] = 32'b11111111111111110111111100111000;
assign LUT_1[17190] = 32'b11111111111111111010011001001101;
assign LUT_1[17191] = 32'b11111111111111110011101011001001;
assign LUT_1[17192] = 32'b11111111111111110101111111011010;
assign LUT_1[17193] = 32'b11111111111111101111010001010110;
assign LUT_1[17194] = 32'b11111111111111110001101101101011;
assign LUT_1[17195] = 32'b11111111111111101010111111100111;
assign LUT_1[17196] = 32'b11111111111111111101111000110001;
assign LUT_1[17197] = 32'b11111111111111110111001010101101;
assign LUT_1[17198] = 32'b11111111111111111001100111000010;
assign LUT_1[17199] = 32'b11111111111111110010111000111110;
assign LUT_1[17200] = 32'b11111111111111111000101101000111;
assign LUT_1[17201] = 32'b11111111111111110001111111000011;
assign LUT_1[17202] = 32'b11111111111111110100011011011000;
assign LUT_1[17203] = 32'b11111111111111101101101101010100;
assign LUT_1[17204] = 32'b00000000000000000000100110011110;
assign LUT_1[17205] = 32'b11111111111111111001111000011010;
assign LUT_1[17206] = 32'b11111111111111111100010100101111;
assign LUT_1[17207] = 32'b11111111111111110101100110101011;
assign LUT_1[17208] = 32'b11111111111111110111111010111100;
assign LUT_1[17209] = 32'b11111111111111110001001100111000;
assign LUT_1[17210] = 32'b11111111111111110011101001001101;
assign LUT_1[17211] = 32'b11111111111111101100111011001001;
assign LUT_1[17212] = 32'b11111111111111111111110100010011;
assign LUT_1[17213] = 32'b11111111111111111001000110001111;
assign LUT_1[17214] = 32'b11111111111111111011100010100100;
assign LUT_1[17215] = 32'b11111111111111110100110100100000;
assign LUT_1[17216] = 32'b11111111111111110111110100001110;
assign LUT_1[17217] = 32'b11111111111111110001000110001010;
assign LUT_1[17218] = 32'b11111111111111110011100010011111;
assign LUT_1[17219] = 32'b11111111111111101100110100011011;
assign LUT_1[17220] = 32'b11111111111111111111101101100101;
assign LUT_1[17221] = 32'b11111111111111111000111111100001;
assign LUT_1[17222] = 32'b11111111111111111011011011110110;
assign LUT_1[17223] = 32'b11111111111111110100101101110010;
assign LUT_1[17224] = 32'b11111111111111110111000010000011;
assign LUT_1[17225] = 32'b11111111111111110000010011111111;
assign LUT_1[17226] = 32'b11111111111111110010110000010100;
assign LUT_1[17227] = 32'b11111111111111101100000010010000;
assign LUT_1[17228] = 32'b11111111111111111110111011011010;
assign LUT_1[17229] = 32'b11111111111111111000001101010110;
assign LUT_1[17230] = 32'b11111111111111111010101001101011;
assign LUT_1[17231] = 32'b11111111111111110011111011100111;
assign LUT_1[17232] = 32'b11111111111111111001101111110000;
assign LUT_1[17233] = 32'b11111111111111110011000001101100;
assign LUT_1[17234] = 32'b11111111111111110101011110000001;
assign LUT_1[17235] = 32'b11111111111111101110101111111101;
assign LUT_1[17236] = 32'b00000000000000000001101001000111;
assign LUT_1[17237] = 32'b11111111111111111010111011000011;
assign LUT_1[17238] = 32'b11111111111111111101010111011000;
assign LUT_1[17239] = 32'b11111111111111110110101001010100;
assign LUT_1[17240] = 32'b11111111111111111000111101100101;
assign LUT_1[17241] = 32'b11111111111111110010001111100001;
assign LUT_1[17242] = 32'b11111111111111110100101011110110;
assign LUT_1[17243] = 32'b11111111111111101101111101110010;
assign LUT_1[17244] = 32'b00000000000000000000110110111100;
assign LUT_1[17245] = 32'b11111111111111111010001000111000;
assign LUT_1[17246] = 32'b11111111111111111100100101001101;
assign LUT_1[17247] = 32'b11111111111111110101110111001001;
assign LUT_1[17248] = 32'b11111111111111111000101111001101;
assign LUT_1[17249] = 32'b11111111111111110010000001001001;
assign LUT_1[17250] = 32'b11111111111111110100011101011110;
assign LUT_1[17251] = 32'b11111111111111101101101111011010;
assign LUT_1[17252] = 32'b00000000000000000000101000100100;
assign LUT_1[17253] = 32'b11111111111111111001111010100000;
assign LUT_1[17254] = 32'b11111111111111111100010110110101;
assign LUT_1[17255] = 32'b11111111111111110101101000110001;
assign LUT_1[17256] = 32'b11111111111111110111111101000010;
assign LUT_1[17257] = 32'b11111111111111110001001110111110;
assign LUT_1[17258] = 32'b11111111111111110011101011010011;
assign LUT_1[17259] = 32'b11111111111111101100111101001111;
assign LUT_1[17260] = 32'b11111111111111111111110110011001;
assign LUT_1[17261] = 32'b11111111111111111001001000010101;
assign LUT_1[17262] = 32'b11111111111111111011100100101010;
assign LUT_1[17263] = 32'b11111111111111110100110110100110;
assign LUT_1[17264] = 32'b11111111111111111010101010101111;
assign LUT_1[17265] = 32'b11111111111111110011111100101011;
assign LUT_1[17266] = 32'b11111111111111110110011001000000;
assign LUT_1[17267] = 32'b11111111111111101111101010111100;
assign LUT_1[17268] = 32'b00000000000000000010100100000110;
assign LUT_1[17269] = 32'b11111111111111111011110110000010;
assign LUT_1[17270] = 32'b11111111111111111110010010010111;
assign LUT_1[17271] = 32'b11111111111111110111100100010011;
assign LUT_1[17272] = 32'b11111111111111111001111000100100;
assign LUT_1[17273] = 32'b11111111111111110011001010100000;
assign LUT_1[17274] = 32'b11111111111111110101100110110101;
assign LUT_1[17275] = 32'b11111111111111101110111000110001;
assign LUT_1[17276] = 32'b00000000000000000001110001111011;
assign LUT_1[17277] = 32'b11111111111111111011000011110111;
assign LUT_1[17278] = 32'b11111111111111111101100000001100;
assign LUT_1[17279] = 32'b11111111111111110110110010001000;
assign LUT_1[17280] = 32'b11111111111111111000110110101001;
assign LUT_1[17281] = 32'b11111111111111110010001000100101;
assign LUT_1[17282] = 32'b11111111111111110100100100111010;
assign LUT_1[17283] = 32'b11111111111111101101110110110110;
assign LUT_1[17284] = 32'b00000000000000000000110000000000;
assign LUT_1[17285] = 32'b11111111111111111010000001111100;
assign LUT_1[17286] = 32'b11111111111111111100011110010001;
assign LUT_1[17287] = 32'b11111111111111110101110000001101;
assign LUT_1[17288] = 32'b11111111111111111000000100011110;
assign LUT_1[17289] = 32'b11111111111111110001010110011010;
assign LUT_1[17290] = 32'b11111111111111110011110010101111;
assign LUT_1[17291] = 32'b11111111111111101101000100101011;
assign LUT_1[17292] = 32'b11111111111111111111111101110101;
assign LUT_1[17293] = 32'b11111111111111111001001111110001;
assign LUT_1[17294] = 32'b11111111111111111011101100000110;
assign LUT_1[17295] = 32'b11111111111111110100111110000010;
assign LUT_1[17296] = 32'b11111111111111111010110010001011;
assign LUT_1[17297] = 32'b11111111111111110100000100000111;
assign LUT_1[17298] = 32'b11111111111111110110100000011100;
assign LUT_1[17299] = 32'b11111111111111101111110010011000;
assign LUT_1[17300] = 32'b00000000000000000010101011100010;
assign LUT_1[17301] = 32'b11111111111111111011111101011110;
assign LUT_1[17302] = 32'b11111111111111111110011001110011;
assign LUT_1[17303] = 32'b11111111111111110111101011101111;
assign LUT_1[17304] = 32'b11111111111111111010000000000000;
assign LUT_1[17305] = 32'b11111111111111110011010001111100;
assign LUT_1[17306] = 32'b11111111111111110101101110010001;
assign LUT_1[17307] = 32'b11111111111111101111000000001101;
assign LUT_1[17308] = 32'b00000000000000000001111001010111;
assign LUT_1[17309] = 32'b11111111111111111011001011010011;
assign LUT_1[17310] = 32'b11111111111111111101100111101000;
assign LUT_1[17311] = 32'b11111111111111110110111001100100;
assign LUT_1[17312] = 32'b11111111111111111001110001101000;
assign LUT_1[17313] = 32'b11111111111111110011000011100100;
assign LUT_1[17314] = 32'b11111111111111110101011111111001;
assign LUT_1[17315] = 32'b11111111111111101110110001110101;
assign LUT_1[17316] = 32'b00000000000000000001101010111111;
assign LUT_1[17317] = 32'b11111111111111111010111100111011;
assign LUT_1[17318] = 32'b11111111111111111101011001010000;
assign LUT_1[17319] = 32'b11111111111111110110101011001100;
assign LUT_1[17320] = 32'b11111111111111111000111111011101;
assign LUT_1[17321] = 32'b11111111111111110010010001011001;
assign LUT_1[17322] = 32'b11111111111111110100101101101110;
assign LUT_1[17323] = 32'b11111111111111101101111111101010;
assign LUT_1[17324] = 32'b00000000000000000000111000110100;
assign LUT_1[17325] = 32'b11111111111111111010001010110000;
assign LUT_1[17326] = 32'b11111111111111111100100111000101;
assign LUT_1[17327] = 32'b11111111111111110101111001000001;
assign LUT_1[17328] = 32'b11111111111111111011101101001010;
assign LUT_1[17329] = 32'b11111111111111110100111111000110;
assign LUT_1[17330] = 32'b11111111111111110111011011011011;
assign LUT_1[17331] = 32'b11111111111111110000101101010111;
assign LUT_1[17332] = 32'b00000000000000000011100110100001;
assign LUT_1[17333] = 32'b11111111111111111100111000011101;
assign LUT_1[17334] = 32'b11111111111111111111010100110010;
assign LUT_1[17335] = 32'b11111111111111111000100110101110;
assign LUT_1[17336] = 32'b11111111111111111010111010111111;
assign LUT_1[17337] = 32'b11111111111111110100001100111011;
assign LUT_1[17338] = 32'b11111111111111110110101001010000;
assign LUT_1[17339] = 32'b11111111111111101111111011001100;
assign LUT_1[17340] = 32'b00000000000000000010110100010110;
assign LUT_1[17341] = 32'b11111111111111111100000110010010;
assign LUT_1[17342] = 32'b11111111111111111110100010100111;
assign LUT_1[17343] = 32'b11111111111111110111110100100011;
assign LUT_1[17344] = 32'b11111111111111111010110100010001;
assign LUT_1[17345] = 32'b11111111111111110100000110001101;
assign LUT_1[17346] = 32'b11111111111111110110100010100010;
assign LUT_1[17347] = 32'b11111111111111101111110100011110;
assign LUT_1[17348] = 32'b00000000000000000010101101101000;
assign LUT_1[17349] = 32'b11111111111111111011111111100100;
assign LUT_1[17350] = 32'b11111111111111111110011011111001;
assign LUT_1[17351] = 32'b11111111111111110111101101110101;
assign LUT_1[17352] = 32'b11111111111111111010000010000110;
assign LUT_1[17353] = 32'b11111111111111110011010100000010;
assign LUT_1[17354] = 32'b11111111111111110101110000010111;
assign LUT_1[17355] = 32'b11111111111111101111000010010011;
assign LUT_1[17356] = 32'b00000000000000000001111011011101;
assign LUT_1[17357] = 32'b11111111111111111011001101011001;
assign LUT_1[17358] = 32'b11111111111111111101101001101110;
assign LUT_1[17359] = 32'b11111111111111110110111011101010;
assign LUT_1[17360] = 32'b11111111111111111100101111110011;
assign LUT_1[17361] = 32'b11111111111111110110000001101111;
assign LUT_1[17362] = 32'b11111111111111111000011110000100;
assign LUT_1[17363] = 32'b11111111111111110001110000000000;
assign LUT_1[17364] = 32'b00000000000000000100101001001010;
assign LUT_1[17365] = 32'b11111111111111111101111011000110;
assign LUT_1[17366] = 32'b00000000000000000000010111011011;
assign LUT_1[17367] = 32'b11111111111111111001101001010111;
assign LUT_1[17368] = 32'b11111111111111111011111101101000;
assign LUT_1[17369] = 32'b11111111111111110101001111100100;
assign LUT_1[17370] = 32'b11111111111111110111101011111001;
assign LUT_1[17371] = 32'b11111111111111110000111101110101;
assign LUT_1[17372] = 32'b00000000000000000011110110111111;
assign LUT_1[17373] = 32'b11111111111111111101001000111011;
assign LUT_1[17374] = 32'b11111111111111111111100101010000;
assign LUT_1[17375] = 32'b11111111111111111000110111001100;
assign LUT_1[17376] = 32'b11111111111111111011101111010000;
assign LUT_1[17377] = 32'b11111111111111110101000001001100;
assign LUT_1[17378] = 32'b11111111111111110111011101100001;
assign LUT_1[17379] = 32'b11111111111111110000101111011101;
assign LUT_1[17380] = 32'b00000000000000000011101000100111;
assign LUT_1[17381] = 32'b11111111111111111100111010100011;
assign LUT_1[17382] = 32'b11111111111111111111010110111000;
assign LUT_1[17383] = 32'b11111111111111111000101000110100;
assign LUT_1[17384] = 32'b11111111111111111010111101000101;
assign LUT_1[17385] = 32'b11111111111111110100001111000001;
assign LUT_1[17386] = 32'b11111111111111110110101011010110;
assign LUT_1[17387] = 32'b11111111111111101111111101010010;
assign LUT_1[17388] = 32'b00000000000000000010110110011100;
assign LUT_1[17389] = 32'b11111111111111111100001000011000;
assign LUT_1[17390] = 32'b11111111111111111110100100101101;
assign LUT_1[17391] = 32'b11111111111111110111110110101001;
assign LUT_1[17392] = 32'b11111111111111111101101010110010;
assign LUT_1[17393] = 32'b11111111111111110110111100101110;
assign LUT_1[17394] = 32'b11111111111111111001011001000011;
assign LUT_1[17395] = 32'b11111111111111110010101010111111;
assign LUT_1[17396] = 32'b00000000000000000101100100001001;
assign LUT_1[17397] = 32'b11111111111111111110110110000101;
assign LUT_1[17398] = 32'b00000000000000000001010010011010;
assign LUT_1[17399] = 32'b11111111111111111010100100010110;
assign LUT_1[17400] = 32'b11111111111111111100111000100111;
assign LUT_1[17401] = 32'b11111111111111110110001010100011;
assign LUT_1[17402] = 32'b11111111111111111000100110111000;
assign LUT_1[17403] = 32'b11111111111111110001111000110100;
assign LUT_1[17404] = 32'b00000000000000000100110001111110;
assign LUT_1[17405] = 32'b11111111111111111110000011111010;
assign LUT_1[17406] = 32'b00000000000000000000100000001111;
assign LUT_1[17407] = 32'b11111111111111111001110010001011;
assign LUT_1[17408] = 32'b00000000000000000100101010101101;
assign LUT_1[17409] = 32'b11111111111111111101111100101001;
assign LUT_1[17410] = 32'b00000000000000000000011000111110;
assign LUT_1[17411] = 32'b11111111111111111001101010111010;
assign LUT_1[17412] = 32'b00000000000000001100100100000100;
assign LUT_1[17413] = 32'b00000000000000000101110110000000;
assign LUT_1[17414] = 32'b00000000000000001000010010010101;
assign LUT_1[17415] = 32'b00000000000000000001100100010001;
assign LUT_1[17416] = 32'b00000000000000000011111000100010;
assign LUT_1[17417] = 32'b11111111111111111101001010011110;
assign LUT_1[17418] = 32'b11111111111111111111100110110011;
assign LUT_1[17419] = 32'b11111111111111111000111000101111;
assign LUT_1[17420] = 32'b00000000000000001011110001111001;
assign LUT_1[17421] = 32'b00000000000000000101000011110101;
assign LUT_1[17422] = 32'b00000000000000000111100000001010;
assign LUT_1[17423] = 32'b00000000000000000000110010000110;
assign LUT_1[17424] = 32'b00000000000000000110100110001111;
assign LUT_1[17425] = 32'b11111111111111111111111000001011;
assign LUT_1[17426] = 32'b00000000000000000010010100100000;
assign LUT_1[17427] = 32'b11111111111111111011100110011100;
assign LUT_1[17428] = 32'b00000000000000001110011111100110;
assign LUT_1[17429] = 32'b00000000000000000111110001100010;
assign LUT_1[17430] = 32'b00000000000000001010001101110111;
assign LUT_1[17431] = 32'b00000000000000000011011111110011;
assign LUT_1[17432] = 32'b00000000000000000101110100000100;
assign LUT_1[17433] = 32'b11111111111111111111000110000000;
assign LUT_1[17434] = 32'b00000000000000000001100010010101;
assign LUT_1[17435] = 32'b11111111111111111010110100010001;
assign LUT_1[17436] = 32'b00000000000000001101101101011011;
assign LUT_1[17437] = 32'b00000000000000000110111111010111;
assign LUT_1[17438] = 32'b00000000000000001001011011101100;
assign LUT_1[17439] = 32'b00000000000000000010101101101000;
assign LUT_1[17440] = 32'b00000000000000000101100101101100;
assign LUT_1[17441] = 32'b11111111111111111110110111101000;
assign LUT_1[17442] = 32'b00000000000000000001010011111101;
assign LUT_1[17443] = 32'b11111111111111111010100101111001;
assign LUT_1[17444] = 32'b00000000000000001101011111000011;
assign LUT_1[17445] = 32'b00000000000000000110110000111111;
assign LUT_1[17446] = 32'b00000000000000001001001101010100;
assign LUT_1[17447] = 32'b00000000000000000010011111010000;
assign LUT_1[17448] = 32'b00000000000000000100110011100001;
assign LUT_1[17449] = 32'b11111111111111111110000101011101;
assign LUT_1[17450] = 32'b00000000000000000000100001110010;
assign LUT_1[17451] = 32'b11111111111111111001110011101110;
assign LUT_1[17452] = 32'b00000000000000001100101100111000;
assign LUT_1[17453] = 32'b00000000000000000101111110110100;
assign LUT_1[17454] = 32'b00000000000000001000011011001001;
assign LUT_1[17455] = 32'b00000000000000000001101101000101;
assign LUT_1[17456] = 32'b00000000000000000111100001001110;
assign LUT_1[17457] = 32'b00000000000000000000110011001010;
assign LUT_1[17458] = 32'b00000000000000000011001111011111;
assign LUT_1[17459] = 32'b11111111111111111100100001011011;
assign LUT_1[17460] = 32'b00000000000000001111011010100101;
assign LUT_1[17461] = 32'b00000000000000001000101100100001;
assign LUT_1[17462] = 32'b00000000000000001011001000110110;
assign LUT_1[17463] = 32'b00000000000000000100011010110010;
assign LUT_1[17464] = 32'b00000000000000000110101111000011;
assign LUT_1[17465] = 32'b00000000000000000000000000111111;
assign LUT_1[17466] = 32'b00000000000000000010011101010100;
assign LUT_1[17467] = 32'b11111111111111111011101111010000;
assign LUT_1[17468] = 32'b00000000000000001110101000011010;
assign LUT_1[17469] = 32'b00000000000000000111111010010110;
assign LUT_1[17470] = 32'b00000000000000001010010110101011;
assign LUT_1[17471] = 32'b00000000000000000011101000100111;
assign LUT_1[17472] = 32'b00000000000000000110101000010101;
assign LUT_1[17473] = 32'b11111111111111111111111010010001;
assign LUT_1[17474] = 32'b00000000000000000010010110100110;
assign LUT_1[17475] = 32'b11111111111111111011101000100010;
assign LUT_1[17476] = 32'b00000000000000001110100001101100;
assign LUT_1[17477] = 32'b00000000000000000111110011101000;
assign LUT_1[17478] = 32'b00000000000000001010001111111101;
assign LUT_1[17479] = 32'b00000000000000000011100001111001;
assign LUT_1[17480] = 32'b00000000000000000101110110001010;
assign LUT_1[17481] = 32'b11111111111111111111001000000110;
assign LUT_1[17482] = 32'b00000000000000000001100100011011;
assign LUT_1[17483] = 32'b11111111111111111010110110010111;
assign LUT_1[17484] = 32'b00000000000000001101101111100001;
assign LUT_1[17485] = 32'b00000000000000000111000001011101;
assign LUT_1[17486] = 32'b00000000000000001001011101110010;
assign LUT_1[17487] = 32'b00000000000000000010101111101110;
assign LUT_1[17488] = 32'b00000000000000001000100011110111;
assign LUT_1[17489] = 32'b00000000000000000001110101110011;
assign LUT_1[17490] = 32'b00000000000000000100010010001000;
assign LUT_1[17491] = 32'b11111111111111111101100100000100;
assign LUT_1[17492] = 32'b00000000000000010000011101001110;
assign LUT_1[17493] = 32'b00000000000000001001101111001010;
assign LUT_1[17494] = 32'b00000000000000001100001011011111;
assign LUT_1[17495] = 32'b00000000000000000101011101011011;
assign LUT_1[17496] = 32'b00000000000000000111110001101100;
assign LUT_1[17497] = 32'b00000000000000000001000011101000;
assign LUT_1[17498] = 32'b00000000000000000011011111111101;
assign LUT_1[17499] = 32'b11111111111111111100110001111001;
assign LUT_1[17500] = 32'b00000000000000001111101011000011;
assign LUT_1[17501] = 32'b00000000000000001000111100111111;
assign LUT_1[17502] = 32'b00000000000000001011011001010100;
assign LUT_1[17503] = 32'b00000000000000000100101011010000;
assign LUT_1[17504] = 32'b00000000000000000111100011010100;
assign LUT_1[17505] = 32'b00000000000000000000110101010000;
assign LUT_1[17506] = 32'b00000000000000000011010001100101;
assign LUT_1[17507] = 32'b11111111111111111100100011100001;
assign LUT_1[17508] = 32'b00000000000000001111011100101011;
assign LUT_1[17509] = 32'b00000000000000001000101110100111;
assign LUT_1[17510] = 32'b00000000000000001011001010111100;
assign LUT_1[17511] = 32'b00000000000000000100011100111000;
assign LUT_1[17512] = 32'b00000000000000000110110001001001;
assign LUT_1[17513] = 32'b00000000000000000000000011000101;
assign LUT_1[17514] = 32'b00000000000000000010011111011010;
assign LUT_1[17515] = 32'b11111111111111111011110001010110;
assign LUT_1[17516] = 32'b00000000000000001110101010100000;
assign LUT_1[17517] = 32'b00000000000000000111111100011100;
assign LUT_1[17518] = 32'b00000000000000001010011000110001;
assign LUT_1[17519] = 32'b00000000000000000011101010101101;
assign LUT_1[17520] = 32'b00000000000000001001011110110110;
assign LUT_1[17521] = 32'b00000000000000000010110000110010;
assign LUT_1[17522] = 32'b00000000000000000101001101000111;
assign LUT_1[17523] = 32'b11111111111111111110011111000011;
assign LUT_1[17524] = 32'b00000000000000010001011000001101;
assign LUT_1[17525] = 32'b00000000000000001010101010001001;
assign LUT_1[17526] = 32'b00000000000000001101000110011110;
assign LUT_1[17527] = 32'b00000000000000000110011000011010;
assign LUT_1[17528] = 32'b00000000000000001000101100101011;
assign LUT_1[17529] = 32'b00000000000000000001111110100111;
assign LUT_1[17530] = 32'b00000000000000000100011010111100;
assign LUT_1[17531] = 32'b11111111111111111101101100111000;
assign LUT_1[17532] = 32'b00000000000000010000100110000010;
assign LUT_1[17533] = 32'b00000000000000001001110111111110;
assign LUT_1[17534] = 32'b00000000000000001100010100010011;
assign LUT_1[17535] = 32'b00000000000000000101100110001111;
assign LUT_1[17536] = 32'b00000000000000000111101010110000;
assign LUT_1[17537] = 32'b00000000000000000000111100101100;
assign LUT_1[17538] = 32'b00000000000000000011011001000001;
assign LUT_1[17539] = 32'b11111111111111111100101010111101;
assign LUT_1[17540] = 32'b00000000000000001111100100000111;
assign LUT_1[17541] = 32'b00000000000000001000110110000011;
assign LUT_1[17542] = 32'b00000000000000001011010010011000;
assign LUT_1[17543] = 32'b00000000000000000100100100010100;
assign LUT_1[17544] = 32'b00000000000000000110111000100101;
assign LUT_1[17545] = 32'b00000000000000000000001010100001;
assign LUT_1[17546] = 32'b00000000000000000010100110110110;
assign LUT_1[17547] = 32'b11111111111111111011111000110010;
assign LUT_1[17548] = 32'b00000000000000001110110001111100;
assign LUT_1[17549] = 32'b00000000000000001000000011111000;
assign LUT_1[17550] = 32'b00000000000000001010100000001101;
assign LUT_1[17551] = 32'b00000000000000000011110010001001;
assign LUT_1[17552] = 32'b00000000000000001001100110010010;
assign LUT_1[17553] = 32'b00000000000000000010111000001110;
assign LUT_1[17554] = 32'b00000000000000000101010100100011;
assign LUT_1[17555] = 32'b11111111111111111110100110011111;
assign LUT_1[17556] = 32'b00000000000000010001011111101001;
assign LUT_1[17557] = 32'b00000000000000001010110001100101;
assign LUT_1[17558] = 32'b00000000000000001101001101111010;
assign LUT_1[17559] = 32'b00000000000000000110011111110110;
assign LUT_1[17560] = 32'b00000000000000001000110100000111;
assign LUT_1[17561] = 32'b00000000000000000010000110000011;
assign LUT_1[17562] = 32'b00000000000000000100100010011000;
assign LUT_1[17563] = 32'b11111111111111111101110100010100;
assign LUT_1[17564] = 32'b00000000000000010000101101011110;
assign LUT_1[17565] = 32'b00000000000000001001111111011010;
assign LUT_1[17566] = 32'b00000000000000001100011011101111;
assign LUT_1[17567] = 32'b00000000000000000101101101101011;
assign LUT_1[17568] = 32'b00000000000000001000100101101111;
assign LUT_1[17569] = 32'b00000000000000000001110111101011;
assign LUT_1[17570] = 32'b00000000000000000100010100000000;
assign LUT_1[17571] = 32'b11111111111111111101100101111100;
assign LUT_1[17572] = 32'b00000000000000010000011111000110;
assign LUT_1[17573] = 32'b00000000000000001001110001000010;
assign LUT_1[17574] = 32'b00000000000000001100001101010111;
assign LUT_1[17575] = 32'b00000000000000000101011111010011;
assign LUT_1[17576] = 32'b00000000000000000111110011100100;
assign LUT_1[17577] = 32'b00000000000000000001000101100000;
assign LUT_1[17578] = 32'b00000000000000000011100001110101;
assign LUT_1[17579] = 32'b11111111111111111100110011110001;
assign LUT_1[17580] = 32'b00000000000000001111101100111011;
assign LUT_1[17581] = 32'b00000000000000001000111110110111;
assign LUT_1[17582] = 32'b00000000000000001011011011001100;
assign LUT_1[17583] = 32'b00000000000000000100101101001000;
assign LUT_1[17584] = 32'b00000000000000001010100001010001;
assign LUT_1[17585] = 32'b00000000000000000011110011001101;
assign LUT_1[17586] = 32'b00000000000000000110001111100010;
assign LUT_1[17587] = 32'b11111111111111111111100001011110;
assign LUT_1[17588] = 32'b00000000000000010010011010101000;
assign LUT_1[17589] = 32'b00000000000000001011101100100100;
assign LUT_1[17590] = 32'b00000000000000001110001000111001;
assign LUT_1[17591] = 32'b00000000000000000111011010110101;
assign LUT_1[17592] = 32'b00000000000000001001101111000110;
assign LUT_1[17593] = 32'b00000000000000000011000001000010;
assign LUT_1[17594] = 32'b00000000000000000101011101010111;
assign LUT_1[17595] = 32'b11111111111111111110101111010011;
assign LUT_1[17596] = 32'b00000000000000010001101000011101;
assign LUT_1[17597] = 32'b00000000000000001010111010011001;
assign LUT_1[17598] = 32'b00000000000000001101010110101110;
assign LUT_1[17599] = 32'b00000000000000000110101000101010;
assign LUT_1[17600] = 32'b00000000000000001001101000011000;
assign LUT_1[17601] = 32'b00000000000000000010111010010100;
assign LUT_1[17602] = 32'b00000000000000000101010110101001;
assign LUT_1[17603] = 32'b11111111111111111110101000100101;
assign LUT_1[17604] = 32'b00000000000000010001100001101111;
assign LUT_1[17605] = 32'b00000000000000001010110011101011;
assign LUT_1[17606] = 32'b00000000000000001101010000000000;
assign LUT_1[17607] = 32'b00000000000000000110100001111100;
assign LUT_1[17608] = 32'b00000000000000001000110110001101;
assign LUT_1[17609] = 32'b00000000000000000010001000001001;
assign LUT_1[17610] = 32'b00000000000000000100100100011110;
assign LUT_1[17611] = 32'b11111111111111111101110110011010;
assign LUT_1[17612] = 32'b00000000000000010000101111100100;
assign LUT_1[17613] = 32'b00000000000000001010000001100000;
assign LUT_1[17614] = 32'b00000000000000001100011101110101;
assign LUT_1[17615] = 32'b00000000000000000101101111110001;
assign LUT_1[17616] = 32'b00000000000000001011100011111010;
assign LUT_1[17617] = 32'b00000000000000000100110101110110;
assign LUT_1[17618] = 32'b00000000000000000111010010001011;
assign LUT_1[17619] = 32'b00000000000000000000100100000111;
assign LUT_1[17620] = 32'b00000000000000010011011101010001;
assign LUT_1[17621] = 32'b00000000000000001100101111001101;
assign LUT_1[17622] = 32'b00000000000000001111001011100010;
assign LUT_1[17623] = 32'b00000000000000001000011101011110;
assign LUT_1[17624] = 32'b00000000000000001010110001101111;
assign LUT_1[17625] = 32'b00000000000000000100000011101011;
assign LUT_1[17626] = 32'b00000000000000000110100000000000;
assign LUT_1[17627] = 32'b11111111111111111111110001111100;
assign LUT_1[17628] = 32'b00000000000000010010101011000110;
assign LUT_1[17629] = 32'b00000000000000001011111101000010;
assign LUT_1[17630] = 32'b00000000000000001110011001010111;
assign LUT_1[17631] = 32'b00000000000000000111101011010011;
assign LUT_1[17632] = 32'b00000000000000001010100011010111;
assign LUT_1[17633] = 32'b00000000000000000011110101010011;
assign LUT_1[17634] = 32'b00000000000000000110010001101000;
assign LUT_1[17635] = 32'b11111111111111111111100011100100;
assign LUT_1[17636] = 32'b00000000000000010010011100101110;
assign LUT_1[17637] = 32'b00000000000000001011101110101010;
assign LUT_1[17638] = 32'b00000000000000001110001010111111;
assign LUT_1[17639] = 32'b00000000000000000111011100111011;
assign LUT_1[17640] = 32'b00000000000000001001110001001100;
assign LUT_1[17641] = 32'b00000000000000000011000011001000;
assign LUT_1[17642] = 32'b00000000000000000101011111011101;
assign LUT_1[17643] = 32'b11111111111111111110110001011001;
assign LUT_1[17644] = 32'b00000000000000010001101010100011;
assign LUT_1[17645] = 32'b00000000000000001010111100011111;
assign LUT_1[17646] = 32'b00000000000000001101011000110100;
assign LUT_1[17647] = 32'b00000000000000000110101010110000;
assign LUT_1[17648] = 32'b00000000000000001100011110111001;
assign LUT_1[17649] = 32'b00000000000000000101110000110101;
assign LUT_1[17650] = 32'b00000000000000001000001101001010;
assign LUT_1[17651] = 32'b00000000000000000001011111000110;
assign LUT_1[17652] = 32'b00000000000000010100011000010000;
assign LUT_1[17653] = 32'b00000000000000001101101010001100;
assign LUT_1[17654] = 32'b00000000000000010000000110100001;
assign LUT_1[17655] = 32'b00000000000000001001011000011101;
assign LUT_1[17656] = 32'b00000000000000001011101100101110;
assign LUT_1[17657] = 32'b00000000000000000100111110101010;
assign LUT_1[17658] = 32'b00000000000000000111011010111111;
assign LUT_1[17659] = 32'b00000000000000000000101100111011;
assign LUT_1[17660] = 32'b00000000000000010011100110000101;
assign LUT_1[17661] = 32'b00000000000000001100111000000001;
assign LUT_1[17662] = 32'b00000000000000001111010100010110;
assign LUT_1[17663] = 32'b00000000000000001000100110010010;
assign LUT_1[17664] = 32'b00000000000000000010011110111001;
assign LUT_1[17665] = 32'b11111111111111111011110000110101;
assign LUT_1[17666] = 32'b11111111111111111110001101001010;
assign LUT_1[17667] = 32'b11111111111111110111011111000110;
assign LUT_1[17668] = 32'b00000000000000001010011000010000;
assign LUT_1[17669] = 32'b00000000000000000011101010001100;
assign LUT_1[17670] = 32'b00000000000000000110000110100001;
assign LUT_1[17671] = 32'b11111111111111111111011000011101;
assign LUT_1[17672] = 32'b00000000000000000001101100101110;
assign LUT_1[17673] = 32'b11111111111111111010111110101010;
assign LUT_1[17674] = 32'b11111111111111111101011010111111;
assign LUT_1[17675] = 32'b11111111111111110110101100111011;
assign LUT_1[17676] = 32'b00000000000000001001100110000101;
assign LUT_1[17677] = 32'b00000000000000000010111000000001;
assign LUT_1[17678] = 32'b00000000000000000101010100010110;
assign LUT_1[17679] = 32'b11111111111111111110100110010010;
assign LUT_1[17680] = 32'b00000000000000000100011010011011;
assign LUT_1[17681] = 32'b11111111111111111101101100010111;
assign LUT_1[17682] = 32'b00000000000000000000001000101100;
assign LUT_1[17683] = 32'b11111111111111111001011010101000;
assign LUT_1[17684] = 32'b00000000000000001100010011110010;
assign LUT_1[17685] = 32'b00000000000000000101100101101110;
assign LUT_1[17686] = 32'b00000000000000001000000010000011;
assign LUT_1[17687] = 32'b00000000000000000001010011111111;
assign LUT_1[17688] = 32'b00000000000000000011101000010000;
assign LUT_1[17689] = 32'b11111111111111111100111010001100;
assign LUT_1[17690] = 32'b11111111111111111111010110100001;
assign LUT_1[17691] = 32'b11111111111111111000101000011101;
assign LUT_1[17692] = 32'b00000000000000001011100001100111;
assign LUT_1[17693] = 32'b00000000000000000100110011100011;
assign LUT_1[17694] = 32'b00000000000000000111001111111000;
assign LUT_1[17695] = 32'b00000000000000000000100001110100;
assign LUT_1[17696] = 32'b00000000000000000011011001111000;
assign LUT_1[17697] = 32'b11111111111111111100101011110100;
assign LUT_1[17698] = 32'b11111111111111111111001000001001;
assign LUT_1[17699] = 32'b11111111111111111000011010000101;
assign LUT_1[17700] = 32'b00000000000000001011010011001111;
assign LUT_1[17701] = 32'b00000000000000000100100101001011;
assign LUT_1[17702] = 32'b00000000000000000111000001100000;
assign LUT_1[17703] = 32'b00000000000000000000010011011100;
assign LUT_1[17704] = 32'b00000000000000000010100111101101;
assign LUT_1[17705] = 32'b11111111111111111011111001101001;
assign LUT_1[17706] = 32'b11111111111111111110010101111110;
assign LUT_1[17707] = 32'b11111111111111110111100111111010;
assign LUT_1[17708] = 32'b00000000000000001010100001000100;
assign LUT_1[17709] = 32'b00000000000000000011110011000000;
assign LUT_1[17710] = 32'b00000000000000000110001111010101;
assign LUT_1[17711] = 32'b11111111111111111111100001010001;
assign LUT_1[17712] = 32'b00000000000000000101010101011010;
assign LUT_1[17713] = 32'b11111111111111111110100111010110;
assign LUT_1[17714] = 32'b00000000000000000001000011101011;
assign LUT_1[17715] = 32'b11111111111111111010010101100111;
assign LUT_1[17716] = 32'b00000000000000001101001110110001;
assign LUT_1[17717] = 32'b00000000000000000110100000101101;
assign LUT_1[17718] = 32'b00000000000000001000111101000010;
assign LUT_1[17719] = 32'b00000000000000000010001110111110;
assign LUT_1[17720] = 32'b00000000000000000100100011001111;
assign LUT_1[17721] = 32'b11111111111111111101110101001011;
assign LUT_1[17722] = 32'b00000000000000000000010001100000;
assign LUT_1[17723] = 32'b11111111111111111001100011011100;
assign LUT_1[17724] = 32'b00000000000000001100011100100110;
assign LUT_1[17725] = 32'b00000000000000000101101110100010;
assign LUT_1[17726] = 32'b00000000000000001000001010110111;
assign LUT_1[17727] = 32'b00000000000000000001011100110011;
assign LUT_1[17728] = 32'b00000000000000000100011100100001;
assign LUT_1[17729] = 32'b11111111111111111101101110011101;
assign LUT_1[17730] = 32'b00000000000000000000001010110010;
assign LUT_1[17731] = 32'b11111111111111111001011100101110;
assign LUT_1[17732] = 32'b00000000000000001100010101111000;
assign LUT_1[17733] = 32'b00000000000000000101100111110100;
assign LUT_1[17734] = 32'b00000000000000001000000100001001;
assign LUT_1[17735] = 32'b00000000000000000001010110000101;
assign LUT_1[17736] = 32'b00000000000000000011101010010110;
assign LUT_1[17737] = 32'b11111111111111111100111100010010;
assign LUT_1[17738] = 32'b11111111111111111111011000100111;
assign LUT_1[17739] = 32'b11111111111111111000101010100011;
assign LUT_1[17740] = 32'b00000000000000001011100011101101;
assign LUT_1[17741] = 32'b00000000000000000100110101101001;
assign LUT_1[17742] = 32'b00000000000000000111010001111110;
assign LUT_1[17743] = 32'b00000000000000000000100011111010;
assign LUT_1[17744] = 32'b00000000000000000110011000000011;
assign LUT_1[17745] = 32'b11111111111111111111101001111111;
assign LUT_1[17746] = 32'b00000000000000000010000110010100;
assign LUT_1[17747] = 32'b11111111111111111011011000010000;
assign LUT_1[17748] = 32'b00000000000000001110010001011010;
assign LUT_1[17749] = 32'b00000000000000000111100011010110;
assign LUT_1[17750] = 32'b00000000000000001001111111101011;
assign LUT_1[17751] = 32'b00000000000000000011010001100111;
assign LUT_1[17752] = 32'b00000000000000000101100101111000;
assign LUT_1[17753] = 32'b11111111111111111110110111110100;
assign LUT_1[17754] = 32'b00000000000000000001010100001001;
assign LUT_1[17755] = 32'b11111111111111111010100110000101;
assign LUT_1[17756] = 32'b00000000000000001101011111001111;
assign LUT_1[17757] = 32'b00000000000000000110110001001011;
assign LUT_1[17758] = 32'b00000000000000001001001101100000;
assign LUT_1[17759] = 32'b00000000000000000010011111011100;
assign LUT_1[17760] = 32'b00000000000000000101010111100000;
assign LUT_1[17761] = 32'b11111111111111111110101001011100;
assign LUT_1[17762] = 32'b00000000000000000001000101110001;
assign LUT_1[17763] = 32'b11111111111111111010010111101101;
assign LUT_1[17764] = 32'b00000000000000001101010000110111;
assign LUT_1[17765] = 32'b00000000000000000110100010110011;
assign LUT_1[17766] = 32'b00000000000000001000111111001000;
assign LUT_1[17767] = 32'b00000000000000000010010001000100;
assign LUT_1[17768] = 32'b00000000000000000100100101010101;
assign LUT_1[17769] = 32'b11111111111111111101110111010001;
assign LUT_1[17770] = 32'b00000000000000000000010011100110;
assign LUT_1[17771] = 32'b11111111111111111001100101100010;
assign LUT_1[17772] = 32'b00000000000000001100011110101100;
assign LUT_1[17773] = 32'b00000000000000000101110000101000;
assign LUT_1[17774] = 32'b00000000000000001000001100111101;
assign LUT_1[17775] = 32'b00000000000000000001011110111001;
assign LUT_1[17776] = 32'b00000000000000000111010011000010;
assign LUT_1[17777] = 32'b00000000000000000000100100111110;
assign LUT_1[17778] = 32'b00000000000000000011000001010011;
assign LUT_1[17779] = 32'b11111111111111111100010011001111;
assign LUT_1[17780] = 32'b00000000000000001111001100011001;
assign LUT_1[17781] = 32'b00000000000000001000011110010101;
assign LUT_1[17782] = 32'b00000000000000001010111010101010;
assign LUT_1[17783] = 32'b00000000000000000100001100100110;
assign LUT_1[17784] = 32'b00000000000000000110100000110111;
assign LUT_1[17785] = 32'b11111111111111111111110010110011;
assign LUT_1[17786] = 32'b00000000000000000010001111001000;
assign LUT_1[17787] = 32'b11111111111111111011100001000100;
assign LUT_1[17788] = 32'b00000000000000001110011010001110;
assign LUT_1[17789] = 32'b00000000000000000111101100001010;
assign LUT_1[17790] = 32'b00000000000000001010001000011111;
assign LUT_1[17791] = 32'b00000000000000000011011010011011;
assign LUT_1[17792] = 32'b00000000000000000101011110111100;
assign LUT_1[17793] = 32'b11111111111111111110110000111000;
assign LUT_1[17794] = 32'b00000000000000000001001101001101;
assign LUT_1[17795] = 32'b11111111111111111010011111001001;
assign LUT_1[17796] = 32'b00000000000000001101011000010011;
assign LUT_1[17797] = 32'b00000000000000000110101010001111;
assign LUT_1[17798] = 32'b00000000000000001001000110100100;
assign LUT_1[17799] = 32'b00000000000000000010011000100000;
assign LUT_1[17800] = 32'b00000000000000000100101100110001;
assign LUT_1[17801] = 32'b11111111111111111101111110101101;
assign LUT_1[17802] = 32'b00000000000000000000011011000010;
assign LUT_1[17803] = 32'b11111111111111111001101100111110;
assign LUT_1[17804] = 32'b00000000000000001100100110001000;
assign LUT_1[17805] = 32'b00000000000000000101111000000100;
assign LUT_1[17806] = 32'b00000000000000001000010100011001;
assign LUT_1[17807] = 32'b00000000000000000001100110010101;
assign LUT_1[17808] = 32'b00000000000000000111011010011110;
assign LUT_1[17809] = 32'b00000000000000000000101100011010;
assign LUT_1[17810] = 32'b00000000000000000011001000101111;
assign LUT_1[17811] = 32'b11111111111111111100011010101011;
assign LUT_1[17812] = 32'b00000000000000001111010011110101;
assign LUT_1[17813] = 32'b00000000000000001000100101110001;
assign LUT_1[17814] = 32'b00000000000000001011000010000110;
assign LUT_1[17815] = 32'b00000000000000000100010100000010;
assign LUT_1[17816] = 32'b00000000000000000110101000010011;
assign LUT_1[17817] = 32'b11111111111111111111111010001111;
assign LUT_1[17818] = 32'b00000000000000000010010110100100;
assign LUT_1[17819] = 32'b11111111111111111011101000100000;
assign LUT_1[17820] = 32'b00000000000000001110100001101010;
assign LUT_1[17821] = 32'b00000000000000000111110011100110;
assign LUT_1[17822] = 32'b00000000000000001010001111111011;
assign LUT_1[17823] = 32'b00000000000000000011100001110111;
assign LUT_1[17824] = 32'b00000000000000000110011001111011;
assign LUT_1[17825] = 32'b11111111111111111111101011110111;
assign LUT_1[17826] = 32'b00000000000000000010001000001100;
assign LUT_1[17827] = 32'b11111111111111111011011010001000;
assign LUT_1[17828] = 32'b00000000000000001110010011010010;
assign LUT_1[17829] = 32'b00000000000000000111100101001110;
assign LUT_1[17830] = 32'b00000000000000001010000001100011;
assign LUT_1[17831] = 32'b00000000000000000011010011011111;
assign LUT_1[17832] = 32'b00000000000000000101100111110000;
assign LUT_1[17833] = 32'b11111111111111111110111001101100;
assign LUT_1[17834] = 32'b00000000000000000001010110000001;
assign LUT_1[17835] = 32'b11111111111111111010100111111101;
assign LUT_1[17836] = 32'b00000000000000001101100001000111;
assign LUT_1[17837] = 32'b00000000000000000110110011000011;
assign LUT_1[17838] = 32'b00000000000000001001001111011000;
assign LUT_1[17839] = 32'b00000000000000000010100001010100;
assign LUT_1[17840] = 32'b00000000000000001000010101011101;
assign LUT_1[17841] = 32'b00000000000000000001100111011001;
assign LUT_1[17842] = 32'b00000000000000000100000011101110;
assign LUT_1[17843] = 32'b11111111111111111101010101101010;
assign LUT_1[17844] = 32'b00000000000000010000001110110100;
assign LUT_1[17845] = 32'b00000000000000001001100000110000;
assign LUT_1[17846] = 32'b00000000000000001011111101000101;
assign LUT_1[17847] = 32'b00000000000000000101001111000001;
assign LUT_1[17848] = 32'b00000000000000000111100011010010;
assign LUT_1[17849] = 32'b00000000000000000000110101001110;
assign LUT_1[17850] = 32'b00000000000000000011010001100011;
assign LUT_1[17851] = 32'b11111111111111111100100011011111;
assign LUT_1[17852] = 32'b00000000000000001111011100101001;
assign LUT_1[17853] = 32'b00000000000000001000101110100101;
assign LUT_1[17854] = 32'b00000000000000001011001010111010;
assign LUT_1[17855] = 32'b00000000000000000100011100110110;
assign LUT_1[17856] = 32'b00000000000000000111011100100100;
assign LUT_1[17857] = 32'b00000000000000000000101110100000;
assign LUT_1[17858] = 32'b00000000000000000011001010110101;
assign LUT_1[17859] = 32'b11111111111111111100011100110001;
assign LUT_1[17860] = 32'b00000000000000001111010101111011;
assign LUT_1[17861] = 32'b00000000000000001000100111110111;
assign LUT_1[17862] = 32'b00000000000000001011000100001100;
assign LUT_1[17863] = 32'b00000000000000000100010110001000;
assign LUT_1[17864] = 32'b00000000000000000110101010011001;
assign LUT_1[17865] = 32'b11111111111111111111111100010101;
assign LUT_1[17866] = 32'b00000000000000000010011000101010;
assign LUT_1[17867] = 32'b11111111111111111011101010100110;
assign LUT_1[17868] = 32'b00000000000000001110100011110000;
assign LUT_1[17869] = 32'b00000000000000000111110101101100;
assign LUT_1[17870] = 32'b00000000000000001010010010000001;
assign LUT_1[17871] = 32'b00000000000000000011100011111101;
assign LUT_1[17872] = 32'b00000000000000001001011000000110;
assign LUT_1[17873] = 32'b00000000000000000010101010000010;
assign LUT_1[17874] = 32'b00000000000000000101000110010111;
assign LUT_1[17875] = 32'b11111111111111111110011000010011;
assign LUT_1[17876] = 32'b00000000000000010001010001011101;
assign LUT_1[17877] = 32'b00000000000000001010100011011001;
assign LUT_1[17878] = 32'b00000000000000001100111111101110;
assign LUT_1[17879] = 32'b00000000000000000110010001101010;
assign LUT_1[17880] = 32'b00000000000000001000100101111011;
assign LUT_1[17881] = 32'b00000000000000000001110111110111;
assign LUT_1[17882] = 32'b00000000000000000100010100001100;
assign LUT_1[17883] = 32'b11111111111111111101100110001000;
assign LUT_1[17884] = 32'b00000000000000010000011111010010;
assign LUT_1[17885] = 32'b00000000000000001001110001001110;
assign LUT_1[17886] = 32'b00000000000000001100001101100011;
assign LUT_1[17887] = 32'b00000000000000000101011111011111;
assign LUT_1[17888] = 32'b00000000000000001000010111100011;
assign LUT_1[17889] = 32'b00000000000000000001101001011111;
assign LUT_1[17890] = 32'b00000000000000000100000101110100;
assign LUT_1[17891] = 32'b11111111111111111101010111110000;
assign LUT_1[17892] = 32'b00000000000000010000010000111010;
assign LUT_1[17893] = 32'b00000000000000001001100010110110;
assign LUT_1[17894] = 32'b00000000000000001011111111001011;
assign LUT_1[17895] = 32'b00000000000000000101010001000111;
assign LUT_1[17896] = 32'b00000000000000000111100101011000;
assign LUT_1[17897] = 32'b00000000000000000000110111010100;
assign LUT_1[17898] = 32'b00000000000000000011010011101001;
assign LUT_1[17899] = 32'b11111111111111111100100101100101;
assign LUT_1[17900] = 32'b00000000000000001111011110101111;
assign LUT_1[17901] = 32'b00000000000000001000110000101011;
assign LUT_1[17902] = 32'b00000000000000001011001101000000;
assign LUT_1[17903] = 32'b00000000000000000100011110111100;
assign LUT_1[17904] = 32'b00000000000000001010010011000101;
assign LUT_1[17905] = 32'b00000000000000000011100101000001;
assign LUT_1[17906] = 32'b00000000000000000110000001010110;
assign LUT_1[17907] = 32'b11111111111111111111010011010010;
assign LUT_1[17908] = 32'b00000000000000010010001100011100;
assign LUT_1[17909] = 32'b00000000000000001011011110011000;
assign LUT_1[17910] = 32'b00000000000000001101111010101101;
assign LUT_1[17911] = 32'b00000000000000000111001100101001;
assign LUT_1[17912] = 32'b00000000000000001001100000111010;
assign LUT_1[17913] = 32'b00000000000000000010110010110110;
assign LUT_1[17914] = 32'b00000000000000000101001111001011;
assign LUT_1[17915] = 32'b11111111111111111110100001000111;
assign LUT_1[17916] = 32'b00000000000000010001011010010001;
assign LUT_1[17917] = 32'b00000000000000001010101100001101;
assign LUT_1[17918] = 32'b00000000000000001101001000100010;
assign LUT_1[17919] = 32'b00000000000000000110011010011110;
assign LUT_1[17920] = 32'b11111111111111111110011001001010;
assign LUT_1[17921] = 32'b11111111111111110111101011000110;
assign LUT_1[17922] = 32'b11111111111111111010000111011011;
assign LUT_1[17923] = 32'b11111111111111110011011001010111;
assign LUT_1[17924] = 32'b00000000000000000110010010100001;
assign LUT_1[17925] = 32'b11111111111111111111100100011101;
assign LUT_1[17926] = 32'b00000000000000000010000000110010;
assign LUT_1[17927] = 32'b11111111111111111011010010101110;
assign LUT_1[17928] = 32'b11111111111111111101100110111111;
assign LUT_1[17929] = 32'b11111111111111110110111000111011;
assign LUT_1[17930] = 32'b11111111111111111001010101010000;
assign LUT_1[17931] = 32'b11111111111111110010100111001100;
assign LUT_1[17932] = 32'b00000000000000000101100000010110;
assign LUT_1[17933] = 32'b11111111111111111110110010010010;
assign LUT_1[17934] = 32'b00000000000000000001001110100111;
assign LUT_1[17935] = 32'b11111111111111111010100000100011;
assign LUT_1[17936] = 32'b00000000000000000000010100101100;
assign LUT_1[17937] = 32'b11111111111111111001100110101000;
assign LUT_1[17938] = 32'b11111111111111111100000010111101;
assign LUT_1[17939] = 32'b11111111111111110101010100111001;
assign LUT_1[17940] = 32'b00000000000000001000001110000011;
assign LUT_1[17941] = 32'b00000000000000000001011111111111;
assign LUT_1[17942] = 32'b00000000000000000011111100010100;
assign LUT_1[17943] = 32'b11111111111111111101001110010000;
assign LUT_1[17944] = 32'b11111111111111111111100010100001;
assign LUT_1[17945] = 32'b11111111111111111000110100011101;
assign LUT_1[17946] = 32'b11111111111111111011010000110010;
assign LUT_1[17947] = 32'b11111111111111110100100010101110;
assign LUT_1[17948] = 32'b00000000000000000111011011111000;
assign LUT_1[17949] = 32'b00000000000000000000101101110100;
assign LUT_1[17950] = 32'b00000000000000000011001010001001;
assign LUT_1[17951] = 32'b11111111111111111100011100000101;
assign LUT_1[17952] = 32'b11111111111111111111010100001001;
assign LUT_1[17953] = 32'b11111111111111111000100110000101;
assign LUT_1[17954] = 32'b11111111111111111011000010011010;
assign LUT_1[17955] = 32'b11111111111111110100010100010110;
assign LUT_1[17956] = 32'b00000000000000000111001101100000;
assign LUT_1[17957] = 32'b00000000000000000000011111011100;
assign LUT_1[17958] = 32'b00000000000000000010111011110001;
assign LUT_1[17959] = 32'b11111111111111111100001101101101;
assign LUT_1[17960] = 32'b11111111111111111110100001111110;
assign LUT_1[17961] = 32'b11111111111111110111110011111010;
assign LUT_1[17962] = 32'b11111111111111111010010000001111;
assign LUT_1[17963] = 32'b11111111111111110011100010001011;
assign LUT_1[17964] = 32'b00000000000000000110011011010101;
assign LUT_1[17965] = 32'b11111111111111111111101101010001;
assign LUT_1[17966] = 32'b00000000000000000010001001100110;
assign LUT_1[17967] = 32'b11111111111111111011011011100010;
assign LUT_1[17968] = 32'b00000000000000000001001111101011;
assign LUT_1[17969] = 32'b11111111111111111010100001100111;
assign LUT_1[17970] = 32'b11111111111111111100111101111100;
assign LUT_1[17971] = 32'b11111111111111110110001111111000;
assign LUT_1[17972] = 32'b00000000000000001001001001000010;
assign LUT_1[17973] = 32'b00000000000000000010011010111110;
assign LUT_1[17974] = 32'b00000000000000000100110111010011;
assign LUT_1[17975] = 32'b11111111111111111110001001001111;
assign LUT_1[17976] = 32'b00000000000000000000011101100000;
assign LUT_1[17977] = 32'b11111111111111111001101111011100;
assign LUT_1[17978] = 32'b11111111111111111100001011110001;
assign LUT_1[17979] = 32'b11111111111111110101011101101101;
assign LUT_1[17980] = 32'b00000000000000001000010110110111;
assign LUT_1[17981] = 32'b00000000000000000001101000110011;
assign LUT_1[17982] = 32'b00000000000000000100000101001000;
assign LUT_1[17983] = 32'b11111111111111111101010111000100;
assign LUT_1[17984] = 32'b00000000000000000000010110110010;
assign LUT_1[17985] = 32'b11111111111111111001101000101110;
assign LUT_1[17986] = 32'b11111111111111111100000101000011;
assign LUT_1[17987] = 32'b11111111111111110101010110111111;
assign LUT_1[17988] = 32'b00000000000000001000010000001001;
assign LUT_1[17989] = 32'b00000000000000000001100010000101;
assign LUT_1[17990] = 32'b00000000000000000011111110011010;
assign LUT_1[17991] = 32'b11111111111111111101010000010110;
assign LUT_1[17992] = 32'b11111111111111111111100100100111;
assign LUT_1[17993] = 32'b11111111111111111000110110100011;
assign LUT_1[17994] = 32'b11111111111111111011010010111000;
assign LUT_1[17995] = 32'b11111111111111110100100100110100;
assign LUT_1[17996] = 32'b00000000000000000111011101111110;
assign LUT_1[17997] = 32'b00000000000000000000101111111010;
assign LUT_1[17998] = 32'b00000000000000000011001100001111;
assign LUT_1[17999] = 32'b11111111111111111100011110001011;
assign LUT_1[18000] = 32'b00000000000000000010010010010100;
assign LUT_1[18001] = 32'b11111111111111111011100100010000;
assign LUT_1[18002] = 32'b11111111111111111110000000100101;
assign LUT_1[18003] = 32'b11111111111111110111010010100001;
assign LUT_1[18004] = 32'b00000000000000001010001011101011;
assign LUT_1[18005] = 32'b00000000000000000011011101100111;
assign LUT_1[18006] = 32'b00000000000000000101111001111100;
assign LUT_1[18007] = 32'b11111111111111111111001011111000;
assign LUT_1[18008] = 32'b00000000000000000001100000001001;
assign LUT_1[18009] = 32'b11111111111111111010110010000101;
assign LUT_1[18010] = 32'b11111111111111111101001110011010;
assign LUT_1[18011] = 32'b11111111111111110110100000010110;
assign LUT_1[18012] = 32'b00000000000000001001011001100000;
assign LUT_1[18013] = 32'b00000000000000000010101011011100;
assign LUT_1[18014] = 32'b00000000000000000101000111110001;
assign LUT_1[18015] = 32'b11111111111111111110011001101101;
assign LUT_1[18016] = 32'b00000000000000000001010001110001;
assign LUT_1[18017] = 32'b11111111111111111010100011101101;
assign LUT_1[18018] = 32'b11111111111111111101000000000010;
assign LUT_1[18019] = 32'b11111111111111110110010001111110;
assign LUT_1[18020] = 32'b00000000000000001001001011001000;
assign LUT_1[18021] = 32'b00000000000000000010011101000100;
assign LUT_1[18022] = 32'b00000000000000000100111001011001;
assign LUT_1[18023] = 32'b11111111111111111110001011010101;
assign LUT_1[18024] = 32'b00000000000000000000011111100110;
assign LUT_1[18025] = 32'b11111111111111111001110001100010;
assign LUT_1[18026] = 32'b11111111111111111100001101110111;
assign LUT_1[18027] = 32'b11111111111111110101011111110011;
assign LUT_1[18028] = 32'b00000000000000001000011000111101;
assign LUT_1[18029] = 32'b00000000000000000001101010111001;
assign LUT_1[18030] = 32'b00000000000000000100000111001110;
assign LUT_1[18031] = 32'b11111111111111111101011001001010;
assign LUT_1[18032] = 32'b00000000000000000011001101010011;
assign LUT_1[18033] = 32'b11111111111111111100011111001111;
assign LUT_1[18034] = 32'b11111111111111111110111011100100;
assign LUT_1[18035] = 32'b11111111111111111000001101100000;
assign LUT_1[18036] = 32'b00000000000000001011000110101010;
assign LUT_1[18037] = 32'b00000000000000000100011000100110;
assign LUT_1[18038] = 32'b00000000000000000110110100111011;
assign LUT_1[18039] = 32'b00000000000000000000000110110111;
assign LUT_1[18040] = 32'b00000000000000000010011011001000;
assign LUT_1[18041] = 32'b11111111111111111011101101000100;
assign LUT_1[18042] = 32'b11111111111111111110001001011001;
assign LUT_1[18043] = 32'b11111111111111110111011011010101;
assign LUT_1[18044] = 32'b00000000000000001010010100011111;
assign LUT_1[18045] = 32'b00000000000000000011100110011011;
assign LUT_1[18046] = 32'b00000000000000000110000010110000;
assign LUT_1[18047] = 32'b11111111111111111111010100101100;
assign LUT_1[18048] = 32'b00000000000000000001011001001101;
assign LUT_1[18049] = 32'b11111111111111111010101011001001;
assign LUT_1[18050] = 32'b11111111111111111101000111011110;
assign LUT_1[18051] = 32'b11111111111111110110011001011010;
assign LUT_1[18052] = 32'b00000000000000001001010010100100;
assign LUT_1[18053] = 32'b00000000000000000010100100100000;
assign LUT_1[18054] = 32'b00000000000000000101000000110101;
assign LUT_1[18055] = 32'b11111111111111111110010010110001;
assign LUT_1[18056] = 32'b00000000000000000000100111000010;
assign LUT_1[18057] = 32'b11111111111111111001111000111110;
assign LUT_1[18058] = 32'b11111111111111111100010101010011;
assign LUT_1[18059] = 32'b11111111111111110101100111001111;
assign LUT_1[18060] = 32'b00000000000000001000100000011001;
assign LUT_1[18061] = 32'b00000000000000000001110010010101;
assign LUT_1[18062] = 32'b00000000000000000100001110101010;
assign LUT_1[18063] = 32'b11111111111111111101100000100110;
assign LUT_1[18064] = 32'b00000000000000000011010100101111;
assign LUT_1[18065] = 32'b11111111111111111100100110101011;
assign LUT_1[18066] = 32'b11111111111111111111000011000000;
assign LUT_1[18067] = 32'b11111111111111111000010100111100;
assign LUT_1[18068] = 32'b00000000000000001011001110000110;
assign LUT_1[18069] = 32'b00000000000000000100100000000010;
assign LUT_1[18070] = 32'b00000000000000000110111100010111;
assign LUT_1[18071] = 32'b00000000000000000000001110010011;
assign LUT_1[18072] = 32'b00000000000000000010100010100100;
assign LUT_1[18073] = 32'b11111111111111111011110100100000;
assign LUT_1[18074] = 32'b11111111111111111110010000110101;
assign LUT_1[18075] = 32'b11111111111111110111100010110001;
assign LUT_1[18076] = 32'b00000000000000001010011011111011;
assign LUT_1[18077] = 32'b00000000000000000011101101110111;
assign LUT_1[18078] = 32'b00000000000000000110001010001100;
assign LUT_1[18079] = 32'b11111111111111111111011100001000;
assign LUT_1[18080] = 32'b00000000000000000010010100001100;
assign LUT_1[18081] = 32'b11111111111111111011100110001000;
assign LUT_1[18082] = 32'b11111111111111111110000010011101;
assign LUT_1[18083] = 32'b11111111111111110111010100011001;
assign LUT_1[18084] = 32'b00000000000000001010001101100011;
assign LUT_1[18085] = 32'b00000000000000000011011111011111;
assign LUT_1[18086] = 32'b00000000000000000101111011110100;
assign LUT_1[18087] = 32'b11111111111111111111001101110000;
assign LUT_1[18088] = 32'b00000000000000000001100010000001;
assign LUT_1[18089] = 32'b11111111111111111010110011111101;
assign LUT_1[18090] = 32'b11111111111111111101010000010010;
assign LUT_1[18091] = 32'b11111111111111110110100010001110;
assign LUT_1[18092] = 32'b00000000000000001001011011011000;
assign LUT_1[18093] = 32'b00000000000000000010101101010100;
assign LUT_1[18094] = 32'b00000000000000000101001001101001;
assign LUT_1[18095] = 32'b11111111111111111110011011100101;
assign LUT_1[18096] = 32'b00000000000000000100001111101110;
assign LUT_1[18097] = 32'b11111111111111111101100001101010;
assign LUT_1[18098] = 32'b11111111111111111111111101111111;
assign LUT_1[18099] = 32'b11111111111111111001001111111011;
assign LUT_1[18100] = 32'b00000000000000001100001001000101;
assign LUT_1[18101] = 32'b00000000000000000101011011000001;
assign LUT_1[18102] = 32'b00000000000000000111110111010110;
assign LUT_1[18103] = 32'b00000000000000000001001001010010;
assign LUT_1[18104] = 32'b00000000000000000011011101100011;
assign LUT_1[18105] = 32'b11111111111111111100101111011111;
assign LUT_1[18106] = 32'b11111111111111111111001011110100;
assign LUT_1[18107] = 32'b11111111111111111000011101110000;
assign LUT_1[18108] = 32'b00000000000000001011010110111010;
assign LUT_1[18109] = 32'b00000000000000000100101000110110;
assign LUT_1[18110] = 32'b00000000000000000111000101001011;
assign LUT_1[18111] = 32'b00000000000000000000010111000111;
assign LUT_1[18112] = 32'b00000000000000000011010110110101;
assign LUT_1[18113] = 32'b11111111111111111100101000110001;
assign LUT_1[18114] = 32'b11111111111111111111000101000110;
assign LUT_1[18115] = 32'b11111111111111111000010111000010;
assign LUT_1[18116] = 32'b00000000000000001011010000001100;
assign LUT_1[18117] = 32'b00000000000000000100100010001000;
assign LUT_1[18118] = 32'b00000000000000000110111110011101;
assign LUT_1[18119] = 32'b00000000000000000000010000011001;
assign LUT_1[18120] = 32'b00000000000000000010100100101010;
assign LUT_1[18121] = 32'b11111111111111111011110110100110;
assign LUT_1[18122] = 32'b11111111111111111110010010111011;
assign LUT_1[18123] = 32'b11111111111111110111100100110111;
assign LUT_1[18124] = 32'b00000000000000001010011110000001;
assign LUT_1[18125] = 32'b00000000000000000011101111111101;
assign LUT_1[18126] = 32'b00000000000000000110001100010010;
assign LUT_1[18127] = 32'b11111111111111111111011110001110;
assign LUT_1[18128] = 32'b00000000000000000101010010010111;
assign LUT_1[18129] = 32'b11111111111111111110100100010011;
assign LUT_1[18130] = 32'b00000000000000000001000000101000;
assign LUT_1[18131] = 32'b11111111111111111010010010100100;
assign LUT_1[18132] = 32'b00000000000000001101001011101110;
assign LUT_1[18133] = 32'b00000000000000000110011101101010;
assign LUT_1[18134] = 32'b00000000000000001000111001111111;
assign LUT_1[18135] = 32'b00000000000000000010001011111011;
assign LUT_1[18136] = 32'b00000000000000000100100000001100;
assign LUT_1[18137] = 32'b11111111111111111101110010001000;
assign LUT_1[18138] = 32'b00000000000000000000001110011101;
assign LUT_1[18139] = 32'b11111111111111111001100000011001;
assign LUT_1[18140] = 32'b00000000000000001100011001100011;
assign LUT_1[18141] = 32'b00000000000000000101101011011111;
assign LUT_1[18142] = 32'b00000000000000001000000111110100;
assign LUT_1[18143] = 32'b00000000000000000001011001110000;
assign LUT_1[18144] = 32'b00000000000000000100010001110100;
assign LUT_1[18145] = 32'b11111111111111111101100011110000;
assign LUT_1[18146] = 32'b00000000000000000000000000000101;
assign LUT_1[18147] = 32'b11111111111111111001010010000001;
assign LUT_1[18148] = 32'b00000000000000001100001011001011;
assign LUT_1[18149] = 32'b00000000000000000101011101000111;
assign LUT_1[18150] = 32'b00000000000000000111111001011100;
assign LUT_1[18151] = 32'b00000000000000000001001011011000;
assign LUT_1[18152] = 32'b00000000000000000011011111101001;
assign LUT_1[18153] = 32'b11111111111111111100110001100101;
assign LUT_1[18154] = 32'b11111111111111111111001101111010;
assign LUT_1[18155] = 32'b11111111111111111000011111110110;
assign LUT_1[18156] = 32'b00000000000000001011011001000000;
assign LUT_1[18157] = 32'b00000000000000000100101010111100;
assign LUT_1[18158] = 32'b00000000000000000111000111010001;
assign LUT_1[18159] = 32'b00000000000000000000011001001101;
assign LUT_1[18160] = 32'b00000000000000000110001101010110;
assign LUT_1[18161] = 32'b11111111111111111111011111010010;
assign LUT_1[18162] = 32'b00000000000000000001111011100111;
assign LUT_1[18163] = 32'b11111111111111111011001101100011;
assign LUT_1[18164] = 32'b00000000000000001110000110101101;
assign LUT_1[18165] = 32'b00000000000000000111011000101001;
assign LUT_1[18166] = 32'b00000000000000001001110100111110;
assign LUT_1[18167] = 32'b00000000000000000011000110111010;
assign LUT_1[18168] = 32'b00000000000000000101011011001011;
assign LUT_1[18169] = 32'b11111111111111111110101101000111;
assign LUT_1[18170] = 32'b00000000000000000001001001011100;
assign LUT_1[18171] = 32'b11111111111111111010011011011000;
assign LUT_1[18172] = 32'b00000000000000001101010100100010;
assign LUT_1[18173] = 32'b00000000000000000110100110011110;
assign LUT_1[18174] = 32'b00000000000000001001000010110011;
assign LUT_1[18175] = 32'b00000000000000000010010100101111;
assign LUT_1[18176] = 32'b11111111111111111100001101010110;
assign LUT_1[18177] = 32'b11111111111111110101011111010010;
assign LUT_1[18178] = 32'b11111111111111110111111011100111;
assign LUT_1[18179] = 32'b11111111111111110001001101100011;
assign LUT_1[18180] = 32'b00000000000000000100000110101101;
assign LUT_1[18181] = 32'b11111111111111111101011000101001;
assign LUT_1[18182] = 32'b11111111111111111111110100111110;
assign LUT_1[18183] = 32'b11111111111111111001000110111010;
assign LUT_1[18184] = 32'b11111111111111111011011011001011;
assign LUT_1[18185] = 32'b11111111111111110100101101000111;
assign LUT_1[18186] = 32'b11111111111111110111001001011100;
assign LUT_1[18187] = 32'b11111111111111110000011011011000;
assign LUT_1[18188] = 32'b00000000000000000011010100100010;
assign LUT_1[18189] = 32'b11111111111111111100100110011110;
assign LUT_1[18190] = 32'b11111111111111111111000010110011;
assign LUT_1[18191] = 32'b11111111111111111000010100101111;
assign LUT_1[18192] = 32'b11111111111111111110001000111000;
assign LUT_1[18193] = 32'b11111111111111110111011010110100;
assign LUT_1[18194] = 32'b11111111111111111001110111001001;
assign LUT_1[18195] = 32'b11111111111111110011001001000101;
assign LUT_1[18196] = 32'b00000000000000000110000010001111;
assign LUT_1[18197] = 32'b11111111111111111111010100001011;
assign LUT_1[18198] = 32'b00000000000000000001110000100000;
assign LUT_1[18199] = 32'b11111111111111111011000010011100;
assign LUT_1[18200] = 32'b11111111111111111101010110101101;
assign LUT_1[18201] = 32'b11111111111111110110101000101001;
assign LUT_1[18202] = 32'b11111111111111111001000100111110;
assign LUT_1[18203] = 32'b11111111111111110010010110111010;
assign LUT_1[18204] = 32'b00000000000000000101010000000100;
assign LUT_1[18205] = 32'b11111111111111111110100010000000;
assign LUT_1[18206] = 32'b00000000000000000000111110010101;
assign LUT_1[18207] = 32'b11111111111111111010010000010001;
assign LUT_1[18208] = 32'b11111111111111111101001000010101;
assign LUT_1[18209] = 32'b11111111111111110110011010010001;
assign LUT_1[18210] = 32'b11111111111111111000110110100110;
assign LUT_1[18211] = 32'b11111111111111110010001000100010;
assign LUT_1[18212] = 32'b00000000000000000101000001101100;
assign LUT_1[18213] = 32'b11111111111111111110010011101000;
assign LUT_1[18214] = 32'b00000000000000000000101111111101;
assign LUT_1[18215] = 32'b11111111111111111010000001111001;
assign LUT_1[18216] = 32'b11111111111111111100010110001010;
assign LUT_1[18217] = 32'b11111111111111110101101000000110;
assign LUT_1[18218] = 32'b11111111111111111000000100011011;
assign LUT_1[18219] = 32'b11111111111111110001010110010111;
assign LUT_1[18220] = 32'b00000000000000000100001111100001;
assign LUT_1[18221] = 32'b11111111111111111101100001011101;
assign LUT_1[18222] = 32'b11111111111111111111111101110010;
assign LUT_1[18223] = 32'b11111111111111111001001111101110;
assign LUT_1[18224] = 32'b11111111111111111111000011110111;
assign LUT_1[18225] = 32'b11111111111111111000010101110011;
assign LUT_1[18226] = 32'b11111111111111111010110010001000;
assign LUT_1[18227] = 32'b11111111111111110100000100000100;
assign LUT_1[18228] = 32'b00000000000000000110111101001110;
assign LUT_1[18229] = 32'b00000000000000000000001111001010;
assign LUT_1[18230] = 32'b00000000000000000010101011011111;
assign LUT_1[18231] = 32'b11111111111111111011111101011011;
assign LUT_1[18232] = 32'b11111111111111111110010001101100;
assign LUT_1[18233] = 32'b11111111111111110111100011101000;
assign LUT_1[18234] = 32'b11111111111111111001111111111101;
assign LUT_1[18235] = 32'b11111111111111110011010001111001;
assign LUT_1[18236] = 32'b00000000000000000110001011000011;
assign LUT_1[18237] = 32'b11111111111111111111011100111111;
assign LUT_1[18238] = 32'b00000000000000000001111001010100;
assign LUT_1[18239] = 32'b11111111111111111011001011010000;
assign LUT_1[18240] = 32'b11111111111111111110001010111110;
assign LUT_1[18241] = 32'b11111111111111110111011100111010;
assign LUT_1[18242] = 32'b11111111111111111001111001001111;
assign LUT_1[18243] = 32'b11111111111111110011001011001011;
assign LUT_1[18244] = 32'b00000000000000000110000100010101;
assign LUT_1[18245] = 32'b11111111111111111111010110010001;
assign LUT_1[18246] = 32'b00000000000000000001110010100110;
assign LUT_1[18247] = 32'b11111111111111111011000100100010;
assign LUT_1[18248] = 32'b11111111111111111101011000110011;
assign LUT_1[18249] = 32'b11111111111111110110101010101111;
assign LUT_1[18250] = 32'b11111111111111111001000111000100;
assign LUT_1[18251] = 32'b11111111111111110010011001000000;
assign LUT_1[18252] = 32'b00000000000000000101010010001010;
assign LUT_1[18253] = 32'b11111111111111111110100100000110;
assign LUT_1[18254] = 32'b00000000000000000001000000011011;
assign LUT_1[18255] = 32'b11111111111111111010010010010111;
assign LUT_1[18256] = 32'b00000000000000000000000110100000;
assign LUT_1[18257] = 32'b11111111111111111001011000011100;
assign LUT_1[18258] = 32'b11111111111111111011110100110001;
assign LUT_1[18259] = 32'b11111111111111110101000110101101;
assign LUT_1[18260] = 32'b00000000000000000111111111110111;
assign LUT_1[18261] = 32'b00000000000000000001010001110011;
assign LUT_1[18262] = 32'b00000000000000000011101110001000;
assign LUT_1[18263] = 32'b11111111111111111101000000000100;
assign LUT_1[18264] = 32'b11111111111111111111010100010101;
assign LUT_1[18265] = 32'b11111111111111111000100110010001;
assign LUT_1[18266] = 32'b11111111111111111011000010100110;
assign LUT_1[18267] = 32'b11111111111111110100010100100010;
assign LUT_1[18268] = 32'b00000000000000000111001101101100;
assign LUT_1[18269] = 32'b00000000000000000000011111101000;
assign LUT_1[18270] = 32'b00000000000000000010111011111101;
assign LUT_1[18271] = 32'b11111111111111111100001101111001;
assign LUT_1[18272] = 32'b11111111111111111111000101111101;
assign LUT_1[18273] = 32'b11111111111111111000010111111001;
assign LUT_1[18274] = 32'b11111111111111111010110100001110;
assign LUT_1[18275] = 32'b11111111111111110100000110001010;
assign LUT_1[18276] = 32'b00000000000000000110111111010100;
assign LUT_1[18277] = 32'b00000000000000000000010001010000;
assign LUT_1[18278] = 32'b00000000000000000010101101100101;
assign LUT_1[18279] = 32'b11111111111111111011111111100001;
assign LUT_1[18280] = 32'b11111111111111111110010011110010;
assign LUT_1[18281] = 32'b11111111111111110111100101101110;
assign LUT_1[18282] = 32'b11111111111111111010000010000011;
assign LUT_1[18283] = 32'b11111111111111110011010011111111;
assign LUT_1[18284] = 32'b00000000000000000110001101001001;
assign LUT_1[18285] = 32'b11111111111111111111011111000101;
assign LUT_1[18286] = 32'b00000000000000000001111011011010;
assign LUT_1[18287] = 32'b11111111111111111011001101010110;
assign LUT_1[18288] = 32'b00000000000000000001000001011111;
assign LUT_1[18289] = 32'b11111111111111111010010011011011;
assign LUT_1[18290] = 32'b11111111111111111100101111110000;
assign LUT_1[18291] = 32'b11111111111111110110000001101100;
assign LUT_1[18292] = 32'b00000000000000001000111010110110;
assign LUT_1[18293] = 32'b00000000000000000010001100110010;
assign LUT_1[18294] = 32'b00000000000000000100101001000111;
assign LUT_1[18295] = 32'b11111111111111111101111011000011;
assign LUT_1[18296] = 32'b00000000000000000000001111010100;
assign LUT_1[18297] = 32'b11111111111111111001100001010000;
assign LUT_1[18298] = 32'b11111111111111111011111101100101;
assign LUT_1[18299] = 32'b11111111111111110101001111100001;
assign LUT_1[18300] = 32'b00000000000000001000001000101011;
assign LUT_1[18301] = 32'b00000000000000000001011010100111;
assign LUT_1[18302] = 32'b00000000000000000011110110111100;
assign LUT_1[18303] = 32'b11111111111111111101001000111000;
assign LUT_1[18304] = 32'b11111111111111111111001101011001;
assign LUT_1[18305] = 32'b11111111111111111000011111010101;
assign LUT_1[18306] = 32'b11111111111111111010111011101010;
assign LUT_1[18307] = 32'b11111111111111110100001101100110;
assign LUT_1[18308] = 32'b00000000000000000111000110110000;
assign LUT_1[18309] = 32'b00000000000000000000011000101100;
assign LUT_1[18310] = 32'b00000000000000000010110101000001;
assign LUT_1[18311] = 32'b11111111111111111100000110111101;
assign LUT_1[18312] = 32'b11111111111111111110011011001110;
assign LUT_1[18313] = 32'b11111111111111110111101101001010;
assign LUT_1[18314] = 32'b11111111111111111010001001011111;
assign LUT_1[18315] = 32'b11111111111111110011011011011011;
assign LUT_1[18316] = 32'b00000000000000000110010100100101;
assign LUT_1[18317] = 32'b11111111111111111111100110100001;
assign LUT_1[18318] = 32'b00000000000000000010000010110110;
assign LUT_1[18319] = 32'b11111111111111111011010100110010;
assign LUT_1[18320] = 32'b00000000000000000001001000111011;
assign LUT_1[18321] = 32'b11111111111111111010011010110111;
assign LUT_1[18322] = 32'b11111111111111111100110111001100;
assign LUT_1[18323] = 32'b11111111111111110110001001001000;
assign LUT_1[18324] = 32'b00000000000000001001000010010010;
assign LUT_1[18325] = 32'b00000000000000000010010100001110;
assign LUT_1[18326] = 32'b00000000000000000100110000100011;
assign LUT_1[18327] = 32'b11111111111111111110000010011111;
assign LUT_1[18328] = 32'b00000000000000000000010110110000;
assign LUT_1[18329] = 32'b11111111111111111001101000101100;
assign LUT_1[18330] = 32'b11111111111111111100000101000001;
assign LUT_1[18331] = 32'b11111111111111110101010110111101;
assign LUT_1[18332] = 32'b00000000000000001000010000000111;
assign LUT_1[18333] = 32'b00000000000000000001100010000011;
assign LUT_1[18334] = 32'b00000000000000000011111110011000;
assign LUT_1[18335] = 32'b11111111111111111101010000010100;
assign LUT_1[18336] = 32'b00000000000000000000001000011000;
assign LUT_1[18337] = 32'b11111111111111111001011010010100;
assign LUT_1[18338] = 32'b11111111111111111011110110101001;
assign LUT_1[18339] = 32'b11111111111111110101001000100101;
assign LUT_1[18340] = 32'b00000000000000001000000001101111;
assign LUT_1[18341] = 32'b00000000000000000001010011101011;
assign LUT_1[18342] = 32'b00000000000000000011110000000000;
assign LUT_1[18343] = 32'b11111111111111111101000001111100;
assign LUT_1[18344] = 32'b11111111111111111111010110001101;
assign LUT_1[18345] = 32'b11111111111111111000101000001001;
assign LUT_1[18346] = 32'b11111111111111111011000100011110;
assign LUT_1[18347] = 32'b11111111111111110100010110011010;
assign LUT_1[18348] = 32'b00000000000000000111001111100100;
assign LUT_1[18349] = 32'b00000000000000000000100001100000;
assign LUT_1[18350] = 32'b00000000000000000010111101110101;
assign LUT_1[18351] = 32'b11111111111111111100001111110001;
assign LUT_1[18352] = 32'b00000000000000000010000011111010;
assign LUT_1[18353] = 32'b11111111111111111011010101110110;
assign LUT_1[18354] = 32'b11111111111111111101110010001011;
assign LUT_1[18355] = 32'b11111111111111110111000100000111;
assign LUT_1[18356] = 32'b00000000000000001001111101010001;
assign LUT_1[18357] = 32'b00000000000000000011001111001101;
assign LUT_1[18358] = 32'b00000000000000000101101011100010;
assign LUT_1[18359] = 32'b11111111111111111110111101011110;
assign LUT_1[18360] = 32'b00000000000000000001010001101111;
assign LUT_1[18361] = 32'b11111111111111111010100011101011;
assign LUT_1[18362] = 32'b11111111111111111101000000000000;
assign LUT_1[18363] = 32'b11111111111111110110010001111100;
assign LUT_1[18364] = 32'b00000000000000001001001011000110;
assign LUT_1[18365] = 32'b00000000000000000010011101000010;
assign LUT_1[18366] = 32'b00000000000000000100111001010111;
assign LUT_1[18367] = 32'b11111111111111111110001011010011;
assign LUT_1[18368] = 32'b00000000000000000001001011000001;
assign LUT_1[18369] = 32'b11111111111111111010011100111101;
assign LUT_1[18370] = 32'b11111111111111111100111001010010;
assign LUT_1[18371] = 32'b11111111111111110110001011001110;
assign LUT_1[18372] = 32'b00000000000000001001000100011000;
assign LUT_1[18373] = 32'b00000000000000000010010110010100;
assign LUT_1[18374] = 32'b00000000000000000100110010101001;
assign LUT_1[18375] = 32'b11111111111111111110000100100101;
assign LUT_1[18376] = 32'b00000000000000000000011000110110;
assign LUT_1[18377] = 32'b11111111111111111001101010110010;
assign LUT_1[18378] = 32'b11111111111111111100000111000111;
assign LUT_1[18379] = 32'b11111111111111110101011001000011;
assign LUT_1[18380] = 32'b00000000000000001000010010001101;
assign LUT_1[18381] = 32'b00000000000000000001100100001001;
assign LUT_1[18382] = 32'b00000000000000000100000000011110;
assign LUT_1[18383] = 32'b11111111111111111101010010011010;
assign LUT_1[18384] = 32'b00000000000000000011000110100011;
assign LUT_1[18385] = 32'b11111111111111111100011000011111;
assign LUT_1[18386] = 32'b11111111111111111110110100110100;
assign LUT_1[18387] = 32'b11111111111111111000000110110000;
assign LUT_1[18388] = 32'b00000000000000001010111111111010;
assign LUT_1[18389] = 32'b00000000000000000100010001110110;
assign LUT_1[18390] = 32'b00000000000000000110101110001011;
assign LUT_1[18391] = 32'b00000000000000000000000000000111;
assign LUT_1[18392] = 32'b00000000000000000010010100011000;
assign LUT_1[18393] = 32'b11111111111111111011100110010100;
assign LUT_1[18394] = 32'b11111111111111111110000010101001;
assign LUT_1[18395] = 32'b11111111111111110111010100100101;
assign LUT_1[18396] = 32'b00000000000000001010001101101111;
assign LUT_1[18397] = 32'b00000000000000000011011111101011;
assign LUT_1[18398] = 32'b00000000000000000101111100000000;
assign LUT_1[18399] = 32'b11111111111111111111001101111100;
assign LUT_1[18400] = 32'b00000000000000000010000110000000;
assign LUT_1[18401] = 32'b11111111111111111011010111111100;
assign LUT_1[18402] = 32'b11111111111111111101110100010001;
assign LUT_1[18403] = 32'b11111111111111110111000110001101;
assign LUT_1[18404] = 32'b00000000000000001001111111010111;
assign LUT_1[18405] = 32'b00000000000000000011010001010011;
assign LUT_1[18406] = 32'b00000000000000000101101101101000;
assign LUT_1[18407] = 32'b11111111111111111110111111100100;
assign LUT_1[18408] = 32'b00000000000000000001010011110101;
assign LUT_1[18409] = 32'b11111111111111111010100101110001;
assign LUT_1[18410] = 32'b11111111111111111101000010000110;
assign LUT_1[18411] = 32'b11111111111111110110010100000010;
assign LUT_1[18412] = 32'b00000000000000001001001101001100;
assign LUT_1[18413] = 32'b00000000000000000010011111001000;
assign LUT_1[18414] = 32'b00000000000000000100111011011101;
assign LUT_1[18415] = 32'b11111111111111111110001101011001;
assign LUT_1[18416] = 32'b00000000000000000100000001100010;
assign LUT_1[18417] = 32'b11111111111111111101010011011110;
assign LUT_1[18418] = 32'b11111111111111111111101111110011;
assign LUT_1[18419] = 32'b11111111111111111001000001101111;
assign LUT_1[18420] = 32'b00000000000000001011111010111001;
assign LUT_1[18421] = 32'b00000000000000000101001100110101;
assign LUT_1[18422] = 32'b00000000000000000111101001001010;
assign LUT_1[18423] = 32'b00000000000000000000111011000110;
assign LUT_1[18424] = 32'b00000000000000000011001111010111;
assign LUT_1[18425] = 32'b11111111111111111100100001010011;
assign LUT_1[18426] = 32'b11111111111111111110111101101000;
assign LUT_1[18427] = 32'b11111111111111111000001111100100;
assign LUT_1[18428] = 32'b00000000000000001011001000101110;
assign LUT_1[18429] = 32'b00000000000000000100011010101010;
assign LUT_1[18430] = 32'b00000000000000000110110110111111;
assign LUT_1[18431] = 32'b00000000000000000000001000111011;
assign LUT_1[18432] = 32'b11111111111111111111010101111000;
assign LUT_1[18433] = 32'b11111111111111111000100111110100;
assign LUT_1[18434] = 32'b11111111111111111011000100001001;
assign LUT_1[18435] = 32'b11111111111111110100010110000101;
assign LUT_1[18436] = 32'b00000000000000000111001111001111;
assign LUT_1[18437] = 32'b00000000000000000000100001001011;
assign LUT_1[18438] = 32'b00000000000000000010111101100000;
assign LUT_1[18439] = 32'b11111111111111111100001111011100;
assign LUT_1[18440] = 32'b11111111111111111110100011101101;
assign LUT_1[18441] = 32'b11111111111111110111110101101001;
assign LUT_1[18442] = 32'b11111111111111111010010001111110;
assign LUT_1[18443] = 32'b11111111111111110011100011111010;
assign LUT_1[18444] = 32'b00000000000000000110011101000100;
assign LUT_1[18445] = 32'b11111111111111111111101111000000;
assign LUT_1[18446] = 32'b00000000000000000010001011010101;
assign LUT_1[18447] = 32'b11111111111111111011011101010001;
assign LUT_1[18448] = 32'b00000000000000000001010001011010;
assign LUT_1[18449] = 32'b11111111111111111010100011010110;
assign LUT_1[18450] = 32'b11111111111111111100111111101011;
assign LUT_1[18451] = 32'b11111111111111110110010001100111;
assign LUT_1[18452] = 32'b00000000000000001001001010110001;
assign LUT_1[18453] = 32'b00000000000000000010011100101101;
assign LUT_1[18454] = 32'b00000000000000000100111001000010;
assign LUT_1[18455] = 32'b11111111111111111110001010111110;
assign LUT_1[18456] = 32'b00000000000000000000011111001111;
assign LUT_1[18457] = 32'b11111111111111111001110001001011;
assign LUT_1[18458] = 32'b11111111111111111100001101100000;
assign LUT_1[18459] = 32'b11111111111111110101011111011100;
assign LUT_1[18460] = 32'b00000000000000001000011000100110;
assign LUT_1[18461] = 32'b00000000000000000001101010100010;
assign LUT_1[18462] = 32'b00000000000000000100000110110111;
assign LUT_1[18463] = 32'b11111111111111111101011000110011;
assign LUT_1[18464] = 32'b00000000000000000000010000110111;
assign LUT_1[18465] = 32'b11111111111111111001100010110011;
assign LUT_1[18466] = 32'b11111111111111111011111111001000;
assign LUT_1[18467] = 32'b11111111111111110101010001000100;
assign LUT_1[18468] = 32'b00000000000000001000001010001110;
assign LUT_1[18469] = 32'b00000000000000000001011100001010;
assign LUT_1[18470] = 32'b00000000000000000011111000011111;
assign LUT_1[18471] = 32'b11111111111111111101001010011011;
assign LUT_1[18472] = 32'b11111111111111111111011110101100;
assign LUT_1[18473] = 32'b11111111111111111000110000101000;
assign LUT_1[18474] = 32'b11111111111111111011001100111101;
assign LUT_1[18475] = 32'b11111111111111110100011110111001;
assign LUT_1[18476] = 32'b00000000000000000111011000000011;
assign LUT_1[18477] = 32'b00000000000000000000101001111111;
assign LUT_1[18478] = 32'b00000000000000000011000110010100;
assign LUT_1[18479] = 32'b11111111111111111100011000010000;
assign LUT_1[18480] = 32'b00000000000000000010001100011001;
assign LUT_1[18481] = 32'b11111111111111111011011110010101;
assign LUT_1[18482] = 32'b11111111111111111101111010101010;
assign LUT_1[18483] = 32'b11111111111111110111001100100110;
assign LUT_1[18484] = 32'b00000000000000001010000101110000;
assign LUT_1[18485] = 32'b00000000000000000011010111101100;
assign LUT_1[18486] = 32'b00000000000000000101110100000001;
assign LUT_1[18487] = 32'b11111111111111111111000101111101;
assign LUT_1[18488] = 32'b00000000000000000001011010001110;
assign LUT_1[18489] = 32'b11111111111111111010101100001010;
assign LUT_1[18490] = 32'b11111111111111111101001000011111;
assign LUT_1[18491] = 32'b11111111111111110110011010011011;
assign LUT_1[18492] = 32'b00000000000000001001010011100101;
assign LUT_1[18493] = 32'b00000000000000000010100101100001;
assign LUT_1[18494] = 32'b00000000000000000101000001110110;
assign LUT_1[18495] = 32'b11111111111111111110010011110010;
assign LUT_1[18496] = 32'b00000000000000000001010011100000;
assign LUT_1[18497] = 32'b11111111111111111010100101011100;
assign LUT_1[18498] = 32'b11111111111111111101000001110001;
assign LUT_1[18499] = 32'b11111111111111110110010011101101;
assign LUT_1[18500] = 32'b00000000000000001001001100110111;
assign LUT_1[18501] = 32'b00000000000000000010011110110011;
assign LUT_1[18502] = 32'b00000000000000000100111011001000;
assign LUT_1[18503] = 32'b11111111111111111110001101000100;
assign LUT_1[18504] = 32'b00000000000000000000100001010101;
assign LUT_1[18505] = 32'b11111111111111111001110011010001;
assign LUT_1[18506] = 32'b11111111111111111100001111100110;
assign LUT_1[18507] = 32'b11111111111111110101100001100010;
assign LUT_1[18508] = 32'b00000000000000001000011010101100;
assign LUT_1[18509] = 32'b00000000000000000001101100101000;
assign LUT_1[18510] = 32'b00000000000000000100001000111101;
assign LUT_1[18511] = 32'b11111111111111111101011010111001;
assign LUT_1[18512] = 32'b00000000000000000011001111000010;
assign LUT_1[18513] = 32'b11111111111111111100100000111110;
assign LUT_1[18514] = 32'b11111111111111111110111101010011;
assign LUT_1[18515] = 32'b11111111111111111000001111001111;
assign LUT_1[18516] = 32'b00000000000000001011001000011001;
assign LUT_1[18517] = 32'b00000000000000000100011010010101;
assign LUT_1[18518] = 32'b00000000000000000110110110101010;
assign LUT_1[18519] = 32'b00000000000000000000001000100110;
assign LUT_1[18520] = 32'b00000000000000000010011100110111;
assign LUT_1[18521] = 32'b11111111111111111011101110110011;
assign LUT_1[18522] = 32'b11111111111111111110001011001000;
assign LUT_1[18523] = 32'b11111111111111110111011101000100;
assign LUT_1[18524] = 32'b00000000000000001010010110001110;
assign LUT_1[18525] = 32'b00000000000000000011101000001010;
assign LUT_1[18526] = 32'b00000000000000000110000100011111;
assign LUT_1[18527] = 32'b11111111111111111111010110011011;
assign LUT_1[18528] = 32'b00000000000000000010001110011111;
assign LUT_1[18529] = 32'b11111111111111111011100000011011;
assign LUT_1[18530] = 32'b11111111111111111101111100110000;
assign LUT_1[18531] = 32'b11111111111111110111001110101100;
assign LUT_1[18532] = 32'b00000000000000001010000111110110;
assign LUT_1[18533] = 32'b00000000000000000011011001110010;
assign LUT_1[18534] = 32'b00000000000000000101110110000111;
assign LUT_1[18535] = 32'b11111111111111111111001000000011;
assign LUT_1[18536] = 32'b00000000000000000001011100010100;
assign LUT_1[18537] = 32'b11111111111111111010101110010000;
assign LUT_1[18538] = 32'b11111111111111111101001010100101;
assign LUT_1[18539] = 32'b11111111111111110110011100100001;
assign LUT_1[18540] = 32'b00000000000000001001010101101011;
assign LUT_1[18541] = 32'b00000000000000000010100111100111;
assign LUT_1[18542] = 32'b00000000000000000101000011111100;
assign LUT_1[18543] = 32'b11111111111111111110010101111000;
assign LUT_1[18544] = 32'b00000000000000000100001010000001;
assign LUT_1[18545] = 32'b11111111111111111101011011111101;
assign LUT_1[18546] = 32'b11111111111111111111111000010010;
assign LUT_1[18547] = 32'b11111111111111111001001010001110;
assign LUT_1[18548] = 32'b00000000000000001100000011011000;
assign LUT_1[18549] = 32'b00000000000000000101010101010100;
assign LUT_1[18550] = 32'b00000000000000000111110001101001;
assign LUT_1[18551] = 32'b00000000000000000001000011100101;
assign LUT_1[18552] = 32'b00000000000000000011010111110110;
assign LUT_1[18553] = 32'b11111111111111111100101001110010;
assign LUT_1[18554] = 32'b11111111111111111111000110000111;
assign LUT_1[18555] = 32'b11111111111111111000011000000011;
assign LUT_1[18556] = 32'b00000000000000001011010001001101;
assign LUT_1[18557] = 32'b00000000000000000100100011001001;
assign LUT_1[18558] = 32'b00000000000000000110111111011110;
assign LUT_1[18559] = 32'b00000000000000000000010001011010;
assign LUT_1[18560] = 32'b00000000000000000010010101111011;
assign LUT_1[18561] = 32'b11111111111111111011100111110111;
assign LUT_1[18562] = 32'b11111111111111111110000100001100;
assign LUT_1[18563] = 32'b11111111111111110111010110001000;
assign LUT_1[18564] = 32'b00000000000000001010001111010010;
assign LUT_1[18565] = 32'b00000000000000000011100001001110;
assign LUT_1[18566] = 32'b00000000000000000101111101100011;
assign LUT_1[18567] = 32'b11111111111111111111001111011111;
assign LUT_1[18568] = 32'b00000000000000000001100011110000;
assign LUT_1[18569] = 32'b11111111111111111010110101101100;
assign LUT_1[18570] = 32'b11111111111111111101010010000001;
assign LUT_1[18571] = 32'b11111111111111110110100011111101;
assign LUT_1[18572] = 32'b00000000000000001001011101000111;
assign LUT_1[18573] = 32'b00000000000000000010101111000011;
assign LUT_1[18574] = 32'b00000000000000000101001011011000;
assign LUT_1[18575] = 32'b11111111111111111110011101010100;
assign LUT_1[18576] = 32'b00000000000000000100010001011101;
assign LUT_1[18577] = 32'b11111111111111111101100011011001;
assign LUT_1[18578] = 32'b11111111111111111111111111101110;
assign LUT_1[18579] = 32'b11111111111111111001010001101010;
assign LUT_1[18580] = 32'b00000000000000001100001010110100;
assign LUT_1[18581] = 32'b00000000000000000101011100110000;
assign LUT_1[18582] = 32'b00000000000000000111111001000101;
assign LUT_1[18583] = 32'b00000000000000000001001011000001;
assign LUT_1[18584] = 32'b00000000000000000011011111010010;
assign LUT_1[18585] = 32'b11111111111111111100110001001110;
assign LUT_1[18586] = 32'b11111111111111111111001101100011;
assign LUT_1[18587] = 32'b11111111111111111000011111011111;
assign LUT_1[18588] = 32'b00000000000000001011011000101001;
assign LUT_1[18589] = 32'b00000000000000000100101010100101;
assign LUT_1[18590] = 32'b00000000000000000111000110111010;
assign LUT_1[18591] = 32'b00000000000000000000011000110110;
assign LUT_1[18592] = 32'b00000000000000000011010000111010;
assign LUT_1[18593] = 32'b11111111111111111100100010110110;
assign LUT_1[18594] = 32'b11111111111111111110111111001011;
assign LUT_1[18595] = 32'b11111111111111111000010001000111;
assign LUT_1[18596] = 32'b00000000000000001011001010010001;
assign LUT_1[18597] = 32'b00000000000000000100011100001101;
assign LUT_1[18598] = 32'b00000000000000000110111000100010;
assign LUT_1[18599] = 32'b00000000000000000000001010011110;
assign LUT_1[18600] = 32'b00000000000000000010011110101111;
assign LUT_1[18601] = 32'b11111111111111111011110000101011;
assign LUT_1[18602] = 32'b11111111111111111110001101000000;
assign LUT_1[18603] = 32'b11111111111111110111011110111100;
assign LUT_1[18604] = 32'b00000000000000001010011000000110;
assign LUT_1[18605] = 32'b00000000000000000011101010000010;
assign LUT_1[18606] = 32'b00000000000000000110000110010111;
assign LUT_1[18607] = 32'b11111111111111111111011000010011;
assign LUT_1[18608] = 32'b00000000000000000101001100011100;
assign LUT_1[18609] = 32'b11111111111111111110011110011000;
assign LUT_1[18610] = 32'b00000000000000000000111010101101;
assign LUT_1[18611] = 32'b11111111111111111010001100101001;
assign LUT_1[18612] = 32'b00000000000000001101000101110011;
assign LUT_1[18613] = 32'b00000000000000000110010111101111;
assign LUT_1[18614] = 32'b00000000000000001000110100000100;
assign LUT_1[18615] = 32'b00000000000000000010000110000000;
assign LUT_1[18616] = 32'b00000000000000000100011010010001;
assign LUT_1[18617] = 32'b11111111111111111101101100001101;
assign LUT_1[18618] = 32'b00000000000000000000001000100010;
assign LUT_1[18619] = 32'b11111111111111111001011010011110;
assign LUT_1[18620] = 32'b00000000000000001100010011101000;
assign LUT_1[18621] = 32'b00000000000000000101100101100100;
assign LUT_1[18622] = 32'b00000000000000001000000001111001;
assign LUT_1[18623] = 32'b00000000000000000001010011110101;
assign LUT_1[18624] = 32'b00000000000000000100010011100011;
assign LUT_1[18625] = 32'b11111111111111111101100101011111;
assign LUT_1[18626] = 32'b00000000000000000000000001110100;
assign LUT_1[18627] = 32'b11111111111111111001010011110000;
assign LUT_1[18628] = 32'b00000000000000001100001100111010;
assign LUT_1[18629] = 32'b00000000000000000101011110110110;
assign LUT_1[18630] = 32'b00000000000000000111111011001011;
assign LUT_1[18631] = 32'b00000000000000000001001101000111;
assign LUT_1[18632] = 32'b00000000000000000011100001011000;
assign LUT_1[18633] = 32'b11111111111111111100110011010100;
assign LUT_1[18634] = 32'b11111111111111111111001111101001;
assign LUT_1[18635] = 32'b11111111111111111000100001100101;
assign LUT_1[18636] = 32'b00000000000000001011011010101111;
assign LUT_1[18637] = 32'b00000000000000000100101100101011;
assign LUT_1[18638] = 32'b00000000000000000111001001000000;
assign LUT_1[18639] = 32'b00000000000000000000011010111100;
assign LUT_1[18640] = 32'b00000000000000000110001111000101;
assign LUT_1[18641] = 32'b11111111111111111111100001000001;
assign LUT_1[18642] = 32'b00000000000000000001111101010110;
assign LUT_1[18643] = 32'b11111111111111111011001111010010;
assign LUT_1[18644] = 32'b00000000000000001110001000011100;
assign LUT_1[18645] = 32'b00000000000000000111011010011000;
assign LUT_1[18646] = 32'b00000000000000001001110110101101;
assign LUT_1[18647] = 32'b00000000000000000011001000101001;
assign LUT_1[18648] = 32'b00000000000000000101011100111010;
assign LUT_1[18649] = 32'b11111111111111111110101110110110;
assign LUT_1[18650] = 32'b00000000000000000001001011001011;
assign LUT_1[18651] = 32'b11111111111111111010011101000111;
assign LUT_1[18652] = 32'b00000000000000001101010110010001;
assign LUT_1[18653] = 32'b00000000000000000110101000001101;
assign LUT_1[18654] = 32'b00000000000000001001000100100010;
assign LUT_1[18655] = 32'b00000000000000000010010110011110;
assign LUT_1[18656] = 32'b00000000000000000101001110100010;
assign LUT_1[18657] = 32'b11111111111111111110100000011110;
assign LUT_1[18658] = 32'b00000000000000000000111100110011;
assign LUT_1[18659] = 32'b11111111111111111010001110101111;
assign LUT_1[18660] = 32'b00000000000000001101000111111001;
assign LUT_1[18661] = 32'b00000000000000000110011001110101;
assign LUT_1[18662] = 32'b00000000000000001000110110001010;
assign LUT_1[18663] = 32'b00000000000000000010001000000110;
assign LUT_1[18664] = 32'b00000000000000000100011100010111;
assign LUT_1[18665] = 32'b11111111111111111101101110010011;
assign LUT_1[18666] = 32'b00000000000000000000001010101000;
assign LUT_1[18667] = 32'b11111111111111111001011100100100;
assign LUT_1[18668] = 32'b00000000000000001100010101101110;
assign LUT_1[18669] = 32'b00000000000000000101100111101010;
assign LUT_1[18670] = 32'b00000000000000001000000011111111;
assign LUT_1[18671] = 32'b00000000000000000001010101111011;
assign LUT_1[18672] = 32'b00000000000000000111001010000100;
assign LUT_1[18673] = 32'b00000000000000000000011100000000;
assign LUT_1[18674] = 32'b00000000000000000010111000010101;
assign LUT_1[18675] = 32'b11111111111111111100001010010001;
assign LUT_1[18676] = 32'b00000000000000001111000011011011;
assign LUT_1[18677] = 32'b00000000000000001000010101010111;
assign LUT_1[18678] = 32'b00000000000000001010110001101100;
assign LUT_1[18679] = 32'b00000000000000000100000011101000;
assign LUT_1[18680] = 32'b00000000000000000110010111111001;
assign LUT_1[18681] = 32'b11111111111111111111101001110101;
assign LUT_1[18682] = 32'b00000000000000000010000110001010;
assign LUT_1[18683] = 32'b11111111111111111011011000000110;
assign LUT_1[18684] = 32'b00000000000000001110010001010000;
assign LUT_1[18685] = 32'b00000000000000000111100011001100;
assign LUT_1[18686] = 32'b00000000000000001001111111100001;
assign LUT_1[18687] = 32'b00000000000000000011010001011101;
assign LUT_1[18688] = 32'b11111111111111111101001010000100;
assign LUT_1[18689] = 32'b11111111111111110110011100000000;
assign LUT_1[18690] = 32'b11111111111111111000111000010101;
assign LUT_1[18691] = 32'b11111111111111110010001010010001;
assign LUT_1[18692] = 32'b00000000000000000101000011011011;
assign LUT_1[18693] = 32'b11111111111111111110010101010111;
assign LUT_1[18694] = 32'b00000000000000000000110001101100;
assign LUT_1[18695] = 32'b11111111111111111010000011101000;
assign LUT_1[18696] = 32'b11111111111111111100010111111001;
assign LUT_1[18697] = 32'b11111111111111110101101001110101;
assign LUT_1[18698] = 32'b11111111111111111000000110001010;
assign LUT_1[18699] = 32'b11111111111111110001011000000110;
assign LUT_1[18700] = 32'b00000000000000000100010001010000;
assign LUT_1[18701] = 32'b11111111111111111101100011001100;
assign LUT_1[18702] = 32'b11111111111111111111111111100001;
assign LUT_1[18703] = 32'b11111111111111111001010001011101;
assign LUT_1[18704] = 32'b11111111111111111111000101100110;
assign LUT_1[18705] = 32'b11111111111111111000010111100010;
assign LUT_1[18706] = 32'b11111111111111111010110011110111;
assign LUT_1[18707] = 32'b11111111111111110100000101110011;
assign LUT_1[18708] = 32'b00000000000000000110111110111101;
assign LUT_1[18709] = 32'b00000000000000000000010000111001;
assign LUT_1[18710] = 32'b00000000000000000010101101001110;
assign LUT_1[18711] = 32'b11111111111111111011111111001010;
assign LUT_1[18712] = 32'b11111111111111111110010011011011;
assign LUT_1[18713] = 32'b11111111111111110111100101010111;
assign LUT_1[18714] = 32'b11111111111111111010000001101100;
assign LUT_1[18715] = 32'b11111111111111110011010011101000;
assign LUT_1[18716] = 32'b00000000000000000110001100110010;
assign LUT_1[18717] = 32'b11111111111111111111011110101110;
assign LUT_1[18718] = 32'b00000000000000000001111011000011;
assign LUT_1[18719] = 32'b11111111111111111011001100111111;
assign LUT_1[18720] = 32'b11111111111111111110000101000011;
assign LUT_1[18721] = 32'b11111111111111110111010110111111;
assign LUT_1[18722] = 32'b11111111111111111001110011010100;
assign LUT_1[18723] = 32'b11111111111111110011000101010000;
assign LUT_1[18724] = 32'b00000000000000000101111110011010;
assign LUT_1[18725] = 32'b11111111111111111111010000010110;
assign LUT_1[18726] = 32'b00000000000000000001101100101011;
assign LUT_1[18727] = 32'b11111111111111111010111110100111;
assign LUT_1[18728] = 32'b11111111111111111101010010111000;
assign LUT_1[18729] = 32'b11111111111111110110100100110100;
assign LUT_1[18730] = 32'b11111111111111111001000001001001;
assign LUT_1[18731] = 32'b11111111111111110010010011000101;
assign LUT_1[18732] = 32'b00000000000000000101001100001111;
assign LUT_1[18733] = 32'b11111111111111111110011110001011;
assign LUT_1[18734] = 32'b00000000000000000000111010100000;
assign LUT_1[18735] = 32'b11111111111111111010001100011100;
assign LUT_1[18736] = 32'b00000000000000000000000000100101;
assign LUT_1[18737] = 32'b11111111111111111001010010100001;
assign LUT_1[18738] = 32'b11111111111111111011101110110110;
assign LUT_1[18739] = 32'b11111111111111110101000000110010;
assign LUT_1[18740] = 32'b00000000000000000111111001111100;
assign LUT_1[18741] = 32'b00000000000000000001001011111000;
assign LUT_1[18742] = 32'b00000000000000000011101000001101;
assign LUT_1[18743] = 32'b11111111111111111100111010001001;
assign LUT_1[18744] = 32'b11111111111111111111001110011010;
assign LUT_1[18745] = 32'b11111111111111111000100000010110;
assign LUT_1[18746] = 32'b11111111111111111010111100101011;
assign LUT_1[18747] = 32'b11111111111111110100001110100111;
assign LUT_1[18748] = 32'b00000000000000000111000111110001;
assign LUT_1[18749] = 32'b00000000000000000000011001101101;
assign LUT_1[18750] = 32'b00000000000000000010110110000010;
assign LUT_1[18751] = 32'b11111111111111111100000111111110;
assign LUT_1[18752] = 32'b11111111111111111111000111101100;
assign LUT_1[18753] = 32'b11111111111111111000011001101000;
assign LUT_1[18754] = 32'b11111111111111111010110101111101;
assign LUT_1[18755] = 32'b11111111111111110100000111111001;
assign LUT_1[18756] = 32'b00000000000000000111000001000011;
assign LUT_1[18757] = 32'b00000000000000000000010010111111;
assign LUT_1[18758] = 32'b00000000000000000010101111010100;
assign LUT_1[18759] = 32'b11111111111111111100000001010000;
assign LUT_1[18760] = 32'b11111111111111111110010101100001;
assign LUT_1[18761] = 32'b11111111111111110111100111011101;
assign LUT_1[18762] = 32'b11111111111111111010000011110010;
assign LUT_1[18763] = 32'b11111111111111110011010101101110;
assign LUT_1[18764] = 32'b00000000000000000110001110111000;
assign LUT_1[18765] = 32'b11111111111111111111100000110100;
assign LUT_1[18766] = 32'b00000000000000000001111101001001;
assign LUT_1[18767] = 32'b11111111111111111011001111000101;
assign LUT_1[18768] = 32'b00000000000000000001000011001110;
assign LUT_1[18769] = 32'b11111111111111111010010101001010;
assign LUT_1[18770] = 32'b11111111111111111100110001011111;
assign LUT_1[18771] = 32'b11111111111111110110000011011011;
assign LUT_1[18772] = 32'b00000000000000001000111100100101;
assign LUT_1[18773] = 32'b00000000000000000010001110100001;
assign LUT_1[18774] = 32'b00000000000000000100101010110110;
assign LUT_1[18775] = 32'b11111111111111111101111100110010;
assign LUT_1[18776] = 32'b00000000000000000000010001000011;
assign LUT_1[18777] = 32'b11111111111111111001100010111111;
assign LUT_1[18778] = 32'b11111111111111111011111111010100;
assign LUT_1[18779] = 32'b11111111111111110101010001010000;
assign LUT_1[18780] = 32'b00000000000000001000001010011010;
assign LUT_1[18781] = 32'b00000000000000000001011100010110;
assign LUT_1[18782] = 32'b00000000000000000011111000101011;
assign LUT_1[18783] = 32'b11111111111111111101001010100111;
assign LUT_1[18784] = 32'b00000000000000000000000010101011;
assign LUT_1[18785] = 32'b11111111111111111001010100100111;
assign LUT_1[18786] = 32'b11111111111111111011110000111100;
assign LUT_1[18787] = 32'b11111111111111110101000010111000;
assign LUT_1[18788] = 32'b00000000000000000111111100000010;
assign LUT_1[18789] = 32'b00000000000000000001001101111110;
assign LUT_1[18790] = 32'b00000000000000000011101010010011;
assign LUT_1[18791] = 32'b11111111111111111100111100001111;
assign LUT_1[18792] = 32'b11111111111111111111010000100000;
assign LUT_1[18793] = 32'b11111111111111111000100010011100;
assign LUT_1[18794] = 32'b11111111111111111010111110110001;
assign LUT_1[18795] = 32'b11111111111111110100010000101101;
assign LUT_1[18796] = 32'b00000000000000000111001001110111;
assign LUT_1[18797] = 32'b00000000000000000000011011110011;
assign LUT_1[18798] = 32'b00000000000000000010111000001000;
assign LUT_1[18799] = 32'b11111111111111111100001010000100;
assign LUT_1[18800] = 32'b00000000000000000001111110001101;
assign LUT_1[18801] = 32'b11111111111111111011010000001001;
assign LUT_1[18802] = 32'b11111111111111111101101100011110;
assign LUT_1[18803] = 32'b11111111111111110110111110011010;
assign LUT_1[18804] = 32'b00000000000000001001110111100100;
assign LUT_1[18805] = 32'b00000000000000000011001001100000;
assign LUT_1[18806] = 32'b00000000000000000101100101110101;
assign LUT_1[18807] = 32'b11111111111111111110110111110001;
assign LUT_1[18808] = 32'b00000000000000000001001100000010;
assign LUT_1[18809] = 32'b11111111111111111010011101111110;
assign LUT_1[18810] = 32'b11111111111111111100111010010011;
assign LUT_1[18811] = 32'b11111111111111110110001100001111;
assign LUT_1[18812] = 32'b00000000000000001001000101011001;
assign LUT_1[18813] = 32'b00000000000000000010010111010101;
assign LUT_1[18814] = 32'b00000000000000000100110011101010;
assign LUT_1[18815] = 32'b11111111111111111110000101100110;
assign LUT_1[18816] = 32'b00000000000000000000001010000111;
assign LUT_1[18817] = 32'b11111111111111111001011100000011;
assign LUT_1[18818] = 32'b11111111111111111011111000011000;
assign LUT_1[18819] = 32'b11111111111111110101001010010100;
assign LUT_1[18820] = 32'b00000000000000001000000011011110;
assign LUT_1[18821] = 32'b00000000000000000001010101011010;
assign LUT_1[18822] = 32'b00000000000000000011110001101111;
assign LUT_1[18823] = 32'b11111111111111111101000011101011;
assign LUT_1[18824] = 32'b11111111111111111111010111111100;
assign LUT_1[18825] = 32'b11111111111111111000101001111000;
assign LUT_1[18826] = 32'b11111111111111111011000110001101;
assign LUT_1[18827] = 32'b11111111111111110100011000001001;
assign LUT_1[18828] = 32'b00000000000000000111010001010011;
assign LUT_1[18829] = 32'b00000000000000000000100011001111;
assign LUT_1[18830] = 32'b00000000000000000010111111100100;
assign LUT_1[18831] = 32'b11111111111111111100010001100000;
assign LUT_1[18832] = 32'b00000000000000000010000101101001;
assign LUT_1[18833] = 32'b11111111111111111011010111100101;
assign LUT_1[18834] = 32'b11111111111111111101110011111010;
assign LUT_1[18835] = 32'b11111111111111110111000101110110;
assign LUT_1[18836] = 32'b00000000000000001001111111000000;
assign LUT_1[18837] = 32'b00000000000000000011010000111100;
assign LUT_1[18838] = 32'b00000000000000000101101101010001;
assign LUT_1[18839] = 32'b11111111111111111110111111001101;
assign LUT_1[18840] = 32'b00000000000000000001010011011110;
assign LUT_1[18841] = 32'b11111111111111111010100101011010;
assign LUT_1[18842] = 32'b11111111111111111101000001101111;
assign LUT_1[18843] = 32'b11111111111111110110010011101011;
assign LUT_1[18844] = 32'b00000000000000001001001100110101;
assign LUT_1[18845] = 32'b00000000000000000010011110110001;
assign LUT_1[18846] = 32'b00000000000000000100111011000110;
assign LUT_1[18847] = 32'b11111111111111111110001101000010;
assign LUT_1[18848] = 32'b00000000000000000001000101000110;
assign LUT_1[18849] = 32'b11111111111111111010010111000010;
assign LUT_1[18850] = 32'b11111111111111111100110011010111;
assign LUT_1[18851] = 32'b11111111111111110110000101010011;
assign LUT_1[18852] = 32'b00000000000000001000111110011101;
assign LUT_1[18853] = 32'b00000000000000000010010000011001;
assign LUT_1[18854] = 32'b00000000000000000100101100101110;
assign LUT_1[18855] = 32'b11111111111111111101111110101010;
assign LUT_1[18856] = 32'b00000000000000000000010010111011;
assign LUT_1[18857] = 32'b11111111111111111001100100110111;
assign LUT_1[18858] = 32'b11111111111111111100000001001100;
assign LUT_1[18859] = 32'b11111111111111110101010011001000;
assign LUT_1[18860] = 32'b00000000000000001000001100010010;
assign LUT_1[18861] = 32'b00000000000000000001011110001110;
assign LUT_1[18862] = 32'b00000000000000000011111010100011;
assign LUT_1[18863] = 32'b11111111111111111101001100011111;
assign LUT_1[18864] = 32'b00000000000000000011000000101000;
assign LUT_1[18865] = 32'b11111111111111111100010010100100;
assign LUT_1[18866] = 32'b11111111111111111110101110111001;
assign LUT_1[18867] = 32'b11111111111111111000000000110101;
assign LUT_1[18868] = 32'b00000000000000001010111001111111;
assign LUT_1[18869] = 32'b00000000000000000100001011111011;
assign LUT_1[18870] = 32'b00000000000000000110101000010000;
assign LUT_1[18871] = 32'b11111111111111111111111010001100;
assign LUT_1[18872] = 32'b00000000000000000010001110011101;
assign LUT_1[18873] = 32'b11111111111111111011100000011001;
assign LUT_1[18874] = 32'b11111111111111111101111100101110;
assign LUT_1[18875] = 32'b11111111111111110111001110101010;
assign LUT_1[18876] = 32'b00000000000000001010000111110100;
assign LUT_1[18877] = 32'b00000000000000000011011001110000;
assign LUT_1[18878] = 32'b00000000000000000101110110000101;
assign LUT_1[18879] = 32'b11111111111111111111001000000001;
assign LUT_1[18880] = 32'b00000000000000000010000111101111;
assign LUT_1[18881] = 32'b11111111111111111011011001101011;
assign LUT_1[18882] = 32'b11111111111111111101110110000000;
assign LUT_1[18883] = 32'b11111111111111110111000111111100;
assign LUT_1[18884] = 32'b00000000000000001010000001000110;
assign LUT_1[18885] = 32'b00000000000000000011010011000010;
assign LUT_1[18886] = 32'b00000000000000000101101111010111;
assign LUT_1[18887] = 32'b11111111111111111111000001010011;
assign LUT_1[18888] = 32'b00000000000000000001010101100100;
assign LUT_1[18889] = 32'b11111111111111111010100111100000;
assign LUT_1[18890] = 32'b11111111111111111101000011110101;
assign LUT_1[18891] = 32'b11111111111111110110010101110001;
assign LUT_1[18892] = 32'b00000000000000001001001110111011;
assign LUT_1[18893] = 32'b00000000000000000010100000110111;
assign LUT_1[18894] = 32'b00000000000000000100111101001100;
assign LUT_1[18895] = 32'b11111111111111111110001111001000;
assign LUT_1[18896] = 32'b00000000000000000100000011010001;
assign LUT_1[18897] = 32'b11111111111111111101010101001101;
assign LUT_1[18898] = 32'b11111111111111111111110001100010;
assign LUT_1[18899] = 32'b11111111111111111001000011011110;
assign LUT_1[18900] = 32'b00000000000000001011111100101000;
assign LUT_1[18901] = 32'b00000000000000000101001110100100;
assign LUT_1[18902] = 32'b00000000000000000111101010111001;
assign LUT_1[18903] = 32'b00000000000000000000111100110101;
assign LUT_1[18904] = 32'b00000000000000000011010001000110;
assign LUT_1[18905] = 32'b11111111111111111100100011000010;
assign LUT_1[18906] = 32'b11111111111111111110111111010111;
assign LUT_1[18907] = 32'b11111111111111111000010001010011;
assign LUT_1[18908] = 32'b00000000000000001011001010011101;
assign LUT_1[18909] = 32'b00000000000000000100011100011001;
assign LUT_1[18910] = 32'b00000000000000000110111000101110;
assign LUT_1[18911] = 32'b00000000000000000000001010101010;
assign LUT_1[18912] = 32'b00000000000000000011000010101110;
assign LUT_1[18913] = 32'b11111111111111111100010100101010;
assign LUT_1[18914] = 32'b11111111111111111110110000111111;
assign LUT_1[18915] = 32'b11111111111111111000000010111011;
assign LUT_1[18916] = 32'b00000000000000001010111100000101;
assign LUT_1[18917] = 32'b00000000000000000100001110000001;
assign LUT_1[18918] = 32'b00000000000000000110101010010110;
assign LUT_1[18919] = 32'b11111111111111111111111100010010;
assign LUT_1[18920] = 32'b00000000000000000010010000100011;
assign LUT_1[18921] = 32'b11111111111111111011100010011111;
assign LUT_1[18922] = 32'b11111111111111111101111110110100;
assign LUT_1[18923] = 32'b11111111111111110111010000110000;
assign LUT_1[18924] = 32'b00000000000000001010001001111010;
assign LUT_1[18925] = 32'b00000000000000000011011011110110;
assign LUT_1[18926] = 32'b00000000000000000101111000001011;
assign LUT_1[18927] = 32'b11111111111111111111001010000111;
assign LUT_1[18928] = 32'b00000000000000000100111110010000;
assign LUT_1[18929] = 32'b11111111111111111110010000001100;
assign LUT_1[18930] = 32'b00000000000000000000101100100001;
assign LUT_1[18931] = 32'b11111111111111111001111110011101;
assign LUT_1[18932] = 32'b00000000000000001100110111100111;
assign LUT_1[18933] = 32'b00000000000000000110001001100011;
assign LUT_1[18934] = 32'b00000000000000001000100101111000;
assign LUT_1[18935] = 32'b00000000000000000001110111110100;
assign LUT_1[18936] = 32'b00000000000000000100001100000101;
assign LUT_1[18937] = 32'b11111111111111111101011110000001;
assign LUT_1[18938] = 32'b11111111111111111111111010010110;
assign LUT_1[18939] = 32'b11111111111111111001001100010010;
assign LUT_1[18940] = 32'b00000000000000001100000101011100;
assign LUT_1[18941] = 32'b00000000000000000101010111011000;
assign LUT_1[18942] = 32'b00000000000000000111110011101101;
assign LUT_1[18943] = 32'b00000000000000000001000101101001;
assign LUT_1[18944] = 32'b11111111111111111001000100010101;
assign LUT_1[18945] = 32'b11111111111111110010010110010001;
assign LUT_1[18946] = 32'b11111111111111110100110010100110;
assign LUT_1[18947] = 32'b11111111111111101110000100100010;
assign LUT_1[18948] = 32'b00000000000000000000111101101100;
assign LUT_1[18949] = 32'b11111111111111111010001111101000;
assign LUT_1[18950] = 32'b11111111111111111100101011111101;
assign LUT_1[18951] = 32'b11111111111111110101111101111001;
assign LUT_1[18952] = 32'b11111111111111111000010010001010;
assign LUT_1[18953] = 32'b11111111111111110001100100000110;
assign LUT_1[18954] = 32'b11111111111111110100000000011011;
assign LUT_1[18955] = 32'b11111111111111101101010010010111;
assign LUT_1[18956] = 32'b00000000000000000000001011100001;
assign LUT_1[18957] = 32'b11111111111111111001011101011101;
assign LUT_1[18958] = 32'b11111111111111111011111001110010;
assign LUT_1[18959] = 32'b11111111111111110101001011101110;
assign LUT_1[18960] = 32'b11111111111111111010111111110111;
assign LUT_1[18961] = 32'b11111111111111110100010001110011;
assign LUT_1[18962] = 32'b11111111111111110110101110001000;
assign LUT_1[18963] = 32'b11111111111111110000000000000100;
assign LUT_1[18964] = 32'b00000000000000000010111001001110;
assign LUT_1[18965] = 32'b11111111111111111100001011001010;
assign LUT_1[18966] = 32'b11111111111111111110100111011111;
assign LUT_1[18967] = 32'b11111111111111110111111001011011;
assign LUT_1[18968] = 32'b11111111111111111010001101101100;
assign LUT_1[18969] = 32'b11111111111111110011011111101000;
assign LUT_1[18970] = 32'b11111111111111110101111011111101;
assign LUT_1[18971] = 32'b11111111111111101111001101111001;
assign LUT_1[18972] = 32'b00000000000000000010000111000011;
assign LUT_1[18973] = 32'b11111111111111111011011000111111;
assign LUT_1[18974] = 32'b11111111111111111101110101010100;
assign LUT_1[18975] = 32'b11111111111111110111000111010000;
assign LUT_1[18976] = 32'b11111111111111111001111111010100;
assign LUT_1[18977] = 32'b11111111111111110011010001010000;
assign LUT_1[18978] = 32'b11111111111111110101101101100101;
assign LUT_1[18979] = 32'b11111111111111101110111111100001;
assign LUT_1[18980] = 32'b00000000000000000001111000101011;
assign LUT_1[18981] = 32'b11111111111111111011001010100111;
assign LUT_1[18982] = 32'b11111111111111111101100110111100;
assign LUT_1[18983] = 32'b11111111111111110110111000111000;
assign LUT_1[18984] = 32'b11111111111111111001001101001001;
assign LUT_1[18985] = 32'b11111111111111110010011111000101;
assign LUT_1[18986] = 32'b11111111111111110100111011011010;
assign LUT_1[18987] = 32'b11111111111111101110001101010110;
assign LUT_1[18988] = 32'b00000000000000000001000110100000;
assign LUT_1[18989] = 32'b11111111111111111010011000011100;
assign LUT_1[18990] = 32'b11111111111111111100110100110001;
assign LUT_1[18991] = 32'b11111111111111110110000110101101;
assign LUT_1[18992] = 32'b11111111111111111011111010110110;
assign LUT_1[18993] = 32'b11111111111111110101001100110010;
assign LUT_1[18994] = 32'b11111111111111110111101001000111;
assign LUT_1[18995] = 32'b11111111111111110000111011000011;
assign LUT_1[18996] = 32'b00000000000000000011110100001101;
assign LUT_1[18997] = 32'b11111111111111111101000110001001;
assign LUT_1[18998] = 32'b11111111111111111111100010011110;
assign LUT_1[18999] = 32'b11111111111111111000110100011010;
assign LUT_1[19000] = 32'b11111111111111111011001000101011;
assign LUT_1[19001] = 32'b11111111111111110100011010100111;
assign LUT_1[19002] = 32'b11111111111111110110110110111100;
assign LUT_1[19003] = 32'b11111111111111110000001000111000;
assign LUT_1[19004] = 32'b00000000000000000011000010000010;
assign LUT_1[19005] = 32'b11111111111111111100010011111110;
assign LUT_1[19006] = 32'b11111111111111111110110000010011;
assign LUT_1[19007] = 32'b11111111111111111000000010001111;
assign LUT_1[19008] = 32'b11111111111111111011000001111101;
assign LUT_1[19009] = 32'b11111111111111110100010011111001;
assign LUT_1[19010] = 32'b11111111111111110110110000001110;
assign LUT_1[19011] = 32'b11111111111111110000000010001010;
assign LUT_1[19012] = 32'b00000000000000000010111011010100;
assign LUT_1[19013] = 32'b11111111111111111100001101010000;
assign LUT_1[19014] = 32'b11111111111111111110101001100101;
assign LUT_1[19015] = 32'b11111111111111110111111011100001;
assign LUT_1[19016] = 32'b11111111111111111010001111110010;
assign LUT_1[19017] = 32'b11111111111111110011100001101110;
assign LUT_1[19018] = 32'b11111111111111110101111110000011;
assign LUT_1[19019] = 32'b11111111111111101111001111111111;
assign LUT_1[19020] = 32'b00000000000000000010001001001001;
assign LUT_1[19021] = 32'b11111111111111111011011011000101;
assign LUT_1[19022] = 32'b11111111111111111101110111011010;
assign LUT_1[19023] = 32'b11111111111111110111001001010110;
assign LUT_1[19024] = 32'b11111111111111111100111101011111;
assign LUT_1[19025] = 32'b11111111111111110110001111011011;
assign LUT_1[19026] = 32'b11111111111111111000101011110000;
assign LUT_1[19027] = 32'b11111111111111110001111101101100;
assign LUT_1[19028] = 32'b00000000000000000100110110110110;
assign LUT_1[19029] = 32'b11111111111111111110001000110010;
assign LUT_1[19030] = 32'b00000000000000000000100101000111;
assign LUT_1[19031] = 32'b11111111111111111001110111000011;
assign LUT_1[19032] = 32'b11111111111111111100001011010100;
assign LUT_1[19033] = 32'b11111111111111110101011101010000;
assign LUT_1[19034] = 32'b11111111111111110111111001100101;
assign LUT_1[19035] = 32'b11111111111111110001001011100001;
assign LUT_1[19036] = 32'b00000000000000000100000100101011;
assign LUT_1[19037] = 32'b11111111111111111101010110100111;
assign LUT_1[19038] = 32'b11111111111111111111110010111100;
assign LUT_1[19039] = 32'b11111111111111111001000100111000;
assign LUT_1[19040] = 32'b11111111111111111011111100111100;
assign LUT_1[19041] = 32'b11111111111111110101001110111000;
assign LUT_1[19042] = 32'b11111111111111110111101011001101;
assign LUT_1[19043] = 32'b11111111111111110000111101001001;
assign LUT_1[19044] = 32'b00000000000000000011110110010011;
assign LUT_1[19045] = 32'b11111111111111111101001000001111;
assign LUT_1[19046] = 32'b11111111111111111111100100100100;
assign LUT_1[19047] = 32'b11111111111111111000110110100000;
assign LUT_1[19048] = 32'b11111111111111111011001010110001;
assign LUT_1[19049] = 32'b11111111111111110100011100101101;
assign LUT_1[19050] = 32'b11111111111111110110111001000010;
assign LUT_1[19051] = 32'b11111111111111110000001010111110;
assign LUT_1[19052] = 32'b00000000000000000011000100001000;
assign LUT_1[19053] = 32'b11111111111111111100010110000100;
assign LUT_1[19054] = 32'b11111111111111111110110010011001;
assign LUT_1[19055] = 32'b11111111111111111000000100010101;
assign LUT_1[19056] = 32'b11111111111111111101111000011110;
assign LUT_1[19057] = 32'b11111111111111110111001010011010;
assign LUT_1[19058] = 32'b11111111111111111001100110101111;
assign LUT_1[19059] = 32'b11111111111111110010111000101011;
assign LUT_1[19060] = 32'b00000000000000000101110001110101;
assign LUT_1[19061] = 32'b11111111111111111111000011110001;
assign LUT_1[19062] = 32'b00000000000000000001100000000110;
assign LUT_1[19063] = 32'b11111111111111111010110010000010;
assign LUT_1[19064] = 32'b11111111111111111101000110010011;
assign LUT_1[19065] = 32'b11111111111111110110011000001111;
assign LUT_1[19066] = 32'b11111111111111111000110100100100;
assign LUT_1[19067] = 32'b11111111111111110010000110100000;
assign LUT_1[19068] = 32'b00000000000000000100111111101010;
assign LUT_1[19069] = 32'b11111111111111111110010001100110;
assign LUT_1[19070] = 32'b00000000000000000000101101111011;
assign LUT_1[19071] = 32'b11111111111111111001111111110111;
assign LUT_1[19072] = 32'b11111111111111111100000100011000;
assign LUT_1[19073] = 32'b11111111111111110101010110010100;
assign LUT_1[19074] = 32'b11111111111111110111110010101001;
assign LUT_1[19075] = 32'b11111111111111110001000100100101;
assign LUT_1[19076] = 32'b00000000000000000011111101101111;
assign LUT_1[19077] = 32'b11111111111111111101001111101011;
assign LUT_1[19078] = 32'b11111111111111111111101100000000;
assign LUT_1[19079] = 32'b11111111111111111000111101111100;
assign LUT_1[19080] = 32'b11111111111111111011010010001101;
assign LUT_1[19081] = 32'b11111111111111110100100100001001;
assign LUT_1[19082] = 32'b11111111111111110111000000011110;
assign LUT_1[19083] = 32'b11111111111111110000010010011010;
assign LUT_1[19084] = 32'b00000000000000000011001011100100;
assign LUT_1[19085] = 32'b11111111111111111100011101100000;
assign LUT_1[19086] = 32'b11111111111111111110111001110101;
assign LUT_1[19087] = 32'b11111111111111111000001011110001;
assign LUT_1[19088] = 32'b11111111111111111101111111111010;
assign LUT_1[19089] = 32'b11111111111111110111010001110110;
assign LUT_1[19090] = 32'b11111111111111111001101110001011;
assign LUT_1[19091] = 32'b11111111111111110011000000000111;
assign LUT_1[19092] = 32'b00000000000000000101111001010001;
assign LUT_1[19093] = 32'b11111111111111111111001011001101;
assign LUT_1[19094] = 32'b00000000000000000001100111100010;
assign LUT_1[19095] = 32'b11111111111111111010111001011110;
assign LUT_1[19096] = 32'b11111111111111111101001101101111;
assign LUT_1[19097] = 32'b11111111111111110110011111101011;
assign LUT_1[19098] = 32'b11111111111111111000111100000000;
assign LUT_1[19099] = 32'b11111111111111110010001101111100;
assign LUT_1[19100] = 32'b00000000000000000101000111000110;
assign LUT_1[19101] = 32'b11111111111111111110011001000010;
assign LUT_1[19102] = 32'b00000000000000000000110101010111;
assign LUT_1[19103] = 32'b11111111111111111010000111010011;
assign LUT_1[19104] = 32'b11111111111111111100111111010111;
assign LUT_1[19105] = 32'b11111111111111110110010001010011;
assign LUT_1[19106] = 32'b11111111111111111000101101101000;
assign LUT_1[19107] = 32'b11111111111111110001111111100100;
assign LUT_1[19108] = 32'b00000000000000000100111000101110;
assign LUT_1[19109] = 32'b11111111111111111110001010101010;
assign LUT_1[19110] = 32'b00000000000000000000100110111111;
assign LUT_1[19111] = 32'b11111111111111111001111000111011;
assign LUT_1[19112] = 32'b11111111111111111100001101001100;
assign LUT_1[19113] = 32'b11111111111111110101011111001000;
assign LUT_1[19114] = 32'b11111111111111110111111011011101;
assign LUT_1[19115] = 32'b11111111111111110001001101011001;
assign LUT_1[19116] = 32'b00000000000000000100000110100011;
assign LUT_1[19117] = 32'b11111111111111111101011000011111;
assign LUT_1[19118] = 32'b11111111111111111111110100110100;
assign LUT_1[19119] = 32'b11111111111111111001000110110000;
assign LUT_1[19120] = 32'b11111111111111111110111010111001;
assign LUT_1[19121] = 32'b11111111111111111000001100110101;
assign LUT_1[19122] = 32'b11111111111111111010101001001010;
assign LUT_1[19123] = 32'b11111111111111110011111011000110;
assign LUT_1[19124] = 32'b00000000000000000110110100010000;
assign LUT_1[19125] = 32'b00000000000000000000000110001100;
assign LUT_1[19126] = 32'b00000000000000000010100010100001;
assign LUT_1[19127] = 32'b11111111111111111011110100011101;
assign LUT_1[19128] = 32'b11111111111111111110001000101110;
assign LUT_1[19129] = 32'b11111111111111110111011010101010;
assign LUT_1[19130] = 32'b11111111111111111001110110111111;
assign LUT_1[19131] = 32'b11111111111111110011001000111011;
assign LUT_1[19132] = 32'b00000000000000000110000010000101;
assign LUT_1[19133] = 32'b11111111111111111111010100000001;
assign LUT_1[19134] = 32'b00000000000000000001110000010110;
assign LUT_1[19135] = 32'b11111111111111111011000010010010;
assign LUT_1[19136] = 32'b11111111111111111110000010000000;
assign LUT_1[19137] = 32'b11111111111111110111010011111100;
assign LUT_1[19138] = 32'b11111111111111111001110000010001;
assign LUT_1[19139] = 32'b11111111111111110011000010001101;
assign LUT_1[19140] = 32'b00000000000000000101111011010111;
assign LUT_1[19141] = 32'b11111111111111111111001101010011;
assign LUT_1[19142] = 32'b00000000000000000001101001101000;
assign LUT_1[19143] = 32'b11111111111111111010111011100100;
assign LUT_1[19144] = 32'b11111111111111111101001111110101;
assign LUT_1[19145] = 32'b11111111111111110110100001110001;
assign LUT_1[19146] = 32'b11111111111111111000111110000110;
assign LUT_1[19147] = 32'b11111111111111110010010000000010;
assign LUT_1[19148] = 32'b00000000000000000101001001001100;
assign LUT_1[19149] = 32'b11111111111111111110011011001000;
assign LUT_1[19150] = 32'b00000000000000000000110111011101;
assign LUT_1[19151] = 32'b11111111111111111010001001011001;
assign LUT_1[19152] = 32'b11111111111111111111111101100010;
assign LUT_1[19153] = 32'b11111111111111111001001111011110;
assign LUT_1[19154] = 32'b11111111111111111011101011110011;
assign LUT_1[19155] = 32'b11111111111111110100111101101111;
assign LUT_1[19156] = 32'b00000000000000000111110110111001;
assign LUT_1[19157] = 32'b00000000000000000001001000110101;
assign LUT_1[19158] = 32'b00000000000000000011100101001010;
assign LUT_1[19159] = 32'b11111111111111111100110111000110;
assign LUT_1[19160] = 32'b11111111111111111111001011010111;
assign LUT_1[19161] = 32'b11111111111111111000011101010011;
assign LUT_1[19162] = 32'b11111111111111111010111001101000;
assign LUT_1[19163] = 32'b11111111111111110100001011100100;
assign LUT_1[19164] = 32'b00000000000000000111000100101110;
assign LUT_1[19165] = 32'b00000000000000000000010110101010;
assign LUT_1[19166] = 32'b00000000000000000010110010111111;
assign LUT_1[19167] = 32'b11111111111111111100000100111011;
assign LUT_1[19168] = 32'b11111111111111111110111100111111;
assign LUT_1[19169] = 32'b11111111111111111000001110111011;
assign LUT_1[19170] = 32'b11111111111111111010101011010000;
assign LUT_1[19171] = 32'b11111111111111110011111101001100;
assign LUT_1[19172] = 32'b00000000000000000110110110010110;
assign LUT_1[19173] = 32'b00000000000000000000001000010010;
assign LUT_1[19174] = 32'b00000000000000000010100100100111;
assign LUT_1[19175] = 32'b11111111111111111011110110100011;
assign LUT_1[19176] = 32'b11111111111111111110001010110100;
assign LUT_1[19177] = 32'b11111111111111110111011100110000;
assign LUT_1[19178] = 32'b11111111111111111001111001000101;
assign LUT_1[19179] = 32'b11111111111111110011001011000001;
assign LUT_1[19180] = 32'b00000000000000000110000100001011;
assign LUT_1[19181] = 32'b11111111111111111111010110000111;
assign LUT_1[19182] = 32'b00000000000000000001110010011100;
assign LUT_1[19183] = 32'b11111111111111111011000100011000;
assign LUT_1[19184] = 32'b00000000000000000000111000100001;
assign LUT_1[19185] = 32'b11111111111111111010001010011101;
assign LUT_1[19186] = 32'b11111111111111111100100110110010;
assign LUT_1[19187] = 32'b11111111111111110101111000101110;
assign LUT_1[19188] = 32'b00000000000000001000110001111000;
assign LUT_1[19189] = 32'b00000000000000000010000011110100;
assign LUT_1[19190] = 32'b00000000000000000100100000001001;
assign LUT_1[19191] = 32'b11111111111111111101110010000101;
assign LUT_1[19192] = 32'b00000000000000000000000110010110;
assign LUT_1[19193] = 32'b11111111111111111001011000010010;
assign LUT_1[19194] = 32'b11111111111111111011110100100111;
assign LUT_1[19195] = 32'b11111111111111110101000110100011;
assign LUT_1[19196] = 32'b00000000000000000111111111101101;
assign LUT_1[19197] = 32'b00000000000000000001010001101001;
assign LUT_1[19198] = 32'b00000000000000000011101101111110;
assign LUT_1[19199] = 32'b11111111111111111100111111111010;
assign LUT_1[19200] = 32'b11111111111111110110111000100001;
assign LUT_1[19201] = 32'b11111111111111110000001010011101;
assign LUT_1[19202] = 32'b11111111111111110010100110110010;
assign LUT_1[19203] = 32'b11111111111111101011111000101110;
assign LUT_1[19204] = 32'b11111111111111111110110001111000;
assign LUT_1[19205] = 32'b11111111111111111000000011110100;
assign LUT_1[19206] = 32'b11111111111111111010100000001001;
assign LUT_1[19207] = 32'b11111111111111110011110010000101;
assign LUT_1[19208] = 32'b11111111111111110110000110010110;
assign LUT_1[19209] = 32'b11111111111111101111011000010010;
assign LUT_1[19210] = 32'b11111111111111110001110100100111;
assign LUT_1[19211] = 32'b11111111111111101011000110100011;
assign LUT_1[19212] = 32'b11111111111111111101111111101101;
assign LUT_1[19213] = 32'b11111111111111110111010001101001;
assign LUT_1[19214] = 32'b11111111111111111001101101111110;
assign LUT_1[19215] = 32'b11111111111111110010111111111010;
assign LUT_1[19216] = 32'b11111111111111111000110100000011;
assign LUT_1[19217] = 32'b11111111111111110010000101111111;
assign LUT_1[19218] = 32'b11111111111111110100100010010100;
assign LUT_1[19219] = 32'b11111111111111101101110100010000;
assign LUT_1[19220] = 32'b00000000000000000000101101011010;
assign LUT_1[19221] = 32'b11111111111111111001111111010110;
assign LUT_1[19222] = 32'b11111111111111111100011011101011;
assign LUT_1[19223] = 32'b11111111111111110101101101100111;
assign LUT_1[19224] = 32'b11111111111111111000000001111000;
assign LUT_1[19225] = 32'b11111111111111110001010011110100;
assign LUT_1[19226] = 32'b11111111111111110011110000001001;
assign LUT_1[19227] = 32'b11111111111111101101000010000101;
assign LUT_1[19228] = 32'b11111111111111111111111011001111;
assign LUT_1[19229] = 32'b11111111111111111001001101001011;
assign LUT_1[19230] = 32'b11111111111111111011101001100000;
assign LUT_1[19231] = 32'b11111111111111110100111011011100;
assign LUT_1[19232] = 32'b11111111111111110111110011100000;
assign LUT_1[19233] = 32'b11111111111111110001000101011100;
assign LUT_1[19234] = 32'b11111111111111110011100001110001;
assign LUT_1[19235] = 32'b11111111111111101100110011101101;
assign LUT_1[19236] = 32'b11111111111111111111101100110111;
assign LUT_1[19237] = 32'b11111111111111111000111110110011;
assign LUT_1[19238] = 32'b11111111111111111011011011001000;
assign LUT_1[19239] = 32'b11111111111111110100101101000100;
assign LUT_1[19240] = 32'b11111111111111110111000001010101;
assign LUT_1[19241] = 32'b11111111111111110000010011010001;
assign LUT_1[19242] = 32'b11111111111111110010101111100110;
assign LUT_1[19243] = 32'b11111111111111101100000001100010;
assign LUT_1[19244] = 32'b11111111111111111110111010101100;
assign LUT_1[19245] = 32'b11111111111111111000001100101000;
assign LUT_1[19246] = 32'b11111111111111111010101000111101;
assign LUT_1[19247] = 32'b11111111111111110011111010111001;
assign LUT_1[19248] = 32'b11111111111111111001101111000010;
assign LUT_1[19249] = 32'b11111111111111110011000000111110;
assign LUT_1[19250] = 32'b11111111111111110101011101010011;
assign LUT_1[19251] = 32'b11111111111111101110101111001111;
assign LUT_1[19252] = 32'b00000000000000000001101000011001;
assign LUT_1[19253] = 32'b11111111111111111010111010010101;
assign LUT_1[19254] = 32'b11111111111111111101010110101010;
assign LUT_1[19255] = 32'b11111111111111110110101000100110;
assign LUT_1[19256] = 32'b11111111111111111000111100110111;
assign LUT_1[19257] = 32'b11111111111111110010001110110011;
assign LUT_1[19258] = 32'b11111111111111110100101011001000;
assign LUT_1[19259] = 32'b11111111111111101101111101000100;
assign LUT_1[19260] = 32'b00000000000000000000110110001110;
assign LUT_1[19261] = 32'b11111111111111111010001000001010;
assign LUT_1[19262] = 32'b11111111111111111100100100011111;
assign LUT_1[19263] = 32'b11111111111111110101110110011011;
assign LUT_1[19264] = 32'b11111111111111111000110110001001;
assign LUT_1[19265] = 32'b11111111111111110010001000000101;
assign LUT_1[19266] = 32'b11111111111111110100100100011010;
assign LUT_1[19267] = 32'b11111111111111101101110110010110;
assign LUT_1[19268] = 32'b00000000000000000000101111100000;
assign LUT_1[19269] = 32'b11111111111111111010000001011100;
assign LUT_1[19270] = 32'b11111111111111111100011101110001;
assign LUT_1[19271] = 32'b11111111111111110101101111101101;
assign LUT_1[19272] = 32'b11111111111111111000000011111110;
assign LUT_1[19273] = 32'b11111111111111110001010101111010;
assign LUT_1[19274] = 32'b11111111111111110011110010001111;
assign LUT_1[19275] = 32'b11111111111111101101000100001011;
assign LUT_1[19276] = 32'b11111111111111111111111101010101;
assign LUT_1[19277] = 32'b11111111111111111001001111010001;
assign LUT_1[19278] = 32'b11111111111111111011101011100110;
assign LUT_1[19279] = 32'b11111111111111110100111101100010;
assign LUT_1[19280] = 32'b11111111111111111010110001101011;
assign LUT_1[19281] = 32'b11111111111111110100000011100111;
assign LUT_1[19282] = 32'b11111111111111110110011111111100;
assign LUT_1[19283] = 32'b11111111111111101111110001111000;
assign LUT_1[19284] = 32'b00000000000000000010101011000010;
assign LUT_1[19285] = 32'b11111111111111111011111100111110;
assign LUT_1[19286] = 32'b11111111111111111110011001010011;
assign LUT_1[19287] = 32'b11111111111111110111101011001111;
assign LUT_1[19288] = 32'b11111111111111111001111111100000;
assign LUT_1[19289] = 32'b11111111111111110011010001011100;
assign LUT_1[19290] = 32'b11111111111111110101101101110001;
assign LUT_1[19291] = 32'b11111111111111101110111111101101;
assign LUT_1[19292] = 32'b00000000000000000001111000110111;
assign LUT_1[19293] = 32'b11111111111111111011001010110011;
assign LUT_1[19294] = 32'b11111111111111111101100111001000;
assign LUT_1[19295] = 32'b11111111111111110110111001000100;
assign LUT_1[19296] = 32'b11111111111111111001110001001000;
assign LUT_1[19297] = 32'b11111111111111110011000011000100;
assign LUT_1[19298] = 32'b11111111111111110101011111011001;
assign LUT_1[19299] = 32'b11111111111111101110110001010101;
assign LUT_1[19300] = 32'b00000000000000000001101010011111;
assign LUT_1[19301] = 32'b11111111111111111010111100011011;
assign LUT_1[19302] = 32'b11111111111111111101011000110000;
assign LUT_1[19303] = 32'b11111111111111110110101010101100;
assign LUT_1[19304] = 32'b11111111111111111000111110111101;
assign LUT_1[19305] = 32'b11111111111111110010010000111001;
assign LUT_1[19306] = 32'b11111111111111110100101101001110;
assign LUT_1[19307] = 32'b11111111111111101101111111001010;
assign LUT_1[19308] = 32'b00000000000000000000111000010100;
assign LUT_1[19309] = 32'b11111111111111111010001010010000;
assign LUT_1[19310] = 32'b11111111111111111100100110100101;
assign LUT_1[19311] = 32'b11111111111111110101111000100001;
assign LUT_1[19312] = 32'b11111111111111111011101100101010;
assign LUT_1[19313] = 32'b11111111111111110100111110100110;
assign LUT_1[19314] = 32'b11111111111111110111011010111011;
assign LUT_1[19315] = 32'b11111111111111110000101100110111;
assign LUT_1[19316] = 32'b00000000000000000011100110000001;
assign LUT_1[19317] = 32'b11111111111111111100110111111101;
assign LUT_1[19318] = 32'b11111111111111111111010100010010;
assign LUT_1[19319] = 32'b11111111111111111000100110001110;
assign LUT_1[19320] = 32'b11111111111111111010111010011111;
assign LUT_1[19321] = 32'b11111111111111110100001100011011;
assign LUT_1[19322] = 32'b11111111111111110110101000110000;
assign LUT_1[19323] = 32'b11111111111111101111111010101100;
assign LUT_1[19324] = 32'b00000000000000000010110011110110;
assign LUT_1[19325] = 32'b11111111111111111100000101110010;
assign LUT_1[19326] = 32'b11111111111111111110100010000111;
assign LUT_1[19327] = 32'b11111111111111110111110100000011;
assign LUT_1[19328] = 32'b11111111111111111001111000100100;
assign LUT_1[19329] = 32'b11111111111111110011001010100000;
assign LUT_1[19330] = 32'b11111111111111110101100110110101;
assign LUT_1[19331] = 32'b11111111111111101110111000110001;
assign LUT_1[19332] = 32'b00000000000000000001110001111011;
assign LUT_1[19333] = 32'b11111111111111111011000011110111;
assign LUT_1[19334] = 32'b11111111111111111101100000001100;
assign LUT_1[19335] = 32'b11111111111111110110110010001000;
assign LUT_1[19336] = 32'b11111111111111111001000110011001;
assign LUT_1[19337] = 32'b11111111111111110010011000010101;
assign LUT_1[19338] = 32'b11111111111111110100110100101010;
assign LUT_1[19339] = 32'b11111111111111101110000110100110;
assign LUT_1[19340] = 32'b00000000000000000000111111110000;
assign LUT_1[19341] = 32'b11111111111111111010010001101100;
assign LUT_1[19342] = 32'b11111111111111111100101110000001;
assign LUT_1[19343] = 32'b11111111111111110101111111111101;
assign LUT_1[19344] = 32'b11111111111111111011110100000110;
assign LUT_1[19345] = 32'b11111111111111110101000110000010;
assign LUT_1[19346] = 32'b11111111111111110111100010010111;
assign LUT_1[19347] = 32'b11111111111111110000110100010011;
assign LUT_1[19348] = 32'b00000000000000000011101101011101;
assign LUT_1[19349] = 32'b11111111111111111100111111011001;
assign LUT_1[19350] = 32'b11111111111111111111011011101110;
assign LUT_1[19351] = 32'b11111111111111111000101101101010;
assign LUT_1[19352] = 32'b11111111111111111011000001111011;
assign LUT_1[19353] = 32'b11111111111111110100010011110111;
assign LUT_1[19354] = 32'b11111111111111110110110000001100;
assign LUT_1[19355] = 32'b11111111111111110000000010001000;
assign LUT_1[19356] = 32'b00000000000000000010111011010010;
assign LUT_1[19357] = 32'b11111111111111111100001101001110;
assign LUT_1[19358] = 32'b11111111111111111110101001100011;
assign LUT_1[19359] = 32'b11111111111111110111111011011111;
assign LUT_1[19360] = 32'b11111111111111111010110011100011;
assign LUT_1[19361] = 32'b11111111111111110100000101011111;
assign LUT_1[19362] = 32'b11111111111111110110100001110100;
assign LUT_1[19363] = 32'b11111111111111101111110011110000;
assign LUT_1[19364] = 32'b00000000000000000010101100111010;
assign LUT_1[19365] = 32'b11111111111111111011111110110110;
assign LUT_1[19366] = 32'b11111111111111111110011011001011;
assign LUT_1[19367] = 32'b11111111111111110111101101000111;
assign LUT_1[19368] = 32'b11111111111111111010000001011000;
assign LUT_1[19369] = 32'b11111111111111110011010011010100;
assign LUT_1[19370] = 32'b11111111111111110101101111101001;
assign LUT_1[19371] = 32'b11111111111111101111000001100101;
assign LUT_1[19372] = 32'b00000000000000000001111010101111;
assign LUT_1[19373] = 32'b11111111111111111011001100101011;
assign LUT_1[19374] = 32'b11111111111111111101101001000000;
assign LUT_1[19375] = 32'b11111111111111110110111010111100;
assign LUT_1[19376] = 32'b11111111111111111100101111000101;
assign LUT_1[19377] = 32'b11111111111111110110000001000001;
assign LUT_1[19378] = 32'b11111111111111111000011101010110;
assign LUT_1[19379] = 32'b11111111111111110001101111010010;
assign LUT_1[19380] = 32'b00000000000000000100101000011100;
assign LUT_1[19381] = 32'b11111111111111111101111010011000;
assign LUT_1[19382] = 32'b00000000000000000000010110101101;
assign LUT_1[19383] = 32'b11111111111111111001101000101001;
assign LUT_1[19384] = 32'b11111111111111111011111100111010;
assign LUT_1[19385] = 32'b11111111111111110101001110110110;
assign LUT_1[19386] = 32'b11111111111111110111101011001011;
assign LUT_1[19387] = 32'b11111111111111110000111101000111;
assign LUT_1[19388] = 32'b00000000000000000011110110010001;
assign LUT_1[19389] = 32'b11111111111111111101001000001101;
assign LUT_1[19390] = 32'b11111111111111111111100100100010;
assign LUT_1[19391] = 32'b11111111111111111000110110011110;
assign LUT_1[19392] = 32'b11111111111111111011110110001100;
assign LUT_1[19393] = 32'b11111111111111110101001000001000;
assign LUT_1[19394] = 32'b11111111111111110111100100011101;
assign LUT_1[19395] = 32'b11111111111111110000110110011001;
assign LUT_1[19396] = 32'b00000000000000000011101111100011;
assign LUT_1[19397] = 32'b11111111111111111101000001011111;
assign LUT_1[19398] = 32'b11111111111111111111011101110100;
assign LUT_1[19399] = 32'b11111111111111111000101111110000;
assign LUT_1[19400] = 32'b11111111111111111011000100000001;
assign LUT_1[19401] = 32'b11111111111111110100010101111101;
assign LUT_1[19402] = 32'b11111111111111110110110010010010;
assign LUT_1[19403] = 32'b11111111111111110000000100001110;
assign LUT_1[19404] = 32'b00000000000000000010111101011000;
assign LUT_1[19405] = 32'b11111111111111111100001111010100;
assign LUT_1[19406] = 32'b11111111111111111110101011101001;
assign LUT_1[19407] = 32'b11111111111111110111111101100101;
assign LUT_1[19408] = 32'b11111111111111111101110001101110;
assign LUT_1[19409] = 32'b11111111111111110111000011101010;
assign LUT_1[19410] = 32'b11111111111111111001011111111111;
assign LUT_1[19411] = 32'b11111111111111110010110001111011;
assign LUT_1[19412] = 32'b00000000000000000101101011000101;
assign LUT_1[19413] = 32'b11111111111111111110111101000001;
assign LUT_1[19414] = 32'b00000000000000000001011001010110;
assign LUT_1[19415] = 32'b11111111111111111010101011010010;
assign LUT_1[19416] = 32'b11111111111111111100111111100011;
assign LUT_1[19417] = 32'b11111111111111110110010001011111;
assign LUT_1[19418] = 32'b11111111111111111000101101110100;
assign LUT_1[19419] = 32'b11111111111111110001111111110000;
assign LUT_1[19420] = 32'b00000000000000000100111000111010;
assign LUT_1[19421] = 32'b11111111111111111110001010110110;
assign LUT_1[19422] = 32'b00000000000000000000100111001011;
assign LUT_1[19423] = 32'b11111111111111111001111001000111;
assign LUT_1[19424] = 32'b11111111111111111100110001001011;
assign LUT_1[19425] = 32'b11111111111111110110000011000111;
assign LUT_1[19426] = 32'b11111111111111111000011111011100;
assign LUT_1[19427] = 32'b11111111111111110001110001011000;
assign LUT_1[19428] = 32'b00000000000000000100101010100010;
assign LUT_1[19429] = 32'b11111111111111111101111100011110;
assign LUT_1[19430] = 32'b00000000000000000000011000110011;
assign LUT_1[19431] = 32'b11111111111111111001101010101111;
assign LUT_1[19432] = 32'b11111111111111111011111111000000;
assign LUT_1[19433] = 32'b11111111111111110101010000111100;
assign LUT_1[19434] = 32'b11111111111111110111101101010001;
assign LUT_1[19435] = 32'b11111111111111110000111111001101;
assign LUT_1[19436] = 32'b00000000000000000011111000010111;
assign LUT_1[19437] = 32'b11111111111111111101001010010011;
assign LUT_1[19438] = 32'b11111111111111111111100110101000;
assign LUT_1[19439] = 32'b11111111111111111000111000100100;
assign LUT_1[19440] = 32'b11111111111111111110101100101101;
assign LUT_1[19441] = 32'b11111111111111110111111110101001;
assign LUT_1[19442] = 32'b11111111111111111010011010111110;
assign LUT_1[19443] = 32'b11111111111111110011101100111010;
assign LUT_1[19444] = 32'b00000000000000000110100110000100;
assign LUT_1[19445] = 32'b11111111111111111111111000000000;
assign LUT_1[19446] = 32'b00000000000000000010010100010101;
assign LUT_1[19447] = 32'b11111111111111111011100110010001;
assign LUT_1[19448] = 32'b11111111111111111101111010100010;
assign LUT_1[19449] = 32'b11111111111111110111001100011110;
assign LUT_1[19450] = 32'b11111111111111111001101000110011;
assign LUT_1[19451] = 32'b11111111111111110010111010101111;
assign LUT_1[19452] = 32'b00000000000000000101110011111001;
assign LUT_1[19453] = 32'b11111111111111111111000101110101;
assign LUT_1[19454] = 32'b00000000000000000001100010001010;
assign LUT_1[19455] = 32'b11111111111111111010110100000110;
assign LUT_1[19456] = 32'b00000000000000000101101100101000;
assign LUT_1[19457] = 32'b11111111111111111110111110100100;
assign LUT_1[19458] = 32'b00000000000000000001011010111001;
assign LUT_1[19459] = 32'b11111111111111111010101100110101;
assign LUT_1[19460] = 32'b00000000000000001101100101111111;
assign LUT_1[19461] = 32'b00000000000000000110110111111011;
assign LUT_1[19462] = 32'b00000000000000001001010100010000;
assign LUT_1[19463] = 32'b00000000000000000010100110001100;
assign LUT_1[19464] = 32'b00000000000000000100111010011101;
assign LUT_1[19465] = 32'b11111111111111111110001100011001;
assign LUT_1[19466] = 32'b00000000000000000000101000101110;
assign LUT_1[19467] = 32'b11111111111111111001111010101010;
assign LUT_1[19468] = 32'b00000000000000001100110011110100;
assign LUT_1[19469] = 32'b00000000000000000110000101110000;
assign LUT_1[19470] = 32'b00000000000000001000100010000101;
assign LUT_1[19471] = 32'b00000000000000000001110100000001;
assign LUT_1[19472] = 32'b00000000000000000111101000001010;
assign LUT_1[19473] = 32'b00000000000000000000111010000110;
assign LUT_1[19474] = 32'b00000000000000000011010110011011;
assign LUT_1[19475] = 32'b11111111111111111100101000010111;
assign LUT_1[19476] = 32'b00000000000000001111100001100001;
assign LUT_1[19477] = 32'b00000000000000001000110011011101;
assign LUT_1[19478] = 32'b00000000000000001011001111110010;
assign LUT_1[19479] = 32'b00000000000000000100100001101110;
assign LUT_1[19480] = 32'b00000000000000000110110101111111;
assign LUT_1[19481] = 32'b00000000000000000000000111111011;
assign LUT_1[19482] = 32'b00000000000000000010100100010000;
assign LUT_1[19483] = 32'b11111111111111111011110110001100;
assign LUT_1[19484] = 32'b00000000000000001110101111010110;
assign LUT_1[19485] = 32'b00000000000000001000000001010010;
assign LUT_1[19486] = 32'b00000000000000001010011101100111;
assign LUT_1[19487] = 32'b00000000000000000011101111100011;
assign LUT_1[19488] = 32'b00000000000000000110100111100111;
assign LUT_1[19489] = 32'b11111111111111111111111001100011;
assign LUT_1[19490] = 32'b00000000000000000010010101111000;
assign LUT_1[19491] = 32'b11111111111111111011100111110100;
assign LUT_1[19492] = 32'b00000000000000001110100000111110;
assign LUT_1[19493] = 32'b00000000000000000111110010111010;
assign LUT_1[19494] = 32'b00000000000000001010001111001111;
assign LUT_1[19495] = 32'b00000000000000000011100001001011;
assign LUT_1[19496] = 32'b00000000000000000101110101011100;
assign LUT_1[19497] = 32'b11111111111111111111000111011000;
assign LUT_1[19498] = 32'b00000000000000000001100011101101;
assign LUT_1[19499] = 32'b11111111111111111010110101101001;
assign LUT_1[19500] = 32'b00000000000000001101101110110011;
assign LUT_1[19501] = 32'b00000000000000000111000000101111;
assign LUT_1[19502] = 32'b00000000000000001001011101000100;
assign LUT_1[19503] = 32'b00000000000000000010101111000000;
assign LUT_1[19504] = 32'b00000000000000001000100011001001;
assign LUT_1[19505] = 32'b00000000000000000001110101000101;
assign LUT_1[19506] = 32'b00000000000000000100010001011010;
assign LUT_1[19507] = 32'b11111111111111111101100011010110;
assign LUT_1[19508] = 32'b00000000000000010000011100100000;
assign LUT_1[19509] = 32'b00000000000000001001101110011100;
assign LUT_1[19510] = 32'b00000000000000001100001010110001;
assign LUT_1[19511] = 32'b00000000000000000101011100101101;
assign LUT_1[19512] = 32'b00000000000000000111110000111110;
assign LUT_1[19513] = 32'b00000000000000000001000010111010;
assign LUT_1[19514] = 32'b00000000000000000011011111001111;
assign LUT_1[19515] = 32'b11111111111111111100110001001011;
assign LUT_1[19516] = 32'b00000000000000001111101010010101;
assign LUT_1[19517] = 32'b00000000000000001000111100010001;
assign LUT_1[19518] = 32'b00000000000000001011011000100110;
assign LUT_1[19519] = 32'b00000000000000000100101010100010;
assign LUT_1[19520] = 32'b00000000000000000111101010010000;
assign LUT_1[19521] = 32'b00000000000000000000111100001100;
assign LUT_1[19522] = 32'b00000000000000000011011000100001;
assign LUT_1[19523] = 32'b11111111111111111100101010011101;
assign LUT_1[19524] = 32'b00000000000000001111100011100111;
assign LUT_1[19525] = 32'b00000000000000001000110101100011;
assign LUT_1[19526] = 32'b00000000000000001011010001111000;
assign LUT_1[19527] = 32'b00000000000000000100100011110100;
assign LUT_1[19528] = 32'b00000000000000000110111000000101;
assign LUT_1[19529] = 32'b00000000000000000000001010000001;
assign LUT_1[19530] = 32'b00000000000000000010100110010110;
assign LUT_1[19531] = 32'b11111111111111111011111000010010;
assign LUT_1[19532] = 32'b00000000000000001110110001011100;
assign LUT_1[19533] = 32'b00000000000000001000000011011000;
assign LUT_1[19534] = 32'b00000000000000001010011111101101;
assign LUT_1[19535] = 32'b00000000000000000011110001101001;
assign LUT_1[19536] = 32'b00000000000000001001100101110010;
assign LUT_1[19537] = 32'b00000000000000000010110111101110;
assign LUT_1[19538] = 32'b00000000000000000101010100000011;
assign LUT_1[19539] = 32'b11111111111111111110100101111111;
assign LUT_1[19540] = 32'b00000000000000010001011111001001;
assign LUT_1[19541] = 32'b00000000000000001010110001000101;
assign LUT_1[19542] = 32'b00000000000000001101001101011010;
assign LUT_1[19543] = 32'b00000000000000000110011111010110;
assign LUT_1[19544] = 32'b00000000000000001000110011100111;
assign LUT_1[19545] = 32'b00000000000000000010000101100011;
assign LUT_1[19546] = 32'b00000000000000000100100001111000;
assign LUT_1[19547] = 32'b11111111111111111101110011110100;
assign LUT_1[19548] = 32'b00000000000000010000101100111110;
assign LUT_1[19549] = 32'b00000000000000001001111110111010;
assign LUT_1[19550] = 32'b00000000000000001100011011001111;
assign LUT_1[19551] = 32'b00000000000000000101101101001011;
assign LUT_1[19552] = 32'b00000000000000001000100101001111;
assign LUT_1[19553] = 32'b00000000000000000001110111001011;
assign LUT_1[19554] = 32'b00000000000000000100010011100000;
assign LUT_1[19555] = 32'b11111111111111111101100101011100;
assign LUT_1[19556] = 32'b00000000000000010000011110100110;
assign LUT_1[19557] = 32'b00000000000000001001110000100010;
assign LUT_1[19558] = 32'b00000000000000001100001100110111;
assign LUT_1[19559] = 32'b00000000000000000101011110110011;
assign LUT_1[19560] = 32'b00000000000000000111110011000100;
assign LUT_1[19561] = 32'b00000000000000000001000101000000;
assign LUT_1[19562] = 32'b00000000000000000011100001010101;
assign LUT_1[19563] = 32'b11111111111111111100110011010001;
assign LUT_1[19564] = 32'b00000000000000001111101100011011;
assign LUT_1[19565] = 32'b00000000000000001000111110010111;
assign LUT_1[19566] = 32'b00000000000000001011011010101100;
assign LUT_1[19567] = 32'b00000000000000000100101100101000;
assign LUT_1[19568] = 32'b00000000000000001010100000110001;
assign LUT_1[19569] = 32'b00000000000000000011110010101101;
assign LUT_1[19570] = 32'b00000000000000000110001111000010;
assign LUT_1[19571] = 32'b11111111111111111111100000111110;
assign LUT_1[19572] = 32'b00000000000000010010011010001000;
assign LUT_1[19573] = 32'b00000000000000001011101100000100;
assign LUT_1[19574] = 32'b00000000000000001110001000011001;
assign LUT_1[19575] = 32'b00000000000000000111011010010101;
assign LUT_1[19576] = 32'b00000000000000001001101110100110;
assign LUT_1[19577] = 32'b00000000000000000011000000100010;
assign LUT_1[19578] = 32'b00000000000000000101011100110111;
assign LUT_1[19579] = 32'b11111111111111111110101110110011;
assign LUT_1[19580] = 32'b00000000000000010001100111111101;
assign LUT_1[19581] = 32'b00000000000000001010111001111001;
assign LUT_1[19582] = 32'b00000000000000001101010110001110;
assign LUT_1[19583] = 32'b00000000000000000110101000001010;
assign LUT_1[19584] = 32'b00000000000000001000101100101011;
assign LUT_1[19585] = 32'b00000000000000000001111110100111;
assign LUT_1[19586] = 32'b00000000000000000100011010111100;
assign LUT_1[19587] = 32'b11111111111111111101101100111000;
assign LUT_1[19588] = 32'b00000000000000010000100110000010;
assign LUT_1[19589] = 32'b00000000000000001001110111111110;
assign LUT_1[19590] = 32'b00000000000000001100010100010011;
assign LUT_1[19591] = 32'b00000000000000000101100110001111;
assign LUT_1[19592] = 32'b00000000000000000111111010100000;
assign LUT_1[19593] = 32'b00000000000000000001001100011100;
assign LUT_1[19594] = 32'b00000000000000000011101000110001;
assign LUT_1[19595] = 32'b11111111111111111100111010101101;
assign LUT_1[19596] = 32'b00000000000000001111110011110111;
assign LUT_1[19597] = 32'b00000000000000001001000101110011;
assign LUT_1[19598] = 32'b00000000000000001011100010001000;
assign LUT_1[19599] = 32'b00000000000000000100110100000100;
assign LUT_1[19600] = 32'b00000000000000001010101000001101;
assign LUT_1[19601] = 32'b00000000000000000011111010001001;
assign LUT_1[19602] = 32'b00000000000000000110010110011110;
assign LUT_1[19603] = 32'b11111111111111111111101000011010;
assign LUT_1[19604] = 32'b00000000000000010010100001100100;
assign LUT_1[19605] = 32'b00000000000000001011110011100000;
assign LUT_1[19606] = 32'b00000000000000001110001111110101;
assign LUT_1[19607] = 32'b00000000000000000111100001110001;
assign LUT_1[19608] = 32'b00000000000000001001110110000010;
assign LUT_1[19609] = 32'b00000000000000000011000111111110;
assign LUT_1[19610] = 32'b00000000000000000101100100010011;
assign LUT_1[19611] = 32'b11111111111111111110110110001111;
assign LUT_1[19612] = 32'b00000000000000010001101111011001;
assign LUT_1[19613] = 32'b00000000000000001011000001010101;
assign LUT_1[19614] = 32'b00000000000000001101011101101010;
assign LUT_1[19615] = 32'b00000000000000000110101111100110;
assign LUT_1[19616] = 32'b00000000000000001001100111101010;
assign LUT_1[19617] = 32'b00000000000000000010111001100110;
assign LUT_1[19618] = 32'b00000000000000000101010101111011;
assign LUT_1[19619] = 32'b11111111111111111110100111110111;
assign LUT_1[19620] = 32'b00000000000000010001100001000001;
assign LUT_1[19621] = 32'b00000000000000001010110010111101;
assign LUT_1[19622] = 32'b00000000000000001101001111010010;
assign LUT_1[19623] = 32'b00000000000000000110100001001110;
assign LUT_1[19624] = 32'b00000000000000001000110101011111;
assign LUT_1[19625] = 32'b00000000000000000010000111011011;
assign LUT_1[19626] = 32'b00000000000000000100100011110000;
assign LUT_1[19627] = 32'b11111111111111111101110101101100;
assign LUT_1[19628] = 32'b00000000000000010000101110110110;
assign LUT_1[19629] = 32'b00000000000000001010000000110010;
assign LUT_1[19630] = 32'b00000000000000001100011101000111;
assign LUT_1[19631] = 32'b00000000000000000101101111000011;
assign LUT_1[19632] = 32'b00000000000000001011100011001100;
assign LUT_1[19633] = 32'b00000000000000000100110101001000;
assign LUT_1[19634] = 32'b00000000000000000111010001011101;
assign LUT_1[19635] = 32'b00000000000000000000100011011001;
assign LUT_1[19636] = 32'b00000000000000010011011100100011;
assign LUT_1[19637] = 32'b00000000000000001100101110011111;
assign LUT_1[19638] = 32'b00000000000000001111001010110100;
assign LUT_1[19639] = 32'b00000000000000001000011100110000;
assign LUT_1[19640] = 32'b00000000000000001010110001000001;
assign LUT_1[19641] = 32'b00000000000000000100000010111101;
assign LUT_1[19642] = 32'b00000000000000000110011111010010;
assign LUT_1[19643] = 32'b11111111111111111111110001001110;
assign LUT_1[19644] = 32'b00000000000000010010101010011000;
assign LUT_1[19645] = 32'b00000000000000001011111100010100;
assign LUT_1[19646] = 32'b00000000000000001110011000101001;
assign LUT_1[19647] = 32'b00000000000000000111101010100101;
assign LUT_1[19648] = 32'b00000000000000001010101010010011;
assign LUT_1[19649] = 32'b00000000000000000011111100001111;
assign LUT_1[19650] = 32'b00000000000000000110011000100100;
assign LUT_1[19651] = 32'b11111111111111111111101010100000;
assign LUT_1[19652] = 32'b00000000000000010010100011101010;
assign LUT_1[19653] = 32'b00000000000000001011110101100110;
assign LUT_1[19654] = 32'b00000000000000001110010001111011;
assign LUT_1[19655] = 32'b00000000000000000111100011110111;
assign LUT_1[19656] = 32'b00000000000000001001111000001000;
assign LUT_1[19657] = 32'b00000000000000000011001010000100;
assign LUT_1[19658] = 32'b00000000000000000101100110011001;
assign LUT_1[19659] = 32'b11111111111111111110111000010101;
assign LUT_1[19660] = 32'b00000000000000010001110001011111;
assign LUT_1[19661] = 32'b00000000000000001011000011011011;
assign LUT_1[19662] = 32'b00000000000000001101011111110000;
assign LUT_1[19663] = 32'b00000000000000000110110001101100;
assign LUT_1[19664] = 32'b00000000000000001100100101110101;
assign LUT_1[19665] = 32'b00000000000000000101110111110001;
assign LUT_1[19666] = 32'b00000000000000001000010100000110;
assign LUT_1[19667] = 32'b00000000000000000001100110000010;
assign LUT_1[19668] = 32'b00000000000000010100011111001100;
assign LUT_1[19669] = 32'b00000000000000001101110001001000;
assign LUT_1[19670] = 32'b00000000000000010000001101011101;
assign LUT_1[19671] = 32'b00000000000000001001011111011001;
assign LUT_1[19672] = 32'b00000000000000001011110011101010;
assign LUT_1[19673] = 32'b00000000000000000101000101100110;
assign LUT_1[19674] = 32'b00000000000000000111100001111011;
assign LUT_1[19675] = 32'b00000000000000000000110011110111;
assign LUT_1[19676] = 32'b00000000000000010011101101000001;
assign LUT_1[19677] = 32'b00000000000000001100111110111101;
assign LUT_1[19678] = 32'b00000000000000001111011011010010;
assign LUT_1[19679] = 32'b00000000000000001000101101001110;
assign LUT_1[19680] = 32'b00000000000000001011100101010010;
assign LUT_1[19681] = 32'b00000000000000000100110111001110;
assign LUT_1[19682] = 32'b00000000000000000111010011100011;
assign LUT_1[19683] = 32'b00000000000000000000100101011111;
assign LUT_1[19684] = 32'b00000000000000010011011110101001;
assign LUT_1[19685] = 32'b00000000000000001100110000100101;
assign LUT_1[19686] = 32'b00000000000000001111001100111010;
assign LUT_1[19687] = 32'b00000000000000001000011110110110;
assign LUT_1[19688] = 32'b00000000000000001010110011000111;
assign LUT_1[19689] = 32'b00000000000000000100000101000011;
assign LUT_1[19690] = 32'b00000000000000000110100001011000;
assign LUT_1[19691] = 32'b11111111111111111111110011010100;
assign LUT_1[19692] = 32'b00000000000000010010101100011110;
assign LUT_1[19693] = 32'b00000000000000001011111110011010;
assign LUT_1[19694] = 32'b00000000000000001110011010101111;
assign LUT_1[19695] = 32'b00000000000000000111101100101011;
assign LUT_1[19696] = 32'b00000000000000001101100000110100;
assign LUT_1[19697] = 32'b00000000000000000110110010110000;
assign LUT_1[19698] = 32'b00000000000000001001001111000101;
assign LUT_1[19699] = 32'b00000000000000000010100001000001;
assign LUT_1[19700] = 32'b00000000000000010101011010001011;
assign LUT_1[19701] = 32'b00000000000000001110101100000111;
assign LUT_1[19702] = 32'b00000000000000010001001000011100;
assign LUT_1[19703] = 32'b00000000000000001010011010011000;
assign LUT_1[19704] = 32'b00000000000000001100101110101001;
assign LUT_1[19705] = 32'b00000000000000000110000000100101;
assign LUT_1[19706] = 32'b00000000000000001000011100111010;
assign LUT_1[19707] = 32'b00000000000000000001101110110110;
assign LUT_1[19708] = 32'b00000000000000010100101000000000;
assign LUT_1[19709] = 32'b00000000000000001101111001111100;
assign LUT_1[19710] = 32'b00000000000000010000010110010001;
assign LUT_1[19711] = 32'b00000000000000001001101000001101;
assign LUT_1[19712] = 32'b00000000000000000011100000110100;
assign LUT_1[19713] = 32'b11111111111111111100110010110000;
assign LUT_1[19714] = 32'b11111111111111111111001111000101;
assign LUT_1[19715] = 32'b11111111111111111000100001000001;
assign LUT_1[19716] = 32'b00000000000000001011011010001011;
assign LUT_1[19717] = 32'b00000000000000000100101100000111;
assign LUT_1[19718] = 32'b00000000000000000111001000011100;
assign LUT_1[19719] = 32'b00000000000000000000011010011000;
assign LUT_1[19720] = 32'b00000000000000000010101110101001;
assign LUT_1[19721] = 32'b11111111111111111100000000100101;
assign LUT_1[19722] = 32'b11111111111111111110011100111010;
assign LUT_1[19723] = 32'b11111111111111110111101110110110;
assign LUT_1[19724] = 32'b00000000000000001010101000000000;
assign LUT_1[19725] = 32'b00000000000000000011111001111100;
assign LUT_1[19726] = 32'b00000000000000000110010110010001;
assign LUT_1[19727] = 32'b11111111111111111111101000001101;
assign LUT_1[19728] = 32'b00000000000000000101011100010110;
assign LUT_1[19729] = 32'b11111111111111111110101110010010;
assign LUT_1[19730] = 32'b00000000000000000001001010100111;
assign LUT_1[19731] = 32'b11111111111111111010011100100011;
assign LUT_1[19732] = 32'b00000000000000001101010101101101;
assign LUT_1[19733] = 32'b00000000000000000110100111101001;
assign LUT_1[19734] = 32'b00000000000000001001000011111110;
assign LUT_1[19735] = 32'b00000000000000000010010101111010;
assign LUT_1[19736] = 32'b00000000000000000100101010001011;
assign LUT_1[19737] = 32'b11111111111111111101111100000111;
assign LUT_1[19738] = 32'b00000000000000000000011000011100;
assign LUT_1[19739] = 32'b11111111111111111001101010011000;
assign LUT_1[19740] = 32'b00000000000000001100100011100010;
assign LUT_1[19741] = 32'b00000000000000000101110101011110;
assign LUT_1[19742] = 32'b00000000000000001000010001110011;
assign LUT_1[19743] = 32'b00000000000000000001100011101111;
assign LUT_1[19744] = 32'b00000000000000000100011011110011;
assign LUT_1[19745] = 32'b11111111111111111101101101101111;
assign LUT_1[19746] = 32'b00000000000000000000001010000100;
assign LUT_1[19747] = 32'b11111111111111111001011100000000;
assign LUT_1[19748] = 32'b00000000000000001100010101001010;
assign LUT_1[19749] = 32'b00000000000000000101100111000110;
assign LUT_1[19750] = 32'b00000000000000001000000011011011;
assign LUT_1[19751] = 32'b00000000000000000001010101010111;
assign LUT_1[19752] = 32'b00000000000000000011101001101000;
assign LUT_1[19753] = 32'b11111111111111111100111011100100;
assign LUT_1[19754] = 32'b11111111111111111111010111111001;
assign LUT_1[19755] = 32'b11111111111111111000101001110101;
assign LUT_1[19756] = 32'b00000000000000001011100010111111;
assign LUT_1[19757] = 32'b00000000000000000100110100111011;
assign LUT_1[19758] = 32'b00000000000000000111010001010000;
assign LUT_1[19759] = 32'b00000000000000000000100011001100;
assign LUT_1[19760] = 32'b00000000000000000110010111010101;
assign LUT_1[19761] = 32'b11111111111111111111101001010001;
assign LUT_1[19762] = 32'b00000000000000000010000101100110;
assign LUT_1[19763] = 32'b11111111111111111011010111100010;
assign LUT_1[19764] = 32'b00000000000000001110010000101100;
assign LUT_1[19765] = 32'b00000000000000000111100010101000;
assign LUT_1[19766] = 32'b00000000000000001001111110111101;
assign LUT_1[19767] = 32'b00000000000000000011010000111001;
assign LUT_1[19768] = 32'b00000000000000000101100101001010;
assign LUT_1[19769] = 32'b11111111111111111110110111000110;
assign LUT_1[19770] = 32'b00000000000000000001010011011011;
assign LUT_1[19771] = 32'b11111111111111111010100101010111;
assign LUT_1[19772] = 32'b00000000000000001101011110100001;
assign LUT_1[19773] = 32'b00000000000000000110110000011101;
assign LUT_1[19774] = 32'b00000000000000001001001100110010;
assign LUT_1[19775] = 32'b00000000000000000010011110101110;
assign LUT_1[19776] = 32'b00000000000000000101011110011100;
assign LUT_1[19777] = 32'b11111111111111111110110000011000;
assign LUT_1[19778] = 32'b00000000000000000001001100101101;
assign LUT_1[19779] = 32'b11111111111111111010011110101001;
assign LUT_1[19780] = 32'b00000000000000001101010111110011;
assign LUT_1[19781] = 32'b00000000000000000110101001101111;
assign LUT_1[19782] = 32'b00000000000000001001000110000100;
assign LUT_1[19783] = 32'b00000000000000000010011000000000;
assign LUT_1[19784] = 32'b00000000000000000100101100010001;
assign LUT_1[19785] = 32'b11111111111111111101111110001101;
assign LUT_1[19786] = 32'b00000000000000000000011010100010;
assign LUT_1[19787] = 32'b11111111111111111001101100011110;
assign LUT_1[19788] = 32'b00000000000000001100100101101000;
assign LUT_1[19789] = 32'b00000000000000000101110111100100;
assign LUT_1[19790] = 32'b00000000000000001000010011111001;
assign LUT_1[19791] = 32'b00000000000000000001100101110101;
assign LUT_1[19792] = 32'b00000000000000000111011001111110;
assign LUT_1[19793] = 32'b00000000000000000000101011111010;
assign LUT_1[19794] = 32'b00000000000000000011001000001111;
assign LUT_1[19795] = 32'b11111111111111111100011010001011;
assign LUT_1[19796] = 32'b00000000000000001111010011010101;
assign LUT_1[19797] = 32'b00000000000000001000100101010001;
assign LUT_1[19798] = 32'b00000000000000001011000001100110;
assign LUT_1[19799] = 32'b00000000000000000100010011100010;
assign LUT_1[19800] = 32'b00000000000000000110100111110011;
assign LUT_1[19801] = 32'b11111111111111111111111001101111;
assign LUT_1[19802] = 32'b00000000000000000010010110000100;
assign LUT_1[19803] = 32'b11111111111111111011101000000000;
assign LUT_1[19804] = 32'b00000000000000001110100001001010;
assign LUT_1[19805] = 32'b00000000000000000111110011000110;
assign LUT_1[19806] = 32'b00000000000000001010001111011011;
assign LUT_1[19807] = 32'b00000000000000000011100001010111;
assign LUT_1[19808] = 32'b00000000000000000110011001011011;
assign LUT_1[19809] = 32'b11111111111111111111101011010111;
assign LUT_1[19810] = 32'b00000000000000000010000111101100;
assign LUT_1[19811] = 32'b11111111111111111011011001101000;
assign LUT_1[19812] = 32'b00000000000000001110010010110010;
assign LUT_1[19813] = 32'b00000000000000000111100100101110;
assign LUT_1[19814] = 32'b00000000000000001010000001000011;
assign LUT_1[19815] = 32'b00000000000000000011010010111111;
assign LUT_1[19816] = 32'b00000000000000000101100111010000;
assign LUT_1[19817] = 32'b11111111111111111110111001001100;
assign LUT_1[19818] = 32'b00000000000000000001010101100001;
assign LUT_1[19819] = 32'b11111111111111111010100111011101;
assign LUT_1[19820] = 32'b00000000000000001101100000100111;
assign LUT_1[19821] = 32'b00000000000000000110110010100011;
assign LUT_1[19822] = 32'b00000000000000001001001110111000;
assign LUT_1[19823] = 32'b00000000000000000010100000110100;
assign LUT_1[19824] = 32'b00000000000000001000010100111101;
assign LUT_1[19825] = 32'b00000000000000000001100110111001;
assign LUT_1[19826] = 32'b00000000000000000100000011001110;
assign LUT_1[19827] = 32'b11111111111111111101010101001010;
assign LUT_1[19828] = 32'b00000000000000010000001110010100;
assign LUT_1[19829] = 32'b00000000000000001001100000010000;
assign LUT_1[19830] = 32'b00000000000000001011111100100101;
assign LUT_1[19831] = 32'b00000000000000000101001110100001;
assign LUT_1[19832] = 32'b00000000000000000111100010110010;
assign LUT_1[19833] = 32'b00000000000000000000110100101110;
assign LUT_1[19834] = 32'b00000000000000000011010001000011;
assign LUT_1[19835] = 32'b11111111111111111100100010111111;
assign LUT_1[19836] = 32'b00000000000000001111011100001001;
assign LUT_1[19837] = 32'b00000000000000001000101110000101;
assign LUT_1[19838] = 32'b00000000000000001011001010011010;
assign LUT_1[19839] = 32'b00000000000000000100011100010110;
assign LUT_1[19840] = 32'b00000000000000000110100000110111;
assign LUT_1[19841] = 32'b11111111111111111111110010110011;
assign LUT_1[19842] = 32'b00000000000000000010001111001000;
assign LUT_1[19843] = 32'b11111111111111111011100001000100;
assign LUT_1[19844] = 32'b00000000000000001110011010001110;
assign LUT_1[19845] = 32'b00000000000000000111101100001010;
assign LUT_1[19846] = 32'b00000000000000001010001000011111;
assign LUT_1[19847] = 32'b00000000000000000011011010011011;
assign LUT_1[19848] = 32'b00000000000000000101101110101100;
assign LUT_1[19849] = 32'b11111111111111111111000000101000;
assign LUT_1[19850] = 32'b00000000000000000001011100111101;
assign LUT_1[19851] = 32'b11111111111111111010101110111001;
assign LUT_1[19852] = 32'b00000000000000001101101000000011;
assign LUT_1[19853] = 32'b00000000000000000110111001111111;
assign LUT_1[19854] = 32'b00000000000000001001010110010100;
assign LUT_1[19855] = 32'b00000000000000000010101000010000;
assign LUT_1[19856] = 32'b00000000000000001000011100011001;
assign LUT_1[19857] = 32'b00000000000000000001101110010101;
assign LUT_1[19858] = 32'b00000000000000000100001010101010;
assign LUT_1[19859] = 32'b11111111111111111101011100100110;
assign LUT_1[19860] = 32'b00000000000000010000010101110000;
assign LUT_1[19861] = 32'b00000000000000001001100111101100;
assign LUT_1[19862] = 32'b00000000000000001100000100000001;
assign LUT_1[19863] = 32'b00000000000000000101010101111101;
assign LUT_1[19864] = 32'b00000000000000000111101010001110;
assign LUT_1[19865] = 32'b00000000000000000000111100001010;
assign LUT_1[19866] = 32'b00000000000000000011011000011111;
assign LUT_1[19867] = 32'b11111111111111111100101010011011;
assign LUT_1[19868] = 32'b00000000000000001111100011100101;
assign LUT_1[19869] = 32'b00000000000000001000110101100001;
assign LUT_1[19870] = 32'b00000000000000001011010001110110;
assign LUT_1[19871] = 32'b00000000000000000100100011110010;
assign LUT_1[19872] = 32'b00000000000000000111011011110110;
assign LUT_1[19873] = 32'b00000000000000000000101101110010;
assign LUT_1[19874] = 32'b00000000000000000011001010000111;
assign LUT_1[19875] = 32'b11111111111111111100011100000011;
assign LUT_1[19876] = 32'b00000000000000001111010101001101;
assign LUT_1[19877] = 32'b00000000000000001000100111001001;
assign LUT_1[19878] = 32'b00000000000000001011000011011110;
assign LUT_1[19879] = 32'b00000000000000000100010101011010;
assign LUT_1[19880] = 32'b00000000000000000110101001101011;
assign LUT_1[19881] = 32'b11111111111111111111111011100111;
assign LUT_1[19882] = 32'b00000000000000000010010111111100;
assign LUT_1[19883] = 32'b11111111111111111011101001111000;
assign LUT_1[19884] = 32'b00000000000000001110100011000010;
assign LUT_1[19885] = 32'b00000000000000000111110100111110;
assign LUT_1[19886] = 32'b00000000000000001010010001010011;
assign LUT_1[19887] = 32'b00000000000000000011100011001111;
assign LUT_1[19888] = 32'b00000000000000001001010111011000;
assign LUT_1[19889] = 32'b00000000000000000010101001010100;
assign LUT_1[19890] = 32'b00000000000000000101000101101001;
assign LUT_1[19891] = 32'b11111111111111111110010111100101;
assign LUT_1[19892] = 32'b00000000000000010001010000101111;
assign LUT_1[19893] = 32'b00000000000000001010100010101011;
assign LUT_1[19894] = 32'b00000000000000001100111111000000;
assign LUT_1[19895] = 32'b00000000000000000110010000111100;
assign LUT_1[19896] = 32'b00000000000000001000100101001101;
assign LUT_1[19897] = 32'b00000000000000000001110111001001;
assign LUT_1[19898] = 32'b00000000000000000100010011011110;
assign LUT_1[19899] = 32'b11111111111111111101100101011010;
assign LUT_1[19900] = 32'b00000000000000010000011110100100;
assign LUT_1[19901] = 32'b00000000000000001001110000100000;
assign LUT_1[19902] = 32'b00000000000000001100001100110101;
assign LUT_1[19903] = 32'b00000000000000000101011110110001;
assign LUT_1[19904] = 32'b00000000000000001000011110011111;
assign LUT_1[19905] = 32'b00000000000000000001110000011011;
assign LUT_1[19906] = 32'b00000000000000000100001100110000;
assign LUT_1[19907] = 32'b11111111111111111101011110101100;
assign LUT_1[19908] = 32'b00000000000000010000010111110110;
assign LUT_1[19909] = 32'b00000000000000001001101001110010;
assign LUT_1[19910] = 32'b00000000000000001100000110000111;
assign LUT_1[19911] = 32'b00000000000000000101011000000011;
assign LUT_1[19912] = 32'b00000000000000000111101100010100;
assign LUT_1[19913] = 32'b00000000000000000000111110010000;
assign LUT_1[19914] = 32'b00000000000000000011011010100101;
assign LUT_1[19915] = 32'b11111111111111111100101100100001;
assign LUT_1[19916] = 32'b00000000000000001111100101101011;
assign LUT_1[19917] = 32'b00000000000000001000110111100111;
assign LUT_1[19918] = 32'b00000000000000001011010011111100;
assign LUT_1[19919] = 32'b00000000000000000100100101111000;
assign LUT_1[19920] = 32'b00000000000000001010011010000001;
assign LUT_1[19921] = 32'b00000000000000000011101011111101;
assign LUT_1[19922] = 32'b00000000000000000110001000010010;
assign LUT_1[19923] = 32'b11111111111111111111011010001110;
assign LUT_1[19924] = 32'b00000000000000010010010011011000;
assign LUT_1[19925] = 32'b00000000000000001011100101010100;
assign LUT_1[19926] = 32'b00000000000000001110000001101001;
assign LUT_1[19927] = 32'b00000000000000000111010011100101;
assign LUT_1[19928] = 32'b00000000000000001001100111110110;
assign LUT_1[19929] = 32'b00000000000000000010111001110010;
assign LUT_1[19930] = 32'b00000000000000000101010110000111;
assign LUT_1[19931] = 32'b11111111111111111110101000000011;
assign LUT_1[19932] = 32'b00000000000000010001100001001101;
assign LUT_1[19933] = 32'b00000000000000001010110011001001;
assign LUT_1[19934] = 32'b00000000000000001101001111011110;
assign LUT_1[19935] = 32'b00000000000000000110100001011010;
assign LUT_1[19936] = 32'b00000000000000001001011001011110;
assign LUT_1[19937] = 32'b00000000000000000010101011011010;
assign LUT_1[19938] = 32'b00000000000000000101000111101111;
assign LUT_1[19939] = 32'b11111111111111111110011001101011;
assign LUT_1[19940] = 32'b00000000000000010001010010110101;
assign LUT_1[19941] = 32'b00000000000000001010100100110001;
assign LUT_1[19942] = 32'b00000000000000001101000001000110;
assign LUT_1[19943] = 32'b00000000000000000110010011000010;
assign LUT_1[19944] = 32'b00000000000000001000100111010011;
assign LUT_1[19945] = 32'b00000000000000000001111001001111;
assign LUT_1[19946] = 32'b00000000000000000100010101100100;
assign LUT_1[19947] = 32'b11111111111111111101100111100000;
assign LUT_1[19948] = 32'b00000000000000010000100000101010;
assign LUT_1[19949] = 32'b00000000000000001001110010100110;
assign LUT_1[19950] = 32'b00000000000000001100001110111011;
assign LUT_1[19951] = 32'b00000000000000000101100000110111;
assign LUT_1[19952] = 32'b00000000000000001011010101000000;
assign LUT_1[19953] = 32'b00000000000000000100100110111100;
assign LUT_1[19954] = 32'b00000000000000000111000011010001;
assign LUT_1[19955] = 32'b00000000000000000000010101001101;
assign LUT_1[19956] = 32'b00000000000000010011001110010111;
assign LUT_1[19957] = 32'b00000000000000001100100000010011;
assign LUT_1[19958] = 32'b00000000000000001110111100101000;
assign LUT_1[19959] = 32'b00000000000000001000001110100100;
assign LUT_1[19960] = 32'b00000000000000001010100010110101;
assign LUT_1[19961] = 32'b00000000000000000011110100110001;
assign LUT_1[19962] = 32'b00000000000000000110010001000110;
assign LUT_1[19963] = 32'b11111111111111111111100011000010;
assign LUT_1[19964] = 32'b00000000000000010010011100001100;
assign LUT_1[19965] = 32'b00000000000000001011101110001000;
assign LUT_1[19966] = 32'b00000000000000001110001010011101;
assign LUT_1[19967] = 32'b00000000000000000111011100011001;
assign LUT_1[19968] = 32'b11111111111111111111011011000101;
assign LUT_1[19969] = 32'b11111111111111111000101101000001;
assign LUT_1[19970] = 32'b11111111111111111011001001010110;
assign LUT_1[19971] = 32'b11111111111111110100011011010010;
assign LUT_1[19972] = 32'b00000000000000000111010100011100;
assign LUT_1[19973] = 32'b00000000000000000000100110011000;
assign LUT_1[19974] = 32'b00000000000000000011000010101101;
assign LUT_1[19975] = 32'b11111111111111111100010100101001;
assign LUT_1[19976] = 32'b11111111111111111110101000111010;
assign LUT_1[19977] = 32'b11111111111111110111111010110110;
assign LUT_1[19978] = 32'b11111111111111111010010111001011;
assign LUT_1[19979] = 32'b11111111111111110011101001000111;
assign LUT_1[19980] = 32'b00000000000000000110100010010001;
assign LUT_1[19981] = 32'b11111111111111111111110100001101;
assign LUT_1[19982] = 32'b00000000000000000010010000100010;
assign LUT_1[19983] = 32'b11111111111111111011100010011110;
assign LUT_1[19984] = 32'b00000000000000000001010110100111;
assign LUT_1[19985] = 32'b11111111111111111010101000100011;
assign LUT_1[19986] = 32'b11111111111111111101000100111000;
assign LUT_1[19987] = 32'b11111111111111110110010110110100;
assign LUT_1[19988] = 32'b00000000000000001001001111111110;
assign LUT_1[19989] = 32'b00000000000000000010100001111010;
assign LUT_1[19990] = 32'b00000000000000000100111110001111;
assign LUT_1[19991] = 32'b11111111111111111110010000001011;
assign LUT_1[19992] = 32'b00000000000000000000100100011100;
assign LUT_1[19993] = 32'b11111111111111111001110110011000;
assign LUT_1[19994] = 32'b11111111111111111100010010101101;
assign LUT_1[19995] = 32'b11111111111111110101100100101001;
assign LUT_1[19996] = 32'b00000000000000001000011101110011;
assign LUT_1[19997] = 32'b00000000000000000001101111101111;
assign LUT_1[19998] = 32'b00000000000000000100001100000100;
assign LUT_1[19999] = 32'b11111111111111111101011110000000;
assign LUT_1[20000] = 32'b00000000000000000000010110000100;
assign LUT_1[20001] = 32'b11111111111111111001101000000000;
assign LUT_1[20002] = 32'b11111111111111111100000100010101;
assign LUT_1[20003] = 32'b11111111111111110101010110010001;
assign LUT_1[20004] = 32'b00000000000000001000001111011011;
assign LUT_1[20005] = 32'b00000000000000000001100001010111;
assign LUT_1[20006] = 32'b00000000000000000011111101101100;
assign LUT_1[20007] = 32'b11111111111111111101001111101000;
assign LUT_1[20008] = 32'b11111111111111111111100011111001;
assign LUT_1[20009] = 32'b11111111111111111000110101110101;
assign LUT_1[20010] = 32'b11111111111111111011010010001010;
assign LUT_1[20011] = 32'b11111111111111110100100100000110;
assign LUT_1[20012] = 32'b00000000000000000111011101010000;
assign LUT_1[20013] = 32'b00000000000000000000101111001100;
assign LUT_1[20014] = 32'b00000000000000000011001011100001;
assign LUT_1[20015] = 32'b11111111111111111100011101011101;
assign LUT_1[20016] = 32'b00000000000000000010010001100110;
assign LUT_1[20017] = 32'b11111111111111111011100011100010;
assign LUT_1[20018] = 32'b11111111111111111101111111110111;
assign LUT_1[20019] = 32'b11111111111111110111010001110011;
assign LUT_1[20020] = 32'b00000000000000001010001010111101;
assign LUT_1[20021] = 32'b00000000000000000011011100111001;
assign LUT_1[20022] = 32'b00000000000000000101111001001110;
assign LUT_1[20023] = 32'b11111111111111111111001011001010;
assign LUT_1[20024] = 32'b00000000000000000001011111011011;
assign LUT_1[20025] = 32'b11111111111111111010110001010111;
assign LUT_1[20026] = 32'b11111111111111111101001101101100;
assign LUT_1[20027] = 32'b11111111111111110110011111101000;
assign LUT_1[20028] = 32'b00000000000000001001011000110010;
assign LUT_1[20029] = 32'b00000000000000000010101010101110;
assign LUT_1[20030] = 32'b00000000000000000101000111000011;
assign LUT_1[20031] = 32'b11111111111111111110011000111111;
assign LUT_1[20032] = 32'b00000000000000000001011000101101;
assign LUT_1[20033] = 32'b11111111111111111010101010101001;
assign LUT_1[20034] = 32'b11111111111111111101000110111110;
assign LUT_1[20035] = 32'b11111111111111110110011000111010;
assign LUT_1[20036] = 32'b00000000000000001001010010000100;
assign LUT_1[20037] = 32'b00000000000000000010100100000000;
assign LUT_1[20038] = 32'b00000000000000000101000000010101;
assign LUT_1[20039] = 32'b11111111111111111110010010010001;
assign LUT_1[20040] = 32'b00000000000000000000100110100010;
assign LUT_1[20041] = 32'b11111111111111111001111000011110;
assign LUT_1[20042] = 32'b11111111111111111100010100110011;
assign LUT_1[20043] = 32'b11111111111111110101100110101111;
assign LUT_1[20044] = 32'b00000000000000001000011111111001;
assign LUT_1[20045] = 32'b00000000000000000001110001110101;
assign LUT_1[20046] = 32'b00000000000000000100001110001010;
assign LUT_1[20047] = 32'b11111111111111111101100000000110;
assign LUT_1[20048] = 32'b00000000000000000011010100001111;
assign LUT_1[20049] = 32'b11111111111111111100100110001011;
assign LUT_1[20050] = 32'b11111111111111111111000010100000;
assign LUT_1[20051] = 32'b11111111111111111000010100011100;
assign LUT_1[20052] = 32'b00000000000000001011001101100110;
assign LUT_1[20053] = 32'b00000000000000000100011111100010;
assign LUT_1[20054] = 32'b00000000000000000110111011110111;
assign LUT_1[20055] = 32'b00000000000000000000001101110011;
assign LUT_1[20056] = 32'b00000000000000000010100010000100;
assign LUT_1[20057] = 32'b11111111111111111011110100000000;
assign LUT_1[20058] = 32'b11111111111111111110010000010101;
assign LUT_1[20059] = 32'b11111111111111110111100010010001;
assign LUT_1[20060] = 32'b00000000000000001010011011011011;
assign LUT_1[20061] = 32'b00000000000000000011101101010111;
assign LUT_1[20062] = 32'b00000000000000000110001001101100;
assign LUT_1[20063] = 32'b11111111111111111111011011101000;
assign LUT_1[20064] = 32'b00000000000000000010010011101100;
assign LUT_1[20065] = 32'b11111111111111111011100101101000;
assign LUT_1[20066] = 32'b11111111111111111110000001111101;
assign LUT_1[20067] = 32'b11111111111111110111010011111001;
assign LUT_1[20068] = 32'b00000000000000001010001101000011;
assign LUT_1[20069] = 32'b00000000000000000011011110111111;
assign LUT_1[20070] = 32'b00000000000000000101111011010100;
assign LUT_1[20071] = 32'b11111111111111111111001101010000;
assign LUT_1[20072] = 32'b00000000000000000001100001100001;
assign LUT_1[20073] = 32'b11111111111111111010110011011101;
assign LUT_1[20074] = 32'b11111111111111111101001111110010;
assign LUT_1[20075] = 32'b11111111111111110110100001101110;
assign LUT_1[20076] = 32'b00000000000000001001011010111000;
assign LUT_1[20077] = 32'b00000000000000000010101100110100;
assign LUT_1[20078] = 32'b00000000000000000101001001001001;
assign LUT_1[20079] = 32'b11111111111111111110011011000101;
assign LUT_1[20080] = 32'b00000000000000000100001111001110;
assign LUT_1[20081] = 32'b11111111111111111101100001001010;
assign LUT_1[20082] = 32'b11111111111111111111111101011111;
assign LUT_1[20083] = 32'b11111111111111111001001111011011;
assign LUT_1[20084] = 32'b00000000000000001100001000100101;
assign LUT_1[20085] = 32'b00000000000000000101011010100001;
assign LUT_1[20086] = 32'b00000000000000000111110110110110;
assign LUT_1[20087] = 32'b00000000000000000001001000110010;
assign LUT_1[20088] = 32'b00000000000000000011011101000011;
assign LUT_1[20089] = 32'b11111111111111111100101110111111;
assign LUT_1[20090] = 32'b11111111111111111111001011010100;
assign LUT_1[20091] = 32'b11111111111111111000011101010000;
assign LUT_1[20092] = 32'b00000000000000001011010110011010;
assign LUT_1[20093] = 32'b00000000000000000100101000010110;
assign LUT_1[20094] = 32'b00000000000000000111000100101011;
assign LUT_1[20095] = 32'b00000000000000000000010110100111;
assign LUT_1[20096] = 32'b00000000000000000010011011001000;
assign LUT_1[20097] = 32'b11111111111111111011101101000100;
assign LUT_1[20098] = 32'b11111111111111111110001001011001;
assign LUT_1[20099] = 32'b11111111111111110111011011010101;
assign LUT_1[20100] = 32'b00000000000000001010010100011111;
assign LUT_1[20101] = 32'b00000000000000000011100110011011;
assign LUT_1[20102] = 32'b00000000000000000110000010110000;
assign LUT_1[20103] = 32'b11111111111111111111010100101100;
assign LUT_1[20104] = 32'b00000000000000000001101000111101;
assign LUT_1[20105] = 32'b11111111111111111010111010111001;
assign LUT_1[20106] = 32'b11111111111111111101010111001110;
assign LUT_1[20107] = 32'b11111111111111110110101001001010;
assign LUT_1[20108] = 32'b00000000000000001001100010010100;
assign LUT_1[20109] = 32'b00000000000000000010110100010000;
assign LUT_1[20110] = 32'b00000000000000000101010000100101;
assign LUT_1[20111] = 32'b11111111111111111110100010100001;
assign LUT_1[20112] = 32'b00000000000000000100010110101010;
assign LUT_1[20113] = 32'b11111111111111111101101000100110;
assign LUT_1[20114] = 32'b00000000000000000000000100111011;
assign LUT_1[20115] = 32'b11111111111111111001010110110111;
assign LUT_1[20116] = 32'b00000000000000001100010000000001;
assign LUT_1[20117] = 32'b00000000000000000101100001111101;
assign LUT_1[20118] = 32'b00000000000000000111111110010010;
assign LUT_1[20119] = 32'b00000000000000000001010000001110;
assign LUT_1[20120] = 32'b00000000000000000011100100011111;
assign LUT_1[20121] = 32'b11111111111111111100110110011011;
assign LUT_1[20122] = 32'b11111111111111111111010010110000;
assign LUT_1[20123] = 32'b11111111111111111000100100101100;
assign LUT_1[20124] = 32'b00000000000000001011011101110110;
assign LUT_1[20125] = 32'b00000000000000000100101111110010;
assign LUT_1[20126] = 32'b00000000000000000111001100000111;
assign LUT_1[20127] = 32'b00000000000000000000011110000011;
assign LUT_1[20128] = 32'b00000000000000000011010110000111;
assign LUT_1[20129] = 32'b11111111111111111100101000000011;
assign LUT_1[20130] = 32'b11111111111111111111000100011000;
assign LUT_1[20131] = 32'b11111111111111111000010110010100;
assign LUT_1[20132] = 32'b00000000000000001011001111011110;
assign LUT_1[20133] = 32'b00000000000000000100100001011010;
assign LUT_1[20134] = 32'b00000000000000000110111101101111;
assign LUT_1[20135] = 32'b00000000000000000000001111101011;
assign LUT_1[20136] = 32'b00000000000000000010100011111100;
assign LUT_1[20137] = 32'b11111111111111111011110101111000;
assign LUT_1[20138] = 32'b11111111111111111110010010001101;
assign LUT_1[20139] = 32'b11111111111111110111100100001001;
assign LUT_1[20140] = 32'b00000000000000001010011101010011;
assign LUT_1[20141] = 32'b00000000000000000011101111001111;
assign LUT_1[20142] = 32'b00000000000000000110001011100100;
assign LUT_1[20143] = 32'b11111111111111111111011101100000;
assign LUT_1[20144] = 32'b00000000000000000101010001101001;
assign LUT_1[20145] = 32'b11111111111111111110100011100101;
assign LUT_1[20146] = 32'b00000000000000000000111111111010;
assign LUT_1[20147] = 32'b11111111111111111010010001110110;
assign LUT_1[20148] = 32'b00000000000000001101001011000000;
assign LUT_1[20149] = 32'b00000000000000000110011100111100;
assign LUT_1[20150] = 32'b00000000000000001000111001010001;
assign LUT_1[20151] = 32'b00000000000000000010001011001101;
assign LUT_1[20152] = 32'b00000000000000000100011111011110;
assign LUT_1[20153] = 32'b11111111111111111101110001011010;
assign LUT_1[20154] = 32'b00000000000000000000001101101111;
assign LUT_1[20155] = 32'b11111111111111111001011111101011;
assign LUT_1[20156] = 32'b00000000000000001100011000110101;
assign LUT_1[20157] = 32'b00000000000000000101101010110001;
assign LUT_1[20158] = 32'b00000000000000001000000111000110;
assign LUT_1[20159] = 32'b00000000000000000001011001000010;
assign LUT_1[20160] = 32'b00000000000000000100011000110000;
assign LUT_1[20161] = 32'b11111111111111111101101010101100;
assign LUT_1[20162] = 32'b00000000000000000000000111000001;
assign LUT_1[20163] = 32'b11111111111111111001011000111101;
assign LUT_1[20164] = 32'b00000000000000001100010010000111;
assign LUT_1[20165] = 32'b00000000000000000101100100000011;
assign LUT_1[20166] = 32'b00000000000000001000000000011000;
assign LUT_1[20167] = 32'b00000000000000000001010010010100;
assign LUT_1[20168] = 32'b00000000000000000011100110100101;
assign LUT_1[20169] = 32'b11111111111111111100111000100001;
assign LUT_1[20170] = 32'b11111111111111111111010100110110;
assign LUT_1[20171] = 32'b11111111111111111000100110110010;
assign LUT_1[20172] = 32'b00000000000000001011011111111100;
assign LUT_1[20173] = 32'b00000000000000000100110001111000;
assign LUT_1[20174] = 32'b00000000000000000111001110001101;
assign LUT_1[20175] = 32'b00000000000000000000100000001001;
assign LUT_1[20176] = 32'b00000000000000000110010100010010;
assign LUT_1[20177] = 32'b11111111111111111111100110001110;
assign LUT_1[20178] = 32'b00000000000000000010000010100011;
assign LUT_1[20179] = 32'b11111111111111111011010100011111;
assign LUT_1[20180] = 32'b00000000000000001110001101101001;
assign LUT_1[20181] = 32'b00000000000000000111011111100101;
assign LUT_1[20182] = 32'b00000000000000001001111011111010;
assign LUT_1[20183] = 32'b00000000000000000011001101110110;
assign LUT_1[20184] = 32'b00000000000000000101100010000111;
assign LUT_1[20185] = 32'b11111111111111111110110100000011;
assign LUT_1[20186] = 32'b00000000000000000001010000011000;
assign LUT_1[20187] = 32'b11111111111111111010100010010100;
assign LUT_1[20188] = 32'b00000000000000001101011011011110;
assign LUT_1[20189] = 32'b00000000000000000110101101011010;
assign LUT_1[20190] = 32'b00000000000000001001001001101111;
assign LUT_1[20191] = 32'b00000000000000000010011011101011;
assign LUT_1[20192] = 32'b00000000000000000101010011101111;
assign LUT_1[20193] = 32'b11111111111111111110100101101011;
assign LUT_1[20194] = 32'b00000000000000000001000010000000;
assign LUT_1[20195] = 32'b11111111111111111010010011111100;
assign LUT_1[20196] = 32'b00000000000000001101001101000110;
assign LUT_1[20197] = 32'b00000000000000000110011111000010;
assign LUT_1[20198] = 32'b00000000000000001000111011010111;
assign LUT_1[20199] = 32'b00000000000000000010001101010011;
assign LUT_1[20200] = 32'b00000000000000000100100001100100;
assign LUT_1[20201] = 32'b11111111111111111101110011100000;
assign LUT_1[20202] = 32'b00000000000000000000001111110101;
assign LUT_1[20203] = 32'b11111111111111111001100001110001;
assign LUT_1[20204] = 32'b00000000000000001100011010111011;
assign LUT_1[20205] = 32'b00000000000000000101101100110111;
assign LUT_1[20206] = 32'b00000000000000001000001001001100;
assign LUT_1[20207] = 32'b00000000000000000001011011001000;
assign LUT_1[20208] = 32'b00000000000000000111001111010001;
assign LUT_1[20209] = 32'b00000000000000000000100001001101;
assign LUT_1[20210] = 32'b00000000000000000010111101100010;
assign LUT_1[20211] = 32'b11111111111111111100001111011110;
assign LUT_1[20212] = 32'b00000000000000001111001000101000;
assign LUT_1[20213] = 32'b00000000000000001000011010100100;
assign LUT_1[20214] = 32'b00000000000000001010110110111001;
assign LUT_1[20215] = 32'b00000000000000000100001000110101;
assign LUT_1[20216] = 32'b00000000000000000110011101000110;
assign LUT_1[20217] = 32'b11111111111111111111101111000010;
assign LUT_1[20218] = 32'b00000000000000000010001011010111;
assign LUT_1[20219] = 32'b11111111111111111011011101010011;
assign LUT_1[20220] = 32'b00000000000000001110010110011101;
assign LUT_1[20221] = 32'b00000000000000000111101000011001;
assign LUT_1[20222] = 32'b00000000000000001010000100101110;
assign LUT_1[20223] = 32'b00000000000000000011010110101010;
assign LUT_1[20224] = 32'b11111111111111111101001111010001;
assign LUT_1[20225] = 32'b11111111111111110110100001001101;
assign LUT_1[20226] = 32'b11111111111111111000111101100010;
assign LUT_1[20227] = 32'b11111111111111110010001111011110;
assign LUT_1[20228] = 32'b00000000000000000101001000101000;
assign LUT_1[20229] = 32'b11111111111111111110011010100100;
assign LUT_1[20230] = 32'b00000000000000000000110110111001;
assign LUT_1[20231] = 32'b11111111111111111010001000110101;
assign LUT_1[20232] = 32'b11111111111111111100011101000110;
assign LUT_1[20233] = 32'b11111111111111110101101111000010;
assign LUT_1[20234] = 32'b11111111111111111000001011010111;
assign LUT_1[20235] = 32'b11111111111111110001011101010011;
assign LUT_1[20236] = 32'b00000000000000000100010110011101;
assign LUT_1[20237] = 32'b11111111111111111101101000011001;
assign LUT_1[20238] = 32'b00000000000000000000000100101110;
assign LUT_1[20239] = 32'b11111111111111111001010110101010;
assign LUT_1[20240] = 32'b11111111111111111111001010110011;
assign LUT_1[20241] = 32'b11111111111111111000011100101111;
assign LUT_1[20242] = 32'b11111111111111111010111001000100;
assign LUT_1[20243] = 32'b11111111111111110100001011000000;
assign LUT_1[20244] = 32'b00000000000000000111000100001010;
assign LUT_1[20245] = 32'b00000000000000000000010110000110;
assign LUT_1[20246] = 32'b00000000000000000010110010011011;
assign LUT_1[20247] = 32'b11111111111111111100000100010111;
assign LUT_1[20248] = 32'b11111111111111111110011000101000;
assign LUT_1[20249] = 32'b11111111111111110111101010100100;
assign LUT_1[20250] = 32'b11111111111111111010000110111001;
assign LUT_1[20251] = 32'b11111111111111110011011000110101;
assign LUT_1[20252] = 32'b00000000000000000110010001111111;
assign LUT_1[20253] = 32'b11111111111111111111100011111011;
assign LUT_1[20254] = 32'b00000000000000000010000000010000;
assign LUT_1[20255] = 32'b11111111111111111011010010001100;
assign LUT_1[20256] = 32'b11111111111111111110001010010000;
assign LUT_1[20257] = 32'b11111111111111110111011100001100;
assign LUT_1[20258] = 32'b11111111111111111001111000100001;
assign LUT_1[20259] = 32'b11111111111111110011001010011101;
assign LUT_1[20260] = 32'b00000000000000000110000011100111;
assign LUT_1[20261] = 32'b11111111111111111111010101100011;
assign LUT_1[20262] = 32'b00000000000000000001110001111000;
assign LUT_1[20263] = 32'b11111111111111111011000011110100;
assign LUT_1[20264] = 32'b11111111111111111101011000000101;
assign LUT_1[20265] = 32'b11111111111111110110101010000001;
assign LUT_1[20266] = 32'b11111111111111111001000110010110;
assign LUT_1[20267] = 32'b11111111111111110010011000010010;
assign LUT_1[20268] = 32'b00000000000000000101010001011100;
assign LUT_1[20269] = 32'b11111111111111111110100011011000;
assign LUT_1[20270] = 32'b00000000000000000000111111101101;
assign LUT_1[20271] = 32'b11111111111111111010010001101001;
assign LUT_1[20272] = 32'b00000000000000000000000101110010;
assign LUT_1[20273] = 32'b11111111111111111001010111101110;
assign LUT_1[20274] = 32'b11111111111111111011110100000011;
assign LUT_1[20275] = 32'b11111111111111110101000101111111;
assign LUT_1[20276] = 32'b00000000000000000111111111001001;
assign LUT_1[20277] = 32'b00000000000000000001010001000101;
assign LUT_1[20278] = 32'b00000000000000000011101101011010;
assign LUT_1[20279] = 32'b11111111111111111100111111010110;
assign LUT_1[20280] = 32'b11111111111111111111010011100111;
assign LUT_1[20281] = 32'b11111111111111111000100101100011;
assign LUT_1[20282] = 32'b11111111111111111011000001111000;
assign LUT_1[20283] = 32'b11111111111111110100010011110100;
assign LUT_1[20284] = 32'b00000000000000000111001100111110;
assign LUT_1[20285] = 32'b00000000000000000000011110111010;
assign LUT_1[20286] = 32'b00000000000000000010111011001111;
assign LUT_1[20287] = 32'b11111111111111111100001101001011;
assign LUT_1[20288] = 32'b11111111111111111111001100111001;
assign LUT_1[20289] = 32'b11111111111111111000011110110101;
assign LUT_1[20290] = 32'b11111111111111111010111011001010;
assign LUT_1[20291] = 32'b11111111111111110100001101000110;
assign LUT_1[20292] = 32'b00000000000000000111000110010000;
assign LUT_1[20293] = 32'b00000000000000000000011000001100;
assign LUT_1[20294] = 32'b00000000000000000010110100100001;
assign LUT_1[20295] = 32'b11111111111111111100000110011101;
assign LUT_1[20296] = 32'b11111111111111111110011010101110;
assign LUT_1[20297] = 32'b11111111111111110111101100101010;
assign LUT_1[20298] = 32'b11111111111111111010001000111111;
assign LUT_1[20299] = 32'b11111111111111110011011010111011;
assign LUT_1[20300] = 32'b00000000000000000110010100000101;
assign LUT_1[20301] = 32'b11111111111111111111100110000001;
assign LUT_1[20302] = 32'b00000000000000000010000010010110;
assign LUT_1[20303] = 32'b11111111111111111011010100010010;
assign LUT_1[20304] = 32'b00000000000000000001001000011011;
assign LUT_1[20305] = 32'b11111111111111111010011010010111;
assign LUT_1[20306] = 32'b11111111111111111100110110101100;
assign LUT_1[20307] = 32'b11111111111111110110001000101000;
assign LUT_1[20308] = 32'b00000000000000001001000001110010;
assign LUT_1[20309] = 32'b00000000000000000010010011101110;
assign LUT_1[20310] = 32'b00000000000000000100110000000011;
assign LUT_1[20311] = 32'b11111111111111111110000001111111;
assign LUT_1[20312] = 32'b00000000000000000000010110010000;
assign LUT_1[20313] = 32'b11111111111111111001101000001100;
assign LUT_1[20314] = 32'b11111111111111111100000100100001;
assign LUT_1[20315] = 32'b11111111111111110101010110011101;
assign LUT_1[20316] = 32'b00000000000000001000001111100111;
assign LUT_1[20317] = 32'b00000000000000000001100001100011;
assign LUT_1[20318] = 32'b00000000000000000011111101111000;
assign LUT_1[20319] = 32'b11111111111111111101001111110100;
assign LUT_1[20320] = 32'b00000000000000000000000111111000;
assign LUT_1[20321] = 32'b11111111111111111001011001110100;
assign LUT_1[20322] = 32'b11111111111111111011110110001001;
assign LUT_1[20323] = 32'b11111111111111110101001000000101;
assign LUT_1[20324] = 32'b00000000000000001000000001001111;
assign LUT_1[20325] = 32'b00000000000000000001010011001011;
assign LUT_1[20326] = 32'b00000000000000000011101111100000;
assign LUT_1[20327] = 32'b11111111111111111101000001011100;
assign LUT_1[20328] = 32'b11111111111111111111010101101101;
assign LUT_1[20329] = 32'b11111111111111111000100111101001;
assign LUT_1[20330] = 32'b11111111111111111011000011111110;
assign LUT_1[20331] = 32'b11111111111111110100010101111010;
assign LUT_1[20332] = 32'b00000000000000000111001111000100;
assign LUT_1[20333] = 32'b00000000000000000000100001000000;
assign LUT_1[20334] = 32'b00000000000000000010111101010101;
assign LUT_1[20335] = 32'b11111111111111111100001111010001;
assign LUT_1[20336] = 32'b00000000000000000010000011011010;
assign LUT_1[20337] = 32'b11111111111111111011010101010110;
assign LUT_1[20338] = 32'b11111111111111111101110001101011;
assign LUT_1[20339] = 32'b11111111111111110111000011100111;
assign LUT_1[20340] = 32'b00000000000000001001111100110001;
assign LUT_1[20341] = 32'b00000000000000000011001110101101;
assign LUT_1[20342] = 32'b00000000000000000101101011000010;
assign LUT_1[20343] = 32'b11111111111111111110111100111110;
assign LUT_1[20344] = 32'b00000000000000000001010001001111;
assign LUT_1[20345] = 32'b11111111111111111010100011001011;
assign LUT_1[20346] = 32'b11111111111111111100111111100000;
assign LUT_1[20347] = 32'b11111111111111110110010001011100;
assign LUT_1[20348] = 32'b00000000000000001001001010100110;
assign LUT_1[20349] = 32'b00000000000000000010011100100010;
assign LUT_1[20350] = 32'b00000000000000000100111000110111;
assign LUT_1[20351] = 32'b11111111111111111110001010110011;
assign LUT_1[20352] = 32'b00000000000000000000001111010100;
assign LUT_1[20353] = 32'b11111111111111111001100001010000;
assign LUT_1[20354] = 32'b11111111111111111011111101100101;
assign LUT_1[20355] = 32'b11111111111111110101001111100001;
assign LUT_1[20356] = 32'b00000000000000001000001000101011;
assign LUT_1[20357] = 32'b00000000000000000001011010100111;
assign LUT_1[20358] = 32'b00000000000000000011110110111100;
assign LUT_1[20359] = 32'b11111111111111111101001000111000;
assign LUT_1[20360] = 32'b11111111111111111111011101001001;
assign LUT_1[20361] = 32'b11111111111111111000101111000101;
assign LUT_1[20362] = 32'b11111111111111111011001011011010;
assign LUT_1[20363] = 32'b11111111111111110100011101010110;
assign LUT_1[20364] = 32'b00000000000000000111010110100000;
assign LUT_1[20365] = 32'b00000000000000000000101000011100;
assign LUT_1[20366] = 32'b00000000000000000011000100110001;
assign LUT_1[20367] = 32'b11111111111111111100010110101101;
assign LUT_1[20368] = 32'b00000000000000000010001010110110;
assign LUT_1[20369] = 32'b11111111111111111011011100110010;
assign LUT_1[20370] = 32'b11111111111111111101111001000111;
assign LUT_1[20371] = 32'b11111111111111110111001011000011;
assign LUT_1[20372] = 32'b00000000000000001010000100001101;
assign LUT_1[20373] = 32'b00000000000000000011010110001001;
assign LUT_1[20374] = 32'b00000000000000000101110010011110;
assign LUT_1[20375] = 32'b11111111111111111111000100011010;
assign LUT_1[20376] = 32'b00000000000000000001011000101011;
assign LUT_1[20377] = 32'b11111111111111111010101010100111;
assign LUT_1[20378] = 32'b11111111111111111101000110111100;
assign LUT_1[20379] = 32'b11111111111111110110011000111000;
assign LUT_1[20380] = 32'b00000000000000001001010010000010;
assign LUT_1[20381] = 32'b00000000000000000010100011111110;
assign LUT_1[20382] = 32'b00000000000000000101000000010011;
assign LUT_1[20383] = 32'b11111111111111111110010010001111;
assign LUT_1[20384] = 32'b00000000000000000001001010010011;
assign LUT_1[20385] = 32'b11111111111111111010011100001111;
assign LUT_1[20386] = 32'b11111111111111111100111000100100;
assign LUT_1[20387] = 32'b11111111111111110110001010100000;
assign LUT_1[20388] = 32'b00000000000000001001000011101010;
assign LUT_1[20389] = 32'b00000000000000000010010101100110;
assign LUT_1[20390] = 32'b00000000000000000100110001111011;
assign LUT_1[20391] = 32'b11111111111111111110000011110111;
assign LUT_1[20392] = 32'b00000000000000000000011000001000;
assign LUT_1[20393] = 32'b11111111111111111001101010000100;
assign LUT_1[20394] = 32'b11111111111111111100000110011001;
assign LUT_1[20395] = 32'b11111111111111110101011000010101;
assign LUT_1[20396] = 32'b00000000000000001000010001011111;
assign LUT_1[20397] = 32'b00000000000000000001100011011011;
assign LUT_1[20398] = 32'b00000000000000000011111111110000;
assign LUT_1[20399] = 32'b11111111111111111101010001101100;
assign LUT_1[20400] = 32'b00000000000000000011000101110101;
assign LUT_1[20401] = 32'b11111111111111111100010111110001;
assign LUT_1[20402] = 32'b11111111111111111110110100000110;
assign LUT_1[20403] = 32'b11111111111111111000000110000010;
assign LUT_1[20404] = 32'b00000000000000001010111111001100;
assign LUT_1[20405] = 32'b00000000000000000100010001001000;
assign LUT_1[20406] = 32'b00000000000000000110101101011101;
assign LUT_1[20407] = 32'b11111111111111111111111111011001;
assign LUT_1[20408] = 32'b00000000000000000010010011101010;
assign LUT_1[20409] = 32'b11111111111111111011100101100110;
assign LUT_1[20410] = 32'b11111111111111111110000001111011;
assign LUT_1[20411] = 32'b11111111111111110111010011110111;
assign LUT_1[20412] = 32'b00000000000000001010001101000001;
assign LUT_1[20413] = 32'b00000000000000000011011110111101;
assign LUT_1[20414] = 32'b00000000000000000101111011010010;
assign LUT_1[20415] = 32'b11111111111111111111001101001110;
assign LUT_1[20416] = 32'b00000000000000000010001100111100;
assign LUT_1[20417] = 32'b11111111111111111011011110111000;
assign LUT_1[20418] = 32'b11111111111111111101111011001101;
assign LUT_1[20419] = 32'b11111111111111110111001101001001;
assign LUT_1[20420] = 32'b00000000000000001010000110010011;
assign LUT_1[20421] = 32'b00000000000000000011011000001111;
assign LUT_1[20422] = 32'b00000000000000000101110100100100;
assign LUT_1[20423] = 32'b11111111111111111111000110100000;
assign LUT_1[20424] = 32'b00000000000000000001011010110001;
assign LUT_1[20425] = 32'b11111111111111111010101100101101;
assign LUT_1[20426] = 32'b11111111111111111101001001000010;
assign LUT_1[20427] = 32'b11111111111111110110011010111110;
assign LUT_1[20428] = 32'b00000000000000001001010100001000;
assign LUT_1[20429] = 32'b00000000000000000010100110000100;
assign LUT_1[20430] = 32'b00000000000000000101000010011001;
assign LUT_1[20431] = 32'b11111111111111111110010100010101;
assign LUT_1[20432] = 32'b00000000000000000100001000011110;
assign LUT_1[20433] = 32'b11111111111111111101011010011010;
assign LUT_1[20434] = 32'b11111111111111111111110110101111;
assign LUT_1[20435] = 32'b11111111111111111001001000101011;
assign LUT_1[20436] = 32'b00000000000000001100000001110101;
assign LUT_1[20437] = 32'b00000000000000000101010011110001;
assign LUT_1[20438] = 32'b00000000000000000111110000000110;
assign LUT_1[20439] = 32'b00000000000000000001000010000010;
assign LUT_1[20440] = 32'b00000000000000000011010110010011;
assign LUT_1[20441] = 32'b11111111111111111100101000001111;
assign LUT_1[20442] = 32'b11111111111111111111000100100100;
assign LUT_1[20443] = 32'b11111111111111111000010110100000;
assign LUT_1[20444] = 32'b00000000000000001011001111101010;
assign LUT_1[20445] = 32'b00000000000000000100100001100110;
assign LUT_1[20446] = 32'b00000000000000000110111101111011;
assign LUT_1[20447] = 32'b00000000000000000000001111110111;
assign LUT_1[20448] = 32'b00000000000000000011000111111011;
assign LUT_1[20449] = 32'b11111111111111111100011001110111;
assign LUT_1[20450] = 32'b11111111111111111110110110001100;
assign LUT_1[20451] = 32'b11111111111111111000001000001000;
assign LUT_1[20452] = 32'b00000000000000001011000001010010;
assign LUT_1[20453] = 32'b00000000000000000100010011001110;
assign LUT_1[20454] = 32'b00000000000000000110101111100011;
assign LUT_1[20455] = 32'b00000000000000000000000001011111;
assign LUT_1[20456] = 32'b00000000000000000010010101110000;
assign LUT_1[20457] = 32'b11111111111111111011100111101100;
assign LUT_1[20458] = 32'b11111111111111111110000100000001;
assign LUT_1[20459] = 32'b11111111111111110111010101111101;
assign LUT_1[20460] = 32'b00000000000000001010001111000111;
assign LUT_1[20461] = 32'b00000000000000000011100001000011;
assign LUT_1[20462] = 32'b00000000000000000101111101011000;
assign LUT_1[20463] = 32'b11111111111111111111001111010100;
assign LUT_1[20464] = 32'b00000000000000000101000011011101;
assign LUT_1[20465] = 32'b11111111111111111110010101011001;
assign LUT_1[20466] = 32'b00000000000000000000110001101110;
assign LUT_1[20467] = 32'b11111111111111111010000011101010;
assign LUT_1[20468] = 32'b00000000000000001100111100110100;
assign LUT_1[20469] = 32'b00000000000000000110001110110000;
assign LUT_1[20470] = 32'b00000000000000001000101011000101;
assign LUT_1[20471] = 32'b00000000000000000001111101000001;
assign LUT_1[20472] = 32'b00000000000000000100010001010010;
assign LUT_1[20473] = 32'b11111111111111111101100011001110;
assign LUT_1[20474] = 32'b11111111111111111111111111100011;
assign LUT_1[20475] = 32'b11111111111111111001010001011111;
assign LUT_1[20476] = 32'b00000000000000001100001010101001;
assign LUT_1[20477] = 32'b00000000000000000101011100100101;
assign LUT_1[20478] = 32'b00000000000000000111111000111010;
assign LUT_1[20479] = 32'b00000000000000000001001010110110;
assign LUT_1[20480] = 32'b11111111111111111110001001000011;
assign LUT_1[20481] = 32'b11111111111111110111011010111111;
assign LUT_1[20482] = 32'b11111111111111111001110111010100;
assign LUT_1[20483] = 32'b11111111111111110011001001010000;
assign LUT_1[20484] = 32'b00000000000000000110000010011010;
assign LUT_1[20485] = 32'b11111111111111111111010100010110;
assign LUT_1[20486] = 32'b00000000000000000001110000101011;
assign LUT_1[20487] = 32'b11111111111111111011000010100111;
assign LUT_1[20488] = 32'b11111111111111111101010110111000;
assign LUT_1[20489] = 32'b11111111111111110110101000110100;
assign LUT_1[20490] = 32'b11111111111111111001000101001001;
assign LUT_1[20491] = 32'b11111111111111110010010111000101;
assign LUT_1[20492] = 32'b00000000000000000101010000001111;
assign LUT_1[20493] = 32'b11111111111111111110100010001011;
assign LUT_1[20494] = 32'b00000000000000000000111110100000;
assign LUT_1[20495] = 32'b11111111111111111010010000011100;
assign LUT_1[20496] = 32'b00000000000000000000000100100101;
assign LUT_1[20497] = 32'b11111111111111111001010110100001;
assign LUT_1[20498] = 32'b11111111111111111011110010110110;
assign LUT_1[20499] = 32'b11111111111111110101000100110010;
assign LUT_1[20500] = 32'b00000000000000000111111101111100;
assign LUT_1[20501] = 32'b00000000000000000001001111111000;
assign LUT_1[20502] = 32'b00000000000000000011101100001101;
assign LUT_1[20503] = 32'b11111111111111111100111110001001;
assign LUT_1[20504] = 32'b11111111111111111111010010011010;
assign LUT_1[20505] = 32'b11111111111111111000100100010110;
assign LUT_1[20506] = 32'b11111111111111111011000000101011;
assign LUT_1[20507] = 32'b11111111111111110100010010100111;
assign LUT_1[20508] = 32'b00000000000000000111001011110001;
assign LUT_1[20509] = 32'b00000000000000000000011101101101;
assign LUT_1[20510] = 32'b00000000000000000010111010000010;
assign LUT_1[20511] = 32'b11111111111111111100001011111110;
assign LUT_1[20512] = 32'b11111111111111111111000100000010;
assign LUT_1[20513] = 32'b11111111111111111000010101111110;
assign LUT_1[20514] = 32'b11111111111111111010110010010011;
assign LUT_1[20515] = 32'b11111111111111110100000100001111;
assign LUT_1[20516] = 32'b00000000000000000110111101011001;
assign LUT_1[20517] = 32'b00000000000000000000001111010101;
assign LUT_1[20518] = 32'b00000000000000000010101011101010;
assign LUT_1[20519] = 32'b11111111111111111011111101100110;
assign LUT_1[20520] = 32'b11111111111111111110010001110111;
assign LUT_1[20521] = 32'b11111111111111110111100011110011;
assign LUT_1[20522] = 32'b11111111111111111010000000001000;
assign LUT_1[20523] = 32'b11111111111111110011010010000100;
assign LUT_1[20524] = 32'b00000000000000000110001011001110;
assign LUT_1[20525] = 32'b11111111111111111111011101001010;
assign LUT_1[20526] = 32'b00000000000000000001111001011111;
assign LUT_1[20527] = 32'b11111111111111111011001011011011;
assign LUT_1[20528] = 32'b00000000000000000000111111100100;
assign LUT_1[20529] = 32'b11111111111111111010010001100000;
assign LUT_1[20530] = 32'b11111111111111111100101101110101;
assign LUT_1[20531] = 32'b11111111111111110101111111110001;
assign LUT_1[20532] = 32'b00000000000000001000111000111011;
assign LUT_1[20533] = 32'b00000000000000000010001010110111;
assign LUT_1[20534] = 32'b00000000000000000100100111001100;
assign LUT_1[20535] = 32'b11111111111111111101111001001000;
assign LUT_1[20536] = 32'b00000000000000000000001101011001;
assign LUT_1[20537] = 32'b11111111111111111001011111010101;
assign LUT_1[20538] = 32'b11111111111111111011111011101010;
assign LUT_1[20539] = 32'b11111111111111110101001101100110;
assign LUT_1[20540] = 32'b00000000000000001000000110110000;
assign LUT_1[20541] = 32'b00000000000000000001011000101100;
assign LUT_1[20542] = 32'b00000000000000000011110101000001;
assign LUT_1[20543] = 32'b11111111111111111101000110111101;
assign LUT_1[20544] = 32'b00000000000000000000000110101011;
assign LUT_1[20545] = 32'b11111111111111111001011000100111;
assign LUT_1[20546] = 32'b11111111111111111011110100111100;
assign LUT_1[20547] = 32'b11111111111111110101000110111000;
assign LUT_1[20548] = 32'b00000000000000001000000000000010;
assign LUT_1[20549] = 32'b00000000000000000001010001111110;
assign LUT_1[20550] = 32'b00000000000000000011101110010011;
assign LUT_1[20551] = 32'b11111111111111111101000000001111;
assign LUT_1[20552] = 32'b11111111111111111111010100100000;
assign LUT_1[20553] = 32'b11111111111111111000100110011100;
assign LUT_1[20554] = 32'b11111111111111111011000010110001;
assign LUT_1[20555] = 32'b11111111111111110100010100101101;
assign LUT_1[20556] = 32'b00000000000000000111001101110111;
assign LUT_1[20557] = 32'b00000000000000000000011111110011;
assign LUT_1[20558] = 32'b00000000000000000010111100001000;
assign LUT_1[20559] = 32'b11111111111111111100001110000100;
assign LUT_1[20560] = 32'b00000000000000000010000010001101;
assign LUT_1[20561] = 32'b11111111111111111011010100001001;
assign LUT_1[20562] = 32'b11111111111111111101110000011110;
assign LUT_1[20563] = 32'b11111111111111110111000010011010;
assign LUT_1[20564] = 32'b00000000000000001001111011100100;
assign LUT_1[20565] = 32'b00000000000000000011001101100000;
assign LUT_1[20566] = 32'b00000000000000000101101001110101;
assign LUT_1[20567] = 32'b11111111111111111110111011110001;
assign LUT_1[20568] = 32'b00000000000000000001010000000010;
assign LUT_1[20569] = 32'b11111111111111111010100001111110;
assign LUT_1[20570] = 32'b11111111111111111100111110010011;
assign LUT_1[20571] = 32'b11111111111111110110010000001111;
assign LUT_1[20572] = 32'b00000000000000001001001001011001;
assign LUT_1[20573] = 32'b00000000000000000010011011010101;
assign LUT_1[20574] = 32'b00000000000000000100110111101010;
assign LUT_1[20575] = 32'b11111111111111111110001001100110;
assign LUT_1[20576] = 32'b00000000000000000001000001101010;
assign LUT_1[20577] = 32'b11111111111111111010010011100110;
assign LUT_1[20578] = 32'b11111111111111111100101111111011;
assign LUT_1[20579] = 32'b11111111111111110110000001110111;
assign LUT_1[20580] = 32'b00000000000000001000111011000001;
assign LUT_1[20581] = 32'b00000000000000000010001100111101;
assign LUT_1[20582] = 32'b00000000000000000100101001010010;
assign LUT_1[20583] = 32'b11111111111111111101111011001110;
assign LUT_1[20584] = 32'b00000000000000000000001111011111;
assign LUT_1[20585] = 32'b11111111111111111001100001011011;
assign LUT_1[20586] = 32'b11111111111111111011111101110000;
assign LUT_1[20587] = 32'b11111111111111110101001111101100;
assign LUT_1[20588] = 32'b00000000000000001000001000110110;
assign LUT_1[20589] = 32'b00000000000000000001011010110010;
assign LUT_1[20590] = 32'b00000000000000000011110111000111;
assign LUT_1[20591] = 32'b11111111111111111101001001000011;
assign LUT_1[20592] = 32'b00000000000000000010111101001100;
assign LUT_1[20593] = 32'b11111111111111111100001111001000;
assign LUT_1[20594] = 32'b11111111111111111110101011011101;
assign LUT_1[20595] = 32'b11111111111111110111111101011001;
assign LUT_1[20596] = 32'b00000000000000001010110110100011;
assign LUT_1[20597] = 32'b00000000000000000100001000011111;
assign LUT_1[20598] = 32'b00000000000000000110100100110100;
assign LUT_1[20599] = 32'b11111111111111111111110110110000;
assign LUT_1[20600] = 32'b00000000000000000010001011000001;
assign LUT_1[20601] = 32'b11111111111111111011011100111101;
assign LUT_1[20602] = 32'b11111111111111111101111001010010;
assign LUT_1[20603] = 32'b11111111111111110111001011001110;
assign LUT_1[20604] = 32'b00000000000000001010000100011000;
assign LUT_1[20605] = 32'b00000000000000000011010110010100;
assign LUT_1[20606] = 32'b00000000000000000101110010101001;
assign LUT_1[20607] = 32'b11111111111111111111000100100101;
assign LUT_1[20608] = 32'b00000000000000000001001001000110;
assign LUT_1[20609] = 32'b11111111111111111010011011000010;
assign LUT_1[20610] = 32'b11111111111111111100110111010111;
assign LUT_1[20611] = 32'b11111111111111110110001001010011;
assign LUT_1[20612] = 32'b00000000000000001001000010011101;
assign LUT_1[20613] = 32'b00000000000000000010010100011001;
assign LUT_1[20614] = 32'b00000000000000000100110000101110;
assign LUT_1[20615] = 32'b11111111111111111110000010101010;
assign LUT_1[20616] = 32'b00000000000000000000010110111011;
assign LUT_1[20617] = 32'b11111111111111111001101000110111;
assign LUT_1[20618] = 32'b11111111111111111100000101001100;
assign LUT_1[20619] = 32'b11111111111111110101010111001000;
assign LUT_1[20620] = 32'b00000000000000001000010000010010;
assign LUT_1[20621] = 32'b00000000000000000001100010001110;
assign LUT_1[20622] = 32'b00000000000000000011111110100011;
assign LUT_1[20623] = 32'b11111111111111111101010000011111;
assign LUT_1[20624] = 32'b00000000000000000011000100101000;
assign LUT_1[20625] = 32'b11111111111111111100010110100100;
assign LUT_1[20626] = 32'b11111111111111111110110010111001;
assign LUT_1[20627] = 32'b11111111111111111000000100110101;
assign LUT_1[20628] = 32'b00000000000000001010111101111111;
assign LUT_1[20629] = 32'b00000000000000000100001111111011;
assign LUT_1[20630] = 32'b00000000000000000110101100010000;
assign LUT_1[20631] = 32'b11111111111111111111111110001100;
assign LUT_1[20632] = 32'b00000000000000000010010010011101;
assign LUT_1[20633] = 32'b11111111111111111011100100011001;
assign LUT_1[20634] = 32'b11111111111111111110000000101110;
assign LUT_1[20635] = 32'b11111111111111110111010010101010;
assign LUT_1[20636] = 32'b00000000000000001010001011110100;
assign LUT_1[20637] = 32'b00000000000000000011011101110000;
assign LUT_1[20638] = 32'b00000000000000000101111010000101;
assign LUT_1[20639] = 32'b11111111111111111111001100000001;
assign LUT_1[20640] = 32'b00000000000000000010000100000101;
assign LUT_1[20641] = 32'b11111111111111111011010110000001;
assign LUT_1[20642] = 32'b11111111111111111101110010010110;
assign LUT_1[20643] = 32'b11111111111111110111000100010010;
assign LUT_1[20644] = 32'b00000000000000001001111101011100;
assign LUT_1[20645] = 32'b00000000000000000011001111011000;
assign LUT_1[20646] = 32'b00000000000000000101101011101101;
assign LUT_1[20647] = 32'b11111111111111111110111101101001;
assign LUT_1[20648] = 32'b00000000000000000001010001111010;
assign LUT_1[20649] = 32'b11111111111111111010100011110110;
assign LUT_1[20650] = 32'b11111111111111111101000000001011;
assign LUT_1[20651] = 32'b11111111111111110110010010000111;
assign LUT_1[20652] = 32'b00000000000000001001001011010001;
assign LUT_1[20653] = 32'b00000000000000000010011101001101;
assign LUT_1[20654] = 32'b00000000000000000100111001100010;
assign LUT_1[20655] = 32'b11111111111111111110001011011110;
assign LUT_1[20656] = 32'b00000000000000000011111111100111;
assign LUT_1[20657] = 32'b11111111111111111101010001100011;
assign LUT_1[20658] = 32'b11111111111111111111101101111000;
assign LUT_1[20659] = 32'b11111111111111111000111111110100;
assign LUT_1[20660] = 32'b00000000000000001011111000111110;
assign LUT_1[20661] = 32'b00000000000000000101001010111010;
assign LUT_1[20662] = 32'b00000000000000000111100111001111;
assign LUT_1[20663] = 32'b00000000000000000000111001001011;
assign LUT_1[20664] = 32'b00000000000000000011001101011100;
assign LUT_1[20665] = 32'b11111111111111111100011111011000;
assign LUT_1[20666] = 32'b11111111111111111110111011101101;
assign LUT_1[20667] = 32'b11111111111111111000001101101001;
assign LUT_1[20668] = 32'b00000000000000001011000110110011;
assign LUT_1[20669] = 32'b00000000000000000100011000101111;
assign LUT_1[20670] = 32'b00000000000000000110110101000100;
assign LUT_1[20671] = 32'b00000000000000000000000111000000;
assign LUT_1[20672] = 32'b00000000000000000011000110101110;
assign LUT_1[20673] = 32'b11111111111111111100011000101010;
assign LUT_1[20674] = 32'b11111111111111111110110100111111;
assign LUT_1[20675] = 32'b11111111111111111000000110111011;
assign LUT_1[20676] = 32'b00000000000000001011000000000101;
assign LUT_1[20677] = 32'b00000000000000000100010010000001;
assign LUT_1[20678] = 32'b00000000000000000110101110010110;
assign LUT_1[20679] = 32'b00000000000000000000000000010010;
assign LUT_1[20680] = 32'b00000000000000000010010100100011;
assign LUT_1[20681] = 32'b11111111111111111011100110011111;
assign LUT_1[20682] = 32'b11111111111111111110000010110100;
assign LUT_1[20683] = 32'b11111111111111110111010100110000;
assign LUT_1[20684] = 32'b00000000000000001010001101111010;
assign LUT_1[20685] = 32'b00000000000000000011011111110110;
assign LUT_1[20686] = 32'b00000000000000000101111100001011;
assign LUT_1[20687] = 32'b11111111111111111111001110000111;
assign LUT_1[20688] = 32'b00000000000000000101000010010000;
assign LUT_1[20689] = 32'b11111111111111111110010100001100;
assign LUT_1[20690] = 32'b00000000000000000000110000100001;
assign LUT_1[20691] = 32'b11111111111111111010000010011101;
assign LUT_1[20692] = 32'b00000000000000001100111011100111;
assign LUT_1[20693] = 32'b00000000000000000110001101100011;
assign LUT_1[20694] = 32'b00000000000000001000101001111000;
assign LUT_1[20695] = 32'b00000000000000000001111011110100;
assign LUT_1[20696] = 32'b00000000000000000100010000000101;
assign LUT_1[20697] = 32'b11111111111111111101100010000001;
assign LUT_1[20698] = 32'b11111111111111111111111110010110;
assign LUT_1[20699] = 32'b11111111111111111001010000010010;
assign LUT_1[20700] = 32'b00000000000000001100001001011100;
assign LUT_1[20701] = 32'b00000000000000000101011011011000;
assign LUT_1[20702] = 32'b00000000000000000111110111101101;
assign LUT_1[20703] = 32'b00000000000000000001001001101001;
assign LUT_1[20704] = 32'b00000000000000000100000001101101;
assign LUT_1[20705] = 32'b11111111111111111101010011101001;
assign LUT_1[20706] = 32'b11111111111111111111101111111110;
assign LUT_1[20707] = 32'b11111111111111111001000001111010;
assign LUT_1[20708] = 32'b00000000000000001011111011000100;
assign LUT_1[20709] = 32'b00000000000000000101001101000000;
assign LUT_1[20710] = 32'b00000000000000000111101001010101;
assign LUT_1[20711] = 32'b00000000000000000000111011010001;
assign LUT_1[20712] = 32'b00000000000000000011001111100010;
assign LUT_1[20713] = 32'b11111111111111111100100001011110;
assign LUT_1[20714] = 32'b11111111111111111110111101110011;
assign LUT_1[20715] = 32'b11111111111111111000001111101111;
assign LUT_1[20716] = 32'b00000000000000001011001000111001;
assign LUT_1[20717] = 32'b00000000000000000100011010110101;
assign LUT_1[20718] = 32'b00000000000000000110110111001010;
assign LUT_1[20719] = 32'b00000000000000000000001001000110;
assign LUT_1[20720] = 32'b00000000000000000101111101001111;
assign LUT_1[20721] = 32'b11111111111111111111001111001011;
assign LUT_1[20722] = 32'b00000000000000000001101011100000;
assign LUT_1[20723] = 32'b11111111111111111010111101011100;
assign LUT_1[20724] = 32'b00000000000000001101110110100110;
assign LUT_1[20725] = 32'b00000000000000000111001000100010;
assign LUT_1[20726] = 32'b00000000000000001001100100110111;
assign LUT_1[20727] = 32'b00000000000000000010110110110011;
assign LUT_1[20728] = 32'b00000000000000000101001011000100;
assign LUT_1[20729] = 32'b11111111111111111110011101000000;
assign LUT_1[20730] = 32'b00000000000000000000111001010101;
assign LUT_1[20731] = 32'b11111111111111111010001011010001;
assign LUT_1[20732] = 32'b00000000000000001101000100011011;
assign LUT_1[20733] = 32'b00000000000000000110010110010111;
assign LUT_1[20734] = 32'b00000000000000001000110010101100;
assign LUT_1[20735] = 32'b00000000000000000010000100101000;
assign LUT_1[20736] = 32'b11111111111111111011111101001111;
assign LUT_1[20737] = 32'b11111111111111110101001111001011;
assign LUT_1[20738] = 32'b11111111111111110111101011100000;
assign LUT_1[20739] = 32'b11111111111111110000111101011100;
assign LUT_1[20740] = 32'b00000000000000000011110110100110;
assign LUT_1[20741] = 32'b11111111111111111101001000100010;
assign LUT_1[20742] = 32'b11111111111111111111100100110111;
assign LUT_1[20743] = 32'b11111111111111111000110110110011;
assign LUT_1[20744] = 32'b11111111111111111011001011000100;
assign LUT_1[20745] = 32'b11111111111111110100011101000000;
assign LUT_1[20746] = 32'b11111111111111110110111001010101;
assign LUT_1[20747] = 32'b11111111111111110000001011010001;
assign LUT_1[20748] = 32'b00000000000000000011000100011011;
assign LUT_1[20749] = 32'b11111111111111111100010110010111;
assign LUT_1[20750] = 32'b11111111111111111110110010101100;
assign LUT_1[20751] = 32'b11111111111111111000000100101000;
assign LUT_1[20752] = 32'b11111111111111111101111000110001;
assign LUT_1[20753] = 32'b11111111111111110111001010101101;
assign LUT_1[20754] = 32'b11111111111111111001100111000010;
assign LUT_1[20755] = 32'b11111111111111110010111000111110;
assign LUT_1[20756] = 32'b00000000000000000101110010001000;
assign LUT_1[20757] = 32'b11111111111111111111000100000100;
assign LUT_1[20758] = 32'b00000000000000000001100000011001;
assign LUT_1[20759] = 32'b11111111111111111010110010010101;
assign LUT_1[20760] = 32'b11111111111111111101000110100110;
assign LUT_1[20761] = 32'b11111111111111110110011000100010;
assign LUT_1[20762] = 32'b11111111111111111000110100110111;
assign LUT_1[20763] = 32'b11111111111111110010000110110011;
assign LUT_1[20764] = 32'b00000000000000000100111111111101;
assign LUT_1[20765] = 32'b11111111111111111110010001111001;
assign LUT_1[20766] = 32'b00000000000000000000101110001110;
assign LUT_1[20767] = 32'b11111111111111111010000000001010;
assign LUT_1[20768] = 32'b11111111111111111100111000001110;
assign LUT_1[20769] = 32'b11111111111111110110001010001010;
assign LUT_1[20770] = 32'b11111111111111111000100110011111;
assign LUT_1[20771] = 32'b11111111111111110001111000011011;
assign LUT_1[20772] = 32'b00000000000000000100110001100101;
assign LUT_1[20773] = 32'b11111111111111111110000011100001;
assign LUT_1[20774] = 32'b00000000000000000000011111110110;
assign LUT_1[20775] = 32'b11111111111111111001110001110010;
assign LUT_1[20776] = 32'b11111111111111111100000110000011;
assign LUT_1[20777] = 32'b11111111111111110101010111111111;
assign LUT_1[20778] = 32'b11111111111111110111110100010100;
assign LUT_1[20779] = 32'b11111111111111110001000110010000;
assign LUT_1[20780] = 32'b00000000000000000011111111011010;
assign LUT_1[20781] = 32'b11111111111111111101010001010110;
assign LUT_1[20782] = 32'b11111111111111111111101101101011;
assign LUT_1[20783] = 32'b11111111111111111000111111100111;
assign LUT_1[20784] = 32'b11111111111111111110110011110000;
assign LUT_1[20785] = 32'b11111111111111111000000101101100;
assign LUT_1[20786] = 32'b11111111111111111010100010000001;
assign LUT_1[20787] = 32'b11111111111111110011110011111101;
assign LUT_1[20788] = 32'b00000000000000000110101101000111;
assign LUT_1[20789] = 32'b11111111111111111111111111000011;
assign LUT_1[20790] = 32'b00000000000000000010011011011000;
assign LUT_1[20791] = 32'b11111111111111111011101101010100;
assign LUT_1[20792] = 32'b11111111111111111110000001100101;
assign LUT_1[20793] = 32'b11111111111111110111010011100001;
assign LUT_1[20794] = 32'b11111111111111111001101111110110;
assign LUT_1[20795] = 32'b11111111111111110011000001110010;
assign LUT_1[20796] = 32'b00000000000000000101111010111100;
assign LUT_1[20797] = 32'b11111111111111111111001100111000;
assign LUT_1[20798] = 32'b00000000000000000001101001001101;
assign LUT_1[20799] = 32'b11111111111111111010111011001001;
assign LUT_1[20800] = 32'b11111111111111111101111010110111;
assign LUT_1[20801] = 32'b11111111111111110111001100110011;
assign LUT_1[20802] = 32'b11111111111111111001101001001000;
assign LUT_1[20803] = 32'b11111111111111110010111011000100;
assign LUT_1[20804] = 32'b00000000000000000101110100001110;
assign LUT_1[20805] = 32'b11111111111111111111000110001010;
assign LUT_1[20806] = 32'b00000000000000000001100010011111;
assign LUT_1[20807] = 32'b11111111111111111010110100011011;
assign LUT_1[20808] = 32'b11111111111111111101001000101100;
assign LUT_1[20809] = 32'b11111111111111110110011010101000;
assign LUT_1[20810] = 32'b11111111111111111000110110111101;
assign LUT_1[20811] = 32'b11111111111111110010001000111001;
assign LUT_1[20812] = 32'b00000000000000000101000010000011;
assign LUT_1[20813] = 32'b11111111111111111110010011111111;
assign LUT_1[20814] = 32'b00000000000000000000110000010100;
assign LUT_1[20815] = 32'b11111111111111111010000010010000;
assign LUT_1[20816] = 32'b11111111111111111111110110011001;
assign LUT_1[20817] = 32'b11111111111111111001001000010101;
assign LUT_1[20818] = 32'b11111111111111111011100100101010;
assign LUT_1[20819] = 32'b11111111111111110100110110100110;
assign LUT_1[20820] = 32'b00000000000000000111101111110000;
assign LUT_1[20821] = 32'b00000000000000000001000001101100;
assign LUT_1[20822] = 32'b00000000000000000011011110000001;
assign LUT_1[20823] = 32'b11111111111111111100101111111101;
assign LUT_1[20824] = 32'b11111111111111111111000100001110;
assign LUT_1[20825] = 32'b11111111111111111000010110001010;
assign LUT_1[20826] = 32'b11111111111111111010110010011111;
assign LUT_1[20827] = 32'b11111111111111110100000100011011;
assign LUT_1[20828] = 32'b00000000000000000110111101100101;
assign LUT_1[20829] = 32'b00000000000000000000001111100001;
assign LUT_1[20830] = 32'b00000000000000000010101011110110;
assign LUT_1[20831] = 32'b11111111111111111011111101110010;
assign LUT_1[20832] = 32'b11111111111111111110110101110110;
assign LUT_1[20833] = 32'b11111111111111111000000111110010;
assign LUT_1[20834] = 32'b11111111111111111010100100000111;
assign LUT_1[20835] = 32'b11111111111111110011110110000011;
assign LUT_1[20836] = 32'b00000000000000000110101111001101;
assign LUT_1[20837] = 32'b00000000000000000000000001001001;
assign LUT_1[20838] = 32'b00000000000000000010011101011110;
assign LUT_1[20839] = 32'b11111111111111111011101111011010;
assign LUT_1[20840] = 32'b11111111111111111110000011101011;
assign LUT_1[20841] = 32'b11111111111111110111010101100111;
assign LUT_1[20842] = 32'b11111111111111111001110001111100;
assign LUT_1[20843] = 32'b11111111111111110011000011111000;
assign LUT_1[20844] = 32'b00000000000000000101111101000010;
assign LUT_1[20845] = 32'b11111111111111111111001110111110;
assign LUT_1[20846] = 32'b00000000000000000001101011010011;
assign LUT_1[20847] = 32'b11111111111111111010111101001111;
assign LUT_1[20848] = 32'b00000000000000000000110001011000;
assign LUT_1[20849] = 32'b11111111111111111010000011010100;
assign LUT_1[20850] = 32'b11111111111111111100011111101001;
assign LUT_1[20851] = 32'b11111111111111110101110001100101;
assign LUT_1[20852] = 32'b00000000000000001000101010101111;
assign LUT_1[20853] = 32'b00000000000000000001111100101011;
assign LUT_1[20854] = 32'b00000000000000000100011001000000;
assign LUT_1[20855] = 32'b11111111111111111101101010111100;
assign LUT_1[20856] = 32'b11111111111111111111111111001101;
assign LUT_1[20857] = 32'b11111111111111111001010001001001;
assign LUT_1[20858] = 32'b11111111111111111011101101011110;
assign LUT_1[20859] = 32'b11111111111111110100111111011010;
assign LUT_1[20860] = 32'b00000000000000000111111000100100;
assign LUT_1[20861] = 32'b00000000000000000001001010100000;
assign LUT_1[20862] = 32'b00000000000000000011100110110101;
assign LUT_1[20863] = 32'b11111111111111111100111000110001;
assign LUT_1[20864] = 32'b11111111111111111110111101010010;
assign LUT_1[20865] = 32'b11111111111111111000001111001110;
assign LUT_1[20866] = 32'b11111111111111111010101011100011;
assign LUT_1[20867] = 32'b11111111111111110011111101011111;
assign LUT_1[20868] = 32'b00000000000000000110110110101001;
assign LUT_1[20869] = 32'b00000000000000000000001000100101;
assign LUT_1[20870] = 32'b00000000000000000010100100111010;
assign LUT_1[20871] = 32'b11111111111111111011110110110110;
assign LUT_1[20872] = 32'b11111111111111111110001011000111;
assign LUT_1[20873] = 32'b11111111111111110111011101000011;
assign LUT_1[20874] = 32'b11111111111111111001111001011000;
assign LUT_1[20875] = 32'b11111111111111110011001011010100;
assign LUT_1[20876] = 32'b00000000000000000110000100011110;
assign LUT_1[20877] = 32'b11111111111111111111010110011010;
assign LUT_1[20878] = 32'b00000000000000000001110010101111;
assign LUT_1[20879] = 32'b11111111111111111011000100101011;
assign LUT_1[20880] = 32'b00000000000000000000111000110100;
assign LUT_1[20881] = 32'b11111111111111111010001010110000;
assign LUT_1[20882] = 32'b11111111111111111100100111000101;
assign LUT_1[20883] = 32'b11111111111111110101111001000001;
assign LUT_1[20884] = 32'b00000000000000001000110010001011;
assign LUT_1[20885] = 32'b00000000000000000010000100000111;
assign LUT_1[20886] = 32'b00000000000000000100100000011100;
assign LUT_1[20887] = 32'b11111111111111111101110010011000;
assign LUT_1[20888] = 32'b00000000000000000000000110101001;
assign LUT_1[20889] = 32'b11111111111111111001011000100101;
assign LUT_1[20890] = 32'b11111111111111111011110100111010;
assign LUT_1[20891] = 32'b11111111111111110101000110110110;
assign LUT_1[20892] = 32'b00000000000000001000000000000000;
assign LUT_1[20893] = 32'b00000000000000000001010001111100;
assign LUT_1[20894] = 32'b00000000000000000011101110010001;
assign LUT_1[20895] = 32'b11111111111111111101000000001101;
assign LUT_1[20896] = 32'b11111111111111111111111000010001;
assign LUT_1[20897] = 32'b11111111111111111001001010001101;
assign LUT_1[20898] = 32'b11111111111111111011100110100010;
assign LUT_1[20899] = 32'b11111111111111110100111000011110;
assign LUT_1[20900] = 32'b00000000000000000111110001101000;
assign LUT_1[20901] = 32'b00000000000000000001000011100100;
assign LUT_1[20902] = 32'b00000000000000000011011111111001;
assign LUT_1[20903] = 32'b11111111111111111100110001110101;
assign LUT_1[20904] = 32'b11111111111111111111000110000110;
assign LUT_1[20905] = 32'b11111111111111111000011000000010;
assign LUT_1[20906] = 32'b11111111111111111010110100010111;
assign LUT_1[20907] = 32'b11111111111111110100000110010011;
assign LUT_1[20908] = 32'b00000000000000000110111111011101;
assign LUT_1[20909] = 32'b00000000000000000000010001011001;
assign LUT_1[20910] = 32'b00000000000000000010101101101110;
assign LUT_1[20911] = 32'b11111111111111111011111111101010;
assign LUT_1[20912] = 32'b00000000000000000001110011110011;
assign LUT_1[20913] = 32'b11111111111111111011000101101111;
assign LUT_1[20914] = 32'b11111111111111111101100010000100;
assign LUT_1[20915] = 32'b11111111111111110110110100000000;
assign LUT_1[20916] = 32'b00000000000000001001101101001010;
assign LUT_1[20917] = 32'b00000000000000000010111111000110;
assign LUT_1[20918] = 32'b00000000000000000101011011011011;
assign LUT_1[20919] = 32'b11111111111111111110101101010111;
assign LUT_1[20920] = 32'b00000000000000000001000001101000;
assign LUT_1[20921] = 32'b11111111111111111010010011100100;
assign LUT_1[20922] = 32'b11111111111111111100101111111001;
assign LUT_1[20923] = 32'b11111111111111110110000001110101;
assign LUT_1[20924] = 32'b00000000000000001000111010111111;
assign LUT_1[20925] = 32'b00000000000000000010001100111011;
assign LUT_1[20926] = 32'b00000000000000000100101001010000;
assign LUT_1[20927] = 32'b11111111111111111101111011001100;
assign LUT_1[20928] = 32'b00000000000000000000111010111010;
assign LUT_1[20929] = 32'b11111111111111111010001100110110;
assign LUT_1[20930] = 32'b11111111111111111100101001001011;
assign LUT_1[20931] = 32'b11111111111111110101111011000111;
assign LUT_1[20932] = 32'b00000000000000001000110100010001;
assign LUT_1[20933] = 32'b00000000000000000010000110001101;
assign LUT_1[20934] = 32'b00000000000000000100100010100010;
assign LUT_1[20935] = 32'b11111111111111111101110100011110;
assign LUT_1[20936] = 32'b00000000000000000000001000101111;
assign LUT_1[20937] = 32'b11111111111111111001011010101011;
assign LUT_1[20938] = 32'b11111111111111111011110111000000;
assign LUT_1[20939] = 32'b11111111111111110101001000111100;
assign LUT_1[20940] = 32'b00000000000000001000000010000110;
assign LUT_1[20941] = 32'b00000000000000000001010100000010;
assign LUT_1[20942] = 32'b00000000000000000011110000010111;
assign LUT_1[20943] = 32'b11111111111111111101000010010011;
assign LUT_1[20944] = 32'b00000000000000000010110110011100;
assign LUT_1[20945] = 32'b11111111111111111100001000011000;
assign LUT_1[20946] = 32'b11111111111111111110100100101101;
assign LUT_1[20947] = 32'b11111111111111110111110110101001;
assign LUT_1[20948] = 32'b00000000000000001010101111110011;
assign LUT_1[20949] = 32'b00000000000000000100000001101111;
assign LUT_1[20950] = 32'b00000000000000000110011110000100;
assign LUT_1[20951] = 32'b11111111111111111111110000000000;
assign LUT_1[20952] = 32'b00000000000000000010000100010001;
assign LUT_1[20953] = 32'b11111111111111111011010110001101;
assign LUT_1[20954] = 32'b11111111111111111101110010100010;
assign LUT_1[20955] = 32'b11111111111111110111000100011110;
assign LUT_1[20956] = 32'b00000000000000001001111101101000;
assign LUT_1[20957] = 32'b00000000000000000011001111100100;
assign LUT_1[20958] = 32'b00000000000000000101101011111001;
assign LUT_1[20959] = 32'b11111111111111111110111101110101;
assign LUT_1[20960] = 32'b00000000000000000001110101111001;
assign LUT_1[20961] = 32'b11111111111111111011000111110101;
assign LUT_1[20962] = 32'b11111111111111111101100100001010;
assign LUT_1[20963] = 32'b11111111111111110110110110000110;
assign LUT_1[20964] = 32'b00000000000000001001101111010000;
assign LUT_1[20965] = 32'b00000000000000000011000001001100;
assign LUT_1[20966] = 32'b00000000000000000101011101100001;
assign LUT_1[20967] = 32'b11111111111111111110101111011101;
assign LUT_1[20968] = 32'b00000000000000000001000011101110;
assign LUT_1[20969] = 32'b11111111111111111010010101101010;
assign LUT_1[20970] = 32'b11111111111111111100110001111111;
assign LUT_1[20971] = 32'b11111111111111110110000011111011;
assign LUT_1[20972] = 32'b00000000000000001000111101000101;
assign LUT_1[20973] = 32'b00000000000000000010001111000001;
assign LUT_1[20974] = 32'b00000000000000000100101011010110;
assign LUT_1[20975] = 32'b11111111111111111101111101010010;
assign LUT_1[20976] = 32'b00000000000000000011110001011011;
assign LUT_1[20977] = 32'b11111111111111111101000011010111;
assign LUT_1[20978] = 32'b11111111111111111111011111101100;
assign LUT_1[20979] = 32'b11111111111111111000110001101000;
assign LUT_1[20980] = 32'b00000000000000001011101010110010;
assign LUT_1[20981] = 32'b00000000000000000100111100101110;
assign LUT_1[20982] = 32'b00000000000000000111011001000011;
assign LUT_1[20983] = 32'b00000000000000000000101010111111;
assign LUT_1[20984] = 32'b00000000000000000010111111010000;
assign LUT_1[20985] = 32'b11111111111111111100010001001100;
assign LUT_1[20986] = 32'b11111111111111111110101101100001;
assign LUT_1[20987] = 32'b11111111111111110111111111011101;
assign LUT_1[20988] = 32'b00000000000000001010111000100111;
assign LUT_1[20989] = 32'b00000000000000000100001010100011;
assign LUT_1[20990] = 32'b00000000000000000110100110111000;
assign LUT_1[20991] = 32'b11111111111111111111111000110100;
assign LUT_1[20992] = 32'b11111111111111110111110111100000;
assign LUT_1[20993] = 32'b11111111111111110001001001011100;
assign LUT_1[20994] = 32'b11111111111111110011100101110001;
assign LUT_1[20995] = 32'b11111111111111101100110111101101;
assign LUT_1[20996] = 32'b11111111111111111111110000110111;
assign LUT_1[20997] = 32'b11111111111111111001000010110011;
assign LUT_1[20998] = 32'b11111111111111111011011111001000;
assign LUT_1[20999] = 32'b11111111111111110100110001000100;
assign LUT_1[21000] = 32'b11111111111111110111000101010101;
assign LUT_1[21001] = 32'b11111111111111110000010111010001;
assign LUT_1[21002] = 32'b11111111111111110010110011100110;
assign LUT_1[21003] = 32'b11111111111111101100000101100010;
assign LUT_1[21004] = 32'b11111111111111111110111110101100;
assign LUT_1[21005] = 32'b11111111111111111000010000101000;
assign LUT_1[21006] = 32'b11111111111111111010101100111101;
assign LUT_1[21007] = 32'b11111111111111110011111110111001;
assign LUT_1[21008] = 32'b11111111111111111001110011000010;
assign LUT_1[21009] = 32'b11111111111111110011000100111110;
assign LUT_1[21010] = 32'b11111111111111110101100001010011;
assign LUT_1[21011] = 32'b11111111111111101110110011001111;
assign LUT_1[21012] = 32'b00000000000000000001101100011001;
assign LUT_1[21013] = 32'b11111111111111111010111110010101;
assign LUT_1[21014] = 32'b11111111111111111101011010101010;
assign LUT_1[21015] = 32'b11111111111111110110101100100110;
assign LUT_1[21016] = 32'b11111111111111111001000000110111;
assign LUT_1[21017] = 32'b11111111111111110010010010110011;
assign LUT_1[21018] = 32'b11111111111111110100101111001000;
assign LUT_1[21019] = 32'b11111111111111101110000001000100;
assign LUT_1[21020] = 32'b00000000000000000000111010001110;
assign LUT_1[21021] = 32'b11111111111111111010001100001010;
assign LUT_1[21022] = 32'b11111111111111111100101000011111;
assign LUT_1[21023] = 32'b11111111111111110101111010011011;
assign LUT_1[21024] = 32'b11111111111111111000110010011111;
assign LUT_1[21025] = 32'b11111111111111110010000100011011;
assign LUT_1[21026] = 32'b11111111111111110100100000110000;
assign LUT_1[21027] = 32'b11111111111111101101110010101100;
assign LUT_1[21028] = 32'b00000000000000000000101011110110;
assign LUT_1[21029] = 32'b11111111111111111001111101110010;
assign LUT_1[21030] = 32'b11111111111111111100011010000111;
assign LUT_1[21031] = 32'b11111111111111110101101100000011;
assign LUT_1[21032] = 32'b11111111111111111000000000010100;
assign LUT_1[21033] = 32'b11111111111111110001010010010000;
assign LUT_1[21034] = 32'b11111111111111110011101110100101;
assign LUT_1[21035] = 32'b11111111111111101101000000100001;
assign LUT_1[21036] = 32'b11111111111111111111111001101011;
assign LUT_1[21037] = 32'b11111111111111111001001011100111;
assign LUT_1[21038] = 32'b11111111111111111011100111111100;
assign LUT_1[21039] = 32'b11111111111111110100111001111000;
assign LUT_1[21040] = 32'b11111111111111111010101110000001;
assign LUT_1[21041] = 32'b11111111111111110011111111111101;
assign LUT_1[21042] = 32'b11111111111111110110011100010010;
assign LUT_1[21043] = 32'b11111111111111101111101110001110;
assign LUT_1[21044] = 32'b00000000000000000010100111011000;
assign LUT_1[21045] = 32'b11111111111111111011111001010100;
assign LUT_1[21046] = 32'b11111111111111111110010101101001;
assign LUT_1[21047] = 32'b11111111111111110111100111100101;
assign LUT_1[21048] = 32'b11111111111111111001111011110110;
assign LUT_1[21049] = 32'b11111111111111110011001101110010;
assign LUT_1[21050] = 32'b11111111111111110101101010000111;
assign LUT_1[21051] = 32'b11111111111111101110111100000011;
assign LUT_1[21052] = 32'b00000000000000000001110101001101;
assign LUT_1[21053] = 32'b11111111111111111011000111001001;
assign LUT_1[21054] = 32'b11111111111111111101100011011110;
assign LUT_1[21055] = 32'b11111111111111110110110101011010;
assign LUT_1[21056] = 32'b11111111111111111001110101001000;
assign LUT_1[21057] = 32'b11111111111111110011000111000100;
assign LUT_1[21058] = 32'b11111111111111110101100011011001;
assign LUT_1[21059] = 32'b11111111111111101110110101010101;
assign LUT_1[21060] = 32'b00000000000000000001101110011111;
assign LUT_1[21061] = 32'b11111111111111111011000000011011;
assign LUT_1[21062] = 32'b11111111111111111101011100110000;
assign LUT_1[21063] = 32'b11111111111111110110101110101100;
assign LUT_1[21064] = 32'b11111111111111111001000010111101;
assign LUT_1[21065] = 32'b11111111111111110010010100111001;
assign LUT_1[21066] = 32'b11111111111111110100110001001110;
assign LUT_1[21067] = 32'b11111111111111101110000011001010;
assign LUT_1[21068] = 32'b00000000000000000000111100010100;
assign LUT_1[21069] = 32'b11111111111111111010001110010000;
assign LUT_1[21070] = 32'b11111111111111111100101010100101;
assign LUT_1[21071] = 32'b11111111111111110101111100100001;
assign LUT_1[21072] = 32'b11111111111111111011110000101010;
assign LUT_1[21073] = 32'b11111111111111110101000010100110;
assign LUT_1[21074] = 32'b11111111111111110111011110111011;
assign LUT_1[21075] = 32'b11111111111111110000110000110111;
assign LUT_1[21076] = 32'b00000000000000000011101010000001;
assign LUT_1[21077] = 32'b11111111111111111100111011111101;
assign LUT_1[21078] = 32'b11111111111111111111011000010010;
assign LUT_1[21079] = 32'b11111111111111111000101010001110;
assign LUT_1[21080] = 32'b11111111111111111010111110011111;
assign LUT_1[21081] = 32'b11111111111111110100010000011011;
assign LUT_1[21082] = 32'b11111111111111110110101100110000;
assign LUT_1[21083] = 32'b11111111111111101111111110101100;
assign LUT_1[21084] = 32'b00000000000000000010110111110110;
assign LUT_1[21085] = 32'b11111111111111111100001001110010;
assign LUT_1[21086] = 32'b11111111111111111110100110000111;
assign LUT_1[21087] = 32'b11111111111111110111111000000011;
assign LUT_1[21088] = 32'b11111111111111111010110000000111;
assign LUT_1[21089] = 32'b11111111111111110100000010000011;
assign LUT_1[21090] = 32'b11111111111111110110011110011000;
assign LUT_1[21091] = 32'b11111111111111101111110000010100;
assign LUT_1[21092] = 32'b00000000000000000010101001011110;
assign LUT_1[21093] = 32'b11111111111111111011111011011010;
assign LUT_1[21094] = 32'b11111111111111111110010111101111;
assign LUT_1[21095] = 32'b11111111111111110111101001101011;
assign LUT_1[21096] = 32'b11111111111111111001111101111100;
assign LUT_1[21097] = 32'b11111111111111110011001111111000;
assign LUT_1[21098] = 32'b11111111111111110101101100001101;
assign LUT_1[21099] = 32'b11111111111111101110111110001001;
assign LUT_1[21100] = 32'b00000000000000000001110111010011;
assign LUT_1[21101] = 32'b11111111111111111011001001001111;
assign LUT_1[21102] = 32'b11111111111111111101100101100100;
assign LUT_1[21103] = 32'b11111111111111110110110111100000;
assign LUT_1[21104] = 32'b11111111111111111100101011101001;
assign LUT_1[21105] = 32'b11111111111111110101111101100101;
assign LUT_1[21106] = 32'b11111111111111111000011001111010;
assign LUT_1[21107] = 32'b11111111111111110001101011110110;
assign LUT_1[21108] = 32'b00000000000000000100100101000000;
assign LUT_1[21109] = 32'b11111111111111111101110110111100;
assign LUT_1[21110] = 32'b00000000000000000000010011010001;
assign LUT_1[21111] = 32'b11111111111111111001100101001101;
assign LUT_1[21112] = 32'b11111111111111111011111001011110;
assign LUT_1[21113] = 32'b11111111111111110101001011011010;
assign LUT_1[21114] = 32'b11111111111111110111100111101111;
assign LUT_1[21115] = 32'b11111111111111110000111001101011;
assign LUT_1[21116] = 32'b00000000000000000011110010110101;
assign LUT_1[21117] = 32'b11111111111111111101000100110001;
assign LUT_1[21118] = 32'b11111111111111111111100001000110;
assign LUT_1[21119] = 32'b11111111111111111000110011000010;
assign LUT_1[21120] = 32'b11111111111111111010110111100011;
assign LUT_1[21121] = 32'b11111111111111110100001001011111;
assign LUT_1[21122] = 32'b11111111111111110110100101110100;
assign LUT_1[21123] = 32'b11111111111111101111110111110000;
assign LUT_1[21124] = 32'b00000000000000000010110000111010;
assign LUT_1[21125] = 32'b11111111111111111100000010110110;
assign LUT_1[21126] = 32'b11111111111111111110011111001011;
assign LUT_1[21127] = 32'b11111111111111110111110001000111;
assign LUT_1[21128] = 32'b11111111111111111010000101011000;
assign LUT_1[21129] = 32'b11111111111111110011010111010100;
assign LUT_1[21130] = 32'b11111111111111110101110011101001;
assign LUT_1[21131] = 32'b11111111111111101111000101100101;
assign LUT_1[21132] = 32'b00000000000000000001111110101111;
assign LUT_1[21133] = 32'b11111111111111111011010000101011;
assign LUT_1[21134] = 32'b11111111111111111101101101000000;
assign LUT_1[21135] = 32'b11111111111111110110111110111100;
assign LUT_1[21136] = 32'b11111111111111111100110011000101;
assign LUT_1[21137] = 32'b11111111111111110110000101000001;
assign LUT_1[21138] = 32'b11111111111111111000100001010110;
assign LUT_1[21139] = 32'b11111111111111110001110011010010;
assign LUT_1[21140] = 32'b00000000000000000100101100011100;
assign LUT_1[21141] = 32'b11111111111111111101111110011000;
assign LUT_1[21142] = 32'b00000000000000000000011010101101;
assign LUT_1[21143] = 32'b11111111111111111001101100101001;
assign LUT_1[21144] = 32'b11111111111111111100000000111010;
assign LUT_1[21145] = 32'b11111111111111110101010010110110;
assign LUT_1[21146] = 32'b11111111111111110111101111001011;
assign LUT_1[21147] = 32'b11111111111111110001000001000111;
assign LUT_1[21148] = 32'b00000000000000000011111010010001;
assign LUT_1[21149] = 32'b11111111111111111101001100001101;
assign LUT_1[21150] = 32'b11111111111111111111101000100010;
assign LUT_1[21151] = 32'b11111111111111111000111010011110;
assign LUT_1[21152] = 32'b11111111111111111011110010100010;
assign LUT_1[21153] = 32'b11111111111111110101000100011110;
assign LUT_1[21154] = 32'b11111111111111110111100000110011;
assign LUT_1[21155] = 32'b11111111111111110000110010101111;
assign LUT_1[21156] = 32'b00000000000000000011101011111001;
assign LUT_1[21157] = 32'b11111111111111111100111101110101;
assign LUT_1[21158] = 32'b11111111111111111111011010001010;
assign LUT_1[21159] = 32'b11111111111111111000101100000110;
assign LUT_1[21160] = 32'b11111111111111111011000000010111;
assign LUT_1[21161] = 32'b11111111111111110100010010010011;
assign LUT_1[21162] = 32'b11111111111111110110101110101000;
assign LUT_1[21163] = 32'b11111111111111110000000000100100;
assign LUT_1[21164] = 32'b00000000000000000010111001101110;
assign LUT_1[21165] = 32'b11111111111111111100001011101010;
assign LUT_1[21166] = 32'b11111111111111111110100111111111;
assign LUT_1[21167] = 32'b11111111111111110111111001111011;
assign LUT_1[21168] = 32'b11111111111111111101101110000100;
assign LUT_1[21169] = 32'b11111111111111110111000000000000;
assign LUT_1[21170] = 32'b11111111111111111001011100010101;
assign LUT_1[21171] = 32'b11111111111111110010101110010001;
assign LUT_1[21172] = 32'b00000000000000000101100111011011;
assign LUT_1[21173] = 32'b11111111111111111110111001010111;
assign LUT_1[21174] = 32'b00000000000000000001010101101100;
assign LUT_1[21175] = 32'b11111111111111111010100111101000;
assign LUT_1[21176] = 32'b11111111111111111100111011111001;
assign LUT_1[21177] = 32'b11111111111111110110001101110101;
assign LUT_1[21178] = 32'b11111111111111111000101010001010;
assign LUT_1[21179] = 32'b11111111111111110001111100000110;
assign LUT_1[21180] = 32'b00000000000000000100110101010000;
assign LUT_1[21181] = 32'b11111111111111111110000111001100;
assign LUT_1[21182] = 32'b00000000000000000000100011100001;
assign LUT_1[21183] = 32'b11111111111111111001110101011101;
assign LUT_1[21184] = 32'b11111111111111111100110101001011;
assign LUT_1[21185] = 32'b11111111111111110110000111000111;
assign LUT_1[21186] = 32'b11111111111111111000100011011100;
assign LUT_1[21187] = 32'b11111111111111110001110101011000;
assign LUT_1[21188] = 32'b00000000000000000100101110100010;
assign LUT_1[21189] = 32'b11111111111111111110000000011110;
assign LUT_1[21190] = 32'b00000000000000000000011100110011;
assign LUT_1[21191] = 32'b11111111111111111001101110101111;
assign LUT_1[21192] = 32'b11111111111111111100000011000000;
assign LUT_1[21193] = 32'b11111111111111110101010100111100;
assign LUT_1[21194] = 32'b11111111111111110111110001010001;
assign LUT_1[21195] = 32'b11111111111111110001000011001101;
assign LUT_1[21196] = 32'b00000000000000000011111100010111;
assign LUT_1[21197] = 32'b11111111111111111101001110010011;
assign LUT_1[21198] = 32'b11111111111111111111101010101000;
assign LUT_1[21199] = 32'b11111111111111111000111100100100;
assign LUT_1[21200] = 32'b11111111111111111110110000101101;
assign LUT_1[21201] = 32'b11111111111111111000000010101001;
assign LUT_1[21202] = 32'b11111111111111111010011110111110;
assign LUT_1[21203] = 32'b11111111111111110011110000111010;
assign LUT_1[21204] = 32'b00000000000000000110101010000100;
assign LUT_1[21205] = 32'b11111111111111111111111100000000;
assign LUT_1[21206] = 32'b00000000000000000010011000010101;
assign LUT_1[21207] = 32'b11111111111111111011101010010001;
assign LUT_1[21208] = 32'b11111111111111111101111110100010;
assign LUT_1[21209] = 32'b11111111111111110111010000011110;
assign LUT_1[21210] = 32'b11111111111111111001101100110011;
assign LUT_1[21211] = 32'b11111111111111110010111110101111;
assign LUT_1[21212] = 32'b00000000000000000101110111111001;
assign LUT_1[21213] = 32'b11111111111111111111001001110101;
assign LUT_1[21214] = 32'b00000000000000000001100110001010;
assign LUT_1[21215] = 32'b11111111111111111010111000000110;
assign LUT_1[21216] = 32'b11111111111111111101110000001010;
assign LUT_1[21217] = 32'b11111111111111110111000010000110;
assign LUT_1[21218] = 32'b11111111111111111001011110011011;
assign LUT_1[21219] = 32'b11111111111111110010110000010111;
assign LUT_1[21220] = 32'b00000000000000000101101001100001;
assign LUT_1[21221] = 32'b11111111111111111110111011011101;
assign LUT_1[21222] = 32'b00000000000000000001010111110010;
assign LUT_1[21223] = 32'b11111111111111111010101001101110;
assign LUT_1[21224] = 32'b11111111111111111100111101111111;
assign LUT_1[21225] = 32'b11111111111111110110001111111011;
assign LUT_1[21226] = 32'b11111111111111111000101100010000;
assign LUT_1[21227] = 32'b11111111111111110001111110001100;
assign LUT_1[21228] = 32'b00000000000000000100110111010110;
assign LUT_1[21229] = 32'b11111111111111111110001001010010;
assign LUT_1[21230] = 32'b00000000000000000000100101100111;
assign LUT_1[21231] = 32'b11111111111111111001110111100011;
assign LUT_1[21232] = 32'b11111111111111111111101011101100;
assign LUT_1[21233] = 32'b11111111111111111000111101101000;
assign LUT_1[21234] = 32'b11111111111111111011011001111101;
assign LUT_1[21235] = 32'b11111111111111110100101011111001;
assign LUT_1[21236] = 32'b00000000000000000111100101000011;
assign LUT_1[21237] = 32'b00000000000000000000110110111111;
assign LUT_1[21238] = 32'b00000000000000000011010011010100;
assign LUT_1[21239] = 32'b11111111111111111100100101010000;
assign LUT_1[21240] = 32'b11111111111111111110111001100001;
assign LUT_1[21241] = 32'b11111111111111111000001011011101;
assign LUT_1[21242] = 32'b11111111111111111010100111110010;
assign LUT_1[21243] = 32'b11111111111111110011111001101110;
assign LUT_1[21244] = 32'b00000000000000000110110010111000;
assign LUT_1[21245] = 32'b00000000000000000000000100110100;
assign LUT_1[21246] = 32'b00000000000000000010100001001001;
assign LUT_1[21247] = 32'b11111111111111111011110011000101;
assign LUT_1[21248] = 32'b11111111111111110101101011101100;
assign LUT_1[21249] = 32'b11111111111111101110111101101000;
assign LUT_1[21250] = 32'b11111111111111110001011001111101;
assign LUT_1[21251] = 32'b11111111111111101010101011111001;
assign LUT_1[21252] = 32'b11111111111111111101100101000011;
assign LUT_1[21253] = 32'b11111111111111110110110110111111;
assign LUT_1[21254] = 32'b11111111111111111001010011010100;
assign LUT_1[21255] = 32'b11111111111111110010100101010000;
assign LUT_1[21256] = 32'b11111111111111110100111001100001;
assign LUT_1[21257] = 32'b11111111111111101110001011011101;
assign LUT_1[21258] = 32'b11111111111111110000100111110010;
assign LUT_1[21259] = 32'b11111111111111101001111001101110;
assign LUT_1[21260] = 32'b11111111111111111100110010111000;
assign LUT_1[21261] = 32'b11111111111111110110000100110100;
assign LUT_1[21262] = 32'b11111111111111111000100001001001;
assign LUT_1[21263] = 32'b11111111111111110001110011000101;
assign LUT_1[21264] = 32'b11111111111111110111100111001110;
assign LUT_1[21265] = 32'b11111111111111110000111001001010;
assign LUT_1[21266] = 32'b11111111111111110011010101011111;
assign LUT_1[21267] = 32'b11111111111111101100100111011011;
assign LUT_1[21268] = 32'b11111111111111111111100000100101;
assign LUT_1[21269] = 32'b11111111111111111000110010100001;
assign LUT_1[21270] = 32'b11111111111111111011001110110110;
assign LUT_1[21271] = 32'b11111111111111110100100000110010;
assign LUT_1[21272] = 32'b11111111111111110110110101000011;
assign LUT_1[21273] = 32'b11111111111111110000000110111111;
assign LUT_1[21274] = 32'b11111111111111110010100011010100;
assign LUT_1[21275] = 32'b11111111111111101011110101010000;
assign LUT_1[21276] = 32'b11111111111111111110101110011010;
assign LUT_1[21277] = 32'b11111111111111111000000000010110;
assign LUT_1[21278] = 32'b11111111111111111010011100101011;
assign LUT_1[21279] = 32'b11111111111111110011101110100111;
assign LUT_1[21280] = 32'b11111111111111110110100110101011;
assign LUT_1[21281] = 32'b11111111111111101111111000100111;
assign LUT_1[21282] = 32'b11111111111111110010010100111100;
assign LUT_1[21283] = 32'b11111111111111101011100110111000;
assign LUT_1[21284] = 32'b11111111111111111110100000000010;
assign LUT_1[21285] = 32'b11111111111111110111110001111110;
assign LUT_1[21286] = 32'b11111111111111111010001110010011;
assign LUT_1[21287] = 32'b11111111111111110011100000001111;
assign LUT_1[21288] = 32'b11111111111111110101110100100000;
assign LUT_1[21289] = 32'b11111111111111101111000110011100;
assign LUT_1[21290] = 32'b11111111111111110001100010110001;
assign LUT_1[21291] = 32'b11111111111111101010110100101101;
assign LUT_1[21292] = 32'b11111111111111111101101101110111;
assign LUT_1[21293] = 32'b11111111111111110110111111110011;
assign LUT_1[21294] = 32'b11111111111111111001011100001000;
assign LUT_1[21295] = 32'b11111111111111110010101110000100;
assign LUT_1[21296] = 32'b11111111111111111000100010001101;
assign LUT_1[21297] = 32'b11111111111111110001110100001001;
assign LUT_1[21298] = 32'b11111111111111110100010000011110;
assign LUT_1[21299] = 32'b11111111111111101101100010011010;
assign LUT_1[21300] = 32'b00000000000000000000011011100100;
assign LUT_1[21301] = 32'b11111111111111111001101101100000;
assign LUT_1[21302] = 32'b11111111111111111100001001110101;
assign LUT_1[21303] = 32'b11111111111111110101011011110001;
assign LUT_1[21304] = 32'b11111111111111110111110000000010;
assign LUT_1[21305] = 32'b11111111111111110001000001111110;
assign LUT_1[21306] = 32'b11111111111111110011011110010011;
assign LUT_1[21307] = 32'b11111111111111101100110000001111;
assign LUT_1[21308] = 32'b11111111111111111111101001011001;
assign LUT_1[21309] = 32'b11111111111111111000111011010101;
assign LUT_1[21310] = 32'b11111111111111111011010111101010;
assign LUT_1[21311] = 32'b11111111111111110100101001100110;
assign LUT_1[21312] = 32'b11111111111111110111101001010100;
assign LUT_1[21313] = 32'b11111111111111110000111011010000;
assign LUT_1[21314] = 32'b11111111111111110011010111100101;
assign LUT_1[21315] = 32'b11111111111111101100101001100001;
assign LUT_1[21316] = 32'b11111111111111111111100010101011;
assign LUT_1[21317] = 32'b11111111111111111000110100100111;
assign LUT_1[21318] = 32'b11111111111111111011010000111100;
assign LUT_1[21319] = 32'b11111111111111110100100010111000;
assign LUT_1[21320] = 32'b11111111111111110110110111001001;
assign LUT_1[21321] = 32'b11111111111111110000001001000101;
assign LUT_1[21322] = 32'b11111111111111110010100101011010;
assign LUT_1[21323] = 32'b11111111111111101011110111010110;
assign LUT_1[21324] = 32'b11111111111111111110110000100000;
assign LUT_1[21325] = 32'b11111111111111111000000010011100;
assign LUT_1[21326] = 32'b11111111111111111010011110110001;
assign LUT_1[21327] = 32'b11111111111111110011110000101101;
assign LUT_1[21328] = 32'b11111111111111111001100100110110;
assign LUT_1[21329] = 32'b11111111111111110010110110110010;
assign LUT_1[21330] = 32'b11111111111111110101010011000111;
assign LUT_1[21331] = 32'b11111111111111101110100101000011;
assign LUT_1[21332] = 32'b00000000000000000001011110001101;
assign LUT_1[21333] = 32'b11111111111111111010110000001001;
assign LUT_1[21334] = 32'b11111111111111111101001100011110;
assign LUT_1[21335] = 32'b11111111111111110110011110011010;
assign LUT_1[21336] = 32'b11111111111111111000110010101011;
assign LUT_1[21337] = 32'b11111111111111110010000100100111;
assign LUT_1[21338] = 32'b11111111111111110100100000111100;
assign LUT_1[21339] = 32'b11111111111111101101110010111000;
assign LUT_1[21340] = 32'b00000000000000000000101100000010;
assign LUT_1[21341] = 32'b11111111111111111001111101111110;
assign LUT_1[21342] = 32'b11111111111111111100011010010011;
assign LUT_1[21343] = 32'b11111111111111110101101100001111;
assign LUT_1[21344] = 32'b11111111111111111000100100010011;
assign LUT_1[21345] = 32'b11111111111111110001110110001111;
assign LUT_1[21346] = 32'b11111111111111110100010010100100;
assign LUT_1[21347] = 32'b11111111111111101101100100100000;
assign LUT_1[21348] = 32'b00000000000000000000011101101010;
assign LUT_1[21349] = 32'b11111111111111111001101111100110;
assign LUT_1[21350] = 32'b11111111111111111100001011111011;
assign LUT_1[21351] = 32'b11111111111111110101011101110111;
assign LUT_1[21352] = 32'b11111111111111110111110010001000;
assign LUT_1[21353] = 32'b11111111111111110001000100000100;
assign LUT_1[21354] = 32'b11111111111111110011100000011001;
assign LUT_1[21355] = 32'b11111111111111101100110010010101;
assign LUT_1[21356] = 32'b11111111111111111111101011011111;
assign LUT_1[21357] = 32'b11111111111111111000111101011011;
assign LUT_1[21358] = 32'b11111111111111111011011001110000;
assign LUT_1[21359] = 32'b11111111111111110100101011101100;
assign LUT_1[21360] = 32'b11111111111111111010011111110101;
assign LUT_1[21361] = 32'b11111111111111110011110001110001;
assign LUT_1[21362] = 32'b11111111111111110110001110000110;
assign LUT_1[21363] = 32'b11111111111111101111100000000010;
assign LUT_1[21364] = 32'b00000000000000000010011001001100;
assign LUT_1[21365] = 32'b11111111111111111011101011001000;
assign LUT_1[21366] = 32'b11111111111111111110000111011101;
assign LUT_1[21367] = 32'b11111111111111110111011001011001;
assign LUT_1[21368] = 32'b11111111111111111001101101101010;
assign LUT_1[21369] = 32'b11111111111111110010111111100110;
assign LUT_1[21370] = 32'b11111111111111110101011011111011;
assign LUT_1[21371] = 32'b11111111111111101110101101110111;
assign LUT_1[21372] = 32'b00000000000000000001100111000001;
assign LUT_1[21373] = 32'b11111111111111111010111000111101;
assign LUT_1[21374] = 32'b11111111111111111101010101010010;
assign LUT_1[21375] = 32'b11111111111111110110100111001110;
assign LUT_1[21376] = 32'b11111111111111111000101011101111;
assign LUT_1[21377] = 32'b11111111111111110001111101101011;
assign LUT_1[21378] = 32'b11111111111111110100011010000000;
assign LUT_1[21379] = 32'b11111111111111101101101011111100;
assign LUT_1[21380] = 32'b00000000000000000000100101000110;
assign LUT_1[21381] = 32'b11111111111111111001110111000010;
assign LUT_1[21382] = 32'b11111111111111111100010011010111;
assign LUT_1[21383] = 32'b11111111111111110101100101010011;
assign LUT_1[21384] = 32'b11111111111111110111111001100100;
assign LUT_1[21385] = 32'b11111111111111110001001011100000;
assign LUT_1[21386] = 32'b11111111111111110011100111110101;
assign LUT_1[21387] = 32'b11111111111111101100111001110001;
assign LUT_1[21388] = 32'b11111111111111111111110010111011;
assign LUT_1[21389] = 32'b11111111111111111001000100110111;
assign LUT_1[21390] = 32'b11111111111111111011100001001100;
assign LUT_1[21391] = 32'b11111111111111110100110011001000;
assign LUT_1[21392] = 32'b11111111111111111010100111010001;
assign LUT_1[21393] = 32'b11111111111111110011111001001101;
assign LUT_1[21394] = 32'b11111111111111110110010101100010;
assign LUT_1[21395] = 32'b11111111111111101111100111011110;
assign LUT_1[21396] = 32'b00000000000000000010100000101000;
assign LUT_1[21397] = 32'b11111111111111111011110010100100;
assign LUT_1[21398] = 32'b11111111111111111110001110111001;
assign LUT_1[21399] = 32'b11111111111111110111100000110101;
assign LUT_1[21400] = 32'b11111111111111111001110101000110;
assign LUT_1[21401] = 32'b11111111111111110011000111000010;
assign LUT_1[21402] = 32'b11111111111111110101100011010111;
assign LUT_1[21403] = 32'b11111111111111101110110101010011;
assign LUT_1[21404] = 32'b00000000000000000001101110011101;
assign LUT_1[21405] = 32'b11111111111111111011000000011001;
assign LUT_1[21406] = 32'b11111111111111111101011100101110;
assign LUT_1[21407] = 32'b11111111111111110110101110101010;
assign LUT_1[21408] = 32'b11111111111111111001100110101110;
assign LUT_1[21409] = 32'b11111111111111110010111000101010;
assign LUT_1[21410] = 32'b11111111111111110101010100111111;
assign LUT_1[21411] = 32'b11111111111111101110100110111011;
assign LUT_1[21412] = 32'b00000000000000000001100000000101;
assign LUT_1[21413] = 32'b11111111111111111010110010000001;
assign LUT_1[21414] = 32'b11111111111111111101001110010110;
assign LUT_1[21415] = 32'b11111111111111110110100000010010;
assign LUT_1[21416] = 32'b11111111111111111000110100100011;
assign LUT_1[21417] = 32'b11111111111111110010000110011111;
assign LUT_1[21418] = 32'b11111111111111110100100010110100;
assign LUT_1[21419] = 32'b11111111111111101101110100110000;
assign LUT_1[21420] = 32'b00000000000000000000101101111010;
assign LUT_1[21421] = 32'b11111111111111111001111111110110;
assign LUT_1[21422] = 32'b11111111111111111100011100001011;
assign LUT_1[21423] = 32'b11111111111111110101101110000111;
assign LUT_1[21424] = 32'b11111111111111111011100010010000;
assign LUT_1[21425] = 32'b11111111111111110100110100001100;
assign LUT_1[21426] = 32'b11111111111111110111010000100001;
assign LUT_1[21427] = 32'b11111111111111110000100010011101;
assign LUT_1[21428] = 32'b00000000000000000011011011100111;
assign LUT_1[21429] = 32'b11111111111111111100101101100011;
assign LUT_1[21430] = 32'b11111111111111111111001001111000;
assign LUT_1[21431] = 32'b11111111111111111000011011110100;
assign LUT_1[21432] = 32'b11111111111111111010110000000101;
assign LUT_1[21433] = 32'b11111111111111110100000010000001;
assign LUT_1[21434] = 32'b11111111111111110110011110010110;
assign LUT_1[21435] = 32'b11111111111111101111110000010010;
assign LUT_1[21436] = 32'b00000000000000000010101001011100;
assign LUT_1[21437] = 32'b11111111111111111011111011011000;
assign LUT_1[21438] = 32'b11111111111111111110010111101101;
assign LUT_1[21439] = 32'b11111111111111110111101001101001;
assign LUT_1[21440] = 32'b11111111111111111010101001010111;
assign LUT_1[21441] = 32'b11111111111111110011111011010011;
assign LUT_1[21442] = 32'b11111111111111110110010111101000;
assign LUT_1[21443] = 32'b11111111111111101111101001100100;
assign LUT_1[21444] = 32'b00000000000000000010100010101110;
assign LUT_1[21445] = 32'b11111111111111111011110100101010;
assign LUT_1[21446] = 32'b11111111111111111110010000111111;
assign LUT_1[21447] = 32'b11111111111111110111100010111011;
assign LUT_1[21448] = 32'b11111111111111111001110111001100;
assign LUT_1[21449] = 32'b11111111111111110011001001001000;
assign LUT_1[21450] = 32'b11111111111111110101100101011101;
assign LUT_1[21451] = 32'b11111111111111101110110111011001;
assign LUT_1[21452] = 32'b00000000000000000001110000100011;
assign LUT_1[21453] = 32'b11111111111111111011000010011111;
assign LUT_1[21454] = 32'b11111111111111111101011110110100;
assign LUT_1[21455] = 32'b11111111111111110110110000110000;
assign LUT_1[21456] = 32'b11111111111111111100100100111001;
assign LUT_1[21457] = 32'b11111111111111110101110110110101;
assign LUT_1[21458] = 32'b11111111111111111000010011001010;
assign LUT_1[21459] = 32'b11111111111111110001100101000110;
assign LUT_1[21460] = 32'b00000000000000000100011110010000;
assign LUT_1[21461] = 32'b11111111111111111101110000001100;
assign LUT_1[21462] = 32'b00000000000000000000001100100001;
assign LUT_1[21463] = 32'b11111111111111111001011110011101;
assign LUT_1[21464] = 32'b11111111111111111011110010101110;
assign LUT_1[21465] = 32'b11111111111111110101000100101010;
assign LUT_1[21466] = 32'b11111111111111110111100000111111;
assign LUT_1[21467] = 32'b11111111111111110000110010111011;
assign LUT_1[21468] = 32'b00000000000000000011101100000101;
assign LUT_1[21469] = 32'b11111111111111111100111110000001;
assign LUT_1[21470] = 32'b11111111111111111111011010010110;
assign LUT_1[21471] = 32'b11111111111111111000101100010010;
assign LUT_1[21472] = 32'b11111111111111111011100100010110;
assign LUT_1[21473] = 32'b11111111111111110100110110010010;
assign LUT_1[21474] = 32'b11111111111111110111010010100111;
assign LUT_1[21475] = 32'b11111111111111110000100100100011;
assign LUT_1[21476] = 32'b00000000000000000011011101101101;
assign LUT_1[21477] = 32'b11111111111111111100101111101001;
assign LUT_1[21478] = 32'b11111111111111111111001011111110;
assign LUT_1[21479] = 32'b11111111111111111000011101111010;
assign LUT_1[21480] = 32'b11111111111111111010110010001011;
assign LUT_1[21481] = 32'b11111111111111110100000100000111;
assign LUT_1[21482] = 32'b11111111111111110110100000011100;
assign LUT_1[21483] = 32'b11111111111111101111110010011000;
assign LUT_1[21484] = 32'b00000000000000000010101011100010;
assign LUT_1[21485] = 32'b11111111111111111011111101011110;
assign LUT_1[21486] = 32'b11111111111111111110011001110011;
assign LUT_1[21487] = 32'b11111111111111110111101011101111;
assign LUT_1[21488] = 32'b11111111111111111101011111111000;
assign LUT_1[21489] = 32'b11111111111111110110110001110100;
assign LUT_1[21490] = 32'b11111111111111111001001110001001;
assign LUT_1[21491] = 32'b11111111111111110010100000000101;
assign LUT_1[21492] = 32'b00000000000000000101011001001111;
assign LUT_1[21493] = 32'b11111111111111111110101011001011;
assign LUT_1[21494] = 32'b00000000000000000001000111100000;
assign LUT_1[21495] = 32'b11111111111111111010011001011100;
assign LUT_1[21496] = 32'b11111111111111111100101101101101;
assign LUT_1[21497] = 32'b11111111111111110101111111101001;
assign LUT_1[21498] = 32'b11111111111111111000011011111110;
assign LUT_1[21499] = 32'b11111111111111110001101101111010;
assign LUT_1[21500] = 32'b00000000000000000100100111000100;
assign LUT_1[21501] = 32'b11111111111111111101111001000000;
assign LUT_1[21502] = 32'b00000000000000000000010101010101;
assign LUT_1[21503] = 32'b11111111111111111001100111010001;
assign LUT_1[21504] = 32'b00000000000000000100011111110011;
assign LUT_1[21505] = 32'b11111111111111111101110001101111;
assign LUT_1[21506] = 32'b00000000000000000000001110000100;
assign LUT_1[21507] = 32'b11111111111111111001100000000000;
assign LUT_1[21508] = 32'b00000000000000001100011001001010;
assign LUT_1[21509] = 32'b00000000000000000101101011000110;
assign LUT_1[21510] = 32'b00000000000000001000000111011011;
assign LUT_1[21511] = 32'b00000000000000000001011001010111;
assign LUT_1[21512] = 32'b00000000000000000011101101101000;
assign LUT_1[21513] = 32'b11111111111111111100111111100100;
assign LUT_1[21514] = 32'b11111111111111111111011011111001;
assign LUT_1[21515] = 32'b11111111111111111000101101110101;
assign LUT_1[21516] = 32'b00000000000000001011100110111111;
assign LUT_1[21517] = 32'b00000000000000000100111000111011;
assign LUT_1[21518] = 32'b00000000000000000111010101010000;
assign LUT_1[21519] = 32'b00000000000000000000100111001100;
assign LUT_1[21520] = 32'b00000000000000000110011011010101;
assign LUT_1[21521] = 32'b11111111111111111111101101010001;
assign LUT_1[21522] = 32'b00000000000000000010001001100110;
assign LUT_1[21523] = 32'b11111111111111111011011011100010;
assign LUT_1[21524] = 32'b00000000000000001110010100101100;
assign LUT_1[21525] = 32'b00000000000000000111100110101000;
assign LUT_1[21526] = 32'b00000000000000001010000010111101;
assign LUT_1[21527] = 32'b00000000000000000011010100111001;
assign LUT_1[21528] = 32'b00000000000000000101101001001010;
assign LUT_1[21529] = 32'b11111111111111111110111011000110;
assign LUT_1[21530] = 32'b00000000000000000001010111011011;
assign LUT_1[21531] = 32'b11111111111111111010101001010111;
assign LUT_1[21532] = 32'b00000000000000001101100010100001;
assign LUT_1[21533] = 32'b00000000000000000110110100011101;
assign LUT_1[21534] = 32'b00000000000000001001010000110010;
assign LUT_1[21535] = 32'b00000000000000000010100010101110;
assign LUT_1[21536] = 32'b00000000000000000101011010110010;
assign LUT_1[21537] = 32'b11111111111111111110101100101110;
assign LUT_1[21538] = 32'b00000000000000000001001001000011;
assign LUT_1[21539] = 32'b11111111111111111010011010111111;
assign LUT_1[21540] = 32'b00000000000000001101010100001001;
assign LUT_1[21541] = 32'b00000000000000000110100110000101;
assign LUT_1[21542] = 32'b00000000000000001001000010011010;
assign LUT_1[21543] = 32'b00000000000000000010010100010110;
assign LUT_1[21544] = 32'b00000000000000000100101000100111;
assign LUT_1[21545] = 32'b11111111111111111101111010100011;
assign LUT_1[21546] = 32'b00000000000000000000010110111000;
assign LUT_1[21547] = 32'b11111111111111111001101000110100;
assign LUT_1[21548] = 32'b00000000000000001100100001111110;
assign LUT_1[21549] = 32'b00000000000000000101110011111010;
assign LUT_1[21550] = 32'b00000000000000001000010000001111;
assign LUT_1[21551] = 32'b00000000000000000001100010001011;
assign LUT_1[21552] = 32'b00000000000000000111010110010100;
assign LUT_1[21553] = 32'b00000000000000000000101000010000;
assign LUT_1[21554] = 32'b00000000000000000011000100100101;
assign LUT_1[21555] = 32'b11111111111111111100010110100001;
assign LUT_1[21556] = 32'b00000000000000001111001111101011;
assign LUT_1[21557] = 32'b00000000000000001000100001100111;
assign LUT_1[21558] = 32'b00000000000000001010111101111100;
assign LUT_1[21559] = 32'b00000000000000000100001111111000;
assign LUT_1[21560] = 32'b00000000000000000110100100001001;
assign LUT_1[21561] = 32'b11111111111111111111110110000101;
assign LUT_1[21562] = 32'b00000000000000000010010010011010;
assign LUT_1[21563] = 32'b11111111111111111011100100010110;
assign LUT_1[21564] = 32'b00000000000000001110011101100000;
assign LUT_1[21565] = 32'b00000000000000000111101111011100;
assign LUT_1[21566] = 32'b00000000000000001010001011110001;
assign LUT_1[21567] = 32'b00000000000000000011011101101101;
assign LUT_1[21568] = 32'b00000000000000000110011101011011;
assign LUT_1[21569] = 32'b11111111111111111111101111010111;
assign LUT_1[21570] = 32'b00000000000000000010001011101100;
assign LUT_1[21571] = 32'b11111111111111111011011101101000;
assign LUT_1[21572] = 32'b00000000000000001110010110110010;
assign LUT_1[21573] = 32'b00000000000000000111101000101110;
assign LUT_1[21574] = 32'b00000000000000001010000101000011;
assign LUT_1[21575] = 32'b00000000000000000011010110111111;
assign LUT_1[21576] = 32'b00000000000000000101101011010000;
assign LUT_1[21577] = 32'b11111111111111111110111101001100;
assign LUT_1[21578] = 32'b00000000000000000001011001100001;
assign LUT_1[21579] = 32'b11111111111111111010101011011101;
assign LUT_1[21580] = 32'b00000000000000001101100100100111;
assign LUT_1[21581] = 32'b00000000000000000110110110100011;
assign LUT_1[21582] = 32'b00000000000000001001010010111000;
assign LUT_1[21583] = 32'b00000000000000000010100100110100;
assign LUT_1[21584] = 32'b00000000000000001000011000111101;
assign LUT_1[21585] = 32'b00000000000000000001101010111001;
assign LUT_1[21586] = 32'b00000000000000000100000111001110;
assign LUT_1[21587] = 32'b11111111111111111101011001001010;
assign LUT_1[21588] = 32'b00000000000000010000010010010100;
assign LUT_1[21589] = 32'b00000000000000001001100100010000;
assign LUT_1[21590] = 32'b00000000000000001100000000100101;
assign LUT_1[21591] = 32'b00000000000000000101010010100001;
assign LUT_1[21592] = 32'b00000000000000000111100110110010;
assign LUT_1[21593] = 32'b00000000000000000000111000101110;
assign LUT_1[21594] = 32'b00000000000000000011010101000011;
assign LUT_1[21595] = 32'b11111111111111111100100110111111;
assign LUT_1[21596] = 32'b00000000000000001111100000001001;
assign LUT_1[21597] = 32'b00000000000000001000110010000101;
assign LUT_1[21598] = 32'b00000000000000001011001110011010;
assign LUT_1[21599] = 32'b00000000000000000100100000010110;
assign LUT_1[21600] = 32'b00000000000000000111011000011010;
assign LUT_1[21601] = 32'b00000000000000000000101010010110;
assign LUT_1[21602] = 32'b00000000000000000011000110101011;
assign LUT_1[21603] = 32'b11111111111111111100011000100111;
assign LUT_1[21604] = 32'b00000000000000001111010001110001;
assign LUT_1[21605] = 32'b00000000000000001000100011101101;
assign LUT_1[21606] = 32'b00000000000000001011000000000010;
assign LUT_1[21607] = 32'b00000000000000000100010001111110;
assign LUT_1[21608] = 32'b00000000000000000110100110001111;
assign LUT_1[21609] = 32'b11111111111111111111111000001011;
assign LUT_1[21610] = 32'b00000000000000000010010100100000;
assign LUT_1[21611] = 32'b11111111111111111011100110011100;
assign LUT_1[21612] = 32'b00000000000000001110011111100110;
assign LUT_1[21613] = 32'b00000000000000000111110001100010;
assign LUT_1[21614] = 32'b00000000000000001010001101110111;
assign LUT_1[21615] = 32'b00000000000000000011011111110011;
assign LUT_1[21616] = 32'b00000000000000001001010011111100;
assign LUT_1[21617] = 32'b00000000000000000010100101111000;
assign LUT_1[21618] = 32'b00000000000000000101000010001101;
assign LUT_1[21619] = 32'b11111111111111111110010100001001;
assign LUT_1[21620] = 32'b00000000000000010001001101010011;
assign LUT_1[21621] = 32'b00000000000000001010011111001111;
assign LUT_1[21622] = 32'b00000000000000001100111011100100;
assign LUT_1[21623] = 32'b00000000000000000110001101100000;
assign LUT_1[21624] = 32'b00000000000000001000100001110001;
assign LUT_1[21625] = 32'b00000000000000000001110011101101;
assign LUT_1[21626] = 32'b00000000000000000100010000000010;
assign LUT_1[21627] = 32'b11111111111111111101100001111110;
assign LUT_1[21628] = 32'b00000000000000010000011011001000;
assign LUT_1[21629] = 32'b00000000000000001001101101000100;
assign LUT_1[21630] = 32'b00000000000000001100001001011001;
assign LUT_1[21631] = 32'b00000000000000000101011011010101;
assign LUT_1[21632] = 32'b00000000000000000111011111110110;
assign LUT_1[21633] = 32'b00000000000000000000110001110010;
assign LUT_1[21634] = 32'b00000000000000000011001110000111;
assign LUT_1[21635] = 32'b11111111111111111100100000000011;
assign LUT_1[21636] = 32'b00000000000000001111011001001101;
assign LUT_1[21637] = 32'b00000000000000001000101011001001;
assign LUT_1[21638] = 32'b00000000000000001011000111011110;
assign LUT_1[21639] = 32'b00000000000000000100011001011010;
assign LUT_1[21640] = 32'b00000000000000000110101101101011;
assign LUT_1[21641] = 32'b11111111111111111111111111100111;
assign LUT_1[21642] = 32'b00000000000000000010011011111100;
assign LUT_1[21643] = 32'b11111111111111111011101101111000;
assign LUT_1[21644] = 32'b00000000000000001110100111000010;
assign LUT_1[21645] = 32'b00000000000000000111111000111110;
assign LUT_1[21646] = 32'b00000000000000001010010101010011;
assign LUT_1[21647] = 32'b00000000000000000011100111001111;
assign LUT_1[21648] = 32'b00000000000000001001011011011000;
assign LUT_1[21649] = 32'b00000000000000000010101101010100;
assign LUT_1[21650] = 32'b00000000000000000101001001101001;
assign LUT_1[21651] = 32'b11111111111111111110011011100101;
assign LUT_1[21652] = 32'b00000000000000010001010100101111;
assign LUT_1[21653] = 32'b00000000000000001010100110101011;
assign LUT_1[21654] = 32'b00000000000000001101000011000000;
assign LUT_1[21655] = 32'b00000000000000000110010100111100;
assign LUT_1[21656] = 32'b00000000000000001000101001001101;
assign LUT_1[21657] = 32'b00000000000000000001111011001001;
assign LUT_1[21658] = 32'b00000000000000000100010111011110;
assign LUT_1[21659] = 32'b11111111111111111101101001011010;
assign LUT_1[21660] = 32'b00000000000000010000100010100100;
assign LUT_1[21661] = 32'b00000000000000001001110100100000;
assign LUT_1[21662] = 32'b00000000000000001100010000110101;
assign LUT_1[21663] = 32'b00000000000000000101100010110001;
assign LUT_1[21664] = 32'b00000000000000001000011010110101;
assign LUT_1[21665] = 32'b00000000000000000001101100110001;
assign LUT_1[21666] = 32'b00000000000000000100001001000110;
assign LUT_1[21667] = 32'b11111111111111111101011011000010;
assign LUT_1[21668] = 32'b00000000000000010000010100001100;
assign LUT_1[21669] = 32'b00000000000000001001100110001000;
assign LUT_1[21670] = 32'b00000000000000001100000010011101;
assign LUT_1[21671] = 32'b00000000000000000101010100011001;
assign LUT_1[21672] = 32'b00000000000000000111101000101010;
assign LUT_1[21673] = 32'b00000000000000000000111010100110;
assign LUT_1[21674] = 32'b00000000000000000011010110111011;
assign LUT_1[21675] = 32'b11111111111111111100101000110111;
assign LUT_1[21676] = 32'b00000000000000001111100010000001;
assign LUT_1[21677] = 32'b00000000000000001000110011111101;
assign LUT_1[21678] = 32'b00000000000000001011010000010010;
assign LUT_1[21679] = 32'b00000000000000000100100010001110;
assign LUT_1[21680] = 32'b00000000000000001010010110010111;
assign LUT_1[21681] = 32'b00000000000000000011101000010011;
assign LUT_1[21682] = 32'b00000000000000000110000100101000;
assign LUT_1[21683] = 32'b11111111111111111111010110100100;
assign LUT_1[21684] = 32'b00000000000000010010001111101110;
assign LUT_1[21685] = 32'b00000000000000001011100001101010;
assign LUT_1[21686] = 32'b00000000000000001101111101111111;
assign LUT_1[21687] = 32'b00000000000000000111001111111011;
assign LUT_1[21688] = 32'b00000000000000001001100100001100;
assign LUT_1[21689] = 32'b00000000000000000010110110001000;
assign LUT_1[21690] = 32'b00000000000000000101010010011101;
assign LUT_1[21691] = 32'b11111111111111111110100100011001;
assign LUT_1[21692] = 32'b00000000000000010001011101100011;
assign LUT_1[21693] = 32'b00000000000000001010101111011111;
assign LUT_1[21694] = 32'b00000000000000001101001011110100;
assign LUT_1[21695] = 32'b00000000000000000110011101110000;
assign LUT_1[21696] = 32'b00000000000000001001011101011110;
assign LUT_1[21697] = 32'b00000000000000000010101111011010;
assign LUT_1[21698] = 32'b00000000000000000101001011101111;
assign LUT_1[21699] = 32'b11111111111111111110011101101011;
assign LUT_1[21700] = 32'b00000000000000010001010110110101;
assign LUT_1[21701] = 32'b00000000000000001010101000110001;
assign LUT_1[21702] = 32'b00000000000000001101000101000110;
assign LUT_1[21703] = 32'b00000000000000000110010111000010;
assign LUT_1[21704] = 32'b00000000000000001000101011010011;
assign LUT_1[21705] = 32'b00000000000000000001111101001111;
assign LUT_1[21706] = 32'b00000000000000000100011001100100;
assign LUT_1[21707] = 32'b11111111111111111101101011100000;
assign LUT_1[21708] = 32'b00000000000000010000100100101010;
assign LUT_1[21709] = 32'b00000000000000001001110110100110;
assign LUT_1[21710] = 32'b00000000000000001100010010111011;
assign LUT_1[21711] = 32'b00000000000000000101100100110111;
assign LUT_1[21712] = 32'b00000000000000001011011001000000;
assign LUT_1[21713] = 32'b00000000000000000100101010111100;
assign LUT_1[21714] = 32'b00000000000000000111000111010001;
assign LUT_1[21715] = 32'b00000000000000000000011001001101;
assign LUT_1[21716] = 32'b00000000000000010011010010010111;
assign LUT_1[21717] = 32'b00000000000000001100100100010011;
assign LUT_1[21718] = 32'b00000000000000001111000000101000;
assign LUT_1[21719] = 32'b00000000000000001000010010100100;
assign LUT_1[21720] = 32'b00000000000000001010100110110101;
assign LUT_1[21721] = 32'b00000000000000000011111000110001;
assign LUT_1[21722] = 32'b00000000000000000110010101000110;
assign LUT_1[21723] = 32'b11111111111111111111100111000010;
assign LUT_1[21724] = 32'b00000000000000010010100000001100;
assign LUT_1[21725] = 32'b00000000000000001011110010001000;
assign LUT_1[21726] = 32'b00000000000000001110001110011101;
assign LUT_1[21727] = 32'b00000000000000000111100000011001;
assign LUT_1[21728] = 32'b00000000000000001010011000011101;
assign LUT_1[21729] = 32'b00000000000000000011101010011001;
assign LUT_1[21730] = 32'b00000000000000000110000110101110;
assign LUT_1[21731] = 32'b11111111111111111111011000101010;
assign LUT_1[21732] = 32'b00000000000000010010010001110100;
assign LUT_1[21733] = 32'b00000000000000001011100011110000;
assign LUT_1[21734] = 32'b00000000000000001110000000000101;
assign LUT_1[21735] = 32'b00000000000000000111010010000001;
assign LUT_1[21736] = 32'b00000000000000001001100110010010;
assign LUT_1[21737] = 32'b00000000000000000010111000001110;
assign LUT_1[21738] = 32'b00000000000000000101010100100011;
assign LUT_1[21739] = 32'b11111111111111111110100110011111;
assign LUT_1[21740] = 32'b00000000000000010001011111101001;
assign LUT_1[21741] = 32'b00000000000000001010110001100101;
assign LUT_1[21742] = 32'b00000000000000001101001101111010;
assign LUT_1[21743] = 32'b00000000000000000110011111110110;
assign LUT_1[21744] = 32'b00000000000000001100010011111111;
assign LUT_1[21745] = 32'b00000000000000000101100101111011;
assign LUT_1[21746] = 32'b00000000000000001000000010010000;
assign LUT_1[21747] = 32'b00000000000000000001010100001100;
assign LUT_1[21748] = 32'b00000000000000010100001101010110;
assign LUT_1[21749] = 32'b00000000000000001101011111010010;
assign LUT_1[21750] = 32'b00000000000000001111111011100111;
assign LUT_1[21751] = 32'b00000000000000001001001101100011;
assign LUT_1[21752] = 32'b00000000000000001011100001110100;
assign LUT_1[21753] = 32'b00000000000000000100110011110000;
assign LUT_1[21754] = 32'b00000000000000000111010000000101;
assign LUT_1[21755] = 32'b00000000000000000000100010000001;
assign LUT_1[21756] = 32'b00000000000000010011011011001011;
assign LUT_1[21757] = 32'b00000000000000001100101101000111;
assign LUT_1[21758] = 32'b00000000000000001111001001011100;
assign LUT_1[21759] = 32'b00000000000000001000011011011000;
assign LUT_1[21760] = 32'b00000000000000000010010011111111;
assign LUT_1[21761] = 32'b11111111111111111011100101111011;
assign LUT_1[21762] = 32'b11111111111111111110000010010000;
assign LUT_1[21763] = 32'b11111111111111110111010100001100;
assign LUT_1[21764] = 32'b00000000000000001010001101010110;
assign LUT_1[21765] = 32'b00000000000000000011011111010010;
assign LUT_1[21766] = 32'b00000000000000000101111011100111;
assign LUT_1[21767] = 32'b11111111111111111111001101100011;
assign LUT_1[21768] = 32'b00000000000000000001100001110100;
assign LUT_1[21769] = 32'b11111111111111111010110011110000;
assign LUT_1[21770] = 32'b11111111111111111101010000000101;
assign LUT_1[21771] = 32'b11111111111111110110100010000001;
assign LUT_1[21772] = 32'b00000000000000001001011011001011;
assign LUT_1[21773] = 32'b00000000000000000010101101000111;
assign LUT_1[21774] = 32'b00000000000000000101001001011100;
assign LUT_1[21775] = 32'b11111111111111111110011011011000;
assign LUT_1[21776] = 32'b00000000000000000100001111100001;
assign LUT_1[21777] = 32'b11111111111111111101100001011101;
assign LUT_1[21778] = 32'b11111111111111111111111101110010;
assign LUT_1[21779] = 32'b11111111111111111001001111101110;
assign LUT_1[21780] = 32'b00000000000000001100001000111000;
assign LUT_1[21781] = 32'b00000000000000000101011010110100;
assign LUT_1[21782] = 32'b00000000000000000111110111001001;
assign LUT_1[21783] = 32'b00000000000000000001001001000101;
assign LUT_1[21784] = 32'b00000000000000000011011101010110;
assign LUT_1[21785] = 32'b11111111111111111100101111010010;
assign LUT_1[21786] = 32'b11111111111111111111001011100111;
assign LUT_1[21787] = 32'b11111111111111111000011101100011;
assign LUT_1[21788] = 32'b00000000000000001011010110101101;
assign LUT_1[21789] = 32'b00000000000000000100101000101001;
assign LUT_1[21790] = 32'b00000000000000000111000100111110;
assign LUT_1[21791] = 32'b00000000000000000000010110111010;
assign LUT_1[21792] = 32'b00000000000000000011001110111110;
assign LUT_1[21793] = 32'b11111111111111111100100000111010;
assign LUT_1[21794] = 32'b11111111111111111110111101001111;
assign LUT_1[21795] = 32'b11111111111111111000001111001011;
assign LUT_1[21796] = 32'b00000000000000001011001000010101;
assign LUT_1[21797] = 32'b00000000000000000100011010010001;
assign LUT_1[21798] = 32'b00000000000000000110110110100110;
assign LUT_1[21799] = 32'b00000000000000000000001000100010;
assign LUT_1[21800] = 32'b00000000000000000010011100110011;
assign LUT_1[21801] = 32'b11111111111111111011101110101111;
assign LUT_1[21802] = 32'b11111111111111111110001011000100;
assign LUT_1[21803] = 32'b11111111111111110111011101000000;
assign LUT_1[21804] = 32'b00000000000000001010010110001010;
assign LUT_1[21805] = 32'b00000000000000000011101000000110;
assign LUT_1[21806] = 32'b00000000000000000110000100011011;
assign LUT_1[21807] = 32'b11111111111111111111010110010111;
assign LUT_1[21808] = 32'b00000000000000000101001010100000;
assign LUT_1[21809] = 32'b11111111111111111110011100011100;
assign LUT_1[21810] = 32'b00000000000000000000111000110001;
assign LUT_1[21811] = 32'b11111111111111111010001010101101;
assign LUT_1[21812] = 32'b00000000000000001101000011110111;
assign LUT_1[21813] = 32'b00000000000000000110010101110011;
assign LUT_1[21814] = 32'b00000000000000001000110010001000;
assign LUT_1[21815] = 32'b00000000000000000010000100000100;
assign LUT_1[21816] = 32'b00000000000000000100011000010101;
assign LUT_1[21817] = 32'b11111111111111111101101010010001;
assign LUT_1[21818] = 32'b00000000000000000000000110100110;
assign LUT_1[21819] = 32'b11111111111111111001011000100010;
assign LUT_1[21820] = 32'b00000000000000001100010001101100;
assign LUT_1[21821] = 32'b00000000000000000101100011101000;
assign LUT_1[21822] = 32'b00000000000000000111111111111101;
assign LUT_1[21823] = 32'b00000000000000000001010001111001;
assign LUT_1[21824] = 32'b00000000000000000100010001100111;
assign LUT_1[21825] = 32'b11111111111111111101100011100011;
assign LUT_1[21826] = 32'b11111111111111111111111111111000;
assign LUT_1[21827] = 32'b11111111111111111001010001110100;
assign LUT_1[21828] = 32'b00000000000000001100001010111110;
assign LUT_1[21829] = 32'b00000000000000000101011100111010;
assign LUT_1[21830] = 32'b00000000000000000111111001001111;
assign LUT_1[21831] = 32'b00000000000000000001001011001011;
assign LUT_1[21832] = 32'b00000000000000000011011111011100;
assign LUT_1[21833] = 32'b11111111111111111100110001011000;
assign LUT_1[21834] = 32'b11111111111111111111001101101101;
assign LUT_1[21835] = 32'b11111111111111111000011111101001;
assign LUT_1[21836] = 32'b00000000000000001011011000110011;
assign LUT_1[21837] = 32'b00000000000000000100101010101111;
assign LUT_1[21838] = 32'b00000000000000000111000111000100;
assign LUT_1[21839] = 32'b00000000000000000000011001000000;
assign LUT_1[21840] = 32'b00000000000000000110001101001001;
assign LUT_1[21841] = 32'b11111111111111111111011111000101;
assign LUT_1[21842] = 32'b00000000000000000001111011011010;
assign LUT_1[21843] = 32'b11111111111111111011001101010110;
assign LUT_1[21844] = 32'b00000000000000001110000110100000;
assign LUT_1[21845] = 32'b00000000000000000111011000011100;
assign LUT_1[21846] = 32'b00000000000000001001110100110001;
assign LUT_1[21847] = 32'b00000000000000000011000110101101;
assign LUT_1[21848] = 32'b00000000000000000101011010111110;
assign LUT_1[21849] = 32'b11111111111111111110101100111010;
assign LUT_1[21850] = 32'b00000000000000000001001001001111;
assign LUT_1[21851] = 32'b11111111111111111010011011001011;
assign LUT_1[21852] = 32'b00000000000000001101010100010101;
assign LUT_1[21853] = 32'b00000000000000000110100110010001;
assign LUT_1[21854] = 32'b00000000000000001001000010100110;
assign LUT_1[21855] = 32'b00000000000000000010010100100010;
assign LUT_1[21856] = 32'b00000000000000000101001100100110;
assign LUT_1[21857] = 32'b11111111111111111110011110100010;
assign LUT_1[21858] = 32'b00000000000000000000111010110111;
assign LUT_1[21859] = 32'b11111111111111111010001100110011;
assign LUT_1[21860] = 32'b00000000000000001101000101111101;
assign LUT_1[21861] = 32'b00000000000000000110010111111001;
assign LUT_1[21862] = 32'b00000000000000001000110100001110;
assign LUT_1[21863] = 32'b00000000000000000010000110001010;
assign LUT_1[21864] = 32'b00000000000000000100011010011011;
assign LUT_1[21865] = 32'b11111111111111111101101100010111;
assign LUT_1[21866] = 32'b00000000000000000000001000101100;
assign LUT_1[21867] = 32'b11111111111111111001011010101000;
assign LUT_1[21868] = 32'b00000000000000001100010011110010;
assign LUT_1[21869] = 32'b00000000000000000101100101101110;
assign LUT_1[21870] = 32'b00000000000000001000000010000011;
assign LUT_1[21871] = 32'b00000000000000000001010011111111;
assign LUT_1[21872] = 32'b00000000000000000111001000001000;
assign LUT_1[21873] = 32'b00000000000000000000011010000100;
assign LUT_1[21874] = 32'b00000000000000000010110110011001;
assign LUT_1[21875] = 32'b11111111111111111100001000010101;
assign LUT_1[21876] = 32'b00000000000000001111000001011111;
assign LUT_1[21877] = 32'b00000000000000001000010011011011;
assign LUT_1[21878] = 32'b00000000000000001010101111110000;
assign LUT_1[21879] = 32'b00000000000000000100000001101100;
assign LUT_1[21880] = 32'b00000000000000000110010101111101;
assign LUT_1[21881] = 32'b11111111111111111111100111111001;
assign LUT_1[21882] = 32'b00000000000000000010000100001110;
assign LUT_1[21883] = 32'b11111111111111111011010110001010;
assign LUT_1[21884] = 32'b00000000000000001110001111010100;
assign LUT_1[21885] = 32'b00000000000000000111100001010000;
assign LUT_1[21886] = 32'b00000000000000001001111101100101;
assign LUT_1[21887] = 32'b00000000000000000011001111100001;
assign LUT_1[21888] = 32'b00000000000000000101010100000010;
assign LUT_1[21889] = 32'b11111111111111111110100101111110;
assign LUT_1[21890] = 32'b00000000000000000001000010010011;
assign LUT_1[21891] = 32'b11111111111111111010010100001111;
assign LUT_1[21892] = 32'b00000000000000001101001101011001;
assign LUT_1[21893] = 32'b00000000000000000110011111010101;
assign LUT_1[21894] = 32'b00000000000000001000111011101010;
assign LUT_1[21895] = 32'b00000000000000000010001101100110;
assign LUT_1[21896] = 32'b00000000000000000100100001110111;
assign LUT_1[21897] = 32'b11111111111111111101110011110011;
assign LUT_1[21898] = 32'b00000000000000000000010000001000;
assign LUT_1[21899] = 32'b11111111111111111001100010000100;
assign LUT_1[21900] = 32'b00000000000000001100011011001110;
assign LUT_1[21901] = 32'b00000000000000000101101101001010;
assign LUT_1[21902] = 32'b00000000000000001000001001011111;
assign LUT_1[21903] = 32'b00000000000000000001011011011011;
assign LUT_1[21904] = 32'b00000000000000000111001111100100;
assign LUT_1[21905] = 32'b00000000000000000000100001100000;
assign LUT_1[21906] = 32'b00000000000000000010111101110101;
assign LUT_1[21907] = 32'b11111111111111111100001111110001;
assign LUT_1[21908] = 32'b00000000000000001111001000111011;
assign LUT_1[21909] = 32'b00000000000000001000011010110111;
assign LUT_1[21910] = 32'b00000000000000001010110111001100;
assign LUT_1[21911] = 32'b00000000000000000100001001001000;
assign LUT_1[21912] = 32'b00000000000000000110011101011001;
assign LUT_1[21913] = 32'b11111111111111111111101111010101;
assign LUT_1[21914] = 32'b00000000000000000010001011101010;
assign LUT_1[21915] = 32'b11111111111111111011011101100110;
assign LUT_1[21916] = 32'b00000000000000001110010110110000;
assign LUT_1[21917] = 32'b00000000000000000111101000101100;
assign LUT_1[21918] = 32'b00000000000000001010000101000001;
assign LUT_1[21919] = 32'b00000000000000000011010110111101;
assign LUT_1[21920] = 32'b00000000000000000110001111000001;
assign LUT_1[21921] = 32'b11111111111111111111100000111101;
assign LUT_1[21922] = 32'b00000000000000000001111101010010;
assign LUT_1[21923] = 32'b11111111111111111011001111001110;
assign LUT_1[21924] = 32'b00000000000000001110001000011000;
assign LUT_1[21925] = 32'b00000000000000000111011010010100;
assign LUT_1[21926] = 32'b00000000000000001001110110101001;
assign LUT_1[21927] = 32'b00000000000000000011001000100101;
assign LUT_1[21928] = 32'b00000000000000000101011100110110;
assign LUT_1[21929] = 32'b11111111111111111110101110110010;
assign LUT_1[21930] = 32'b00000000000000000001001011000111;
assign LUT_1[21931] = 32'b11111111111111111010011101000011;
assign LUT_1[21932] = 32'b00000000000000001101010110001101;
assign LUT_1[21933] = 32'b00000000000000000110101000001001;
assign LUT_1[21934] = 32'b00000000000000001001000100011110;
assign LUT_1[21935] = 32'b00000000000000000010010110011010;
assign LUT_1[21936] = 32'b00000000000000001000001010100011;
assign LUT_1[21937] = 32'b00000000000000000001011100011111;
assign LUT_1[21938] = 32'b00000000000000000011111000110100;
assign LUT_1[21939] = 32'b11111111111111111101001010110000;
assign LUT_1[21940] = 32'b00000000000000010000000011111010;
assign LUT_1[21941] = 32'b00000000000000001001010101110110;
assign LUT_1[21942] = 32'b00000000000000001011110010001011;
assign LUT_1[21943] = 32'b00000000000000000101000100000111;
assign LUT_1[21944] = 32'b00000000000000000111011000011000;
assign LUT_1[21945] = 32'b00000000000000000000101010010100;
assign LUT_1[21946] = 32'b00000000000000000011000110101001;
assign LUT_1[21947] = 32'b11111111111111111100011000100101;
assign LUT_1[21948] = 32'b00000000000000001111010001101111;
assign LUT_1[21949] = 32'b00000000000000001000100011101011;
assign LUT_1[21950] = 32'b00000000000000001011000000000000;
assign LUT_1[21951] = 32'b00000000000000000100010001111100;
assign LUT_1[21952] = 32'b00000000000000000111010001101010;
assign LUT_1[21953] = 32'b00000000000000000000100011100110;
assign LUT_1[21954] = 32'b00000000000000000010111111111011;
assign LUT_1[21955] = 32'b11111111111111111100010001110111;
assign LUT_1[21956] = 32'b00000000000000001111001011000001;
assign LUT_1[21957] = 32'b00000000000000001000011100111101;
assign LUT_1[21958] = 32'b00000000000000001010111001010010;
assign LUT_1[21959] = 32'b00000000000000000100001011001110;
assign LUT_1[21960] = 32'b00000000000000000110011111011111;
assign LUT_1[21961] = 32'b11111111111111111111110001011011;
assign LUT_1[21962] = 32'b00000000000000000010001101110000;
assign LUT_1[21963] = 32'b11111111111111111011011111101100;
assign LUT_1[21964] = 32'b00000000000000001110011000110110;
assign LUT_1[21965] = 32'b00000000000000000111101010110010;
assign LUT_1[21966] = 32'b00000000000000001010000111000111;
assign LUT_1[21967] = 32'b00000000000000000011011001000011;
assign LUT_1[21968] = 32'b00000000000000001001001101001100;
assign LUT_1[21969] = 32'b00000000000000000010011111001000;
assign LUT_1[21970] = 32'b00000000000000000100111011011101;
assign LUT_1[21971] = 32'b11111111111111111110001101011001;
assign LUT_1[21972] = 32'b00000000000000010001000110100011;
assign LUT_1[21973] = 32'b00000000000000001010011000011111;
assign LUT_1[21974] = 32'b00000000000000001100110100110100;
assign LUT_1[21975] = 32'b00000000000000000110000110110000;
assign LUT_1[21976] = 32'b00000000000000001000011011000001;
assign LUT_1[21977] = 32'b00000000000000000001101100111101;
assign LUT_1[21978] = 32'b00000000000000000100001001010010;
assign LUT_1[21979] = 32'b11111111111111111101011011001110;
assign LUT_1[21980] = 32'b00000000000000010000010100011000;
assign LUT_1[21981] = 32'b00000000000000001001100110010100;
assign LUT_1[21982] = 32'b00000000000000001100000010101001;
assign LUT_1[21983] = 32'b00000000000000000101010100100101;
assign LUT_1[21984] = 32'b00000000000000001000001100101001;
assign LUT_1[21985] = 32'b00000000000000000001011110100101;
assign LUT_1[21986] = 32'b00000000000000000011111010111010;
assign LUT_1[21987] = 32'b11111111111111111101001100110110;
assign LUT_1[21988] = 32'b00000000000000010000000110000000;
assign LUT_1[21989] = 32'b00000000000000001001010111111100;
assign LUT_1[21990] = 32'b00000000000000001011110100010001;
assign LUT_1[21991] = 32'b00000000000000000101000110001101;
assign LUT_1[21992] = 32'b00000000000000000111011010011110;
assign LUT_1[21993] = 32'b00000000000000000000101100011010;
assign LUT_1[21994] = 32'b00000000000000000011001000101111;
assign LUT_1[21995] = 32'b11111111111111111100011010101011;
assign LUT_1[21996] = 32'b00000000000000001111010011110101;
assign LUT_1[21997] = 32'b00000000000000001000100101110001;
assign LUT_1[21998] = 32'b00000000000000001011000010000110;
assign LUT_1[21999] = 32'b00000000000000000100010100000010;
assign LUT_1[22000] = 32'b00000000000000001010001000001011;
assign LUT_1[22001] = 32'b00000000000000000011011010000111;
assign LUT_1[22002] = 32'b00000000000000000101110110011100;
assign LUT_1[22003] = 32'b11111111111111111111001000011000;
assign LUT_1[22004] = 32'b00000000000000010010000001100010;
assign LUT_1[22005] = 32'b00000000000000001011010011011110;
assign LUT_1[22006] = 32'b00000000000000001101101111110011;
assign LUT_1[22007] = 32'b00000000000000000111000001101111;
assign LUT_1[22008] = 32'b00000000000000001001010110000000;
assign LUT_1[22009] = 32'b00000000000000000010100111111100;
assign LUT_1[22010] = 32'b00000000000000000101000100010001;
assign LUT_1[22011] = 32'b11111111111111111110010110001101;
assign LUT_1[22012] = 32'b00000000000000010001001111010111;
assign LUT_1[22013] = 32'b00000000000000001010100001010011;
assign LUT_1[22014] = 32'b00000000000000001100111101101000;
assign LUT_1[22015] = 32'b00000000000000000110001111100100;
assign LUT_1[22016] = 32'b11111111111111111110001110010000;
assign LUT_1[22017] = 32'b11111111111111110111100000001100;
assign LUT_1[22018] = 32'b11111111111111111001111100100001;
assign LUT_1[22019] = 32'b11111111111111110011001110011101;
assign LUT_1[22020] = 32'b00000000000000000110000111100111;
assign LUT_1[22021] = 32'b11111111111111111111011001100011;
assign LUT_1[22022] = 32'b00000000000000000001110101111000;
assign LUT_1[22023] = 32'b11111111111111111011000111110100;
assign LUT_1[22024] = 32'b11111111111111111101011100000101;
assign LUT_1[22025] = 32'b11111111111111110110101110000001;
assign LUT_1[22026] = 32'b11111111111111111001001010010110;
assign LUT_1[22027] = 32'b11111111111111110010011100010010;
assign LUT_1[22028] = 32'b00000000000000000101010101011100;
assign LUT_1[22029] = 32'b11111111111111111110100111011000;
assign LUT_1[22030] = 32'b00000000000000000001000011101101;
assign LUT_1[22031] = 32'b11111111111111111010010101101001;
assign LUT_1[22032] = 32'b00000000000000000000001001110010;
assign LUT_1[22033] = 32'b11111111111111111001011011101110;
assign LUT_1[22034] = 32'b11111111111111111011111000000011;
assign LUT_1[22035] = 32'b11111111111111110101001001111111;
assign LUT_1[22036] = 32'b00000000000000001000000011001001;
assign LUT_1[22037] = 32'b00000000000000000001010101000101;
assign LUT_1[22038] = 32'b00000000000000000011110001011010;
assign LUT_1[22039] = 32'b11111111111111111101000011010110;
assign LUT_1[22040] = 32'b11111111111111111111010111100111;
assign LUT_1[22041] = 32'b11111111111111111000101001100011;
assign LUT_1[22042] = 32'b11111111111111111011000101111000;
assign LUT_1[22043] = 32'b11111111111111110100010111110100;
assign LUT_1[22044] = 32'b00000000000000000111010000111110;
assign LUT_1[22045] = 32'b00000000000000000000100010111010;
assign LUT_1[22046] = 32'b00000000000000000010111111001111;
assign LUT_1[22047] = 32'b11111111111111111100010001001011;
assign LUT_1[22048] = 32'b11111111111111111111001001001111;
assign LUT_1[22049] = 32'b11111111111111111000011011001011;
assign LUT_1[22050] = 32'b11111111111111111010110111100000;
assign LUT_1[22051] = 32'b11111111111111110100001001011100;
assign LUT_1[22052] = 32'b00000000000000000111000010100110;
assign LUT_1[22053] = 32'b00000000000000000000010100100010;
assign LUT_1[22054] = 32'b00000000000000000010110000110111;
assign LUT_1[22055] = 32'b11111111111111111100000010110011;
assign LUT_1[22056] = 32'b11111111111111111110010111000100;
assign LUT_1[22057] = 32'b11111111111111110111101001000000;
assign LUT_1[22058] = 32'b11111111111111111010000101010101;
assign LUT_1[22059] = 32'b11111111111111110011010111010001;
assign LUT_1[22060] = 32'b00000000000000000110010000011011;
assign LUT_1[22061] = 32'b11111111111111111111100010010111;
assign LUT_1[22062] = 32'b00000000000000000001111110101100;
assign LUT_1[22063] = 32'b11111111111111111011010000101000;
assign LUT_1[22064] = 32'b00000000000000000001000100110001;
assign LUT_1[22065] = 32'b11111111111111111010010110101101;
assign LUT_1[22066] = 32'b11111111111111111100110011000010;
assign LUT_1[22067] = 32'b11111111111111110110000100111110;
assign LUT_1[22068] = 32'b00000000000000001000111110001000;
assign LUT_1[22069] = 32'b00000000000000000010010000000100;
assign LUT_1[22070] = 32'b00000000000000000100101100011001;
assign LUT_1[22071] = 32'b11111111111111111101111110010101;
assign LUT_1[22072] = 32'b00000000000000000000010010100110;
assign LUT_1[22073] = 32'b11111111111111111001100100100010;
assign LUT_1[22074] = 32'b11111111111111111100000000110111;
assign LUT_1[22075] = 32'b11111111111111110101010010110011;
assign LUT_1[22076] = 32'b00000000000000001000001011111101;
assign LUT_1[22077] = 32'b00000000000000000001011101111001;
assign LUT_1[22078] = 32'b00000000000000000011111010001110;
assign LUT_1[22079] = 32'b11111111111111111101001100001010;
assign LUT_1[22080] = 32'b00000000000000000000001011111000;
assign LUT_1[22081] = 32'b11111111111111111001011101110100;
assign LUT_1[22082] = 32'b11111111111111111011111010001001;
assign LUT_1[22083] = 32'b11111111111111110101001100000101;
assign LUT_1[22084] = 32'b00000000000000001000000101001111;
assign LUT_1[22085] = 32'b00000000000000000001010111001011;
assign LUT_1[22086] = 32'b00000000000000000011110011100000;
assign LUT_1[22087] = 32'b11111111111111111101000101011100;
assign LUT_1[22088] = 32'b11111111111111111111011001101101;
assign LUT_1[22089] = 32'b11111111111111111000101011101001;
assign LUT_1[22090] = 32'b11111111111111111011000111111110;
assign LUT_1[22091] = 32'b11111111111111110100011001111010;
assign LUT_1[22092] = 32'b00000000000000000111010011000100;
assign LUT_1[22093] = 32'b00000000000000000000100101000000;
assign LUT_1[22094] = 32'b00000000000000000011000001010101;
assign LUT_1[22095] = 32'b11111111111111111100010011010001;
assign LUT_1[22096] = 32'b00000000000000000010000111011010;
assign LUT_1[22097] = 32'b11111111111111111011011001010110;
assign LUT_1[22098] = 32'b11111111111111111101110101101011;
assign LUT_1[22099] = 32'b11111111111111110111000111100111;
assign LUT_1[22100] = 32'b00000000000000001010000000110001;
assign LUT_1[22101] = 32'b00000000000000000011010010101101;
assign LUT_1[22102] = 32'b00000000000000000101101111000010;
assign LUT_1[22103] = 32'b11111111111111111111000000111110;
assign LUT_1[22104] = 32'b00000000000000000001010101001111;
assign LUT_1[22105] = 32'b11111111111111111010100111001011;
assign LUT_1[22106] = 32'b11111111111111111101000011100000;
assign LUT_1[22107] = 32'b11111111111111110110010101011100;
assign LUT_1[22108] = 32'b00000000000000001001001110100110;
assign LUT_1[22109] = 32'b00000000000000000010100000100010;
assign LUT_1[22110] = 32'b00000000000000000100111100110111;
assign LUT_1[22111] = 32'b11111111111111111110001110110011;
assign LUT_1[22112] = 32'b00000000000000000001000110110111;
assign LUT_1[22113] = 32'b11111111111111111010011000110011;
assign LUT_1[22114] = 32'b11111111111111111100110101001000;
assign LUT_1[22115] = 32'b11111111111111110110000111000100;
assign LUT_1[22116] = 32'b00000000000000001001000000001110;
assign LUT_1[22117] = 32'b00000000000000000010010010001010;
assign LUT_1[22118] = 32'b00000000000000000100101110011111;
assign LUT_1[22119] = 32'b11111111111111111110000000011011;
assign LUT_1[22120] = 32'b00000000000000000000010100101100;
assign LUT_1[22121] = 32'b11111111111111111001100110101000;
assign LUT_1[22122] = 32'b11111111111111111100000010111101;
assign LUT_1[22123] = 32'b11111111111111110101010100111001;
assign LUT_1[22124] = 32'b00000000000000001000001110000011;
assign LUT_1[22125] = 32'b00000000000000000001011111111111;
assign LUT_1[22126] = 32'b00000000000000000011111100010100;
assign LUT_1[22127] = 32'b11111111111111111101001110010000;
assign LUT_1[22128] = 32'b00000000000000000011000010011001;
assign LUT_1[22129] = 32'b11111111111111111100010100010101;
assign LUT_1[22130] = 32'b11111111111111111110110000101010;
assign LUT_1[22131] = 32'b11111111111111111000000010100110;
assign LUT_1[22132] = 32'b00000000000000001010111011110000;
assign LUT_1[22133] = 32'b00000000000000000100001101101100;
assign LUT_1[22134] = 32'b00000000000000000110101010000001;
assign LUT_1[22135] = 32'b11111111111111111111111011111101;
assign LUT_1[22136] = 32'b00000000000000000010010000001110;
assign LUT_1[22137] = 32'b11111111111111111011100010001010;
assign LUT_1[22138] = 32'b11111111111111111101111110011111;
assign LUT_1[22139] = 32'b11111111111111110111010000011011;
assign LUT_1[22140] = 32'b00000000000000001010001001100101;
assign LUT_1[22141] = 32'b00000000000000000011011011100001;
assign LUT_1[22142] = 32'b00000000000000000101110111110110;
assign LUT_1[22143] = 32'b11111111111111111111001001110010;
assign LUT_1[22144] = 32'b00000000000000000001001110010011;
assign LUT_1[22145] = 32'b11111111111111111010100000001111;
assign LUT_1[22146] = 32'b11111111111111111100111100100100;
assign LUT_1[22147] = 32'b11111111111111110110001110100000;
assign LUT_1[22148] = 32'b00000000000000001001000111101010;
assign LUT_1[22149] = 32'b00000000000000000010011001100110;
assign LUT_1[22150] = 32'b00000000000000000100110101111011;
assign LUT_1[22151] = 32'b11111111111111111110000111110111;
assign LUT_1[22152] = 32'b00000000000000000000011100001000;
assign LUT_1[22153] = 32'b11111111111111111001101110000100;
assign LUT_1[22154] = 32'b11111111111111111100001010011001;
assign LUT_1[22155] = 32'b11111111111111110101011100010101;
assign LUT_1[22156] = 32'b00000000000000001000010101011111;
assign LUT_1[22157] = 32'b00000000000000000001100111011011;
assign LUT_1[22158] = 32'b00000000000000000100000011110000;
assign LUT_1[22159] = 32'b11111111111111111101010101101100;
assign LUT_1[22160] = 32'b00000000000000000011001001110101;
assign LUT_1[22161] = 32'b11111111111111111100011011110001;
assign LUT_1[22162] = 32'b11111111111111111110111000000110;
assign LUT_1[22163] = 32'b11111111111111111000001010000010;
assign LUT_1[22164] = 32'b00000000000000001011000011001100;
assign LUT_1[22165] = 32'b00000000000000000100010101001000;
assign LUT_1[22166] = 32'b00000000000000000110110001011101;
assign LUT_1[22167] = 32'b00000000000000000000000011011001;
assign LUT_1[22168] = 32'b00000000000000000010010111101010;
assign LUT_1[22169] = 32'b11111111111111111011101001100110;
assign LUT_1[22170] = 32'b11111111111111111110000101111011;
assign LUT_1[22171] = 32'b11111111111111110111010111110111;
assign LUT_1[22172] = 32'b00000000000000001010010001000001;
assign LUT_1[22173] = 32'b00000000000000000011100010111101;
assign LUT_1[22174] = 32'b00000000000000000101111111010010;
assign LUT_1[22175] = 32'b11111111111111111111010001001110;
assign LUT_1[22176] = 32'b00000000000000000010001001010010;
assign LUT_1[22177] = 32'b11111111111111111011011011001110;
assign LUT_1[22178] = 32'b11111111111111111101110111100011;
assign LUT_1[22179] = 32'b11111111111111110111001001011111;
assign LUT_1[22180] = 32'b00000000000000001010000010101001;
assign LUT_1[22181] = 32'b00000000000000000011010100100101;
assign LUT_1[22182] = 32'b00000000000000000101110000111010;
assign LUT_1[22183] = 32'b11111111111111111111000010110110;
assign LUT_1[22184] = 32'b00000000000000000001010111000111;
assign LUT_1[22185] = 32'b11111111111111111010101001000011;
assign LUT_1[22186] = 32'b11111111111111111101000101011000;
assign LUT_1[22187] = 32'b11111111111111110110010111010100;
assign LUT_1[22188] = 32'b00000000000000001001010000011110;
assign LUT_1[22189] = 32'b00000000000000000010100010011010;
assign LUT_1[22190] = 32'b00000000000000000100111110101111;
assign LUT_1[22191] = 32'b11111111111111111110010000101011;
assign LUT_1[22192] = 32'b00000000000000000100000100110100;
assign LUT_1[22193] = 32'b11111111111111111101010110110000;
assign LUT_1[22194] = 32'b11111111111111111111110011000101;
assign LUT_1[22195] = 32'b11111111111111111001000101000001;
assign LUT_1[22196] = 32'b00000000000000001011111110001011;
assign LUT_1[22197] = 32'b00000000000000000101010000000111;
assign LUT_1[22198] = 32'b00000000000000000111101100011100;
assign LUT_1[22199] = 32'b00000000000000000000111110011000;
assign LUT_1[22200] = 32'b00000000000000000011010010101001;
assign LUT_1[22201] = 32'b11111111111111111100100100100101;
assign LUT_1[22202] = 32'b11111111111111111111000000111010;
assign LUT_1[22203] = 32'b11111111111111111000010010110110;
assign LUT_1[22204] = 32'b00000000000000001011001100000000;
assign LUT_1[22205] = 32'b00000000000000000100011101111100;
assign LUT_1[22206] = 32'b00000000000000000110111010010001;
assign LUT_1[22207] = 32'b00000000000000000000001100001101;
assign LUT_1[22208] = 32'b00000000000000000011001011111011;
assign LUT_1[22209] = 32'b11111111111111111100011101110111;
assign LUT_1[22210] = 32'b11111111111111111110111010001100;
assign LUT_1[22211] = 32'b11111111111111111000001100001000;
assign LUT_1[22212] = 32'b00000000000000001011000101010010;
assign LUT_1[22213] = 32'b00000000000000000100010111001110;
assign LUT_1[22214] = 32'b00000000000000000110110011100011;
assign LUT_1[22215] = 32'b00000000000000000000000101011111;
assign LUT_1[22216] = 32'b00000000000000000010011001110000;
assign LUT_1[22217] = 32'b11111111111111111011101011101100;
assign LUT_1[22218] = 32'b11111111111111111110001000000001;
assign LUT_1[22219] = 32'b11111111111111110111011001111101;
assign LUT_1[22220] = 32'b00000000000000001010010011000111;
assign LUT_1[22221] = 32'b00000000000000000011100101000011;
assign LUT_1[22222] = 32'b00000000000000000110000001011000;
assign LUT_1[22223] = 32'b11111111111111111111010011010100;
assign LUT_1[22224] = 32'b00000000000000000101000111011101;
assign LUT_1[22225] = 32'b11111111111111111110011001011001;
assign LUT_1[22226] = 32'b00000000000000000000110101101110;
assign LUT_1[22227] = 32'b11111111111111111010000111101010;
assign LUT_1[22228] = 32'b00000000000000001101000000110100;
assign LUT_1[22229] = 32'b00000000000000000110010010110000;
assign LUT_1[22230] = 32'b00000000000000001000101111000101;
assign LUT_1[22231] = 32'b00000000000000000010000001000001;
assign LUT_1[22232] = 32'b00000000000000000100010101010010;
assign LUT_1[22233] = 32'b11111111111111111101100111001110;
assign LUT_1[22234] = 32'b00000000000000000000000011100011;
assign LUT_1[22235] = 32'b11111111111111111001010101011111;
assign LUT_1[22236] = 32'b00000000000000001100001110101001;
assign LUT_1[22237] = 32'b00000000000000000101100000100101;
assign LUT_1[22238] = 32'b00000000000000000111111100111010;
assign LUT_1[22239] = 32'b00000000000000000001001110110110;
assign LUT_1[22240] = 32'b00000000000000000100000110111010;
assign LUT_1[22241] = 32'b11111111111111111101011000110110;
assign LUT_1[22242] = 32'b11111111111111111111110101001011;
assign LUT_1[22243] = 32'b11111111111111111001000111000111;
assign LUT_1[22244] = 32'b00000000000000001100000000010001;
assign LUT_1[22245] = 32'b00000000000000000101010010001101;
assign LUT_1[22246] = 32'b00000000000000000111101110100010;
assign LUT_1[22247] = 32'b00000000000000000001000000011110;
assign LUT_1[22248] = 32'b00000000000000000011010100101111;
assign LUT_1[22249] = 32'b11111111111111111100100110101011;
assign LUT_1[22250] = 32'b11111111111111111111000011000000;
assign LUT_1[22251] = 32'b11111111111111111000010100111100;
assign LUT_1[22252] = 32'b00000000000000001011001110000110;
assign LUT_1[22253] = 32'b00000000000000000100100000000010;
assign LUT_1[22254] = 32'b00000000000000000110111100010111;
assign LUT_1[22255] = 32'b00000000000000000000001110010011;
assign LUT_1[22256] = 32'b00000000000000000110000010011100;
assign LUT_1[22257] = 32'b11111111111111111111010100011000;
assign LUT_1[22258] = 32'b00000000000000000001110000101101;
assign LUT_1[22259] = 32'b11111111111111111011000010101001;
assign LUT_1[22260] = 32'b00000000000000001101111011110011;
assign LUT_1[22261] = 32'b00000000000000000111001101101111;
assign LUT_1[22262] = 32'b00000000000000001001101010000100;
assign LUT_1[22263] = 32'b00000000000000000010111100000000;
assign LUT_1[22264] = 32'b00000000000000000101010000010001;
assign LUT_1[22265] = 32'b11111111111111111110100010001101;
assign LUT_1[22266] = 32'b00000000000000000000111110100010;
assign LUT_1[22267] = 32'b11111111111111111010010000011110;
assign LUT_1[22268] = 32'b00000000000000001101001001101000;
assign LUT_1[22269] = 32'b00000000000000000110011011100100;
assign LUT_1[22270] = 32'b00000000000000001000110111111001;
assign LUT_1[22271] = 32'b00000000000000000010001001110101;
assign LUT_1[22272] = 32'b11111111111111111100000010011100;
assign LUT_1[22273] = 32'b11111111111111110101010100011000;
assign LUT_1[22274] = 32'b11111111111111110111110000101101;
assign LUT_1[22275] = 32'b11111111111111110001000010101001;
assign LUT_1[22276] = 32'b00000000000000000011111011110011;
assign LUT_1[22277] = 32'b11111111111111111101001101101111;
assign LUT_1[22278] = 32'b11111111111111111111101010000100;
assign LUT_1[22279] = 32'b11111111111111111000111100000000;
assign LUT_1[22280] = 32'b11111111111111111011010000010001;
assign LUT_1[22281] = 32'b11111111111111110100100010001101;
assign LUT_1[22282] = 32'b11111111111111110110111110100010;
assign LUT_1[22283] = 32'b11111111111111110000010000011110;
assign LUT_1[22284] = 32'b00000000000000000011001001101000;
assign LUT_1[22285] = 32'b11111111111111111100011011100100;
assign LUT_1[22286] = 32'b11111111111111111110110111111001;
assign LUT_1[22287] = 32'b11111111111111111000001001110101;
assign LUT_1[22288] = 32'b11111111111111111101111101111110;
assign LUT_1[22289] = 32'b11111111111111110111001111111010;
assign LUT_1[22290] = 32'b11111111111111111001101100001111;
assign LUT_1[22291] = 32'b11111111111111110010111110001011;
assign LUT_1[22292] = 32'b00000000000000000101110111010101;
assign LUT_1[22293] = 32'b11111111111111111111001001010001;
assign LUT_1[22294] = 32'b00000000000000000001100101100110;
assign LUT_1[22295] = 32'b11111111111111111010110111100010;
assign LUT_1[22296] = 32'b11111111111111111101001011110011;
assign LUT_1[22297] = 32'b11111111111111110110011101101111;
assign LUT_1[22298] = 32'b11111111111111111000111010000100;
assign LUT_1[22299] = 32'b11111111111111110010001100000000;
assign LUT_1[22300] = 32'b00000000000000000101000101001010;
assign LUT_1[22301] = 32'b11111111111111111110010111000110;
assign LUT_1[22302] = 32'b00000000000000000000110011011011;
assign LUT_1[22303] = 32'b11111111111111111010000101010111;
assign LUT_1[22304] = 32'b11111111111111111100111101011011;
assign LUT_1[22305] = 32'b11111111111111110110001111010111;
assign LUT_1[22306] = 32'b11111111111111111000101011101100;
assign LUT_1[22307] = 32'b11111111111111110001111101101000;
assign LUT_1[22308] = 32'b00000000000000000100110110110010;
assign LUT_1[22309] = 32'b11111111111111111110001000101110;
assign LUT_1[22310] = 32'b00000000000000000000100101000011;
assign LUT_1[22311] = 32'b11111111111111111001110110111111;
assign LUT_1[22312] = 32'b11111111111111111100001011010000;
assign LUT_1[22313] = 32'b11111111111111110101011101001100;
assign LUT_1[22314] = 32'b11111111111111110111111001100001;
assign LUT_1[22315] = 32'b11111111111111110001001011011101;
assign LUT_1[22316] = 32'b00000000000000000100000100100111;
assign LUT_1[22317] = 32'b11111111111111111101010110100011;
assign LUT_1[22318] = 32'b11111111111111111111110010111000;
assign LUT_1[22319] = 32'b11111111111111111001000100110100;
assign LUT_1[22320] = 32'b11111111111111111110111000111101;
assign LUT_1[22321] = 32'b11111111111111111000001010111001;
assign LUT_1[22322] = 32'b11111111111111111010100111001110;
assign LUT_1[22323] = 32'b11111111111111110011111001001010;
assign LUT_1[22324] = 32'b00000000000000000110110010010100;
assign LUT_1[22325] = 32'b00000000000000000000000100010000;
assign LUT_1[22326] = 32'b00000000000000000010100000100101;
assign LUT_1[22327] = 32'b11111111111111111011110010100001;
assign LUT_1[22328] = 32'b11111111111111111110000110110010;
assign LUT_1[22329] = 32'b11111111111111110111011000101110;
assign LUT_1[22330] = 32'b11111111111111111001110101000011;
assign LUT_1[22331] = 32'b11111111111111110011000110111111;
assign LUT_1[22332] = 32'b00000000000000000110000000001001;
assign LUT_1[22333] = 32'b11111111111111111111010010000101;
assign LUT_1[22334] = 32'b00000000000000000001101110011010;
assign LUT_1[22335] = 32'b11111111111111111011000000010110;
assign LUT_1[22336] = 32'b11111111111111111110000000000100;
assign LUT_1[22337] = 32'b11111111111111110111010010000000;
assign LUT_1[22338] = 32'b11111111111111111001101110010101;
assign LUT_1[22339] = 32'b11111111111111110011000000010001;
assign LUT_1[22340] = 32'b00000000000000000101111001011011;
assign LUT_1[22341] = 32'b11111111111111111111001011010111;
assign LUT_1[22342] = 32'b00000000000000000001100111101100;
assign LUT_1[22343] = 32'b11111111111111111010111001101000;
assign LUT_1[22344] = 32'b11111111111111111101001101111001;
assign LUT_1[22345] = 32'b11111111111111110110011111110101;
assign LUT_1[22346] = 32'b11111111111111111000111100001010;
assign LUT_1[22347] = 32'b11111111111111110010001110000110;
assign LUT_1[22348] = 32'b00000000000000000101000111010000;
assign LUT_1[22349] = 32'b11111111111111111110011001001100;
assign LUT_1[22350] = 32'b00000000000000000000110101100001;
assign LUT_1[22351] = 32'b11111111111111111010000111011101;
assign LUT_1[22352] = 32'b11111111111111111111111011100110;
assign LUT_1[22353] = 32'b11111111111111111001001101100010;
assign LUT_1[22354] = 32'b11111111111111111011101001110111;
assign LUT_1[22355] = 32'b11111111111111110100111011110011;
assign LUT_1[22356] = 32'b00000000000000000111110100111101;
assign LUT_1[22357] = 32'b00000000000000000001000110111001;
assign LUT_1[22358] = 32'b00000000000000000011100011001110;
assign LUT_1[22359] = 32'b11111111111111111100110101001010;
assign LUT_1[22360] = 32'b11111111111111111111001001011011;
assign LUT_1[22361] = 32'b11111111111111111000011011010111;
assign LUT_1[22362] = 32'b11111111111111111010110111101100;
assign LUT_1[22363] = 32'b11111111111111110100001001101000;
assign LUT_1[22364] = 32'b00000000000000000111000010110010;
assign LUT_1[22365] = 32'b00000000000000000000010100101110;
assign LUT_1[22366] = 32'b00000000000000000010110001000011;
assign LUT_1[22367] = 32'b11111111111111111100000010111111;
assign LUT_1[22368] = 32'b11111111111111111110111011000011;
assign LUT_1[22369] = 32'b11111111111111111000001100111111;
assign LUT_1[22370] = 32'b11111111111111111010101001010100;
assign LUT_1[22371] = 32'b11111111111111110011111011010000;
assign LUT_1[22372] = 32'b00000000000000000110110100011010;
assign LUT_1[22373] = 32'b00000000000000000000000110010110;
assign LUT_1[22374] = 32'b00000000000000000010100010101011;
assign LUT_1[22375] = 32'b11111111111111111011110100100111;
assign LUT_1[22376] = 32'b11111111111111111110001000111000;
assign LUT_1[22377] = 32'b11111111111111110111011010110100;
assign LUT_1[22378] = 32'b11111111111111111001110111001001;
assign LUT_1[22379] = 32'b11111111111111110011001001000101;
assign LUT_1[22380] = 32'b00000000000000000110000010001111;
assign LUT_1[22381] = 32'b11111111111111111111010100001011;
assign LUT_1[22382] = 32'b00000000000000000001110000100000;
assign LUT_1[22383] = 32'b11111111111111111011000010011100;
assign LUT_1[22384] = 32'b00000000000000000000110110100101;
assign LUT_1[22385] = 32'b11111111111111111010001000100001;
assign LUT_1[22386] = 32'b11111111111111111100100100110110;
assign LUT_1[22387] = 32'b11111111111111110101110110110010;
assign LUT_1[22388] = 32'b00000000000000001000101111111100;
assign LUT_1[22389] = 32'b00000000000000000010000001111000;
assign LUT_1[22390] = 32'b00000000000000000100011110001101;
assign LUT_1[22391] = 32'b11111111111111111101110000001001;
assign LUT_1[22392] = 32'b00000000000000000000000100011010;
assign LUT_1[22393] = 32'b11111111111111111001010110010110;
assign LUT_1[22394] = 32'b11111111111111111011110010101011;
assign LUT_1[22395] = 32'b11111111111111110101000100100111;
assign LUT_1[22396] = 32'b00000000000000000111111101110001;
assign LUT_1[22397] = 32'b00000000000000000001001111101101;
assign LUT_1[22398] = 32'b00000000000000000011101100000010;
assign LUT_1[22399] = 32'b11111111111111111100111101111110;
assign LUT_1[22400] = 32'b11111111111111111111000010011111;
assign LUT_1[22401] = 32'b11111111111111111000010100011011;
assign LUT_1[22402] = 32'b11111111111111111010110000110000;
assign LUT_1[22403] = 32'b11111111111111110100000010101100;
assign LUT_1[22404] = 32'b00000000000000000110111011110110;
assign LUT_1[22405] = 32'b00000000000000000000001101110010;
assign LUT_1[22406] = 32'b00000000000000000010101010000111;
assign LUT_1[22407] = 32'b11111111111111111011111100000011;
assign LUT_1[22408] = 32'b11111111111111111110010000010100;
assign LUT_1[22409] = 32'b11111111111111110111100010010000;
assign LUT_1[22410] = 32'b11111111111111111001111110100101;
assign LUT_1[22411] = 32'b11111111111111110011010000100001;
assign LUT_1[22412] = 32'b00000000000000000110001001101011;
assign LUT_1[22413] = 32'b11111111111111111111011011100111;
assign LUT_1[22414] = 32'b00000000000000000001110111111100;
assign LUT_1[22415] = 32'b11111111111111111011001001111000;
assign LUT_1[22416] = 32'b00000000000000000000111110000001;
assign LUT_1[22417] = 32'b11111111111111111010001111111101;
assign LUT_1[22418] = 32'b11111111111111111100101100010010;
assign LUT_1[22419] = 32'b11111111111111110101111110001110;
assign LUT_1[22420] = 32'b00000000000000001000110111011000;
assign LUT_1[22421] = 32'b00000000000000000010001001010100;
assign LUT_1[22422] = 32'b00000000000000000100100101101001;
assign LUT_1[22423] = 32'b11111111111111111101110111100101;
assign LUT_1[22424] = 32'b00000000000000000000001011110110;
assign LUT_1[22425] = 32'b11111111111111111001011101110010;
assign LUT_1[22426] = 32'b11111111111111111011111010000111;
assign LUT_1[22427] = 32'b11111111111111110101001100000011;
assign LUT_1[22428] = 32'b00000000000000001000000101001101;
assign LUT_1[22429] = 32'b00000000000000000001010111001001;
assign LUT_1[22430] = 32'b00000000000000000011110011011110;
assign LUT_1[22431] = 32'b11111111111111111101000101011010;
assign LUT_1[22432] = 32'b11111111111111111111111101011110;
assign LUT_1[22433] = 32'b11111111111111111001001111011010;
assign LUT_1[22434] = 32'b11111111111111111011101011101111;
assign LUT_1[22435] = 32'b11111111111111110100111101101011;
assign LUT_1[22436] = 32'b00000000000000000111110110110101;
assign LUT_1[22437] = 32'b00000000000000000001001000110001;
assign LUT_1[22438] = 32'b00000000000000000011100101000110;
assign LUT_1[22439] = 32'b11111111111111111100110111000010;
assign LUT_1[22440] = 32'b11111111111111111111001011010011;
assign LUT_1[22441] = 32'b11111111111111111000011101001111;
assign LUT_1[22442] = 32'b11111111111111111010111001100100;
assign LUT_1[22443] = 32'b11111111111111110100001011100000;
assign LUT_1[22444] = 32'b00000000000000000111000100101010;
assign LUT_1[22445] = 32'b00000000000000000000010110100110;
assign LUT_1[22446] = 32'b00000000000000000010110010111011;
assign LUT_1[22447] = 32'b11111111111111111100000100110111;
assign LUT_1[22448] = 32'b00000000000000000001111001000000;
assign LUT_1[22449] = 32'b11111111111111111011001010111100;
assign LUT_1[22450] = 32'b11111111111111111101100111010001;
assign LUT_1[22451] = 32'b11111111111111110110111001001101;
assign LUT_1[22452] = 32'b00000000000000001001110010010111;
assign LUT_1[22453] = 32'b00000000000000000011000100010011;
assign LUT_1[22454] = 32'b00000000000000000101100000101000;
assign LUT_1[22455] = 32'b11111111111111111110110010100100;
assign LUT_1[22456] = 32'b00000000000000000001000110110101;
assign LUT_1[22457] = 32'b11111111111111111010011000110001;
assign LUT_1[22458] = 32'b11111111111111111100110101000110;
assign LUT_1[22459] = 32'b11111111111111110110000111000010;
assign LUT_1[22460] = 32'b00000000000000001001000000001100;
assign LUT_1[22461] = 32'b00000000000000000010010010001000;
assign LUT_1[22462] = 32'b00000000000000000100101110011101;
assign LUT_1[22463] = 32'b11111111111111111110000000011001;
assign LUT_1[22464] = 32'b00000000000000000001000000000111;
assign LUT_1[22465] = 32'b11111111111111111010010010000011;
assign LUT_1[22466] = 32'b11111111111111111100101110011000;
assign LUT_1[22467] = 32'b11111111111111110110000000010100;
assign LUT_1[22468] = 32'b00000000000000001000111001011110;
assign LUT_1[22469] = 32'b00000000000000000010001011011010;
assign LUT_1[22470] = 32'b00000000000000000100100111101111;
assign LUT_1[22471] = 32'b11111111111111111101111001101011;
assign LUT_1[22472] = 32'b00000000000000000000001101111100;
assign LUT_1[22473] = 32'b11111111111111111001011111111000;
assign LUT_1[22474] = 32'b11111111111111111011111100001101;
assign LUT_1[22475] = 32'b11111111111111110101001110001001;
assign LUT_1[22476] = 32'b00000000000000001000000111010011;
assign LUT_1[22477] = 32'b00000000000000000001011001001111;
assign LUT_1[22478] = 32'b00000000000000000011110101100100;
assign LUT_1[22479] = 32'b11111111111111111101000111100000;
assign LUT_1[22480] = 32'b00000000000000000010111011101001;
assign LUT_1[22481] = 32'b11111111111111111100001101100101;
assign LUT_1[22482] = 32'b11111111111111111110101001111010;
assign LUT_1[22483] = 32'b11111111111111110111111011110110;
assign LUT_1[22484] = 32'b00000000000000001010110101000000;
assign LUT_1[22485] = 32'b00000000000000000100000110111100;
assign LUT_1[22486] = 32'b00000000000000000110100011010001;
assign LUT_1[22487] = 32'b11111111111111111111110101001101;
assign LUT_1[22488] = 32'b00000000000000000010001001011110;
assign LUT_1[22489] = 32'b11111111111111111011011011011010;
assign LUT_1[22490] = 32'b11111111111111111101110111101111;
assign LUT_1[22491] = 32'b11111111111111110111001001101011;
assign LUT_1[22492] = 32'b00000000000000001010000010110101;
assign LUT_1[22493] = 32'b00000000000000000011010100110001;
assign LUT_1[22494] = 32'b00000000000000000101110001000110;
assign LUT_1[22495] = 32'b11111111111111111111000011000010;
assign LUT_1[22496] = 32'b00000000000000000001111011000110;
assign LUT_1[22497] = 32'b11111111111111111011001101000010;
assign LUT_1[22498] = 32'b11111111111111111101101001010111;
assign LUT_1[22499] = 32'b11111111111111110110111011010011;
assign LUT_1[22500] = 32'b00000000000000001001110100011101;
assign LUT_1[22501] = 32'b00000000000000000011000110011001;
assign LUT_1[22502] = 32'b00000000000000000101100010101110;
assign LUT_1[22503] = 32'b11111111111111111110110100101010;
assign LUT_1[22504] = 32'b00000000000000000001001000111011;
assign LUT_1[22505] = 32'b11111111111111111010011010110111;
assign LUT_1[22506] = 32'b11111111111111111100110111001100;
assign LUT_1[22507] = 32'b11111111111111110110001001001000;
assign LUT_1[22508] = 32'b00000000000000001001000010010010;
assign LUT_1[22509] = 32'b00000000000000000010010100001110;
assign LUT_1[22510] = 32'b00000000000000000100110000100011;
assign LUT_1[22511] = 32'b11111111111111111110000010011111;
assign LUT_1[22512] = 32'b00000000000000000011110110101000;
assign LUT_1[22513] = 32'b11111111111111111101001000100100;
assign LUT_1[22514] = 32'b11111111111111111111100100111001;
assign LUT_1[22515] = 32'b11111111111111111000110110110101;
assign LUT_1[22516] = 32'b00000000000000001011101111111111;
assign LUT_1[22517] = 32'b00000000000000000101000001111011;
assign LUT_1[22518] = 32'b00000000000000000111011110010000;
assign LUT_1[22519] = 32'b00000000000000000000110000001100;
assign LUT_1[22520] = 32'b00000000000000000011000100011101;
assign LUT_1[22521] = 32'b11111111111111111100010110011001;
assign LUT_1[22522] = 32'b11111111111111111110110010101110;
assign LUT_1[22523] = 32'b11111111111111111000000100101010;
assign LUT_1[22524] = 32'b00000000000000001010111101110100;
assign LUT_1[22525] = 32'b00000000000000000100001111110000;
assign LUT_1[22526] = 32'b00000000000000000110101100000101;
assign LUT_1[22527] = 32'b11111111111111111111111110000001;
assign LUT_1[22528] = 32'b11111111111111111111001010111110;
assign LUT_1[22529] = 32'b11111111111111111000011100111010;
assign LUT_1[22530] = 32'b11111111111111111010111001001111;
assign LUT_1[22531] = 32'b11111111111111110100001011001011;
assign LUT_1[22532] = 32'b00000000000000000111000100010101;
assign LUT_1[22533] = 32'b00000000000000000000010110010001;
assign LUT_1[22534] = 32'b00000000000000000010110010100110;
assign LUT_1[22535] = 32'b11111111111111111100000100100010;
assign LUT_1[22536] = 32'b11111111111111111110011000110011;
assign LUT_1[22537] = 32'b11111111111111110111101010101111;
assign LUT_1[22538] = 32'b11111111111111111010000111000100;
assign LUT_1[22539] = 32'b11111111111111110011011001000000;
assign LUT_1[22540] = 32'b00000000000000000110010010001010;
assign LUT_1[22541] = 32'b11111111111111111111100100000110;
assign LUT_1[22542] = 32'b00000000000000000010000000011011;
assign LUT_1[22543] = 32'b11111111111111111011010010010111;
assign LUT_1[22544] = 32'b00000000000000000001000110100000;
assign LUT_1[22545] = 32'b11111111111111111010011000011100;
assign LUT_1[22546] = 32'b11111111111111111100110100110001;
assign LUT_1[22547] = 32'b11111111111111110110000110101101;
assign LUT_1[22548] = 32'b00000000000000001000111111110111;
assign LUT_1[22549] = 32'b00000000000000000010010001110011;
assign LUT_1[22550] = 32'b00000000000000000100101110001000;
assign LUT_1[22551] = 32'b11111111111111111110000000000100;
assign LUT_1[22552] = 32'b00000000000000000000010100010101;
assign LUT_1[22553] = 32'b11111111111111111001100110010001;
assign LUT_1[22554] = 32'b11111111111111111100000010100110;
assign LUT_1[22555] = 32'b11111111111111110101010100100010;
assign LUT_1[22556] = 32'b00000000000000001000001101101100;
assign LUT_1[22557] = 32'b00000000000000000001011111101000;
assign LUT_1[22558] = 32'b00000000000000000011111011111101;
assign LUT_1[22559] = 32'b11111111111111111101001101111001;
assign LUT_1[22560] = 32'b00000000000000000000000101111101;
assign LUT_1[22561] = 32'b11111111111111111001010111111001;
assign LUT_1[22562] = 32'b11111111111111111011110100001110;
assign LUT_1[22563] = 32'b11111111111111110101000110001010;
assign LUT_1[22564] = 32'b00000000000000000111111111010100;
assign LUT_1[22565] = 32'b00000000000000000001010001010000;
assign LUT_1[22566] = 32'b00000000000000000011101101100101;
assign LUT_1[22567] = 32'b11111111111111111100111111100001;
assign LUT_1[22568] = 32'b11111111111111111111010011110010;
assign LUT_1[22569] = 32'b11111111111111111000100101101110;
assign LUT_1[22570] = 32'b11111111111111111011000010000011;
assign LUT_1[22571] = 32'b11111111111111110100010011111111;
assign LUT_1[22572] = 32'b00000000000000000111001101001001;
assign LUT_1[22573] = 32'b00000000000000000000011111000101;
assign LUT_1[22574] = 32'b00000000000000000010111011011010;
assign LUT_1[22575] = 32'b11111111111111111100001101010110;
assign LUT_1[22576] = 32'b00000000000000000010000001011111;
assign LUT_1[22577] = 32'b11111111111111111011010011011011;
assign LUT_1[22578] = 32'b11111111111111111101101111110000;
assign LUT_1[22579] = 32'b11111111111111110111000001101100;
assign LUT_1[22580] = 32'b00000000000000001001111010110110;
assign LUT_1[22581] = 32'b00000000000000000011001100110010;
assign LUT_1[22582] = 32'b00000000000000000101101001000111;
assign LUT_1[22583] = 32'b11111111111111111110111011000011;
assign LUT_1[22584] = 32'b00000000000000000001001111010100;
assign LUT_1[22585] = 32'b11111111111111111010100001010000;
assign LUT_1[22586] = 32'b11111111111111111100111101100101;
assign LUT_1[22587] = 32'b11111111111111110110001111100001;
assign LUT_1[22588] = 32'b00000000000000001001001000101011;
assign LUT_1[22589] = 32'b00000000000000000010011010100111;
assign LUT_1[22590] = 32'b00000000000000000100110110111100;
assign LUT_1[22591] = 32'b11111111111111111110001000111000;
assign LUT_1[22592] = 32'b00000000000000000001001000100110;
assign LUT_1[22593] = 32'b11111111111111111010011010100010;
assign LUT_1[22594] = 32'b11111111111111111100110110110111;
assign LUT_1[22595] = 32'b11111111111111110110001000110011;
assign LUT_1[22596] = 32'b00000000000000001001000001111101;
assign LUT_1[22597] = 32'b00000000000000000010010011111001;
assign LUT_1[22598] = 32'b00000000000000000100110000001110;
assign LUT_1[22599] = 32'b11111111111111111110000010001010;
assign LUT_1[22600] = 32'b00000000000000000000010110011011;
assign LUT_1[22601] = 32'b11111111111111111001101000010111;
assign LUT_1[22602] = 32'b11111111111111111100000100101100;
assign LUT_1[22603] = 32'b11111111111111110101010110101000;
assign LUT_1[22604] = 32'b00000000000000001000001111110010;
assign LUT_1[22605] = 32'b00000000000000000001100001101110;
assign LUT_1[22606] = 32'b00000000000000000011111110000011;
assign LUT_1[22607] = 32'b11111111111111111101001111111111;
assign LUT_1[22608] = 32'b00000000000000000011000100001000;
assign LUT_1[22609] = 32'b11111111111111111100010110000100;
assign LUT_1[22610] = 32'b11111111111111111110110010011001;
assign LUT_1[22611] = 32'b11111111111111111000000100010101;
assign LUT_1[22612] = 32'b00000000000000001010111101011111;
assign LUT_1[22613] = 32'b00000000000000000100001111011011;
assign LUT_1[22614] = 32'b00000000000000000110101011110000;
assign LUT_1[22615] = 32'b11111111111111111111111101101100;
assign LUT_1[22616] = 32'b00000000000000000010010001111101;
assign LUT_1[22617] = 32'b11111111111111111011100011111001;
assign LUT_1[22618] = 32'b11111111111111111110000000001110;
assign LUT_1[22619] = 32'b11111111111111110111010010001010;
assign LUT_1[22620] = 32'b00000000000000001010001011010100;
assign LUT_1[22621] = 32'b00000000000000000011011101010000;
assign LUT_1[22622] = 32'b00000000000000000101111001100101;
assign LUT_1[22623] = 32'b11111111111111111111001011100001;
assign LUT_1[22624] = 32'b00000000000000000010000011100101;
assign LUT_1[22625] = 32'b11111111111111111011010101100001;
assign LUT_1[22626] = 32'b11111111111111111101110001110110;
assign LUT_1[22627] = 32'b11111111111111110111000011110010;
assign LUT_1[22628] = 32'b00000000000000001001111100111100;
assign LUT_1[22629] = 32'b00000000000000000011001110111000;
assign LUT_1[22630] = 32'b00000000000000000101101011001101;
assign LUT_1[22631] = 32'b11111111111111111110111101001001;
assign LUT_1[22632] = 32'b00000000000000000001010001011010;
assign LUT_1[22633] = 32'b11111111111111111010100011010110;
assign LUT_1[22634] = 32'b11111111111111111100111111101011;
assign LUT_1[22635] = 32'b11111111111111110110010001100111;
assign LUT_1[22636] = 32'b00000000000000001001001010110001;
assign LUT_1[22637] = 32'b00000000000000000010011100101101;
assign LUT_1[22638] = 32'b00000000000000000100111001000010;
assign LUT_1[22639] = 32'b11111111111111111110001010111110;
assign LUT_1[22640] = 32'b00000000000000000011111111000111;
assign LUT_1[22641] = 32'b11111111111111111101010001000011;
assign LUT_1[22642] = 32'b11111111111111111111101101011000;
assign LUT_1[22643] = 32'b11111111111111111000111111010100;
assign LUT_1[22644] = 32'b00000000000000001011111000011110;
assign LUT_1[22645] = 32'b00000000000000000101001010011010;
assign LUT_1[22646] = 32'b00000000000000000111100110101111;
assign LUT_1[22647] = 32'b00000000000000000000111000101011;
assign LUT_1[22648] = 32'b00000000000000000011001100111100;
assign LUT_1[22649] = 32'b11111111111111111100011110111000;
assign LUT_1[22650] = 32'b11111111111111111110111011001101;
assign LUT_1[22651] = 32'b11111111111111111000001101001001;
assign LUT_1[22652] = 32'b00000000000000001011000110010011;
assign LUT_1[22653] = 32'b00000000000000000100011000001111;
assign LUT_1[22654] = 32'b00000000000000000110110100100100;
assign LUT_1[22655] = 32'b00000000000000000000000110100000;
assign LUT_1[22656] = 32'b00000000000000000010001011000001;
assign LUT_1[22657] = 32'b11111111111111111011011100111101;
assign LUT_1[22658] = 32'b11111111111111111101111001010010;
assign LUT_1[22659] = 32'b11111111111111110111001011001110;
assign LUT_1[22660] = 32'b00000000000000001010000100011000;
assign LUT_1[22661] = 32'b00000000000000000011010110010100;
assign LUT_1[22662] = 32'b00000000000000000101110010101001;
assign LUT_1[22663] = 32'b11111111111111111111000100100101;
assign LUT_1[22664] = 32'b00000000000000000001011000110110;
assign LUT_1[22665] = 32'b11111111111111111010101010110010;
assign LUT_1[22666] = 32'b11111111111111111101000111000111;
assign LUT_1[22667] = 32'b11111111111111110110011001000011;
assign LUT_1[22668] = 32'b00000000000000001001010010001101;
assign LUT_1[22669] = 32'b00000000000000000010100100001001;
assign LUT_1[22670] = 32'b00000000000000000101000000011110;
assign LUT_1[22671] = 32'b11111111111111111110010010011010;
assign LUT_1[22672] = 32'b00000000000000000100000110100011;
assign LUT_1[22673] = 32'b11111111111111111101011000011111;
assign LUT_1[22674] = 32'b11111111111111111111110100110100;
assign LUT_1[22675] = 32'b11111111111111111001000110110000;
assign LUT_1[22676] = 32'b00000000000000001011111111111010;
assign LUT_1[22677] = 32'b00000000000000000101010001110110;
assign LUT_1[22678] = 32'b00000000000000000111101110001011;
assign LUT_1[22679] = 32'b00000000000000000001000000000111;
assign LUT_1[22680] = 32'b00000000000000000011010100011000;
assign LUT_1[22681] = 32'b11111111111111111100100110010100;
assign LUT_1[22682] = 32'b11111111111111111111000010101001;
assign LUT_1[22683] = 32'b11111111111111111000010100100101;
assign LUT_1[22684] = 32'b00000000000000001011001101101111;
assign LUT_1[22685] = 32'b00000000000000000100011111101011;
assign LUT_1[22686] = 32'b00000000000000000110111100000000;
assign LUT_1[22687] = 32'b00000000000000000000001101111100;
assign LUT_1[22688] = 32'b00000000000000000011000110000000;
assign LUT_1[22689] = 32'b11111111111111111100010111111100;
assign LUT_1[22690] = 32'b11111111111111111110110100010001;
assign LUT_1[22691] = 32'b11111111111111111000000110001101;
assign LUT_1[22692] = 32'b00000000000000001010111111010111;
assign LUT_1[22693] = 32'b00000000000000000100010001010011;
assign LUT_1[22694] = 32'b00000000000000000110101101101000;
assign LUT_1[22695] = 32'b11111111111111111111111111100100;
assign LUT_1[22696] = 32'b00000000000000000010010011110101;
assign LUT_1[22697] = 32'b11111111111111111011100101110001;
assign LUT_1[22698] = 32'b11111111111111111110000010000110;
assign LUT_1[22699] = 32'b11111111111111110111010100000010;
assign LUT_1[22700] = 32'b00000000000000001010001101001100;
assign LUT_1[22701] = 32'b00000000000000000011011111001000;
assign LUT_1[22702] = 32'b00000000000000000101111011011101;
assign LUT_1[22703] = 32'b11111111111111111111001101011001;
assign LUT_1[22704] = 32'b00000000000000000101000001100010;
assign LUT_1[22705] = 32'b11111111111111111110010011011110;
assign LUT_1[22706] = 32'b00000000000000000000101111110011;
assign LUT_1[22707] = 32'b11111111111111111010000001101111;
assign LUT_1[22708] = 32'b00000000000000001100111010111001;
assign LUT_1[22709] = 32'b00000000000000000110001100110101;
assign LUT_1[22710] = 32'b00000000000000001000101001001010;
assign LUT_1[22711] = 32'b00000000000000000001111011000110;
assign LUT_1[22712] = 32'b00000000000000000100001111010111;
assign LUT_1[22713] = 32'b11111111111111111101100001010011;
assign LUT_1[22714] = 32'b11111111111111111111111101101000;
assign LUT_1[22715] = 32'b11111111111111111001001111100100;
assign LUT_1[22716] = 32'b00000000000000001100001000101110;
assign LUT_1[22717] = 32'b00000000000000000101011010101010;
assign LUT_1[22718] = 32'b00000000000000000111110110111111;
assign LUT_1[22719] = 32'b00000000000000000001001000111011;
assign LUT_1[22720] = 32'b00000000000000000100001000101001;
assign LUT_1[22721] = 32'b11111111111111111101011010100101;
assign LUT_1[22722] = 32'b11111111111111111111110110111010;
assign LUT_1[22723] = 32'b11111111111111111001001000110110;
assign LUT_1[22724] = 32'b00000000000000001100000010000000;
assign LUT_1[22725] = 32'b00000000000000000101010011111100;
assign LUT_1[22726] = 32'b00000000000000000111110000010001;
assign LUT_1[22727] = 32'b00000000000000000001000010001101;
assign LUT_1[22728] = 32'b00000000000000000011010110011110;
assign LUT_1[22729] = 32'b11111111111111111100101000011010;
assign LUT_1[22730] = 32'b11111111111111111111000100101111;
assign LUT_1[22731] = 32'b11111111111111111000010110101011;
assign LUT_1[22732] = 32'b00000000000000001011001111110101;
assign LUT_1[22733] = 32'b00000000000000000100100001110001;
assign LUT_1[22734] = 32'b00000000000000000110111110000110;
assign LUT_1[22735] = 32'b00000000000000000000010000000010;
assign LUT_1[22736] = 32'b00000000000000000110000100001011;
assign LUT_1[22737] = 32'b11111111111111111111010110000111;
assign LUT_1[22738] = 32'b00000000000000000001110010011100;
assign LUT_1[22739] = 32'b11111111111111111011000100011000;
assign LUT_1[22740] = 32'b00000000000000001101111101100010;
assign LUT_1[22741] = 32'b00000000000000000111001111011110;
assign LUT_1[22742] = 32'b00000000000000001001101011110011;
assign LUT_1[22743] = 32'b00000000000000000010111101101111;
assign LUT_1[22744] = 32'b00000000000000000101010010000000;
assign LUT_1[22745] = 32'b11111111111111111110100011111100;
assign LUT_1[22746] = 32'b00000000000000000001000000010001;
assign LUT_1[22747] = 32'b11111111111111111010010010001101;
assign LUT_1[22748] = 32'b00000000000000001101001011010111;
assign LUT_1[22749] = 32'b00000000000000000110011101010011;
assign LUT_1[22750] = 32'b00000000000000001000111001101000;
assign LUT_1[22751] = 32'b00000000000000000010001011100100;
assign LUT_1[22752] = 32'b00000000000000000101000011101000;
assign LUT_1[22753] = 32'b11111111111111111110010101100100;
assign LUT_1[22754] = 32'b00000000000000000000110001111001;
assign LUT_1[22755] = 32'b11111111111111111010000011110101;
assign LUT_1[22756] = 32'b00000000000000001100111100111111;
assign LUT_1[22757] = 32'b00000000000000000110001110111011;
assign LUT_1[22758] = 32'b00000000000000001000101011010000;
assign LUT_1[22759] = 32'b00000000000000000001111101001100;
assign LUT_1[22760] = 32'b00000000000000000100010001011101;
assign LUT_1[22761] = 32'b11111111111111111101100011011001;
assign LUT_1[22762] = 32'b11111111111111111111111111101110;
assign LUT_1[22763] = 32'b11111111111111111001010001101010;
assign LUT_1[22764] = 32'b00000000000000001100001010110100;
assign LUT_1[22765] = 32'b00000000000000000101011100110000;
assign LUT_1[22766] = 32'b00000000000000000111111001000101;
assign LUT_1[22767] = 32'b00000000000000000001001011000001;
assign LUT_1[22768] = 32'b00000000000000000110111111001010;
assign LUT_1[22769] = 32'b00000000000000000000010001000110;
assign LUT_1[22770] = 32'b00000000000000000010101101011011;
assign LUT_1[22771] = 32'b11111111111111111011111111010111;
assign LUT_1[22772] = 32'b00000000000000001110111000100001;
assign LUT_1[22773] = 32'b00000000000000001000001010011101;
assign LUT_1[22774] = 32'b00000000000000001010100110110010;
assign LUT_1[22775] = 32'b00000000000000000011111000101110;
assign LUT_1[22776] = 32'b00000000000000000110001100111111;
assign LUT_1[22777] = 32'b11111111111111111111011110111011;
assign LUT_1[22778] = 32'b00000000000000000001111011010000;
assign LUT_1[22779] = 32'b11111111111111111011001101001100;
assign LUT_1[22780] = 32'b00000000000000001110000110010110;
assign LUT_1[22781] = 32'b00000000000000000111011000010010;
assign LUT_1[22782] = 32'b00000000000000001001110100100111;
assign LUT_1[22783] = 32'b00000000000000000011000110100011;
assign LUT_1[22784] = 32'b11111111111111111100111111001010;
assign LUT_1[22785] = 32'b11111111111111110110010001000110;
assign LUT_1[22786] = 32'b11111111111111111000101101011011;
assign LUT_1[22787] = 32'b11111111111111110001111111010111;
assign LUT_1[22788] = 32'b00000000000000000100111000100001;
assign LUT_1[22789] = 32'b11111111111111111110001010011101;
assign LUT_1[22790] = 32'b00000000000000000000100110110010;
assign LUT_1[22791] = 32'b11111111111111111001111000101110;
assign LUT_1[22792] = 32'b11111111111111111100001100111111;
assign LUT_1[22793] = 32'b11111111111111110101011110111011;
assign LUT_1[22794] = 32'b11111111111111110111111011010000;
assign LUT_1[22795] = 32'b11111111111111110001001101001100;
assign LUT_1[22796] = 32'b00000000000000000100000110010110;
assign LUT_1[22797] = 32'b11111111111111111101011000010010;
assign LUT_1[22798] = 32'b11111111111111111111110100100111;
assign LUT_1[22799] = 32'b11111111111111111001000110100011;
assign LUT_1[22800] = 32'b11111111111111111110111010101100;
assign LUT_1[22801] = 32'b11111111111111111000001100101000;
assign LUT_1[22802] = 32'b11111111111111111010101000111101;
assign LUT_1[22803] = 32'b11111111111111110011111010111001;
assign LUT_1[22804] = 32'b00000000000000000110110100000011;
assign LUT_1[22805] = 32'b00000000000000000000000101111111;
assign LUT_1[22806] = 32'b00000000000000000010100010010100;
assign LUT_1[22807] = 32'b11111111111111111011110100010000;
assign LUT_1[22808] = 32'b11111111111111111110001000100001;
assign LUT_1[22809] = 32'b11111111111111110111011010011101;
assign LUT_1[22810] = 32'b11111111111111111001110110110010;
assign LUT_1[22811] = 32'b11111111111111110011001000101110;
assign LUT_1[22812] = 32'b00000000000000000110000001111000;
assign LUT_1[22813] = 32'b11111111111111111111010011110100;
assign LUT_1[22814] = 32'b00000000000000000001110000001001;
assign LUT_1[22815] = 32'b11111111111111111011000010000101;
assign LUT_1[22816] = 32'b11111111111111111101111010001001;
assign LUT_1[22817] = 32'b11111111111111110111001100000101;
assign LUT_1[22818] = 32'b11111111111111111001101000011010;
assign LUT_1[22819] = 32'b11111111111111110010111010010110;
assign LUT_1[22820] = 32'b00000000000000000101110011100000;
assign LUT_1[22821] = 32'b11111111111111111111000101011100;
assign LUT_1[22822] = 32'b00000000000000000001100001110001;
assign LUT_1[22823] = 32'b11111111111111111010110011101101;
assign LUT_1[22824] = 32'b11111111111111111101000111111110;
assign LUT_1[22825] = 32'b11111111111111110110011001111010;
assign LUT_1[22826] = 32'b11111111111111111000110110001111;
assign LUT_1[22827] = 32'b11111111111111110010001000001011;
assign LUT_1[22828] = 32'b00000000000000000101000001010101;
assign LUT_1[22829] = 32'b11111111111111111110010011010001;
assign LUT_1[22830] = 32'b00000000000000000000101111100110;
assign LUT_1[22831] = 32'b11111111111111111010000001100010;
assign LUT_1[22832] = 32'b11111111111111111111110101101011;
assign LUT_1[22833] = 32'b11111111111111111001000111100111;
assign LUT_1[22834] = 32'b11111111111111111011100011111100;
assign LUT_1[22835] = 32'b11111111111111110100110101111000;
assign LUT_1[22836] = 32'b00000000000000000111101111000010;
assign LUT_1[22837] = 32'b00000000000000000001000000111110;
assign LUT_1[22838] = 32'b00000000000000000011011101010011;
assign LUT_1[22839] = 32'b11111111111111111100101111001111;
assign LUT_1[22840] = 32'b11111111111111111111000011100000;
assign LUT_1[22841] = 32'b11111111111111111000010101011100;
assign LUT_1[22842] = 32'b11111111111111111010110001110001;
assign LUT_1[22843] = 32'b11111111111111110100000011101101;
assign LUT_1[22844] = 32'b00000000000000000110111100110111;
assign LUT_1[22845] = 32'b00000000000000000000001110110011;
assign LUT_1[22846] = 32'b00000000000000000010101011001000;
assign LUT_1[22847] = 32'b11111111111111111011111101000100;
assign LUT_1[22848] = 32'b11111111111111111110111100110010;
assign LUT_1[22849] = 32'b11111111111111111000001110101110;
assign LUT_1[22850] = 32'b11111111111111111010101011000011;
assign LUT_1[22851] = 32'b11111111111111110011111100111111;
assign LUT_1[22852] = 32'b00000000000000000110110110001001;
assign LUT_1[22853] = 32'b00000000000000000000001000000101;
assign LUT_1[22854] = 32'b00000000000000000010100100011010;
assign LUT_1[22855] = 32'b11111111111111111011110110010110;
assign LUT_1[22856] = 32'b11111111111111111110001010100111;
assign LUT_1[22857] = 32'b11111111111111110111011100100011;
assign LUT_1[22858] = 32'b11111111111111111001111000111000;
assign LUT_1[22859] = 32'b11111111111111110011001010110100;
assign LUT_1[22860] = 32'b00000000000000000110000011111110;
assign LUT_1[22861] = 32'b11111111111111111111010101111010;
assign LUT_1[22862] = 32'b00000000000000000001110010001111;
assign LUT_1[22863] = 32'b11111111111111111011000100001011;
assign LUT_1[22864] = 32'b00000000000000000000111000010100;
assign LUT_1[22865] = 32'b11111111111111111010001010010000;
assign LUT_1[22866] = 32'b11111111111111111100100110100101;
assign LUT_1[22867] = 32'b11111111111111110101111000100001;
assign LUT_1[22868] = 32'b00000000000000001000110001101011;
assign LUT_1[22869] = 32'b00000000000000000010000011100111;
assign LUT_1[22870] = 32'b00000000000000000100011111111100;
assign LUT_1[22871] = 32'b11111111111111111101110001111000;
assign LUT_1[22872] = 32'b00000000000000000000000110001001;
assign LUT_1[22873] = 32'b11111111111111111001011000000101;
assign LUT_1[22874] = 32'b11111111111111111011110100011010;
assign LUT_1[22875] = 32'b11111111111111110101000110010110;
assign LUT_1[22876] = 32'b00000000000000000111111111100000;
assign LUT_1[22877] = 32'b00000000000000000001010001011100;
assign LUT_1[22878] = 32'b00000000000000000011101101110001;
assign LUT_1[22879] = 32'b11111111111111111100111111101101;
assign LUT_1[22880] = 32'b11111111111111111111110111110001;
assign LUT_1[22881] = 32'b11111111111111111001001001101101;
assign LUT_1[22882] = 32'b11111111111111111011100110000010;
assign LUT_1[22883] = 32'b11111111111111110100110111111110;
assign LUT_1[22884] = 32'b00000000000000000111110001001000;
assign LUT_1[22885] = 32'b00000000000000000001000011000100;
assign LUT_1[22886] = 32'b00000000000000000011011111011001;
assign LUT_1[22887] = 32'b11111111111111111100110001010101;
assign LUT_1[22888] = 32'b11111111111111111111000101100110;
assign LUT_1[22889] = 32'b11111111111111111000010111100010;
assign LUT_1[22890] = 32'b11111111111111111010110011110111;
assign LUT_1[22891] = 32'b11111111111111110100000101110011;
assign LUT_1[22892] = 32'b00000000000000000110111110111101;
assign LUT_1[22893] = 32'b00000000000000000000010000111001;
assign LUT_1[22894] = 32'b00000000000000000010101101001110;
assign LUT_1[22895] = 32'b11111111111111111011111111001010;
assign LUT_1[22896] = 32'b00000000000000000001110011010011;
assign LUT_1[22897] = 32'b11111111111111111011000101001111;
assign LUT_1[22898] = 32'b11111111111111111101100001100100;
assign LUT_1[22899] = 32'b11111111111111110110110011100000;
assign LUT_1[22900] = 32'b00000000000000001001101100101010;
assign LUT_1[22901] = 32'b00000000000000000010111110100110;
assign LUT_1[22902] = 32'b00000000000000000101011010111011;
assign LUT_1[22903] = 32'b11111111111111111110101100110111;
assign LUT_1[22904] = 32'b00000000000000000001000001001000;
assign LUT_1[22905] = 32'b11111111111111111010010011000100;
assign LUT_1[22906] = 32'b11111111111111111100101111011001;
assign LUT_1[22907] = 32'b11111111111111110110000001010101;
assign LUT_1[22908] = 32'b00000000000000001000111010011111;
assign LUT_1[22909] = 32'b00000000000000000010001100011011;
assign LUT_1[22910] = 32'b00000000000000000100101000110000;
assign LUT_1[22911] = 32'b11111111111111111101111010101100;
assign LUT_1[22912] = 32'b11111111111111111111111111001101;
assign LUT_1[22913] = 32'b11111111111111111001010001001001;
assign LUT_1[22914] = 32'b11111111111111111011101101011110;
assign LUT_1[22915] = 32'b11111111111111110100111111011010;
assign LUT_1[22916] = 32'b00000000000000000111111000100100;
assign LUT_1[22917] = 32'b00000000000000000001001010100000;
assign LUT_1[22918] = 32'b00000000000000000011100110110101;
assign LUT_1[22919] = 32'b11111111111111111100111000110001;
assign LUT_1[22920] = 32'b11111111111111111111001101000010;
assign LUT_1[22921] = 32'b11111111111111111000011110111110;
assign LUT_1[22922] = 32'b11111111111111111010111011010011;
assign LUT_1[22923] = 32'b11111111111111110100001101001111;
assign LUT_1[22924] = 32'b00000000000000000111000110011001;
assign LUT_1[22925] = 32'b00000000000000000000011000010101;
assign LUT_1[22926] = 32'b00000000000000000010110100101010;
assign LUT_1[22927] = 32'b11111111111111111100000110100110;
assign LUT_1[22928] = 32'b00000000000000000001111010101111;
assign LUT_1[22929] = 32'b11111111111111111011001100101011;
assign LUT_1[22930] = 32'b11111111111111111101101001000000;
assign LUT_1[22931] = 32'b11111111111111110110111010111100;
assign LUT_1[22932] = 32'b00000000000000001001110100000110;
assign LUT_1[22933] = 32'b00000000000000000011000110000010;
assign LUT_1[22934] = 32'b00000000000000000101100010010111;
assign LUT_1[22935] = 32'b11111111111111111110110100010011;
assign LUT_1[22936] = 32'b00000000000000000001001000100100;
assign LUT_1[22937] = 32'b11111111111111111010011010100000;
assign LUT_1[22938] = 32'b11111111111111111100110110110101;
assign LUT_1[22939] = 32'b11111111111111110110001000110001;
assign LUT_1[22940] = 32'b00000000000000001001000001111011;
assign LUT_1[22941] = 32'b00000000000000000010010011110111;
assign LUT_1[22942] = 32'b00000000000000000100110000001100;
assign LUT_1[22943] = 32'b11111111111111111110000010001000;
assign LUT_1[22944] = 32'b00000000000000000000111010001100;
assign LUT_1[22945] = 32'b11111111111111111010001100001000;
assign LUT_1[22946] = 32'b11111111111111111100101000011101;
assign LUT_1[22947] = 32'b11111111111111110101111010011001;
assign LUT_1[22948] = 32'b00000000000000001000110011100011;
assign LUT_1[22949] = 32'b00000000000000000010000101011111;
assign LUT_1[22950] = 32'b00000000000000000100100001110100;
assign LUT_1[22951] = 32'b11111111111111111101110011110000;
assign LUT_1[22952] = 32'b00000000000000000000001000000001;
assign LUT_1[22953] = 32'b11111111111111111001011001111101;
assign LUT_1[22954] = 32'b11111111111111111011110110010010;
assign LUT_1[22955] = 32'b11111111111111110101001000001110;
assign LUT_1[22956] = 32'b00000000000000001000000001011000;
assign LUT_1[22957] = 32'b00000000000000000001010011010100;
assign LUT_1[22958] = 32'b00000000000000000011101111101001;
assign LUT_1[22959] = 32'b11111111111111111101000001100101;
assign LUT_1[22960] = 32'b00000000000000000010110101101110;
assign LUT_1[22961] = 32'b11111111111111111100000111101010;
assign LUT_1[22962] = 32'b11111111111111111110100011111111;
assign LUT_1[22963] = 32'b11111111111111110111110101111011;
assign LUT_1[22964] = 32'b00000000000000001010101111000101;
assign LUT_1[22965] = 32'b00000000000000000100000001000001;
assign LUT_1[22966] = 32'b00000000000000000110011101010110;
assign LUT_1[22967] = 32'b11111111111111111111101111010010;
assign LUT_1[22968] = 32'b00000000000000000010000011100011;
assign LUT_1[22969] = 32'b11111111111111111011010101011111;
assign LUT_1[22970] = 32'b11111111111111111101110001110100;
assign LUT_1[22971] = 32'b11111111111111110111000011110000;
assign LUT_1[22972] = 32'b00000000000000001001111100111010;
assign LUT_1[22973] = 32'b00000000000000000011001110110110;
assign LUT_1[22974] = 32'b00000000000000000101101011001011;
assign LUT_1[22975] = 32'b11111111111111111110111101000111;
assign LUT_1[22976] = 32'b00000000000000000001111100110101;
assign LUT_1[22977] = 32'b11111111111111111011001110110001;
assign LUT_1[22978] = 32'b11111111111111111101101011000110;
assign LUT_1[22979] = 32'b11111111111111110110111101000010;
assign LUT_1[22980] = 32'b00000000000000001001110110001100;
assign LUT_1[22981] = 32'b00000000000000000011001000001000;
assign LUT_1[22982] = 32'b00000000000000000101100100011101;
assign LUT_1[22983] = 32'b11111111111111111110110110011001;
assign LUT_1[22984] = 32'b00000000000000000001001010101010;
assign LUT_1[22985] = 32'b11111111111111111010011100100110;
assign LUT_1[22986] = 32'b11111111111111111100111000111011;
assign LUT_1[22987] = 32'b11111111111111110110001010110111;
assign LUT_1[22988] = 32'b00000000000000001001000100000001;
assign LUT_1[22989] = 32'b00000000000000000010010101111101;
assign LUT_1[22990] = 32'b00000000000000000100110010010010;
assign LUT_1[22991] = 32'b11111111111111111110000100001110;
assign LUT_1[22992] = 32'b00000000000000000011111000010111;
assign LUT_1[22993] = 32'b11111111111111111101001010010011;
assign LUT_1[22994] = 32'b11111111111111111111100110101000;
assign LUT_1[22995] = 32'b11111111111111111000111000100100;
assign LUT_1[22996] = 32'b00000000000000001011110001101110;
assign LUT_1[22997] = 32'b00000000000000000101000011101010;
assign LUT_1[22998] = 32'b00000000000000000111011111111111;
assign LUT_1[22999] = 32'b00000000000000000000110001111011;
assign LUT_1[23000] = 32'b00000000000000000011000110001100;
assign LUT_1[23001] = 32'b11111111111111111100011000001000;
assign LUT_1[23002] = 32'b11111111111111111110110100011101;
assign LUT_1[23003] = 32'b11111111111111111000000110011001;
assign LUT_1[23004] = 32'b00000000000000001010111111100011;
assign LUT_1[23005] = 32'b00000000000000000100010001011111;
assign LUT_1[23006] = 32'b00000000000000000110101101110100;
assign LUT_1[23007] = 32'b11111111111111111111111111110000;
assign LUT_1[23008] = 32'b00000000000000000010110111110100;
assign LUT_1[23009] = 32'b11111111111111111100001001110000;
assign LUT_1[23010] = 32'b11111111111111111110100110000101;
assign LUT_1[23011] = 32'b11111111111111110111111000000001;
assign LUT_1[23012] = 32'b00000000000000001010110001001011;
assign LUT_1[23013] = 32'b00000000000000000100000011000111;
assign LUT_1[23014] = 32'b00000000000000000110011111011100;
assign LUT_1[23015] = 32'b11111111111111111111110001011000;
assign LUT_1[23016] = 32'b00000000000000000010000101101001;
assign LUT_1[23017] = 32'b11111111111111111011010111100101;
assign LUT_1[23018] = 32'b11111111111111111101110011111010;
assign LUT_1[23019] = 32'b11111111111111110111000101110110;
assign LUT_1[23020] = 32'b00000000000000001001111111000000;
assign LUT_1[23021] = 32'b00000000000000000011010000111100;
assign LUT_1[23022] = 32'b00000000000000000101101101010001;
assign LUT_1[23023] = 32'b11111111111111111110111111001101;
assign LUT_1[23024] = 32'b00000000000000000100110011010110;
assign LUT_1[23025] = 32'b11111111111111111110000101010010;
assign LUT_1[23026] = 32'b00000000000000000000100001100111;
assign LUT_1[23027] = 32'b11111111111111111001110011100011;
assign LUT_1[23028] = 32'b00000000000000001100101100101101;
assign LUT_1[23029] = 32'b00000000000000000101111110101001;
assign LUT_1[23030] = 32'b00000000000000001000011010111110;
assign LUT_1[23031] = 32'b00000000000000000001101100111010;
assign LUT_1[23032] = 32'b00000000000000000100000001001011;
assign LUT_1[23033] = 32'b11111111111111111101010011000111;
assign LUT_1[23034] = 32'b11111111111111111111101111011100;
assign LUT_1[23035] = 32'b11111111111111111001000001011000;
assign LUT_1[23036] = 32'b00000000000000001011111010100010;
assign LUT_1[23037] = 32'b00000000000000000101001100011110;
assign LUT_1[23038] = 32'b00000000000000000111101000110011;
assign LUT_1[23039] = 32'b00000000000000000000111010101111;
assign LUT_1[23040] = 32'b11111111111111111000111001011011;
assign LUT_1[23041] = 32'b11111111111111110010001011010111;
assign LUT_1[23042] = 32'b11111111111111110100100111101100;
assign LUT_1[23043] = 32'b11111111111111101101111001101000;
assign LUT_1[23044] = 32'b00000000000000000000110010110010;
assign LUT_1[23045] = 32'b11111111111111111010000100101110;
assign LUT_1[23046] = 32'b11111111111111111100100001000011;
assign LUT_1[23047] = 32'b11111111111111110101110010111111;
assign LUT_1[23048] = 32'b11111111111111111000000111010000;
assign LUT_1[23049] = 32'b11111111111111110001011001001100;
assign LUT_1[23050] = 32'b11111111111111110011110101100001;
assign LUT_1[23051] = 32'b11111111111111101101000111011101;
assign LUT_1[23052] = 32'b00000000000000000000000000100111;
assign LUT_1[23053] = 32'b11111111111111111001010010100011;
assign LUT_1[23054] = 32'b11111111111111111011101110111000;
assign LUT_1[23055] = 32'b11111111111111110101000000110100;
assign LUT_1[23056] = 32'b11111111111111111010110100111101;
assign LUT_1[23057] = 32'b11111111111111110100000110111001;
assign LUT_1[23058] = 32'b11111111111111110110100011001110;
assign LUT_1[23059] = 32'b11111111111111101111110101001010;
assign LUT_1[23060] = 32'b00000000000000000010101110010100;
assign LUT_1[23061] = 32'b11111111111111111100000000010000;
assign LUT_1[23062] = 32'b11111111111111111110011100100101;
assign LUT_1[23063] = 32'b11111111111111110111101110100001;
assign LUT_1[23064] = 32'b11111111111111111010000010110010;
assign LUT_1[23065] = 32'b11111111111111110011010100101110;
assign LUT_1[23066] = 32'b11111111111111110101110001000011;
assign LUT_1[23067] = 32'b11111111111111101111000010111111;
assign LUT_1[23068] = 32'b00000000000000000001111100001001;
assign LUT_1[23069] = 32'b11111111111111111011001110000101;
assign LUT_1[23070] = 32'b11111111111111111101101010011010;
assign LUT_1[23071] = 32'b11111111111111110110111100010110;
assign LUT_1[23072] = 32'b11111111111111111001110100011010;
assign LUT_1[23073] = 32'b11111111111111110011000110010110;
assign LUT_1[23074] = 32'b11111111111111110101100010101011;
assign LUT_1[23075] = 32'b11111111111111101110110100100111;
assign LUT_1[23076] = 32'b00000000000000000001101101110001;
assign LUT_1[23077] = 32'b11111111111111111010111111101101;
assign LUT_1[23078] = 32'b11111111111111111101011100000010;
assign LUT_1[23079] = 32'b11111111111111110110101101111110;
assign LUT_1[23080] = 32'b11111111111111111001000010001111;
assign LUT_1[23081] = 32'b11111111111111110010010100001011;
assign LUT_1[23082] = 32'b11111111111111110100110000100000;
assign LUT_1[23083] = 32'b11111111111111101110000010011100;
assign LUT_1[23084] = 32'b00000000000000000000111011100110;
assign LUT_1[23085] = 32'b11111111111111111010001101100010;
assign LUT_1[23086] = 32'b11111111111111111100101001110111;
assign LUT_1[23087] = 32'b11111111111111110101111011110011;
assign LUT_1[23088] = 32'b11111111111111111011101111111100;
assign LUT_1[23089] = 32'b11111111111111110101000001111000;
assign LUT_1[23090] = 32'b11111111111111110111011110001101;
assign LUT_1[23091] = 32'b11111111111111110000110000001001;
assign LUT_1[23092] = 32'b00000000000000000011101001010011;
assign LUT_1[23093] = 32'b11111111111111111100111011001111;
assign LUT_1[23094] = 32'b11111111111111111111010111100100;
assign LUT_1[23095] = 32'b11111111111111111000101001100000;
assign LUT_1[23096] = 32'b11111111111111111010111101110001;
assign LUT_1[23097] = 32'b11111111111111110100001111101101;
assign LUT_1[23098] = 32'b11111111111111110110101100000010;
assign LUT_1[23099] = 32'b11111111111111101111111101111110;
assign LUT_1[23100] = 32'b00000000000000000010110111001000;
assign LUT_1[23101] = 32'b11111111111111111100001001000100;
assign LUT_1[23102] = 32'b11111111111111111110100101011001;
assign LUT_1[23103] = 32'b11111111111111110111110111010101;
assign LUT_1[23104] = 32'b11111111111111111010110111000011;
assign LUT_1[23105] = 32'b11111111111111110100001000111111;
assign LUT_1[23106] = 32'b11111111111111110110100101010100;
assign LUT_1[23107] = 32'b11111111111111101111110111010000;
assign LUT_1[23108] = 32'b00000000000000000010110000011010;
assign LUT_1[23109] = 32'b11111111111111111100000010010110;
assign LUT_1[23110] = 32'b11111111111111111110011110101011;
assign LUT_1[23111] = 32'b11111111111111110111110000100111;
assign LUT_1[23112] = 32'b11111111111111111010000100111000;
assign LUT_1[23113] = 32'b11111111111111110011010110110100;
assign LUT_1[23114] = 32'b11111111111111110101110011001001;
assign LUT_1[23115] = 32'b11111111111111101111000101000101;
assign LUT_1[23116] = 32'b00000000000000000001111110001111;
assign LUT_1[23117] = 32'b11111111111111111011010000001011;
assign LUT_1[23118] = 32'b11111111111111111101101100100000;
assign LUT_1[23119] = 32'b11111111111111110110111110011100;
assign LUT_1[23120] = 32'b11111111111111111100110010100101;
assign LUT_1[23121] = 32'b11111111111111110110000100100001;
assign LUT_1[23122] = 32'b11111111111111111000100000110110;
assign LUT_1[23123] = 32'b11111111111111110001110010110010;
assign LUT_1[23124] = 32'b00000000000000000100101011111100;
assign LUT_1[23125] = 32'b11111111111111111101111101111000;
assign LUT_1[23126] = 32'b00000000000000000000011010001101;
assign LUT_1[23127] = 32'b11111111111111111001101100001001;
assign LUT_1[23128] = 32'b11111111111111111100000000011010;
assign LUT_1[23129] = 32'b11111111111111110101010010010110;
assign LUT_1[23130] = 32'b11111111111111110111101110101011;
assign LUT_1[23131] = 32'b11111111111111110001000000100111;
assign LUT_1[23132] = 32'b00000000000000000011111001110001;
assign LUT_1[23133] = 32'b11111111111111111101001011101101;
assign LUT_1[23134] = 32'b11111111111111111111101000000010;
assign LUT_1[23135] = 32'b11111111111111111000111001111110;
assign LUT_1[23136] = 32'b11111111111111111011110010000010;
assign LUT_1[23137] = 32'b11111111111111110101000011111110;
assign LUT_1[23138] = 32'b11111111111111110111100000010011;
assign LUT_1[23139] = 32'b11111111111111110000110010001111;
assign LUT_1[23140] = 32'b00000000000000000011101011011001;
assign LUT_1[23141] = 32'b11111111111111111100111101010101;
assign LUT_1[23142] = 32'b11111111111111111111011001101010;
assign LUT_1[23143] = 32'b11111111111111111000101011100110;
assign LUT_1[23144] = 32'b11111111111111111010111111110111;
assign LUT_1[23145] = 32'b11111111111111110100010001110011;
assign LUT_1[23146] = 32'b11111111111111110110101110001000;
assign LUT_1[23147] = 32'b11111111111111110000000000000100;
assign LUT_1[23148] = 32'b00000000000000000010111001001110;
assign LUT_1[23149] = 32'b11111111111111111100001011001010;
assign LUT_1[23150] = 32'b11111111111111111110100111011111;
assign LUT_1[23151] = 32'b11111111111111110111111001011011;
assign LUT_1[23152] = 32'b11111111111111111101101101100100;
assign LUT_1[23153] = 32'b11111111111111110110111111100000;
assign LUT_1[23154] = 32'b11111111111111111001011011110101;
assign LUT_1[23155] = 32'b11111111111111110010101101110001;
assign LUT_1[23156] = 32'b00000000000000000101100110111011;
assign LUT_1[23157] = 32'b11111111111111111110111000110111;
assign LUT_1[23158] = 32'b00000000000000000001010101001100;
assign LUT_1[23159] = 32'b11111111111111111010100111001000;
assign LUT_1[23160] = 32'b11111111111111111100111011011001;
assign LUT_1[23161] = 32'b11111111111111110110001101010101;
assign LUT_1[23162] = 32'b11111111111111111000101001101010;
assign LUT_1[23163] = 32'b11111111111111110001111011100110;
assign LUT_1[23164] = 32'b00000000000000000100110100110000;
assign LUT_1[23165] = 32'b11111111111111111110000110101100;
assign LUT_1[23166] = 32'b00000000000000000000100011000001;
assign LUT_1[23167] = 32'b11111111111111111001110100111101;
assign LUT_1[23168] = 32'b11111111111111111011111001011110;
assign LUT_1[23169] = 32'b11111111111111110101001011011010;
assign LUT_1[23170] = 32'b11111111111111110111100111101111;
assign LUT_1[23171] = 32'b11111111111111110000111001101011;
assign LUT_1[23172] = 32'b00000000000000000011110010110101;
assign LUT_1[23173] = 32'b11111111111111111101000100110001;
assign LUT_1[23174] = 32'b11111111111111111111100001000110;
assign LUT_1[23175] = 32'b11111111111111111000110011000010;
assign LUT_1[23176] = 32'b11111111111111111011000111010011;
assign LUT_1[23177] = 32'b11111111111111110100011001001111;
assign LUT_1[23178] = 32'b11111111111111110110110101100100;
assign LUT_1[23179] = 32'b11111111111111110000000111100000;
assign LUT_1[23180] = 32'b00000000000000000011000000101010;
assign LUT_1[23181] = 32'b11111111111111111100010010100110;
assign LUT_1[23182] = 32'b11111111111111111110101110111011;
assign LUT_1[23183] = 32'b11111111111111111000000000110111;
assign LUT_1[23184] = 32'b11111111111111111101110101000000;
assign LUT_1[23185] = 32'b11111111111111110111000110111100;
assign LUT_1[23186] = 32'b11111111111111111001100011010001;
assign LUT_1[23187] = 32'b11111111111111110010110101001101;
assign LUT_1[23188] = 32'b00000000000000000101101110010111;
assign LUT_1[23189] = 32'b11111111111111111111000000010011;
assign LUT_1[23190] = 32'b00000000000000000001011100101000;
assign LUT_1[23191] = 32'b11111111111111111010101110100100;
assign LUT_1[23192] = 32'b11111111111111111101000010110101;
assign LUT_1[23193] = 32'b11111111111111110110010100110001;
assign LUT_1[23194] = 32'b11111111111111111000110001000110;
assign LUT_1[23195] = 32'b11111111111111110010000011000010;
assign LUT_1[23196] = 32'b00000000000000000100111100001100;
assign LUT_1[23197] = 32'b11111111111111111110001110001000;
assign LUT_1[23198] = 32'b00000000000000000000101010011101;
assign LUT_1[23199] = 32'b11111111111111111001111100011001;
assign LUT_1[23200] = 32'b11111111111111111100110100011101;
assign LUT_1[23201] = 32'b11111111111111110110000110011001;
assign LUT_1[23202] = 32'b11111111111111111000100010101110;
assign LUT_1[23203] = 32'b11111111111111110001110100101010;
assign LUT_1[23204] = 32'b00000000000000000100101101110100;
assign LUT_1[23205] = 32'b11111111111111111101111111110000;
assign LUT_1[23206] = 32'b00000000000000000000011100000101;
assign LUT_1[23207] = 32'b11111111111111111001101110000001;
assign LUT_1[23208] = 32'b11111111111111111100000010010010;
assign LUT_1[23209] = 32'b11111111111111110101010100001110;
assign LUT_1[23210] = 32'b11111111111111110111110000100011;
assign LUT_1[23211] = 32'b11111111111111110001000010011111;
assign LUT_1[23212] = 32'b00000000000000000011111011101001;
assign LUT_1[23213] = 32'b11111111111111111101001101100101;
assign LUT_1[23214] = 32'b11111111111111111111101001111010;
assign LUT_1[23215] = 32'b11111111111111111000111011110110;
assign LUT_1[23216] = 32'b11111111111111111110101111111111;
assign LUT_1[23217] = 32'b11111111111111111000000001111011;
assign LUT_1[23218] = 32'b11111111111111111010011110010000;
assign LUT_1[23219] = 32'b11111111111111110011110000001100;
assign LUT_1[23220] = 32'b00000000000000000110101001010110;
assign LUT_1[23221] = 32'b11111111111111111111111011010010;
assign LUT_1[23222] = 32'b00000000000000000010010111100111;
assign LUT_1[23223] = 32'b11111111111111111011101001100011;
assign LUT_1[23224] = 32'b11111111111111111101111101110100;
assign LUT_1[23225] = 32'b11111111111111110111001111110000;
assign LUT_1[23226] = 32'b11111111111111111001101100000101;
assign LUT_1[23227] = 32'b11111111111111110010111110000001;
assign LUT_1[23228] = 32'b00000000000000000101110111001011;
assign LUT_1[23229] = 32'b11111111111111111111001001000111;
assign LUT_1[23230] = 32'b00000000000000000001100101011100;
assign LUT_1[23231] = 32'b11111111111111111010110111011000;
assign LUT_1[23232] = 32'b11111111111111111101110111000110;
assign LUT_1[23233] = 32'b11111111111111110111001001000010;
assign LUT_1[23234] = 32'b11111111111111111001100101010111;
assign LUT_1[23235] = 32'b11111111111111110010110111010011;
assign LUT_1[23236] = 32'b00000000000000000101110000011101;
assign LUT_1[23237] = 32'b11111111111111111111000010011001;
assign LUT_1[23238] = 32'b00000000000000000001011110101110;
assign LUT_1[23239] = 32'b11111111111111111010110000101010;
assign LUT_1[23240] = 32'b11111111111111111101000100111011;
assign LUT_1[23241] = 32'b11111111111111110110010110110111;
assign LUT_1[23242] = 32'b11111111111111111000110011001100;
assign LUT_1[23243] = 32'b11111111111111110010000101001000;
assign LUT_1[23244] = 32'b00000000000000000100111110010010;
assign LUT_1[23245] = 32'b11111111111111111110010000001110;
assign LUT_1[23246] = 32'b00000000000000000000101100100011;
assign LUT_1[23247] = 32'b11111111111111111001111110011111;
assign LUT_1[23248] = 32'b11111111111111111111110010101000;
assign LUT_1[23249] = 32'b11111111111111111001000100100100;
assign LUT_1[23250] = 32'b11111111111111111011100000111001;
assign LUT_1[23251] = 32'b11111111111111110100110010110101;
assign LUT_1[23252] = 32'b00000000000000000111101011111111;
assign LUT_1[23253] = 32'b00000000000000000000111101111011;
assign LUT_1[23254] = 32'b00000000000000000011011010010000;
assign LUT_1[23255] = 32'b11111111111111111100101100001100;
assign LUT_1[23256] = 32'b11111111111111111111000000011101;
assign LUT_1[23257] = 32'b11111111111111111000010010011001;
assign LUT_1[23258] = 32'b11111111111111111010101110101110;
assign LUT_1[23259] = 32'b11111111111111110100000000101010;
assign LUT_1[23260] = 32'b00000000000000000110111001110100;
assign LUT_1[23261] = 32'b00000000000000000000001011110000;
assign LUT_1[23262] = 32'b00000000000000000010101000000101;
assign LUT_1[23263] = 32'b11111111111111111011111010000001;
assign LUT_1[23264] = 32'b11111111111111111110110010000101;
assign LUT_1[23265] = 32'b11111111111111111000000100000001;
assign LUT_1[23266] = 32'b11111111111111111010100000010110;
assign LUT_1[23267] = 32'b11111111111111110011110010010010;
assign LUT_1[23268] = 32'b00000000000000000110101011011100;
assign LUT_1[23269] = 32'b11111111111111111111111101011000;
assign LUT_1[23270] = 32'b00000000000000000010011001101101;
assign LUT_1[23271] = 32'b11111111111111111011101011101001;
assign LUT_1[23272] = 32'b11111111111111111101111111111010;
assign LUT_1[23273] = 32'b11111111111111110111010001110110;
assign LUT_1[23274] = 32'b11111111111111111001101110001011;
assign LUT_1[23275] = 32'b11111111111111110011000000000111;
assign LUT_1[23276] = 32'b00000000000000000101111001010001;
assign LUT_1[23277] = 32'b11111111111111111111001011001101;
assign LUT_1[23278] = 32'b00000000000000000001100111100010;
assign LUT_1[23279] = 32'b11111111111111111010111001011110;
assign LUT_1[23280] = 32'b00000000000000000000101101100111;
assign LUT_1[23281] = 32'b11111111111111111001111111100011;
assign LUT_1[23282] = 32'b11111111111111111100011011111000;
assign LUT_1[23283] = 32'b11111111111111110101101101110100;
assign LUT_1[23284] = 32'b00000000000000001000100110111110;
assign LUT_1[23285] = 32'b00000000000000000001111000111010;
assign LUT_1[23286] = 32'b00000000000000000100010101001111;
assign LUT_1[23287] = 32'b11111111111111111101100111001011;
assign LUT_1[23288] = 32'b11111111111111111111111011011100;
assign LUT_1[23289] = 32'b11111111111111111001001101011000;
assign LUT_1[23290] = 32'b11111111111111111011101001101101;
assign LUT_1[23291] = 32'b11111111111111110100111011101001;
assign LUT_1[23292] = 32'b00000000000000000111110100110011;
assign LUT_1[23293] = 32'b00000000000000000001000110101111;
assign LUT_1[23294] = 32'b00000000000000000011100011000100;
assign LUT_1[23295] = 32'b11111111111111111100110101000000;
assign LUT_1[23296] = 32'b11111111111111110110101101100111;
assign LUT_1[23297] = 32'b11111111111111101111111111100011;
assign LUT_1[23298] = 32'b11111111111111110010011011111000;
assign LUT_1[23299] = 32'b11111111111111101011101101110100;
assign LUT_1[23300] = 32'b11111111111111111110100110111110;
assign LUT_1[23301] = 32'b11111111111111110111111000111010;
assign LUT_1[23302] = 32'b11111111111111111010010101001111;
assign LUT_1[23303] = 32'b11111111111111110011100111001011;
assign LUT_1[23304] = 32'b11111111111111110101111011011100;
assign LUT_1[23305] = 32'b11111111111111101111001101011000;
assign LUT_1[23306] = 32'b11111111111111110001101001101101;
assign LUT_1[23307] = 32'b11111111111111101010111011101001;
assign LUT_1[23308] = 32'b11111111111111111101110100110011;
assign LUT_1[23309] = 32'b11111111111111110111000110101111;
assign LUT_1[23310] = 32'b11111111111111111001100011000100;
assign LUT_1[23311] = 32'b11111111111111110010110101000000;
assign LUT_1[23312] = 32'b11111111111111111000101001001001;
assign LUT_1[23313] = 32'b11111111111111110001111011000101;
assign LUT_1[23314] = 32'b11111111111111110100010111011010;
assign LUT_1[23315] = 32'b11111111111111101101101001010110;
assign LUT_1[23316] = 32'b00000000000000000000100010100000;
assign LUT_1[23317] = 32'b11111111111111111001110100011100;
assign LUT_1[23318] = 32'b11111111111111111100010000110001;
assign LUT_1[23319] = 32'b11111111111111110101100010101101;
assign LUT_1[23320] = 32'b11111111111111110111110110111110;
assign LUT_1[23321] = 32'b11111111111111110001001000111010;
assign LUT_1[23322] = 32'b11111111111111110011100101001111;
assign LUT_1[23323] = 32'b11111111111111101100110111001011;
assign LUT_1[23324] = 32'b11111111111111111111110000010101;
assign LUT_1[23325] = 32'b11111111111111111001000010010001;
assign LUT_1[23326] = 32'b11111111111111111011011110100110;
assign LUT_1[23327] = 32'b11111111111111110100110000100010;
assign LUT_1[23328] = 32'b11111111111111110111101000100110;
assign LUT_1[23329] = 32'b11111111111111110000111010100010;
assign LUT_1[23330] = 32'b11111111111111110011010110110111;
assign LUT_1[23331] = 32'b11111111111111101100101000110011;
assign LUT_1[23332] = 32'b11111111111111111111100001111101;
assign LUT_1[23333] = 32'b11111111111111111000110011111001;
assign LUT_1[23334] = 32'b11111111111111111011010000001110;
assign LUT_1[23335] = 32'b11111111111111110100100010001010;
assign LUT_1[23336] = 32'b11111111111111110110110110011011;
assign LUT_1[23337] = 32'b11111111111111110000001000010111;
assign LUT_1[23338] = 32'b11111111111111110010100100101100;
assign LUT_1[23339] = 32'b11111111111111101011110110101000;
assign LUT_1[23340] = 32'b11111111111111111110101111110010;
assign LUT_1[23341] = 32'b11111111111111111000000001101110;
assign LUT_1[23342] = 32'b11111111111111111010011110000011;
assign LUT_1[23343] = 32'b11111111111111110011101111111111;
assign LUT_1[23344] = 32'b11111111111111111001100100001000;
assign LUT_1[23345] = 32'b11111111111111110010110110000100;
assign LUT_1[23346] = 32'b11111111111111110101010010011001;
assign LUT_1[23347] = 32'b11111111111111101110100100010101;
assign LUT_1[23348] = 32'b00000000000000000001011101011111;
assign LUT_1[23349] = 32'b11111111111111111010101111011011;
assign LUT_1[23350] = 32'b11111111111111111101001011110000;
assign LUT_1[23351] = 32'b11111111111111110110011101101100;
assign LUT_1[23352] = 32'b11111111111111111000110001111101;
assign LUT_1[23353] = 32'b11111111111111110010000011111001;
assign LUT_1[23354] = 32'b11111111111111110100100000001110;
assign LUT_1[23355] = 32'b11111111111111101101110010001010;
assign LUT_1[23356] = 32'b00000000000000000000101011010100;
assign LUT_1[23357] = 32'b11111111111111111001111101010000;
assign LUT_1[23358] = 32'b11111111111111111100011001100101;
assign LUT_1[23359] = 32'b11111111111111110101101011100001;
assign LUT_1[23360] = 32'b11111111111111111000101011001111;
assign LUT_1[23361] = 32'b11111111111111110001111101001011;
assign LUT_1[23362] = 32'b11111111111111110100011001100000;
assign LUT_1[23363] = 32'b11111111111111101101101011011100;
assign LUT_1[23364] = 32'b00000000000000000000100100100110;
assign LUT_1[23365] = 32'b11111111111111111001110110100010;
assign LUT_1[23366] = 32'b11111111111111111100010010110111;
assign LUT_1[23367] = 32'b11111111111111110101100100110011;
assign LUT_1[23368] = 32'b11111111111111110111111001000100;
assign LUT_1[23369] = 32'b11111111111111110001001011000000;
assign LUT_1[23370] = 32'b11111111111111110011100111010101;
assign LUT_1[23371] = 32'b11111111111111101100111001010001;
assign LUT_1[23372] = 32'b11111111111111111111110010011011;
assign LUT_1[23373] = 32'b11111111111111111001000100010111;
assign LUT_1[23374] = 32'b11111111111111111011100000101100;
assign LUT_1[23375] = 32'b11111111111111110100110010101000;
assign LUT_1[23376] = 32'b11111111111111111010100110110001;
assign LUT_1[23377] = 32'b11111111111111110011111000101101;
assign LUT_1[23378] = 32'b11111111111111110110010101000010;
assign LUT_1[23379] = 32'b11111111111111101111100110111110;
assign LUT_1[23380] = 32'b00000000000000000010100000001000;
assign LUT_1[23381] = 32'b11111111111111111011110010000100;
assign LUT_1[23382] = 32'b11111111111111111110001110011001;
assign LUT_1[23383] = 32'b11111111111111110111100000010101;
assign LUT_1[23384] = 32'b11111111111111111001110100100110;
assign LUT_1[23385] = 32'b11111111111111110011000110100010;
assign LUT_1[23386] = 32'b11111111111111110101100010110111;
assign LUT_1[23387] = 32'b11111111111111101110110100110011;
assign LUT_1[23388] = 32'b00000000000000000001101101111101;
assign LUT_1[23389] = 32'b11111111111111111010111111111001;
assign LUT_1[23390] = 32'b11111111111111111101011100001110;
assign LUT_1[23391] = 32'b11111111111111110110101110001010;
assign LUT_1[23392] = 32'b11111111111111111001100110001110;
assign LUT_1[23393] = 32'b11111111111111110010111000001010;
assign LUT_1[23394] = 32'b11111111111111110101010100011111;
assign LUT_1[23395] = 32'b11111111111111101110100110011011;
assign LUT_1[23396] = 32'b00000000000000000001011111100101;
assign LUT_1[23397] = 32'b11111111111111111010110001100001;
assign LUT_1[23398] = 32'b11111111111111111101001101110110;
assign LUT_1[23399] = 32'b11111111111111110110011111110010;
assign LUT_1[23400] = 32'b11111111111111111000110100000011;
assign LUT_1[23401] = 32'b11111111111111110010000101111111;
assign LUT_1[23402] = 32'b11111111111111110100100010010100;
assign LUT_1[23403] = 32'b11111111111111101101110100010000;
assign LUT_1[23404] = 32'b00000000000000000000101101011010;
assign LUT_1[23405] = 32'b11111111111111111001111111010110;
assign LUT_1[23406] = 32'b11111111111111111100011011101011;
assign LUT_1[23407] = 32'b11111111111111110101101101100111;
assign LUT_1[23408] = 32'b11111111111111111011100001110000;
assign LUT_1[23409] = 32'b11111111111111110100110011101100;
assign LUT_1[23410] = 32'b11111111111111110111010000000001;
assign LUT_1[23411] = 32'b11111111111111110000100001111101;
assign LUT_1[23412] = 32'b00000000000000000011011011000111;
assign LUT_1[23413] = 32'b11111111111111111100101101000011;
assign LUT_1[23414] = 32'b11111111111111111111001001011000;
assign LUT_1[23415] = 32'b11111111111111111000011011010100;
assign LUT_1[23416] = 32'b11111111111111111010101111100101;
assign LUT_1[23417] = 32'b11111111111111110100000001100001;
assign LUT_1[23418] = 32'b11111111111111110110011101110110;
assign LUT_1[23419] = 32'b11111111111111101111101111110010;
assign LUT_1[23420] = 32'b00000000000000000010101000111100;
assign LUT_1[23421] = 32'b11111111111111111011111010111000;
assign LUT_1[23422] = 32'b11111111111111111110010111001101;
assign LUT_1[23423] = 32'b11111111111111110111101001001001;
assign LUT_1[23424] = 32'b11111111111111111001101101101010;
assign LUT_1[23425] = 32'b11111111111111110010111111100110;
assign LUT_1[23426] = 32'b11111111111111110101011011111011;
assign LUT_1[23427] = 32'b11111111111111101110101101110111;
assign LUT_1[23428] = 32'b00000000000000000001100111000001;
assign LUT_1[23429] = 32'b11111111111111111010111000111101;
assign LUT_1[23430] = 32'b11111111111111111101010101010010;
assign LUT_1[23431] = 32'b11111111111111110110100111001110;
assign LUT_1[23432] = 32'b11111111111111111000111011011111;
assign LUT_1[23433] = 32'b11111111111111110010001101011011;
assign LUT_1[23434] = 32'b11111111111111110100101001110000;
assign LUT_1[23435] = 32'b11111111111111101101111011101100;
assign LUT_1[23436] = 32'b00000000000000000000110100110110;
assign LUT_1[23437] = 32'b11111111111111111010000110110010;
assign LUT_1[23438] = 32'b11111111111111111100100011000111;
assign LUT_1[23439] = 32'b11111111111111110101110101000011;
assign LUT_1[23440] = 32'b11111111111111111011101001001100;
assign LUT_1[23441] = 32'b11111111111111110100111011001000;
assign LUT_1[23442] = 32'b11111111111111110111010111011101;
assign LUT_1[23443] = 32'b11111111111111110000101001011001;
assign LUT_1[23444] = 32'b00000000000000000011100010100011;
assign LUT_1[23445] = 32'b11111111111111111100110100011111;
assign LUT_1[23446] = 32'b11111111111111111111010000110100;
assign LUT_1[23447] = 32'b11111111111111111000100010110000;
assign LUT_1[23448] = 32'b11111111111111111010110111000001;
assign LUT_1[23449] = 32'b11111111111111110100001000111101;
assign LUT_1[23450] = 32'b11111111111111110110100101010010;
assign LUT_1[23451] = 32'b11111111111111101111110111001110;
assign LUT_1[23452] = 32'b00000000000000000010110000011000;
assign LUT_1[23453] = 32'b11111111111111111100000010010100;
assign LUT_1[23454] = 32'b11111111111111111110011110101001;
assign LUT_1[23455] = 32'b11111111111111110111110000100101;
assign LUT_1[23456] = 32'b11111111111111111010101000101001;
assign LUT_1[23457] = 32'b11111111111111110011111010100101;
assign LUT_1[23458] = 32'b11111111111111110110010110111010;
assign LUT_1[23459] = 32'b11111111111111101111101000110110;
assign LUT_1[23460] = 32'b00000000000000000010100010000000;
assign LUT_1[23461] = 32'b11111111111111111011110011111100;
assign LUT_1[23462] = 32'b11111111111111111110010000010001;
assign LUT_1[23463] = 32'b11111111111111110111100010001101;
assign LUT_1[23464] = 32'b11111111111111111001110110011110;
assign LUT_1[23465] = 32'b11111111111111110011001000011010;
assign LUT_1[23466] = 32'b11111111111111110101100100101111;
assign LUT_1[23467] = 32'b11111111111111101110110110101011;
assign LUT_1[23468] = 32'b00000000000000000001101111110101;
assign LUT_1[23469] = 32'b11111111111111111011000001110001;
assign LUT_1[23470] = 32'b11111111111111111101011110000110;
assign LUT_1[23471] = 32'b11111111111111110110110000000010;
assign LUT_1[23472] = 32'b11111111111111111100100100001011;
assign LUT_1[23473] = 32'b11111111111111110101110110000111;
assign LUT_1[23474] = 32'b11111111111111111000010010011100;
assign LUT_1[23475] = 32'b11111111111111110001100100011000;
assign LUT_1[23476] = 32'b00000000000000000100011101100010;
assign LUT_1[23477] = 32'b11111111111111111101101111011110;
assign LUT_1[23478] = 32'b00000000000000000000001011110011;
assign LUT_1[23479] = 32'b11111111111111111001011101101111;
assign LUT_1[23480] = 32'b11111111111111111011110010000000;
assign LUT_1[23481] = 32'b11111111111111110101000011111100;
assign LUT_1[23482] = 32'b11111111111111110111100000010001;
assign LUT_1[23483] = 32'b11111111111111110000110010001101;
assign LUT_1[23484] = 32'b00000000000000000011101011010111;
assign LUT_1[23485] = 32'b11111111111111111100111101010011;
assign LUT_1[23486] = 32'b11111111111111111111011001101000;
assign LUT_1[23487] = 32'b11111111111111111000101011100100;
assign LUT_1[23488] = 32'b11111111111111111011101011010010;
assign LUT_1[23489] = 32'b11111111111111110100111101001110;
assign LUT_1[23490] = 32'b11111111111111110111011001100011;
assign LUT_1[23491] = 32'b11111111111111110000101011011111;
assign LUT_1[23492] = 32'b00000000000000000011100100101001;
assign LUT_1[23493] = 32'b11111111111111111100110110100101;
assign LUT_1[23494] = 32'b11111111111111111111010010111010;
assign LUT_1[23495] = 32'b11111111111111111000100100110110;
assign LUT_1[23496] = 32'b11111111111111111010111001000111;
assign LUT_1[23497] = 32'b11111111111111110100001011000011;
assign LUT_1[23498] = 32'b11111111111111110110100111011000;
assign LUT_1[23499] = 32'b11111111111111101111111001010100;
assign LUT_1[23500] = 32'b00000000000000000010110010011110;
assign LUT_1[23501] = 32'b11111111111111111100000100011010;
assign LUT_1[23502] = 32'b11111111111111111110100000101111;
assign LUT_1[23503] = 32'b11111111111111110111110010101011;
assign LUT_1[23504] = 32'b11111111111111111101100110110100;
assign LUT_1[23505] = 32'b11111111111111110110111000110000;
assign LUT_1[23506] = 32'b11111111111111111001010101000101;
assign LUT_1[23507] = 32'b11111111111111110010100111000001;
assign LUT_1[23508] = 32'b00000000000000000101100000001011;
assign LUT_1[23509] = 32'b11111111111111111110110010000111;
assign LUT_1[23510] = 32'b00000000000000000001001110011100;
assign LUT_1[23511] = 32'b11111111111111111010100000011000;
assign LUT_1[23512] = 32'b11111111111111111100110100101001;
assign LUT_1[23513] = 32'b11111111111111110110000110100101;
assign LUT_1[23514] = 32'b11111111111111111000100010111010;
assign LUT_1[23515] = 32'b11111111111111110001110100110110;
assign LUT_1[23516] = 32'b00000000000000000100101110000000;
assign LUT_1[23517] = 32'b11111111111111111101111111111100;
assign LUT_1[23518] = 32'b00000000000000000000011100010001;
assign LUT_1[23519] = 32'b11111111111111111001101110001101;
assign LUT_1[23520] = 32'b11111111111111111100100110010001;
assign LUT_1[23521] = 32'b11111111111111110101111000001101;
assign LUT_1[23522] = 32'b11111111111111111000010100100010;
assign LUT_1[23523] = 32'b11111111111111110001100110011110;
assign LUT_1[23524] = 32'b00000000000000000100011111101000;
assign LUT_1[23525] = 32'b11111111111111111101110001100100;
assign LUT_1[23526] = 32'b00000000000000000000001101111001;
assign LUT_1[23527] = 32'b11111111111111111001011111110101;
assign LUT_1[23528] = 32'b11111111111111111011110100000110;
assign LUT_1[23529] = 32'b11111111111111110101000110000010;
assign LUT_1[23530] = 32'b11111111111111110111100010010111;
assign LUT_1[23531] = 32'b11111111111111110000110100010011;
assign LUT_1[23532] = 32'b00000000000000000011101101011101;
assign LUT_1[23533] = 32'b11111111111111111100111111011001;
assign LUT_1[23534] = 32'b11111111111111111111011011101110;
assign LUT_1[23535] = 32'b11111111111111111000101101101010;
assign LUT_1[23536] = 32'b11111111111111111110100001110011;
assign LUT_1[23537] = 32'b11111111111111110111110011101111;
assign LUT_1[23538] = 32'b11111111111111111010010000000100;
assign LUT_1[23539] = 32'b11111111111111110011100010000000;
assign LUT_1[23540] = 32'b00000000000000000110011011001010;
assign LUT_1[23541] = 32'b11111111111111111111101101000110;
assign LUT_1[23542] = 32'b00000000000000000010001001011011;
assign LUT_1[23543] = 32'b11111111111111111011011011010111;
assign LUT_1[23544] = 32'b11111111111111111101101111101000;
assign LUT_1[23545] = 32'b11111111111111110111000001100100;
assign LUT_1[23546] = 32'b11111111111111111001011101111001;
assign LUT_1[23547] = 32'b11111111111111110010101111110101;
assign LUT_1[23548] = 32'b00000000000000000101101000111111;
assign LUT_1[23549] = 32'b11111111111111111110111010111011;
assign LUT_1[23550] = 32'b00000000000000000001010111010000;
assign LUT_1[23551] = 32'b11111111111111111010101001001100;
assign LUT_1[23552] = 32'b00000000000000000101100001101110;
assign LUT_1[23553] = 32'b11111111111111111110110011101010;
assign LUT_1[23554] = 32'b00000000000000000001001111111111;
assign LUT_1[23555] = 32'b11111111111111111010100001111011;
assign LUT_1[23556] = 32'b00000000000000001101011011000101;
assign LUT_1[23557] = 32'b00000000000000000110101101000001;
assign LUT_1[23558] = 32'b00000000000000001001001001010110;
assign LUT_1[23559] = 32'b00000000000000000010011011010010;
assign LUT_1[23560] = 32'b00000000000000000100101111100011;
assign LUT_1[23561] = 32'b11111111111111111110000001011111;
assign LUT_1[23562] = 32'b00000000000000000000011101110100;
assign LUT_1[23563] = 32'b11111111111111111001101111110000;
assign LUT_1[23564] = 32'b00000000000000001100101000111010;
assign LUT_1[23565] = 32'b00000000000000000101111010110110;
assign LUT_1[23566] = 32'b00000000000000001000010111001011;
assign LUT_1[23567] = 32'b00000000000000000001101001000111;
assign LUT_1[23568] = 32'b00000000000000000111011101010000;
assign LUT_1[23569] = 32'b00000000000000000000101111001100;
assign LUT_1[23570] = 32'b00000000000000000011001011100001;
assign LUT_1[23571] = 32'b11111111111111111100011101011101;
assign LUT_1[23572] = 32'b00000000000000001111010110100111;
assign LUT_1[23573] = 32'b00000000000000001000101000100011;
assign LUT_1[23574] = 32'b00000000000000001011000100111000;
assign LUT_1[23575] = 32'b00000000000000000100010110110100;
assign LUT_1[23576] = 32'b00000000000000000110101011000101;
assign LUT_1[23577] = 32'b11111111111111111111111101000001;
assign LUT_1[23578] = 32'b00000000000000000010011001010110;
assign LUT_1[23579] = 32'b11111111111111111011101011010010;
assign LUT_1[23580] = 32'b00000000000000001110100100011100;
assign LUT_1[23581] = 32'b00000000000000000111110110011000;
assign LUT_1[23582] = 32'b00000000000000001010010010101101;
assign LUT_1[23583] = 32'b00000000000000000011100100101001;
assign LUT_1[23584] = 32'b00000000000000000110011100101101;
assign LUT_1[23585] = 32'b11111111111111111111101110101001;
assign LUT_1[23586] = 32'b00000000000000000010001010111110;
assign LUT_1[23587] = 32'b11111111111111111011011100111010;
assign LUT_1[23588] = 32'b00000000000000001110010110000100;
assign LUT_1[23589] = 32'b00000000000000000111101000000000;
assign LUT_1[23590] = 32'b00000000000000001010000100010101;
assign LUT_1[23591] = 32'b00000000000000000011010110010001;
assign LUT_1[23592] = 32'b00000000000000000101101010100010;
assign LUT_1[23593] = 32'b11111111111111111110111100011110;
assign LUT_1[23594] = 32'b00000000000000000001011000110011;
assign LUT_1[23595] = 32'b11111111111111111010101010101111;
assign LUT_1[23596] = 32'b00000000000000001101100011111001;
assign LUT_1[23597] = 32'b00000000000000000110110101110101;
assign LUT_1[23598] = 32'b00000000000000001001010010001010;
assign LUT_1[23599] = 32'b00000000000000000010100100000110;
assign LUT_1[23600] = 32'b00000000000000001000011000001111;
assign LUT_1[23601] = 32'b00000000000000000001101010001011;
assign LUT_1[23602] = 32'b00000000000000000100000110100000;
assign LUT_1[23603] = 32'b11111111111111111101011000011100;
assign LUT_1[23604] = 32'b00000000000000010000010001100110;
assign LUT_1[23605] = 32'b00000000000000001001100011100010;
assign LUT_1[23606] = 32'b00000000000000001011111111110111;
assign LUT_1[23607] = 32'b00000000000000000101010001110011;
assign LUT_1[23608] = 32'b00000000000000000111100110000100;
assign LUT_1[23609] = 32'b00000000000000000000111000000000;
assign LUT_1[23610] = 32'b00000000000000000011010100010101;
assign LUT_1[23611] = 32'b11111111111111111100100110010001;
assign LUT_1[23612] = 32'b00000000000000001111011111011011;
assign LUT_1[23613] = 32'b00000000000000001000110001010111;
assign LUT_1[23614] = 32'b00000000000000001011001101101100;
assign LUT_1[23615] = 32'b00000000000000000100011111101000;
assign LUT_1[23616] = 32'b00000000000000000111011111010110;
assign LUT_1[23617] = 32'b00000000000000000000110001010010;
assign LUT_1[23618] = 32'b00000000000000000011001101100111;
assign LUT_1[23619] = 32'b11111111111111111100011111100011;
assign LUT_1[23620] = 32'b00000000000000001111011000101101;
assign LUT_1[23621] = 32'b00000000000000001000101010101001;
assign LUT_1[23622] = 32'b00000000000000001011000110111110;
assign LUT_1[23623] = 32'b00000000000000000100011000111010;
assign LUT_1[23624] = 32'b00000000000000000110101101001011;
assign LUT_1[23625] = 32'b11111111111111111111111111000111;
assign LUT_1[23626] = 32'b00000000000000000010011011011100;
assign LUT_1[23627] = 32'b11111111111111111011101101011000;
assign LUT_1[23628] = 32'b00000000000000001110100110100010;
assign LUT_1[23629] = 32'b00000000000000000111111000011110;
assign LUT_1[23630] = 32'b00000000000000001010010100110011;
assign LUT_1[23631] = 32'b00000000000000000011100110101111;
assign LUT_1[23632] = 32'b00000000000000001001011010111000;
assign LUT_1[23633] = 32'b00000000000000000010101100110100;
assign LUT_1[23634] = 32'b00000000000000000101001001001001;
assign LUT_1[23635] = 32'b11111111111111111110011011000101;
assign LUT_1[23636] = 32'b00000000000000010001010100001111;
assign LUT_1[23637] = 32'b00000000000000001010100110001011;
assign LUT_1[23638] = 32'b00000000000000001101000010100000;
assign LUT_1[23639] = 32'b00000000000000000110010100011100;
assign LUT_1[23640] = 32'b00000000000000001000101000101101;
assign LUT_1[23641] = 32'b00000000000000000001111010101001;
assign LUT_1[23642] = 32'b00000000000000000100010110111110;
assign LUT_1[23643] = 32'b11111111111111111101101000111010;
assign LUT_1[23644] = 32'b00000000000000010000100010000100;
assign LUT_1[23645] = 32'b00000000000000001001110100000000;
assign LUT_1[23646] = 32'b00000000000000001100010000010101;
assign LUT_1[23647] = 32'b00000000000000000101100010010001;
assign LUT_1[23648] = 32'b00000000000000001000011010010101;
assign LUT_1[23649] = 32'b00000000000000000001101100010001;
assign LUT_1[23650] = 32'b00000000000000000100001000100110;
assign LUT_1[23651] = 32'b11111111111111111101011010100010;
assign LUT_1[23652] = 32'b00000000000000010000010011101100;
assign LUT_1[23653] = 32'b00000000000000001001100101101000;
assign LUT_1[23654] = 32'b00000000000000001100000001111101;
assign LUT_1[23655] = 32'b00000000000000000101010011111001;
assign LUT_1[23656] = 32'b00000000000000000111101000001010;
assign LUT_1[23657] = 32'b00000000000000000000111010000110;
assign LUT_1[23658] = 32'b00000000000000000011010110011011;
assign LUT_1[23659] = 32'b11111111111111111100101000010111;
assign LUT_1[23660] = 32'b00000000000000001111100001100001;
assign LUT_1[23661] = 32'b00000000000000001000110011011101;
assign LUT_1[23662] = 32'b00000000000000001011001111110010;
assign LUT_1[23663] = 32'b00000000000000000100100001101110;
assign LUT_1[23664] = 32'b00000000000000001010010101110111;
assign LUT_1[23665] = 32'b00000000000000000011100111110011;
assign LUT_1[23666] = 32'b00000000000000000110000100001000;
assign LUT_1[23667] = 32'b11111111111111111111010110000100;
assign LUT_1[23668] = 32'b00000000000000010010001111001110;
assign LUT_1[23669] = 32'b00000000000000001011100001001010;
assign LUT_1[23670] = 32'b00000000000000001101111101011111;
assign LUT_1[23671] = 32'b00000000000000000111001111011011;
assign LUT_1[23672] = 32'b00000000000000001001100011101100;
assign LUT_1[23673] = 32'b00000000000000000010110101101000;
assign LUT_1[23674] = 32'b00000000000000000101010001111101;
assign LUT_1[23675] = 32'b11111111111111111110100011111001;
assign LUT_1[23676] = 32'b00000000000000010001011101000011;
assign LUT_1[23677] = 32'b00000000000000001010101110111111;
assign LUT_1[23678] = 32'b00000000000000001101001011010100;
assign LUT_1[23679] = 32'b00000000000000000110011101010000;
assign LUT_1[23680] = 32'b00000000000000001000100001110001;
assign LUT_1[23681] = 32'b00000000000000000001110011101101;
assign LUT_1[23682] = 32'b00000000000000000100010000000010;
assign LUT_1[23683] = 32'b11111111111111111101100001111110;
assign LUT_1[23684] = 32'b00000000000000010000011011001000;
assign LUT_1[23685] = 32'b00000000000000001001101101000100;
assign LUT_1[23686] = 32'b00000000000000001100001001011001;
assign LUT_1[23687] = 32'b00000000000000000101011011010101;
assign LUT_1[23688] = 32'b00000000000000000111101111100110;
assign LUT_1[23689] = 32'b00000000000000000001000001100010;
assign LUT_1[23690] = 32'b00000000000000000011011101110111;
assign LUT_1[23691] = 32'b11111111111111111100101111110011;
assign LUT_1[23692] = 32'b00000000000000001111101000111101;
assign LUT_1[23693] = 32'b00000000000000001000111010111001;
assign LUT_1[23694] = 32'b00000000000000001011010111001110;
assign LUT_1[23695] = 32'b00000000000000000100101001001010;
assign LUT_1[23696] = 32'b00000000000000001010011101010011;
assign LUT_1[23697] = 32'b00000000000000000011101111001111;
assign LUT_1[23698] = 32'b00000000000000000110001011100100;
assign LUT_1[23699] = 32'b11111111111111111111011101100000;
assign LUT_1[23700] = 32'b00000000000000010010010110101010;
assign LUT_1[23701] = 32'b00000000000000001011101000100110;
assign LUT_1[23702] = 32'b00000000000000001110000100111011;
assign LUT_1[23703] = 32'b00000000000000000111010110110111;
assign LUT_1[23704] = 32'b00000000000000001001101011001000;
assign LUT_1[23705] = 32'b00000000000000000010111101000100;
assign LUT_1[23706] = 32'b00000000000000000101011001011001;
assign LUT_1[23707] = 32'b11111111111111111110101011010101;
assign LUT_1[23708] = 32'b00000000000000010001100100011111;
assign LUT_1[23709] = 32'b00000000000000001010110110011011;
assign LUT_1[23710] = 32'b00000000000000001101010010110000;
assign LUT_1[23711] = 32'b00000000000000000110100100101100;
assign LUT_1[23712] = 32'b00000000000000001001011100110000;
assign LUT_1[23713] = 32'b00000000000000000010101110101100;
assign LUT_1[23714] = 32'b00000000000000000101001011000001;
assign LUT_1[23715] = 32'b11111111111111111110011100111101;
assign LUT_1[23716] = 32'b00000000000000010001010110000111;
assign LUT_1[23717] = 32'b00000000000000001010101000000011;
assign LUT_1[23718] = 32'b00000000000000001101000100011000;
assign LUT_1[23719] = 32'b00000000000000000110010110010100;
assign LUT_1[23720] = 32'b00000000000000001000101010100101;
assign LUT_1[23721] = 32'b00000000000000000001111100100001;
assign LUT_1[23722] = 32'b00000000000000000100011000110110;
assign LUT_1[23723] = 32'b11111111111111111101101010110010;
assign LUT_1[23724] = 32'b00000000000000010000100011111100;
assign LUT_1[23725] = 32'b00000000000000001001110101111000;
assign LUT_1[23726] = 32'b00000000000000001100010010001101;
assign LUT_1[23727] = 32'b00000000000000000101100100001001;
assign LUT_1[23728] = 32'b00000000000000001011011000010010;
assign LUT_1[23729] = 32'b00000000000000000100101010001110;
assign LUT_1[23730] = 32'b00000000000000000111000110100011;
assign LUT_1[23731] = 32'b00000000000000000000011000011111;
assign LUT_1[23732] = 32'b00000000000000010011010001101001;
assign LUT_1[23733] = 32'b00000000000000001100100011100101;
assign LUT_1[23734] = 32'b00000000000000001110111111111010;
assign LUT_1[23735] = 32'b00000000000000001000010001110110;
assign LUT_1[23736] = 32'b00000000000000001010100110000111;
assign LUT_1[23737] = 32'b00000000000000000011111000000011;
assign LUT_1[23738] = 32'b00000000000000000110010100011000;
assign LUT_1[23739] = 32'b11111111111111111111100110010100;
assign LUT_1[23740] = 32'b00000000000000010010011111011110;
assign LUT_1[23741] = 32'b00000000000000001011110001011010;
assign LUT_1[23742] = 32'b00000000000000001110001101101111;
assign LUT_1[23743] = 32'b00000000000000000111011111101011;
assign LUT_1[23744] = 32'b00000000000000001010011111011001;
assign LUT_1[23745] = 32'b00000000000000000011110001010101;
assign LUT_1[23746] = 32'b00000000000000000110001101101010;
assign LUT_1[23747] = 32'b11111111111111111111011111100110;
assign LUT_1[23748] = 32'b00000000000000010010011000110000;
assign LUT_1[23749] = 32'b00000000000000001011101010101100;
assign LUT_1[23750] = 32'b00000000000000001110000111000001;
assign LUT_1[23751] = 32'b00000000000000000111011000111101;
assign LUT_1[23752] = 32'b00000000000000001001101101001110;
assign LUT_1[23753] = 32'b00000000000000000010111111001010;
assign LUT_1[23754] = 32'b00000000000000000101011011011111;
assign LUT_1[23755] = 32'b11111111111111111110101101011011;
assign LUT_1[23756] = 32'b00000000000000010001100110100101;
assign LUT_1[23757] = 32'b00000000000000001010111000100001;
assign LUT_1[23758] = 32'b00000000000000001101010100110110;
assign LUT_1[23759] = 32'b00000000000000000110100110110010;
assign LUT_1[23760] = 32'b00000000000000001100011010111011;
assign LUT_1[23761] = 32'b00000000000000000101101100110111;
assign LUT_1[23762] = 32'b00000000000000001000001001001100;
assign LUT_1[23763] = 32'b00000000000000000001011011001000;
assign LUT_1[23764] = 32'b00000000000000010100010100010010;
assign LUT_1[23765] = 32'b00000000000000001101100110001110;
assign LUT_1[23766] = 32'b00000000000000010000000010100011;
assign LUT_1[23767] = 32'b00000000000000001001010100011111;
assign LUT_1[23768] = 32'b00000000000000001011101000110000;
assign LUT_1[23769] = 32'b00000000000000000100111010101100;
assign LUT_1[23770] = 32'b00000000000000000111010111000001;
assign LUT_1[23771] = 32'b00000000000000000000101000111101;
assign LUT_1[23772] = 32'b00000000000000010011100010000111;
assign LUT_1[23773] = 32'b00000000000000001100110100000011;
assign LUT_1[23774] = 32'b00000000000000001111010000011000;
assign LUT_1[23775] = 32'b00000000000000001000100010010100;
assign LUT_1[23776] = 32'b00000000000000001011011010011000;
assign LUT_1[23777] = 32'b00000000000000000100101100010100;
assign LUT_1[23778] = 32'b00000000000000000111001000101001;
assign LUT_1[23779] = 32'b00000000000000000000011010100101;
assign LUT_1[23780] = 32'b00000000000000010011010011101111;
assign LUT_1[23781] = 32'b00000000000000001100100101101011;
assign LUT_1[23782] = 32'b00000000000000001111000010000000;
assign LUT_1[23783] = 32'b00000000000000001000010011111100;
assign LUT_1[23784] = 32'b00000000000000001010101000001101;
assign LUT_1[23785] = 32'b00000000000000000011111010001001;
assign LUT_1[23786] = 32'b00000000000000000110010110011110;
assign LUT_1[23787] = 32'b11111111111111111111101000011010;
assign LUT_1[23788] = 32'b00000000000000010010100001100100;
assign LUT_1[23789] = 32'b00000000000000001011110011100000;
assign LUT_1[23790] = 32'b00000000000000001110001111110101;
assign LUT_1[23791] = 32'b00000000000000000111100001110001;
assign LUT_1[23792] = 32'b00000000000000001101010101111010;
assign LUT_1[23793] = 32'b00000000000000000110100111110110;
assign LUT_1[23794] = 32'b00000000000000001001000100001011;
assign LUT_1[23795] = 32'b00000000000000000010010110000111;
assign LUT_1[23796] = 32'b00000000000000010101001111010001;
assign LUT_1[23797] = 32'b00000000000000001110100001001101;
assign LUT_1[23798] = 32'b00000000000000010000111101100010;
assign LUT_1[23799] = 32'b00000000000000001010001111011110;
assign LUT_1[23800] = 32'b00000000000000001100100011101111;
assign LUT_1[23801] = 32'b00000000000000000101110101101011;
assign LUT_1[23802] = 32'b00000000000000001000010010000000;
assign LUT_1[23803] = 32'b00000000000000000001100011111100;
assign LUT_1[23804] = 32'b00000000000000010100011101000110;
assign LUT_1[23805] = 32'b00000000000000001101101111000010;
assign LUT_1[23806] = 32'b00000000000000010000001011010111;
assign LUT_1[23807] = 32'b00000000000000001001011101010011;
assign LUT_1[23808] = 32'b00000000000000000011010101111010;
assign LUT_1[23809] = 32'b11111111111111111100100111110110;
assign LUT_1[23810] = 32'b11111111111111111111000100001011;
assign LUT_1[23811] = 32'b11111111111111111000010110000111;
assign LUT_1[23812] = 32'b00000000000000001011001111010001;
assign LUT_1[23813] = 32'b00000000000000000100100001001101;
assign LUT_1[23814] = 32'b00000000000000000110111101100010;
assign LUT_1[23815] = 32'b00000000000000000000001111011110;
assign LUT_1[23816] = 32'b00000000000000000010100011101111;
assign LUT_1[23817] = 32'b11111111111111111011110101101011;
assign LUT_1[23818] = 32'b11111111111111111110010010000000;
assign LUT_1[23819] = 32'b11111111111111110111100011111100;
assign LUT_1[23820] = 32'b00000000000000001010011101000110;
assign LUT_1[23821] = 32'b00000000000000000011101111000010;
assign LUT_1[23822] = 32'b00000000000000000110001011010111;
assign LUT_1[23823] = 32'b11111111111111111111011101010011;
assign LUT_1[23824] = 32'b00000000000000000101010001011100;
assign LUT_1[23825] = 32'b11111111111111111110100011011000;
assign LUT_1[23826] = 32'b00000000000000000000111111101101;
assign LUT_1[23827] = 32'b11111111111111111010010001101001;
assign LUT_1[23828] = 32'b00000000000000001101001010110011;
assign LUT_1[23829] = 32'b00000000000000000110011100101111;
assign LUT_1[23830] = 32'b00000000000000001000111001000100;
assign LUT_1[23831] = 32'b00000000000000000010001011000000;
assign LUT_1[23832] = 32'b00000000000000000100011111010001;
assign LUT_1[23833] = 32'b11111111111111111101110001001101;
assign LUT_1[23834] = 32'b00000000000000000000001101100010;
assign LUT_1[23835] = 32'b11111111111111111001011111011110;
assign LUT_1[23836] = 32'b00000000000000001100011000101000;
assign LUT_1[23837] = 32'b00000000000000000101101010100100;
assign LUT_1[23838] = 32'b00000000000000001000000110111001;
assign LUT_1[23839] = 32'b00000000000000000001011000110101;
assign LUT_1[23840] = 32'b00000000000000000100010000111001;
assign LUT_1[23841] = 32'b11111111111111111101100010110101;
assign LUT_1[23842] = 32'b11111111111111111111111111001010;
assign LUT_1[23843] = 32'b11111111111111111001010001000110;
assign LUT_1[23844] = 32'b00000000000000001100001010010000;
assign LUT_1[23845] = 32'b00000000000000000101011100001100;
assign LUT_1[23846] = 32'b00000000000000000111111000100001;
assign LUT_1[23847] = 32'b00000000000000000001001010011101;
assign LUT_1[23848] = 32'b00000000000000000011011110101110;
assign LUT_1[23849] = 32'b11111111111111111100110000101010;
assign LUT_1[23850] = 32'b11111111111111111111001100111111;
assign LUT_1[23851] = 32'b11111111111111111000011110111011;
assign LUT_1[23852] = 32'b00000000000000001011011000000101;
assign LUT_1[23853] = 32'b00000000000000000100101010000001;
assign LUT_1[23854] = 32'b00000000000000000111000110010110;
assign LUT_1[23855] = 32'b00000000000000000000011000010010;
assign LUT_1[23856] = 32'b00000000000000000110001100011011;
assign LUT_1[23857] = 32'b11111111111111111111011110010111;
assign LUT_1[23858] = 32'b00000000000000000001111010101100;
assign LUT_1[23859] = 32'b11111111111111111011001100101000;
assign LUT_1[23860] = 32'b00000000000000001110000101110010;
assign LUT_1[23861] = 32'b00000000000000000111010111101110;
assign LUT_1[23862] = 32'b00000000000000001001110100000011;
assign LUT_1[23863] = 32'b00000000000000000011000101111111;
assign LUT_1[23864] = 32'b00000000000000000101011010010000;
assign LUT_1[23865] = 32'b11111111111111111110101100001100;
assign LUT_1[23866] = 32'b00000000000000000001001000100001;
assign LUT_1[23867] = 32'b11111111111111111010011010011101;
assign LUT_1[23868] = 32'b00000000000000001101010011100111;
assign LUT_1[23869] = 32'b00000000000000000110100101100011;
assign LUT_1[23870] = 32'b00000000000000001001000001111000;
assign LUT_1[23871] = 32'b00000000000000000010010011110100;
assign LUT_1[23872] = 32'b00000000000000000101010011100010;
assign LUT_1[23873] = 32'b11111111111111111110100101011110;
assign LUT_1[23874] = 32'b00000000000000000001000001110011;
assign LUT_1[23875] = 32'b11111111111111111010010011101111;
assign LUT_1[23876] = 32'b00000000000000001101001100111001;
assign LUT_1[23877] = 32'b00000000000000000110011110110101;
assign LUT_1[23878] = 32'b00000000000000001000111011001010;
assign LUT_1[23879] = 32'b00000000000000000010001101000110;
assign LUT_1[23880] = 32'b00000000000000000100100001010111;
assign LUT_1[23881] = 32'b11111111111111111101110011010011;
assign LUT_1[23882] = 32'b00000000000000000000001111101000;
assign LUT_1[23883] = 32'b11111111111111111001100001100100;
assign LUT_1[23884] = 32'b00000000000000001100011010101110;
assign LUT_1[23885] = 32'b00000000000000000101101100101010;
assign LUT_1[23886] = 32'b00000000000000001000001000111111;
assign LUT_1[23887] = 32'b00000000000000000001011010111011;
assign LUT_1[23888] = 32'b00000000000000000111001111000100;
assign LUT_1[23889] = 32'b00000000000000000000100001000000;
assign LUT_1[23890] = 32'b00000000000000000010111101010101;
assign LUT_1[23891] = 32'b11111111111111111100001111010001;
assign LUT_1[23892] = 32'b00000000000000001111001000011011;
assign LUT_1[23893] = 32'b00000000000000001000011010010111;
assign LUT_1[23894] = 32'b00000000000000001010110110101100;
assign LUT_1[23895] = 32'b00000000000000000100001000101000;
assign LUT_1[23896] = 32'b00000000000000000110011100111001;
assign LUT_1[23897] = 32'b11111111111111111111101110110101;
assign LUT_1[23898] = 32'b00000000000000000010001011001010;
assign LUT_1[23899] = 32'b11111111111111111011011101000110;
assign LUT_1[23900] = 32'b00000000000000001110010110010000;
assign LUT_1[23901] = 32'b00000000000000000111101000001100;
assign LUT_1[23902] = 32'b00000000000000001010000100100001;
assign LUT_1[23903] = 32'b00000000000000000011010110011101;
assign LUT_1[23904] = 32'b00000000000000000110001110100001;
assign LUT_1[23905] = 32'b11111111111111111111100000011101;
assign LUT_1[23906] = 32'b00000000000000000001111100110010;
assign LUT_1[23907] = 32'b11111111111111111011001110101110;
assign LUT_1[23908] = 32'b00000000000000001110000111111000;
assign LUT_1[23909] = 32'b00000000000000000111011001110100;
assign LUT_1[23910] = 32'b00000000000000001001110110001001;
assign LUT_1[23911] = 32'b00000000000000000011001000000101;
assign LUT_1[23912] = 32'b00000000000000000101011100010110;
assign LUT_1[23913] = 32'b11111111111111111110101110010010;
assign LUT_1[23914] = 32'b00000000000000000001001010100111;
assign LUT_1[23915] = 32'b11111111111111111010011100100011;
assign LUT_1[23916] = 32'b00000000000000001101010101101101;
assign LUT_1[23917] = 32'b00000000000000000110100111101001;
assign LUT_1[23918] = 32'b00000000000000001001000011111110;
assign LUT_1[23919] = 32'b00000000000000000010010101111010;
assign LUT_1[23920] = 32'b00000000000000001000001010000011;
assign LUT_1[23921] = 32'b00000000000000000001011011111111;
assign LUT_1[23922] = 32'b00000000000000000011111000010100;
assign LUT_1[23923] = 32'b11111111111111111101001010010000;
assign LUT_1[23924] = 32'b00000000000000010000000011011010;
assign LUT_1[23925] = 32'b00000000000000001001010101010110;
assign LUT_1[23926] = 32'b00000000000000001011110001101011;
assign LUT_1[23927] = 32'b00000000000000000101000011100111;
assign LUT_1[23928] = 32'b00000000000000000111010111111000;
assign LUT_1[23929] = 32'b00000000000000000000101001110100;
assign LUT_1[23930] = 32'b00000000000000000011000110001001;
assign LUT_1[23931] = 32'b11111111111111111100011000000101;
assign LUT_1[23932] = 32'b00000000000000001111010001001111;
assign LUT_1[23933] = 32'b00000000000000001000100011001011;
assign LUT_1[23934] = 32'b00000000000000001010111111100000;
assign LUT_1[23935] = 32'b00000000000000000100010001011100;
assign LUT_1[23936] = 32'b00000000000000000110010101111101;
assign LUT_1[23937] = 32'b11111111111111111111100111111001;
assign LUT_1[23938] = 32'b00000000000000000010000100001110;
assign LUT_1[23939] = 32'b11111111111111111011010110001010;
assign LUT_1[23940] = 32'b00000000000000001110001111010100;
assign LUT_1[23941] = 32'b00000000000000000111100001010000;
assign LUT_1[23942] = 32'b00000000000000001001111101100101;
assign LUT_1[23943] = 32'b00000000000000000011001111100001;
assign LUT_1[23944] = 32'b00000000000000000101100011110010;
assign LUT_1[23945] = 32'b11111111111111111110110101101110;
assign LUT_1[23946] = 32'b00000000000000000001010010000011;
assign LUT_1[23947] = 32'b11111111111111111010100011111111;
assign LUT_1[23948] = 32'b00000000000000001101011101001001;
assign LUT_1[23949] = 32'b00000000000000000110101111000101;
assign LUT_1[23950] = 32'b00000000000000001001001011011010;
assign LUT_1[23951] = 32'b00000000000000000010011101010110;
assign LUT_1[23952] = 32'b00000000000000001000010001011111;
assign LUT_1[23953] = 32'b00000000000000000001100011011011;
assign LUT_1[23954] = 32'b00000000000000000011111111110000;
assign LUT_1[23955] = 32'b11111111111111111101010001101100;
assign LUT_1[23956] = 32'b00000000000000010000001010110110;
assign LUT_1[23957] = 32'b00000000000000001001011100110010;
assign LUT_1[23958] = 32'b00000000000000001011111001000111;
assign LUT_1[23959] = 32'b00000000000000000101001011000011;
assign LUT_1[23960] = 32'b00000000000000000111011111010100;
assign LUT_1[23961] = 32'b00000000000000000000110001010000;
assign LUT_1[23962] = 32'b00000000000000000011001101100101;
assign LUT_1[23963] = 32'b11111111111111111100011111100001;
assign LUT_1[23964] = 32'b00000000000000001111011000101011;
assign LUT_1[23965] = 32'b00000000000000001000101010100111;
assign LUT_1[23966] = 32'b00000000000000001011000110111100;
assign LUT_1[23967] = 32'b00000000000000000100011000111000;
assign LUT_1[23968] = 32'b00000000000000000111010000111100;
assign LUT_1[23969] = 32'b00000000000000000000100010111000;
assign LUT_1[23970] = 32'b00000000000000000010111111001101;
assign LUT_1[23971] = 32'b11111111111111111100010001001001;
assign LUT_1[23972] = 32'b00000000000000001111001010010011;
assign LUT_1[23973] = 32'b00000000000000001000011100001111;
assign LUT_1[23974] = 32'b00000000000000001010111000100100;
assign LUT_1[23975] = 32'b00000000000000000100001010100000;
assign LUT_1[23976] = 32'b00000000000000000110011110110001;
assign LUT_1[23977] = 32'b11111111111111111111110000101101;
assign LUT_1[23978] = 32'b00000000000000000010001101000010;
assign LUT_1[23979] = 32'b11111111111111111011011110111110;
assign LUT_1[23980] = 32'b00000000000000001110011000001000;
assign LUT_1[23981] = 32'b00000000000000000111101010000100;
assign LUT_1[23982] = 32'b00000000000000001010000110011001;
assign LUT_1[23983] = 32'b00000000000000000011011000010101;
assign LUT_1[23984] = 32'b00000000000000001001001100011110;
assign LUT_1[23985] = 32'b00000000000000000010011110011010;
assign LUT_1[23986] = 32'b00000000000000000100111010101111;
assign LUT_1[23987] = 32'b11111111111111111110001100101011;
assign LUT_1[23988] = 32'b00000000000000010001000101110101;
assign LUT_1[23989] = 32'b00000000000000001010010111110001;
assign LUT_1[23990] = 32'b00000000000000001100110100000110;
assign LUT_1[23991] = 32'b00000000000000000110000110000010;
assign LUT_1[23992] = 32'b00000000000000001000011010010011;
assign LUT_1[23993] = 32'b00000000000000000001101100001111;
assign LUT_1[23994] = 32'b00000000000000000100001000100100;
assign LUT_1[23995] = 32'b11111111111111111101011010100000;
assign LUT_1[23996] = 32'b00000000000000010000010011101010;
assign LUT_1[23997] = 32'b00000000000000001001100101100110;
assign LUT_1[23998] = 32'b00000000000000001100000001111011;
assign LUT_1[23999] = 32'b00000000000000000101010011110111;
assign LUT_1[24000] = 32'b00000000000000001000010011100101;
assign LUT_1[24001] = 32'b00000000000000000001100101100001;
assign LUT_1[24002] = 32'b00000000000000000100000001110110;
assign LUT_1[24003] = 32'b11111111111111111101010011110010;
assign LUT_1[24004] = 32'b00000000000000010000001100111100;
assign LUT_1[24005] = 32'b00000000000000001001011110111000;
assign LUT_1[24006] = 32'b00000000000000001011111011001101;
assign LUT_1[24007] = 32'b00000000000000000101001101001001;
assign LUT_1[24008] = 32'b00000000000000000111100001011010;
assign LUT_1[24009] = 32'b00000000000000000000110011010110;
assign LUT_1[24010] = 32'b00000000000000000011001111101011;
assign LUT_1[24011] = 32'b11111111111111111100100001100111;
assign LUT_1[24012] = 32'b00000000000000001111011010110001;
assign LUT_1[24013] = 32'b00000000000000001000101100101101;
assign LUT_1[24014] = 32'b00000000000000001011001001000010;
assign LUT_1[24015] = 32'b00000000000000000100011010111110;
assign LUT_1[24016] = 32'b00000000000000001010001111000111;
assign LUT_1[24017] = 32'b00000000000000000011100001000011;
assign LUT_1[24018] = 32'b00000000000000000101111101011000;
assign LUT_1[24019] = 32'b11111111111111111111001111010100;
assign LUT_1[24020] = 32'b00000000000000010010001000011110;
assign LUT_1[24021] = 32'b00000000000000001011011010011010;
assign LUT_1[24022] = 32'b00000000000000001101110110101111;
assign LUT_1[24023] = 32'b00000000000000000111001000101011;
assign LUT_1[24024] = 32'b00000000000000001001011100111100;
assign LUT_1[24025] = 32'b00000000000000000010101110111000;
assign LUT_1[24026] = 32'b00000000000000000101001011001101;
assign LUT_1[24027] = 32'b11111111111111111110011101001001;
assign LUT_1[24028] = 32'b00000000000000010001010110010011;
assign LUT_1[24029] = 32'b00000000000000001010101000001111;
assign LUT_1[24030] = 32'b00000000000000001101000100100100;
assign LUT_1[24031] = 32'b00000000000000000110010110100000;
assign LUT_1[24032] = 32'b00000000000000001001001110100100;
assign LUT_1[24033] = 32'b00000000000000000010100000100000;
assign LUT_1[24034] = 32'b00000000000000000100111100110101;
assign LUT_1[24035] = 32'b11111111111111111110001110110001;
assign LUT_1[24036] = 32'b00000000000000010001000111111011;
assign LUT_1[24037] = 32'b00000000000000001010011001110111;
assign LUT_1[24038] = 32'b00000000000000001100110110001100;
assign LUT_1[24039] = 32'b00000000000000000110001000001000;
assign LUT_1[24040] = 32'b00000000000000001000011100011001;
assign LUT_1[24041] = 32'b00000000000000000001101110010101;
assign LUT_1[24042] = 32'b00000000000000000100001010101010;
assign LUT_1[24043] = 32'b11111111111111111101011100100110;
assign LUT_1[24044] = 32'b00000000000000010000010101110000;
assign LUT_1[24045] = 32'b00000000000000001001100111101100;
assign LUT_1[24046] = 32'b00000000000000001100000100000001;
assign LUT_1[24047] = 32'b00000000000000000101010101111101;
assign LUT_1[24048] = 32'b00000000000000001011001010000110;
assign LUT_1[24049] = 32'b00000000000000000100011100000010;
assign LUT_1[24050] = 32'b00000000000000000110111000010111;
assign LUT_1[24051] = 32'b00000000000000000000001010010011;
assign LUT_1[24052] = 32'b00000000000000010011000011011101;
assign LUT_1[24053] = 32'b00000000000000001100010101011001;
assign LUT_1[24054] = 32'b00000000000000001110110001101110;
assign LUT_1[24055] = 32'b00000000000000001000000011101010;
assign LUT_1[24056] = 32'b00000000000000001010010111111011;
assign LUT_1[24057] = 32'b00000000000000000011101001110111;
assign LUT_1[24058] = 32'b00000000000000000110000110001100;
assign LUT_1[24059] = 32'b11111111111111111111011000001000;
assign LUT_1[24060] = 32'b00000000000000010010010001010010;
assign LUT_1[24061] = 32'b00000000000000001011100011001110;
assign LUT_1[24062] = 32'b00000000000000001101111111100011;
assign LUT_1[24063] = 32'b00000000000000000111010001011111;
assign LUT_1[24064] = 32'b11111111111111111111010000001011;
assign LUT_1[24065] = 32'b11111111111111111000100010000111;
assign LUT_1[24066] = 32'b11111111111111111010111110011100;
assign LUT_1[24067] = 32'b11111111111111110100010000011000;
assign LUT_1[24068] = 32'b00000000000000000111001001100010;
assign LUT_1[24069] = 32'b00000000000000000000011011011110;
assign LUT_1[24070] = 32'b00000000000000000010110111110011;
assign LUT_1[24071] = 32'b11111111111111111100001001101111;
assign LUT_1[24072] = 32'b11111111111111111110011110000000;
assign LUT_1[24073] = 32'b11111111111111110111101111111100;
assign LUT_1[24074] = 32'b11111111111111111010001100010001;
assign LUT_1[24075] = 32'b11111111111111110011011110001101;
assign LUT_1[24076] = 32'b00000000000000000110010111010111;
assign LUT_1[24077] = 32'b11111111111111111111101001010011;
assign LUT_1[24078] = 32'b00000000000000000010000101101000;
assign LUT_1[24079] = 32'b11111111111111111011010111100100;
assign LUT_1[24080] = 32'b00000000000000000001001011101101;
assign LUT_1[24081] = 32'b11111111111111111010011101101001;
assign LUT_1[24082] = 32'b11111111111111111100111001111110;
assign LUT_1[24083] = 32'b11111111111111110110001011111010;
assign LUT_1[24084] = 32'b00000000000000001001000101000100;
assign LUT_1[24085] = 32'b00000000000000000010010111000000;
assign LUT_1[24086] = 32'b00000000000000000100110011010101;
assign LUT_1[24087] = 32'b11111111111111111110000101010001;
assign LUT_1[24088] = 32'b00000000000000000000011001100010;
assign LUT_1[24089] = 32'b11111111111111111001101011011110;
assign LUT_1[24090] = 32'b11111111111111111100000111110011;
assign LUT_1[24091] = 32'b11111111111111110101011001101111;
assign LUT_1[24092] = 32'b00000000000000001000010010111001;
assign LUT_1[24093] = 32'b00000000000000000001100100110101;
assign LUT_1[24094] = 32'b00000000000000000100000001001010;
assign LUT_1[24095] = 32'b11111111111111111101010011000110;
assign LUT_1[24096] = 32'b00000000000000000000001011001010;
assign LUT_1[24097] = 32'b11111111111111111001011101000110;
assign LUT_1[24098] = 32'b11111111111111111011111001011011;
assign LUT_1[24099] = 32'b11111111111111110101001011010111;
assign LUT_1[24100] = 32'b00000000000000001000000100100001;
assign LUT_1[24101] = 32'b00000000000000000001010110011101;
assign LUT_1[24102] = 32'b00000000000000000011110010110010;
assign LUT_1[24103] = 32'b11111111111111111101000100101110;
assign LUT_1[24104] = 32'b11111111111111111111011000111111;
assign LUT_1[24105] = 32'b11111111111111111000101010111011;
assign LUT_1[24106] = 32'b11111111111111111011000111010000;
assign LUT_1[24107] = 32'b11111111111111110100011001001100;
assign LUT_1[24108] = 32'b00000000000000000111010010010110;
assign LUT_1[24109] = 32'b00000000000000000000100100010010;
assign LUT_1[24110] = 32'b00000000000000000011000000100111;
assign LUT_1[24111] = 32'b11111111111111111100010010100011;
assign LUT_1[24112] = 32'b00000000000000000010000110101100;
assign LUT_1[24113] = 32'b11111111111111111011011000101000;
assign LUT_1[24114] = 32'b11111111111111111101110100111101;
assign LUT_1[24115] = 32'b11111111111111110111000110111001;
assign LUT_1[24116] = 32'b00000000000000001010000000000011;
assign LUT_1[24117] = 32'b00000000000000000011010001111111;
assign LUT_1[24118] = 32'b00000000000000000101101110010100;
assign LUT_1[24119] = 32'b11111111111111111111000000010000;
assign LUT_1[24120] = 32'b00000000000000000001010100100001;
assign LUT_1[24121] = 32'b11111111111111111010100110011101;
assign LUT_1[24122] = 32'b11111111111111111101000010110010;
assign LUT_1[24123] = 32'b11111111111111110110010100101110;
assign LUT_1[24124] = 32'b00000000000000001001001101111000;
assign LUT_1[24125] = 32'b00000000000000000010011111110100;
assign LUT_1[24126] = 32'b00000000000000000100111100001001;
assign LUT_1[24127] = 32'b11111111111111111110001110000101;
assign LUT_1[24128] = 32'b00000000000000000001001101110011;
assign LUT_1[24129] = 32'b11111111111111111010011111101111;
assign LUT_1[24130] = 32'b11111111111111111100111100000100;
assign LUT_1[24131] = 32'b11111111111111110110001110000000;
assign LUT_1[24132] = 32'b00000000000000001001000111001010;
assign LUT_1[24133] = 32'b00000000000000000010011001000110;
assign LUT_1[24134] = 32'b00000000000000000100110101011011;
assign LUT_1[24135] = 32'b11111111111111111110000111010111;
assign LUT_1[24136] = 32'b00000000000000000000011011101000;
assign LUT_1[24137] = 32'b11111111111111111001101101100100;
assign LUT_1[24138] = 32'b11111111111111111100001001111001;
assign LUT_1[24139] = 32'b11111111111111110101011011110101;
assign LUT_1[24140] = 32'b00000000000000001000010100111111;
assign LUT_1[24141] = 32'b00000000000000000001100110111011;
assign LUT_1[24142] = 32'b00000000000000000100000011010000;
assign LUT_1[24143] = 32'b11111111111111111101010101001100;
assign LUT_1[24144] = 32'b00000000000000000011001001010101;
assign LUT_1[24145] = 32'b11111111111111111100011011010001;
assign LUT_1[24146] = 32'b11111111111111111110110111100110;
assign LUT_1[24147] = 32'b11111111111111111000001001100010;
assign LUT_1[24148] = 32'b00000000000000001011000010101100;
assign LUT_1[24149] = 32'b00000000000000000100010100101000;
assign LUT_1[24150] = 32'b00000000000000000110110000111101;
assign LUT_1[24151] = 32'b00000000000000000000000010111001;
assign LUT_1[24152] = 32'b00000000000000000010010111001010;
assign LUT_1[24153] = 32'b11111111111111111011101001000110;
assign LUT_1[24154] = 32'b11111111111111111110000101011011;
assign LUT_1[24155] = 32'b11111111111111110111010111010111;
assign LUT_1[24156] = 32'b00000000000000001010010000100001;
assign LUT_1[24157] = 32'b00000000000000000011100010011101;
assign LUT_1[24158] = 32'b00000000000000000101111110110010;
assign LUT_1[24159] = 32'b11111111111111111111010000101110;
assign LUT_1[24160] = 32'b00000000000000000010001000110010;
assign LUT_1[24161] = 32'b11111111111111111011011010101110;
assign LUT_1[24162] = 32'b11111111111111111101110111000011;
assign LUT_1[24163] = 32'b11111111111111110111001000111111;
assign LUT_1[24164] = 32'b00000000000000001010000010001001;
assign LUT_1[24165] = 32'b00000000000000000011010100000101;
assign LUT_1[24166] = 32'b00000000000000000101110000011010;
assign LUT_1[24167] = 32'b11111111111111111111000010010110;
assign LUT_1[24168] = 32'b00000000000000000001010110100111;
assign LUT_1[24169] = 32'b11111111111111111010101000100011;
assign LUT_1[24170] = 32'b11111111111111111101000100111000;
assign LUT_1[24171] = 32'b11111111111111110110010110110100;
assign LUT_1[24172] = 32'b00000000000000001001001111111110;
assign LUT_1[24173] = 32'b00000000000000000010100001111010;
assign LUT_1[24174] = 32'b00000000000000000100111110001111;
assign LUT_1[24175] = 32'b11111111111111111110010000001011;
assign LUT_1[24176] = 32'b00000000000000000100000100010100;
assign LUT_1[24177] = 32'b11111111111111111101010110010000;
assign LUT_1[24178] = 32'b11111111111111111111110010100101;
assign LUT_1[24179] = 32'b11111111111111111001000100100001;
assign LUT_1[24180] = 32'b00000000000000001011111101101011;
assign LUT_1[24181] = 32'b00000000000000000101001111100111;
assign LUT_1[24182] = 32'b00000000000000000111101011111100;
assign LUT_1[24183] = 32'b00000000000000000000111101111000;
assign LUT_1[24184] = 32'b00000000000000000011010010001001;
assign LUT_1[24185] = 32'b11111111111111111100100100000101;
assign LUT_1[24186] = 32'b11111111111111111111000000011010;
assign LUT_1[24187] = 32'b11111111111111111000010010010110;
assign LUT_1[24188] = 32'b00000000000000001011001011100000;
assign LUT_1[24189] = 32'b00000000000000000100011101011100;
assign LUT_1[24190] = 32'b00000000000000000110111001110001;
assign LUT_1[24191] = 32'b00000000000000000000001011101101;
assign LUT_1[24192] = 32'b00000000000000000010010000001110;
assign LUT_1[24193] = 32'b11111111111111111011100010001010;
assign LUT_1[24194] = 32'b11111111111111111101111110011111;
assign LUT_1[24195] = 32'b11111111111111110111010000011011;
assign LUT_1[24196] = 32'b00000000000000001010001001100101;
assign LUT_1[24197] = 32'b00000000000000000011011011100001;
assign LUT_1[24198] = 32'b00000000000000000101110111110110;
assign LUT_1[24199] = 32'b11111111111111111111001001110010;
assign LUT_1[24200] = 32'b00000000000000000001011110000011;
assign LUT_1[24201] = 32'b11111111111111111010101111111111;
assign LUT_1[24202] = 32'b11111111111111111101001100010100;
assign LUT_1[24203] = 32'b11111111111111110110011110010000;
assign LUT_1[24204] = 32'b00000000000000001001010111011010;
assign LUT_1[24205] = 32'b00000000000000000010101001010110;
assign LUT_1[24206] = 32'b00000000000000000101000101101011;
assign LUT_1[24207] = 32'b11111111111111111110010111100111;
assign LUT_1[24208] = 32'b00000000000000000100001011110000;
assign LUT_1[24209] = 32'b11111111111111111101011101101100;
assign LUT_1[24210] = 32'b11111111111111111111111010000001;
assign LUT_1[24211] = 32'b11111111111111111001001011111101;
assign LUT_1[24212] = 32'b00000000000000001100000101000111;
assign LUT_1[24213] = 32'b00000000000000000101010111000011;
assign LUT_1[24214] = 32'b00000000000000000111110011011000;
assign LUT_1[24215] = 32'b00000000000000000001000101010100;
assign LUT_1[24216] = 32'b00000000000000000011011001100101;
assign LUT_1[24217] = 32'b11111111111111111100101011100001;
assign LUT_1[24218] = 32'b11111111111111111111000111110110;
assign LUT_1[24219] = 32'b11111111111111111000011001110010;
assign LUT_1[24220] = 32'b00000000000000001011010010111100;
assign LUT_1[24221] = 32'b00000000000000000100100100111000;
assign LUT_1[24222] = 32'b00000000000000000111000001001101;
assign LUT_1[24223] = 32'b00000000000000000000010011001001;
assign LUT_1[24224] = 32'b00000000000000000011001011001101;
assign LUT_1[24225] = 32'b11111111111111111100011101001001;
assign LUT_1[24226] = 32'b11111111111111111110111001011110;
assign LUT_1[24227] = 32'b11111111111111111000001011011010;
assign LUT_1[24228] = 32'b00000000000000001011000100100100;
assign LUT_1[24229] = 32'b00000000000000000100010110100000;
assign LUT_1[24230] = 32'b00000000000000000110110010110101;
assign LUT_1[24231] = 32'b00000000000000000000000100110001;
assign LUT_1[24232] = 32'b00000000000000000010011001000010;
assign LUT_1[24233] = 32'b11111111111111111011101010111110;
assign LUT_1[24234] = 32'b11111111111111111110000111010011;
assign LUT_1[24235] = 32'b11111111111111110111011001001111;
assign LUT_1[24236] = 32'b00000000000000001010010010011001;
assign LUT_1[24237] = 32'b00000000000000000011100100010101;
assign LUT_1[24238] = 32'b00000000000000000110000000101010;
assign LUT_1[24239] = 32'b11111111111111111111010010100110;
assign LUT_1[24240] = 32'b00000000000000000101000110101111;
assign LUT_1[24241] = 32'b11111111111111111110011000101011;
assign LUT_1[24242] = 32'b00000000000000000000110101000000;
assign LUT_1[24243] = 32'b11111111111111111010000110111100;
assign LUT_1[24244] = 32'b00000000000000001101000000000110;
assign LUT_1[24245] = 32'b00000000000000000110010010000010;
assign LUT_1[24246] = 32'b00000000000000001000101110010111;
assign LUT_1[24247] = 32'b00000000000000000010000000010011;
assign LUT_1[24248] = 32'b00000000000000000100010100100100;
assign LUT_1[24249] = 32'b11111111111111111101100110100000;
assign LUT_1[24250] = 32'b00000000000000000000000010110101;
assign LUT_1[24251] = 32'b11111111111111111001010100110001;
assign LUT_1[24252] = 32'b00000000000000001100001101111011;
assign LUT_1[24253] = 32'b00000000000000000101011111110111;
assign LUT_1[24254] = 32'b00000000000000000111111100001100;
assign LUT_1[24255] = 32'b00000000000000000001001110001000;
assign LUT_1[24256] = 32'b00000000000000000100001101110110;
assign LUT_1[24257] = 32'b11111111111111111101011111110010;
assign LUT_1[24258] = 32'b11111111111111111111111100000111;
assign LUT_1[24259] = 32'b11111111111111111001001110000011;
assign LUT_1[24260] = 32'b00000000000000001100000111001101;
assign LUT_1[24261] = 32'b00000000000000000101011001001001;
assign LUT_1[24262] = 32'b00000000000000000111110101011110;
assign LUT_1[24263] = 32'b00000000000000000001000111011010;
assign LUT_1[24264] = 32'b00000000000000000011011011101011;
assign LUT_1[24265] = 32'b11111111111111111100101101100111;
assign LUT_1[24266] = 32'b11111111111111111111001001111100;
assign LUT_1[24267] = 32'b11111111111111111000011011111000;
assign LUT_1[24268] = 32'b00000000000000001011010101000010;
assign LUT_1[24269] = 32'b00000000000000000100100110111110;
assign LUT_1[24270] = 32'b00000000000000000111000011010011;
assign LUT_1[24271] = 32'b00000000000000000000010101001111;
assign LUT_1[24272] = 32'b00000000000000000110001001011000;
assign LUT_1[24273] = 32'b11111111111111111111011011010100;
assign LUT_1[24274] = 32'b00000000000000000001110111101001;
assign LUT_1[24275] = 32'b11111111111111111011001001100101;
assign LUT_1[24276] = 32'b00000000000000001110000010101111;
assign LUT_1[24277] = 32'b00000000000000000111010100101011;
assign LUT_1[24278] = 32'b00000000000000001001110001000000;
assign LUT_1[24279] = 32'b00000000000000000011000010111100;
assign LUT_1[24280] = 32'b00000000000000000101010111001101;
assign LUT_1[24281] = 32'b11111111111111111110101001001001;
assign LUT_1[24282] = 32'b00000000000000000001000101011110;
assign LUT_1[24283] = 32'b11111111111111111010010111011010;
assign LUT_1[24284] = 32'b00000000000000001101010000100100;
assign LUT_1[24285] = 32'b00000000000000000110100010100000;
assign LUT_1[24286] = 32'b00000000000000001000111110110101;
assign LUT_1[24287] = 32'b00000000000000000010010000110001;
assign LUT_1[24288] = 32'b00000000000000000101001000110101;
assign LUT_1[24289] = 32'b11111111111111111110011010110001;
assign LUT_1[24290] = 32'b00000000000000000000110111000110;
assign LUT_1[24291] = 32'b11111111111111111010001001000010;
assign LUT_1[24292] = 32'b00000000000000001101000010001100;
assign LUT_1[24293] = 32'b00000000000000000110010100001000;
assign LUT_1[24294] = 32'b00000000000000001000110000011101;
assign LUT_1[24295] = 32'b00000000000000000010000010011001;
assign LUT_1[24296] = 32'b00000000000000000100010110101010;
assign LUT_1[24297] = 32'b11111111111111111101101000100110;
assign LUT_1[24298] = 32'b00000000000000000000000100111011;
assign LUT_1[24299] = 32'b11111111111111111001010110110111;
assign LUT_1[24300] = 32'b00000000000000001100010000000001;
assign LUT_1[24301] = 32'b00000000000000000101100001111101;
assign LUT_1[24302] = 32'b00000000000000000111111110010010;
assign LUT_1[24303] = 32'b00000000000000000001010000001110;
assign LUT_1[24304] = 32'b00000000000000000111000100010111;
assign LUT_1[24305] = 32'b00000000000000000000010110010011;
assign LUT_1[24306] = 32'b00000000000000000010110010101000;
assign LUT_1[24307] = 32'b11111111111111111100000100100100;
assign LUT_1[24308] = 32'b00000000000000001110111101101110;
assign LUT_1[24309] = 32'b00000000000000001000001111101010;
assign LUT_1[24310] = 32'b00000000000000001010101011111111;
assign LUT_1[24311] = 32'b00000000000000000011111101111011;
assign LUT_1[24312] = 32'b00000000000000000110010010001100;
assign LUT_1[24313] = 32'b11111111111111111111100100001000;
assign LUT_1[24314] = 32'b00000000000000000010000000011101;
assign LUT_1[24315] = 32'b11111111111111111011010010011001;
assign LUT_1[24316] = 32'b00000000000000001110001011100011;
assign LUT_1[24317] = 32'b00000000000000000111011101011111;
assign LUT_1[24318] = 32'b00000000000000001001111001110100;
assign LUT_1[24319] = 32'b00000000000000000011001011110000;
assign LUT_1[24320] = 32'b11111111111111111101000100010111;
assign LUT_1[24321] = 32'b11111111111111110110010110010011;
assign LUT_1[24322] = 32'b11111111111111111000110010101000;
assign LUT_1[24323] = 32'b11111111111111110010000100100100;
assign LUT_1[24324] = 32'b00000000000000000100111101101110;
assign LUT_1[24325] = 32'b11111111111111111110001111101010;
assign LUT_1[24326] = 32'b00000000000000000000101011111111;
assign LUT_1[24327] = 32'b11111111111111111001111101111011;
assign LUT_1[24328] = 32'b11111111111111111100010010001100;
assign LUT_1[24329] = 32'b11111111111111110101100100001000;
assign LUT_1[24330] = 32'b11111111111111111000000000011101;
assign LUT_1[24331] = 32'b11111111111111110001010010011001;
assign LUT_1[24332] = 32'b00000000000000000100001011100011;
assign LUT_1[24333] = 32'b11111111111111111101011101011111;
assign LUT_1[24334] = 32'b11111111111111111111111001110100;
assign LUT_1[24335] = 32'b11111111111111111001001011110000;
assign LUT_1[24336] = 32'b11111111111111111110111111111001;
assign LUT_1[24337] = 32'b11111111111111111000010001110101;
assign LUT_1[24338] = 32'b11111111111111111010101110001010;
assign LUT_1[24339] = 32'b11111111111111110100000000000110;
assign LUT_1[24340] = 32'b00000000000000000110111001010000;
assign LUT_1[24341] = 32'b00000000000000000000001011001100;
assign LUT_1[24342] = 32'b00000000000000000010100111100001;
assign LUT_1[24343] = 32'b11111111111111111011111001011101;
assign LUT_1[24344] = 32'b11111111111111111110001101101110;
assign LUT_1[24345] = 32'b11111111111111110111011111101010;
assign LUT_1[24346] = 32'b11111111111111111001111011111111;
assign LUT_1[24347] = 32'b11111111111111110011001101111011;
assign LUT_1[24348] = 32'b00000000000000000110000111000101;
assign LUT_1[24349] = 32'b11111111111111111111011001000001;
assign LUT_1[24350] = 32'b00000000000000000001110101010110;
assign LUT_1[24351] = 32'b11111111111111111011000111010010;
assign LUT_1[24352] = 32'b11111111111111111101111111010110;
assign LUT_1[24353] = 32'b11111111111111110111010001010010;
assign LUT_1[24354] = 32'b11111111111111111001101101100111;
assign LUT_1[24355] = 32'b11111111111111110010111111100011;
assign LUT_1[24356] = 32'b00000000000000000101111000101101;
assign LUT_1[24357] = 32'b11111111111111111111001010101001;
assign LUT_1[24358] = 32'b00000000000000000001100110111110;
assign LUT_1[24359] = 32'b11111111111111111010111000111010;
assign LUT_1[24360] = 32'b11111111111111111101001101001011;
assign LUT_1[24361] = 32'b11111111111111110110011111000111;
assign LUT_1[24362] = 32'b11111111111111111000111011011100;
assign LUT_1[24363] = 32'b11111111111111110010001101011000;
assign LUT_1[24364] = 32'b00000000000000000101000110100010;
assign LUT_1[24365] = 32'b11111111111111111110011000011110;
assign LUT_1[24366] = 32'b00000000000000000000110100110011;
assign LUT_1[24367] = 32'b11111111111111111010000110101111;
assign LUT_1[24368] = 32'b11111111111111111111111010111000;
assign LUT_1[24369] = 32'b11111111111111111001001100110100;
assign LUT_1[24370] = 32'b11111111111111111011101001001001;
assign LUT_1[24371] = 32'b11111111111111110100111011000101;
assign LUT_1[24372] = 32'b00000000000000000111110100001111;
assign LUT_1[24373] = 32'b00000000000000000001000110001011;
assign LUT_1[24374] = 32'b00000000000000000011100010100000;
assign LUT_1[24375] = 32'b11111111111111111100110100011100;
assign LUT_1[24376] = 32'b11111111111111111111001000101101;
assign LUT_1[24377] = 32'b11111111111111111000011010101001;
assign LUT_1[24378] = 32'b11111111111111111010110110111110;
assign LUT_1[24379] = 32'b11111111111111110100001000111010;
assign LUT_1[24380] = 32'b00000000000000000111000010000100;
assign LUT_1[24381] = 32'b00000000000000000000010100000000;
assign LUT_1[24382] = 32'b00000000000000000010110000010101;
assign LUT_1[24383] = 32'b11111111111111111100000010010001;
assign LUT_1[24384] = 32'b11111111111111111111000001111111;
assign LUT_1[24385] = 32'b11111111111111111000010011111011;
assign LUT_1[24386] = 32'b11111111111111111010110000010000;
assign LUT_1[24387] = 32'b11111111111111110100000010001100;
assign LUT_1[24388] = 32'b00000000000000000110111011010110;
assign LUT_1[24389] = 32'b00000000000000000000001101010010;
assign LUT_1[24390] = 32'b00000000000000000010101001100111;
assign LUT_1[24391] = 32'b11111111111111111011111011100011;
assign LUT_1[24392] = 32'b11111111111111111110001111110100;
assign LUT_1[24393] = 32'b11111111111111110111100001110000;
assign LUT_1[24394] = 32'b11111111111111111001111110000101;
assign LUT_1[24395] = 32'b11111111111111110011010000000001;
assign LUT_1[24396] = 32'b00000000000000000110001001001011;
assign LUT_1[24397] = 32'b11111111111111111111011011000111;
assign LUT_1[24398] = 32'b00000000000000000001110111011100;
assign LUT_1[24399] = 32'b11111111111111111011001001011000;
assign LUT_1[24400] = 32'b00000000000000000000111101100001;
assign LUT_1[24401] = 32'b11111111111111111010001111011101;
assign LUT_1[24402] = 32'b11111111111111111100101011110010;
assign LUT_1[24403] = 32'b11111111111111110101111101101110;
assign LUT_1[24404] = 32'b00000000000000001000110110111000;
assign LUT_1[24405] = 32'b00000000000000000010001000110100;
assign LUT_1[24406] = 32'b00000000000000000100100101001001;
assign LUT_1[24407] = 32'b11111111111111111101110111000101;
assign LUT_1[24408] = 32'b00000000000000000000001011010110;
assign LUT_1[24409] = 32'b11111111111111111001011101010010;
assign LUT_1[24410] = 32'b11111111111111111011111001100111;
assign LUT_1[24411] = 32'b11111111111111110101001011100011;
assign LUT_1[24412] = 32'b00000000000000001000000100101101;
assign LUT_1[24413] = 32'b00000000000000000001010110101001;
assign LUT_1[24414] = 32'b00000000000000000011110010111110;
assign LUT_1[24415] = 32'b11111111111111111101000100111010;
assign LUT_1[24416] = 32'b11111111111111111111111100111110;
assign LUT_1[24417] = 32'b11111111111111111001001110111010;
assign LUT_1[24418] = 32'b11111111111111111011101011001111;
assign LUT_1[24419] = 32'b11111111111111110100111101001011;
assign LUT_1[24420] = 32'b00000000000000000111110110010101;
assign LUT_1[24421] = 32'b00000000000000000001001000010001;
assign LUT_1[24422] = 32'b00000000000000000011100100100110;
assign LUT_1[24423] = 32'b11111111111111111100110110100010;
assign LUT_1[24424] = 32'b11111111111111111111001010110011;
assign LUT_1[24425] = 32'b11111111111111111000011100101111;
assign LUT_1[24426] = 32'b11111111111111111010111001000100;
assign LUT_1[24427] = 32'b11111111111111110100001011000000;
assign LUT_1[24428] = 32'b00000000000000000111000100001010;
assign LUT_1[24429] = 32'b00000000000000000000010110000110;
assign LUT_1[24430] = 32'b00000000000000000010110010011011;
assign LUT_1[24431] = 32'b11111111111111111100000100010111;
assign LUT_1[24432] = 32'b00000000000000000001111000100000;
assign LUT_1[24433] = 32'b11111111111111111011001010011100;
assign LUT_1[24434] = 32'b11111111111111111101100110110001;
assign LUT_1[24435] = 32'b11111111111111110110111000101101;
assign LUT_1[24436] = 32'b00000000000000001001110001110111;
assign LUT_1[24437] = 32'b00000000000000000011000011110011;
assign LUT_1[24438] = 32'b00000000000000000101100000001000;
assign LUT_1[24439] = 32'b11111111111111111110110010000100;
assign LUT_1[24440] = 32'b00000000000000000001000110010101;
assign LUT_1[24441] = 32'b11111111111111111010011000010001;
assign LUT_1[24442] = 32'b11111111111111111100110100100110;
assign LUT_1[24443] = 32'b11111111111111110110000110100010;
assign LUT_1[24444] = 32'b00000000000000001000111111101100;
assign LUT_1[24445] = 32'b00000000000000000010010001101000;
assign LUT_1[24446] = 32'b00000000000000000100101101111101;
assign LUT_1[24447] = 32'b11111111111111111101111111111001;
assign LUT_1[24448] = 32'b00000000000000000000000100011010;
assign LUT_1[24449] = 32'b11111111111111111001010110010110;
assign LUT_1[24450] = 32'b11111111111111111011110010101011;
assign LUT_1[24451] = 32'b11111111111111110101000100100111;
assign LUT_1[24452] = 32'b00000000000000000111111101110001;
assign LUT_1[24453] = 32'b00000000000000000001001111101101;
assign LUT_1[24454] = 32'b00000000000000000011101100000010;
assign LUT_1[24455] = 32'b11111111111111111100111101111110;
assign LUT_1[24456] = 32'b11111111111111111111010010001111;
assign LUT_1[24457] = 32'b11111111111111111000100100001011;
assign LUT_1[24458] = 32'b11111111111111111011000000100000;
assign LUT_1[24459] = 32'b11111111111111110100010010011100;
assign LUT_1[24460] = 32'b00000000000000000111001011100110;
assign LUT_1[24461] = 32'b00000000000000000000011101100010;
assign LUT_1[24462] = 32'b00000000000000000010111001110111;
assign LUT_1[24463] = 32'b11111111111111111100001011110011;
assign LUT_1[24464] = 32'b00000000000000000001111111111100;
assign LUT_1[24465] = 32'b11111111111111111011010001111000;
assign LUT_1[24466] = 32'b11111111111111111101101110001101;
assign LUT_1[24467] = 32'b11111111111111110111000000001001;
assign LUT_1[24468] = 32'b00000000000000001001111001010011;
assign LUT_1[24469] = 32'b00000000000000000011001011001111;
assign LUT_1[24470] = 32'b00000000000000000101100111100100;
assign LUT_1[24471] = 32'b11111111111111111110111001100000;
assign LUT_1[24472] = 32'b00000000000000000001001101110001;
assign LUT_1[24473] = 32'b11111111111111111010011111101101;
assign LUT_1[24474] = 32'b11111111111111111100111100000010;
assign LUT_1[24475] = 32'b11111111111111110110001101111110;
assign LUT_1[24476] = 32'b00000000000000001001000111001000;
assign LUT_1[24477] = 32'b00000000000000000010011001000100;
assign LUT_1[24478] = 32'b00000000000000000100110101011001;
assign LUT_1[24479] = 32'b11111111111111111110000111010101;
assign LUT_1[24480] = 32'b00000000000000000000111111011001;
assign LUT_1[24481] = 32'b11111111111111111010010001010101;
assign LUT_1[24482] = 32'b11111111111111111100101101101010;
assign LUT_1[24483] = 32'b11111111111111110101111111100110;
assign LUT_1[24484] = 32'b00000000000000001000111000110000;
assign LUT_1[24485] = 32'b00000000000000000010001010101100;
assign LUT_1[24486] = 32'b00000000000000000100100111000001;
assign LUT_1[24487] = 32'b11111111111111111101111000111101;
assign LUT_1[24488] = 32'b00000000000000000000001101001110;
assign LUT_1[24489] = 32'b11111111111111111001011111001010;
assign LUT_1[24490] = 32'b11111111111111111011111011011111;
assign LUT_1[24491] = 32'b11111111111111110101001101011011;
assign LUT_1[24492] = 32'b00000000000000001000000110100101;
assign LUT_1[24493] = 32'b00000000000000000001011000100001;
assign LUT_1[24494] = 32'b00000000000000000011110100110110;
assign LUT_1[24495] = 32'b11111111111111111101000110110010;
assign LUT_1[24496] = 32'b00000000000000000010111010111011;
assign LUT_1[24497] = 32'b11111111111111111100001100110111;
assign LUT_1[24498] = 32'b11111111111111111110101001001100;
assign LUT_1[24499] = 32'b11111111111111110111111011001000;
assign LUT_1[24500] = 32'b00000000000000001010110100010010;
assign LUT_1[24501] = 32'b00000000000000000100000110001110;
assign LUT_1[24502] = 32'b00000000000000000110100010100011;
assign LUT_1[24503] = 32'b11111111111111111111110100011111;
assign LUT_1[24504] = 32'b00000000000000000010001000110000;
assign LUT_1[24505] = 32'b11111111111111111011011010101100;
assign LUT_1[24506] = 32'b11111111111111111101110111000001;
assign LUT_1[24507] = 32'b11111111111111110111001000111101;
assign LUT_1[24508] = 32'b00000000000000001010000010000111;
assign LUT_1[24509] = 32'b00000000000000000011010100000011;
assign LUT_1[24510] = 32'b00000000000000000101110000011000;
assign LUT_1[24511] = 32'b11111111111111111111000010010100;
assign LUT_1[24512] = 32'b00000000000000000010000010000010;
assign LUT_1[24513] = 32'b11111111111111111011010011111110;
assign LUT_1[24514] = 32'b11111111111111111101110000010011;
assign LUT_1[24515] = 32'b11111111111111110111000010001111;
assign LUT_1[24516] = 32'b00000000000000001001111011011001;
assign LUT_1[24517] = 32'b00000000000000000011001101010101;
assign LUT_1[24518] = 32'b00000000000000000101101001101010;
assign LUT_1[24519] = 32'b11111111111111111110111011100110;
assign LUT_1[24520] = 32'b00000000000000000001001111110111;
assign LUT_1[24521] = 32'b11111111111111111010100001110011;
assign LUT_1[24522] = 32'b11111111111111111100111110001000;
assign LUT_1[24523] = 32'b11111111111111110110010000000100;
assign LUT_1[24524] = 32'b00000000000000001001001001001110;
assign LUT_1[24525] = 32'b00000000000000000010011011001010;
assign LUT_1[24526] = 32'b00000000000000000100110111011111;
assign LUT_1[24527] = 32'b11111111111111111110001001011011;
assign LUT_1[24528] = 32'b00000000000000000011111101100100;
assign LUT_1[24529] = 32'b11111111111111111101001111100000;
assign LUT_1[24530] = 32'b11111111111111111111101011110101;
assign LUT_1[24531] = 32'b11111111111111111000111101110001;
assign LUT_1[24532] = 32'b00000000000000001011110110111011;
assign LUT_1[24533] = 32'b00000000000000000101001000110111;
assign LUT_1[24534] = 32'b00000000000000000111100101001100;
assign LUT_1[24535] = 32'b00000000000000000000110111001000;
assign LUT_1[24536] = 32'b00000000000000000011001011011001;
assign LUT_1[24537] = 32'b11111111111111111100011101010101;
assign LUT_1[24538] = 32'b11111111111111111110111001101010;
assign LUT_1[24539] = 32'b11111111111111111000001011100110;
assign LUT_1[24540] = 32'b00000000000000001011000100110000;
assign LUT_1[24541] = 32'b00000000000000000100010110101100;
assign LUT_1[24542] = 32'b00000000000000000110110011000001;
assign LUT_1[24543] = 32'b00000000000000000000000100111101;
assign LUT_1[24544] = 32'b00000000000000000010111101000001;
assign LUT_1[24545] = 32'b11111111111111111100001110111101;
assign LUT_1[24546] = 32'b11111111111111111110101011010010;
assign LUT_1[24547] = 32'b11111111111111110111111101001110;
assign LUT_1[24548] = 32'b00000000000000001010110110011000;
assign LUT_1[24549] = 32'b00000000000000000100001000010100;
assign LUT_1[24550] = 32'b00000000000000000110100100101001;
assign LUT_1[24551] = 32'b11111111111111111111110110100101;
assign LUT_1[24552] = 32'b00000000000000000010001010110110;
assign LUT_1[24553] = 32'b11111111111111111011011100110010;
assign LUT_1[24554] = 32'b11111111111111111101111001000111;
assign LUT_1[24555] = 32'b11111111111111110111001011000011;
assign LUT_1[24556] = 32'b00000000000000001010000100001101;
assign LUT_1[24557] = 32'b00000000000000000011010110001001;
assign LUT_1[24558] = 32'b00000000000000000101110010011110;
assign LUT_1[24559] = 32'b11111111111111111111000100011010;
assign LUT_1[24560] = 32'b00000000000000000100111000100011;
assign LUT_1[24561] = 32'b11111111111111111110001010011111;
assign LUT_1[24562] = 32'b00000000000000000000100110110100;
assign LUT_1[24563] = 32'b11111111111111111001111000110000;
assign LUT_1[24564] = 32'b00000000000000001100110001111010;
assign LUT_1[24565] = 32'b00000000000000000110000011110110;
assign LUT_1[24566] = 32'b00000000000000001000100000001011;
assign LUT_1[24567] = 32'b00000000000000000001110010000111;
assign LUT_1[24568] = 32'b00000000000000000100000110011000;
assign LUT_1[24569] = 32'b11111111111111111101011000010100;
assign LUT_1[24570] = 32'b11111111111111111111110100101001;
assign LUT_1[24571] = 32'b11111111111111111001000110100101;
assign LUT_1[24572] = 32'b00000000000000001011111111101111;
assign LUT_1[24573] = 32'b00000000000000000101010001101011;
assign LUT_1[24574] = 32'b00000000000000000111101110000000;
assign LUT_1[24575] = 32'b00000000000000000000111111111100;
assign LUT_1[24576] = 32'b00000000000000000001011100100000;
assign LUT_1[24577] = 32'b11111111111111111010101110011100;
assign LUT_1[24578] = 32'b11111111111111111101001010110001;
assign LUT_1[24579] = 32'b11111111111111110110011100101101;
assign LUT_1[24580] = 32'b00000000000000001001010101110111;
assign LUT_1[24581] = 32'b00000000000000000010100111110011;
assign LUT_1[24582] = 32'b00000000000000000101000100001000;
assign LUT_1[24583] = 32'b11111111111111111110010110000100;
assign LUT_1[24584] = 32'b00000000000000000000101010010101;
assign LUT_1[24585] = 32'b11111111111111111001111100010001;
assign LUT_1[24586] = 32'b11111111111111111100011000100110;
assign LUT_1[24587] = 32'b11111111111111110101101010100010;
assign LUT_1[24588] = 32'b00000000000000001000100011101100;
assign LUT_1[24589] = 32'b00000000000000000001110101101000;
assign LUT_1[24590] = 32'b00000000000000000100010001111101;
assign LUT_1[24591] = 32'b11111111111111111101100011111001;
assign LUT_1[24592] = 32'b00000000000000000011011000000010;
assign LUT_1[24593] = 32'b11111111111111111100101001111110;
assign LUT_1[24594] = 32'b11111111111111111111000110010011;
assign LUT_1[24595] = 32'b11111111111111111000011000001111;
assign LUT_1[24596] = 32'b00000000000000001011010001011001;
assign LUT_1[24597] = 32'b00000000000000000100100011010101;
assign LUT_1[24598] = 32'b00000000000000000110111111101010;
assign LUT_1[24599] = 32'b00000000000000000000010001100110;
assign LUT_1[24600] = 32'b00000000000000000010100101110111;
assign LUT_1[24601] = 32'b11111111111111111011110111110011;
assign LUT_1[24602] = 32'b11111111111111111110010100001000;
assign LUT_1[24603] = 32'b11111111111111110111100110000100;
assign LUT_1[24604] = 32'b00000000000000001010011111001110;
assign LUT_1[24605] = 32'b00000000000000000011110001001010;
assign LUT_1[24606] = 32'b00000000000000000110001101011111;
assign LUT_1[24607] = 32'b11111111111111111111011111011011;
assign LUT_1[24608] = 32'b00000000000000000010010111011111;
assign LUT_1[24609] = 32'b11111111111111111011101001011011;
assign LUT_1[24610] = 32'b11111111111111111110000101110000;
assign LUT_1[24611] = 32'b11111111111111110111010111101100;
assign LUT_1[24612] = 32'b00000000000000001010010000110110;
assign LUT_1[24613] = 32'b00000000000000000011100010110010;
assign LUT_1[24614] = 32'b00000000000000000101111111000111;
assign LUT_1[24615] = 32'b11111111111111111111010001000011;
assign LUT_1[24616] = 32'b00000000000000000001100101010100;
assign LUT_1[24617] = 32'b11111111111111111010110111010000;
assign LUT_1[24618] = 32'b11111111111111111101010011100101;
assign LUT_1[24619] = 32'b11111111111111110110100101100001;
assign LUT_1[24620] = 32'b00000000000000001001011110101011;
assign LUT_1[24621] = 32'b00000000000000000010110000100111;
assign LUT_1[24622] = 32'b00000000000000000101001100111100;
assign LUT_1[24623] = 32'b11111111111111111110011110111000;
assign LUT_1[24624] = 32'b00000000000000000100010011000001;
assign LUT_1[24625] = 32'b11111111111111111101100100111101;
assign LUT_1[24626] = 32'b00000000000000000000000001010010;
assign LUT_1[24627] = 32'b11111111111111111001010011001110;
assign LUT_1[24628] = 32'b00000000000000001100001100011000;
assign LUT_1[24629] = 32'b00000000000000000101011110010100;
assign LUT_1[24630] = 32'b00000000000000000111111010101001;
assign LUT_1[24631] = 32'b00000000000000000001001100100101;
assign LUT_1[24632] = 32'b00000000000000000011100000110110;
assign LUT_1[24633] = 32'b11111111111111111100110010110010;
assign LUT_1[24634] = 32'b11111111111111111111001111000111;
assign LUT_1[24635] = 32'b11111111111111111000100001000011;
assign LUT_1[24636] = 32'b00000000000000001011011010001101;
assign LUT_1[24637] = 32'b00000000000000000100101100001001;
assign LUT_1[24638] = 32'b00000000000000000111001000011110;
assign LUT_1[24639] = 32'b00000000000000000000011010011010;
assign LUT_1[24640] = 32'b00000000000000000011011010001000;
assign LUT_1[24641] = 32'b11111111111111111100101100000100;
assign LUT_1[24642] = 32'b11111111111111111111001000011001;
assign LUT_1[24643] = 32'b11111111111111111000011010010101;
assign LUT_1[24644] = 32'b00000000000000001011010011011111;
assign LUT_1[24645] = 32'b00000000000000000100100101011011;
assign LUT_1[24646] = 32'b00000000000000000111000001110000;
assign LUT_1[24647] = 32'b00000000000000000000010011101100;
assign LUT_1[24648] = 32'b00000000000000000010100111111101;
assign LUT_1[24649] = 32'b11111111111111111011111001111001;
assign LUT_1[24650] = 32'b11111111111111111110010110001110;
assign LUT_1[24651] = 32'b11111111111111110111101000001010;
assign LUT_1[24652] = 32'b00000000000000001010100001010100;
assign LUT_1[24653] = 32'b00000000000000000011110011010000;
assign LUT_1[24654] = 32'b00000000000000000110001111100101;
assign LUT_1[24655] = 32'b11111111111111111111100001100001;
assign LUT_1[24656] = 32'b00000000000000000101010101101010;
assign LUT_1[24657] = 32'b11111111111111111110100111100110;
assign LUT_1[24658] = 32'b00000000000000000001000011111011;
assign LUT_1[24659] = 32'b11111111111111111010010101110111;
assign LUT_1[24660] = 32'b00000000000000001101001111000001;
assign LUT_1[24661] = 32'b00000000000000000110100000111101;
assign LUT_1[24662] = 32'b00000000000000001000111101010010;
assign LUT_1[24663] = 32'b00000000000000000010001111001110;
assign LUT_1[24664] = 32'b00000000000000000100100011011111;
assign LUT_1[24665] = 32'b11111111111111111101110101011011;
assign LUT_1[24666] = 32'b00000000000000000000010001110000;
assign LUT_1[24667] = 32'b11111111111111111001100011101100;
assign LUT_1[24668] = 32'b00000000000000001100011100110110;
assign LUT_1[24669] = 32'b00000000000000000101101110110010;
assign LUT_1[24670] = 32'b00000000000000001000001011000111;
assign LUT_1[24671] = 32'b00000000000000000001011101000011;
assign LUT_1[24672] = 32'b00000000000000000100010101000111;
assign LUT_1[24673] = 32'b11111111111111111101100111000011;
assign LUT_1[24674] = 32'b00000000000000000000000011011000;
assign LUT_1[24675] = 32'b11111111111111111001010101010100;
assign LUT_1[24676] = 32'b00000000000000001100001110011110;
assign LUT_1[24677] = 32'b00000000000000000101100000011010;
assign LUT_1[24678] = 32'b00000000000000000111111100101111;
assign LUT_1[24679] = 32'b00000000000000000001001110101011;
assign LUT_1[24680] = 32'b00000000000000000011100010111100;
assign LUT_1[24681] = 32'b11111111111111111100110100111000;
assign LUT_1[24682] = 32'b11111111111111111111010001001101;
assign LUT_1[24683] = 32'b11111111111111111000100011001001;
assign LUT_1[24684] = 32'b00000000000000001011011100010011;
assign LUT_1[24685] = 32'b00000000000000000100101110001111;
assign LUT_1[24686] = 32'b00000000000000000111001010100100;
assign LUT_1[24687] = 32'b00000000000000000000011100100000;
assign LUT_1[24688] = 32'b00000000000000000110010000101001;
assign LUT_1[24689] = 32'b11111111111111111111100010100101;
assign LUT_1[24690] = 32'b00000000000000000001111110111010;
assign LUT_1[24691] = 32'b11111111111111111011010000110110;
assign LUT_1[24692] = 32'b00000000000000001110001010000000;
assign LUT_1[24693] = 32'b00000000000000000111011011111100;
assign LUT_1[24694] = 32'b00000000000000001001111000010001;
assign LUT_1[24695] = 32'b00000000000000000011001010001101;
assign LUT_1[24696] = 32'b00000000000000000101011110011110;
assign LUT_1[24697] = 32'b11111111111111111110110000011010;
assign LUT_1[24698] = 32'b00000000000000000001001100101111;
assign LUT_1[24699] = 32'b11111111111111111010011110101011;
assign LUT_1[24700] = 32'b00000000000000001101010111110101;
assign LUT_1[24701] = 32'b00000000000000000110101001110001;
assign LUT_1[24702] = 32'b00000000000000001001000110000110;
assign LUT_1[24703] = 32'b00000000000000000010011000000010;
assign LUT_1[24704] = 32'b00000000000000000100011100100011;
assign LUT_1[24705] = 32'b11111111111111111101101110011111;
assign LUT_1[24706] = 32'b00000000000000000000001010110100;
assign LUT_1[24707] = 32'b11111111111111111001011100110000;
assign LUT_1[24708] = 32'b00000000000000001100010101111010;
assign LUT_1[24709] = 32'b00000000000000000101100111110110;
assign LUT_1[24710] = 32'b00000000000000001000000100001011;
assign LUT_1[24711] = 32'b00000000000000000001010110000111;
assign LUT_1[24712] = 32'b00000000000000000011101010011000;
assign LUT_1[24713] = 32'b11111111111111111100111100010100;
assign LUT_1[24714] = 32'b11111111111111111111011000101001;
assign LUT_1[24715] = 32'b11111111111111111000101010100101;
assign LUT_1[24716] = 32'b00000000000000001011100011101111;
assign LUT_1[24717] = 32'b00000000000000000100110101101011;
assign LUT_1[24718] = 32'b00000000000000000111010010000000;
assign LUT_1[24719] = 32'b00000000000000000000100011111100;
assign LUT_1[24720] = 32'b00000000000000000110011000000101;
assign LUT_1[24721] = 32'b11111111111111111111101010000001;
assign LUT_1[24722] = 32'b00000000000000000010000110010110;
assign LUT_1[24723] = 32'b11111111111111111011011000010010;
assign LUT_1[24724] = 32'b00000000000000001110010001011100;
assign LUT_1[24725] = 32'b00000000000000000111100011011000;
assign LUT_1[24726] = 32'b00000000000000001001111111101101;
assign LUT_1[24727] = 32'b00000000000000000011010001101001;
assign LUT_1[24728] = 32'b00000000000000000101100101111010;
assign LUT_1[24729] = 32'b11111111111111111110110111110110;
assign LUT_1[24730] = 32'b00000000000000000001010100001011;
assign LUT_1[24731] = 32'b11111111111111111010100110000111;
assign LUT_1[24732] = 32'b00000000000000001101011111010001;
assign LUT_1[24733] = 32'b00000000000000000110110001001101;
assign LUT_1[24734] = 32'b00000000000000001001001101100010;
assign LUT_1[24735] = 32'b00000000000000000010011111011110;
assign LUT_1[24736] = 32'b00000000000000000101010111100010;
assign LUT_1[24737] = 32'b11111111111111111110101001011110;
assign LUT_1[24738] = 32'b00000000000000000001000101110011;
assign LUT_1[24739] = 32'b11111111111111111010010111101111;
assign LUT_1[24740] = 32'b00000000000000001101010000111001;
assign LUT_1[24741] = 32'b00000000000000000110100010110101;
assign LUT_1[24742] = 32'b00000000000000001000111111001010;
assign LUT_1[24743] = 32'b00000000000000000010010001000110;
assign LUT_1[24744] = 32'b00000000000000000100100101010111;
assign LUT_1[24745] = 32'b11111111111111111101110111010011;
assign LUT_1[24746] = 32'b00000000000000000000010011101000;
assign LUT_1[24747] = 32'b11111111111111111001100101100100;
assign LUT_1[24748] = 32'b00000000000000001100011110101110;
assign LUT_1[24749] = 32'b00000000000000000101110000101010;
assign LUT_1[24750] = 32'b00000000000000001000001100111111;
assign LUT_1[24751] = 32'b00000000000000000001011110111011;
assign LUT_1[24752] = 32'b00000000000000000111010011000100;
assign LUT_1[24753] = 32'b00000000000000000000100101000000;
assign LUT_1[24754] = 32'b00000000000000000011000001010101;
assign LUT_1[24755] = 32'b11111111111111111100010011010001;
assign LUT_1[24756] = 32'b00000000000000001111001100011011;
assign LUT_1[24757] = 32'b00000000000000001000011110010111;
assign LUT_1[24758] = 32'b00000000000000001010111010101100;
assign LUT_1[24759] = 32'b00000000000000000100001100101000;
assign LUT_1[24760] = 32'b00000000000000000110100000111001;
assign LUT_1[24761] = 32'b11111111111111111111110010110101;
assign LUT_1[24762] = 32'b00000000000000000010001111001010;
assign LUT_1[24763] = 32'b11111111111111111011100001000110;
assign LUT_1[24764] = 32'b00000000000000001110011010010000;
assign LUT_1[24765] = 32'b00000000000000000111101100001100;
assign LUT_1[24766] = 32'b00000000000000001010001000100001;
assign LUT_1[24767] = 32'b00000000000000000011011010011101;
assign LUT_1[24768] = 32'b00000000000000000110011010001011;
assign LUT_1[24769] = 32'b11111111111111111111101100000111;
assign LUT_1[24770] = 32'b00000000000000000010001000011100;
assign LUT_1[24771] = 32'b11111111111111111011011010011000;
assign LUT_1[24772] = 32'b00000000000000001110010011100010;
assign LUT_1[24773] = 32'b00000000000000000111100101011110;
assign LUT_1[24774] = 32'b00000000000000001010000001110011;
assign LUT_1[24775] = 32'b00000000000000000011010011101111;
assign LUT_1[24776] = 32'b00000000000000000101101000000000;
assign LUT_1[24777] = 32'b11111111111111111110111001111100;
assign LUT_1[24778] = 32'b00000000000000000001010110010001;
assign LUT_1[24779] = 32'b11111111111111111010101000001101;
assign LUT_1[24780] = 32'b00000000000000001101100001010111;
assign LUT_1[24781] = 32'b00000000000000000110110011010011;
assign LUT_1[24782] = 32'b00000000000000001001001111101000;
assign LUT_1[24783] = 32'b00000000000000000010100001100100;
assign LUT_1[24784] = 32'b00000000000000001000010101101101;
assign LUT_1[24785] = 32'b00000000000000000001100111101001;
assign LUT_1[24786] = 32'b00000000000000000100000011111110;
assign LUT_1[24787] = 32'b11111111111111111101010101111010;
assign LUT_1[24788] = 32'b00000000000000010000001111000100;
assign LUT_1[24789] = 32'b00000000000000001001100001000000;
assign LUT_1[24790] = 32'b00000000000000001011111101010101;
assign LUT_1[24791] = 32'b00000000000000000101001111010001;
assign LUT_1[24792] = 32'b00000000000000000111100011100010;
assign LUT_1[24793] = 32'b00000000000000000000110101011110;
assign LUT_1[24794] = 32'b00000000000000000011010001110011;
assign LUT_1[24795] = 32'b11111111111111111100100011101111;
assign LUT_1[24796] = 32'b00000000000000001111011100111001;
assign LUT_1[24797] = 32'b00000000000000001000101110110101;
assign LUT_1[24798] = 32'b00000000000000001011001011001010;
assign LUT_1[24799] = 32'b00000000000000000100011101000110;
assign LUT_1[24800] = 32'b00000000000000000111010101001010;
assign LUT_1[24801] = 32'b00000000000000000000100111000110;
assign LUT_1[24802] = 32'b00000000000000000011000011011011;
assign LUT_1[24803] = 32'b11111111111111111100010101010111;
assign LUT_1[24804] = 32'b00000000000000001111001110100001;
assign LUT_1[24805] = 32'b00000000000000001000100000011101;
assign LUT_1[24806] = 32'b00000000000000001010111100110010;
assign LUT_1[24807] = 32'b00000000000000000100001110101110;
assign LUT_1[24808] = 32'b00000000000000000110100010111111;
assign LUT_1[24809] = 32'b11111111111111111111110100111011;
assign LUT_1[24810] = 32'b00000000000000000010010001010000;
assign LUT_1[24811] = 32'b11111111111111111011100011001100;
assign LUT_1[24812] = 32'b00000000000000001110011100010110;
assign LUT_1[24813] = 32'b00000000000000000111101110010010;
assign LUT_1[24814] = 32'b00000000000000001010001010100111;
assign LUT_1[24815] = 32'b00000000000000000011011100100011;
assign LUT_1[24816] = 32'b00000000000000001001010000101100;
assign LUT_1[24817] = 32'b00000000000000000010100010101000;
assign LUT_1[24818] = 32'b00000000000000000100111110111101;
assign LUT_1[24819] = 32'b11111111111111111110010000111001;
assign LUT_1[24820] = 32'b00000000000000010001001010000011;
assign LUT_1[24821] = 32'b00000000000000001010011011111111;
assign LUT_1[24822] = 32'b00000000000000001100111000010100;
assign LUT_1[24823] = 32'b00000000000000000110001010010000;
assign LUT_1[24824] = 32'b00000000000000001000011110100001;
assign LUT_1[24825] = 32'b00000000000000000001110000011101;
assign LUT_1[24826] = 32'b00000000000000000100001100110010;
assign LUT_1[24827] = 32'b11111111111111111101011110101110;
assign LUT_1[24828] = 32'b00000000000000010000010111111000;
assign LUT_1[24829] = 32'b00000000000000001001101001110100;
assign LUT_1[24830] = 32'b00000000000000001100000110001001;
assign LUT_1[24831] = 32'b00000000000000000101011000000101;
assign LUT_1[24832] = 32'b11111111111111111111010000101100;
assign LUT_1[24833] = 32'b11111111111111111000100010101000;
assign LUT_1[24834] = 32'b11111111111111111010111110111101;
assign LUT_1[24835] = 32'b11111111111111110100010000111001;
assign LUT_1[24836] = 32'b00000000000000000111001010000011;
assign LUT_1[24837] = 32'b00000000000000000000011011111111;
assign LUT_1[24838] = 32'b00000000000000000010111000010100;
assign LUT_1[24839] = 32'b11111111111111111100001010010000;
assign LUT_1[24840] = 32'b11111111111111111110011110100001;
assign LUT_1[24841] = 32'b11111111111111110111110000011101;
assign LUT_1[24842] = 32'b11111111111111111010001100110010;
assign LUT_1[24843] = 32'b11111111111111110011011110101110;
assign LUT_1[24844] = 32'b00000000000000000110010111111000;
assign LUT_1[24845] = 32'b11111111111111111111101001110100;
assign LUT_1[24846] = 32'b00000000000000000010000110001001;
assign LUT_1[24847] = 32'b11111111111111111011011000000101;
assign LUT_1[24848] = 32'b00000000000000000001001100001110;
assign LUT_1[24849] = 32'b11111111111111111010011110001010;
assign LUT_1[24850] = 32'b11111111111111111100111010011111;
assign LUT_1[24851] = 32'b11111111111111110110001100011011;
assign LUT_1[24852] = 32'b00000000000000001001000101100101;
assign LUT_1[24853] = 32'b00000000000000000010010111100001;
assign LUT_1[24854] = 32'b00000000000000000100110011110110;
assign LUT_1[24855] = 32'b11111111111111111110000101110010;
assign LUT_1[24856] = 32'b00000000000000000000011010000011;
assign LUT_1[24857] = 32'b11111111111111111001101011111111;
assign LUT_1[24858] = 32'b11111111111111111100001000010100;
assign LUT_1[24859] = 32'b11111111111111110101011010010000;
assign LUT_1[24860] = 32'b00000000000000001000010011011010;
assign LUT_1[24861] = 32'b00000000000000000001100101010110;
assign LUT_1[24862] = 32'b00000000000000000100000001101011;
assign LUT_1[24863] = 32'b11111111111111111101010011100111;
assign LUT_1[24864] = 32'b00000000000000000000001011101011;
assign LUT_1[24865] = 32'b11111111111111111001011101100111;
assign LUT_1[24866] = 32'b11111111111111111011111001111100;
assign LUT_1[24867] = 32'b11111111111111110101001011111000;
assign LUT_1[24868] = 32'b00000000000000001000000101000010;
assign LUT_1[24869] = 32'b00000000000000000001010110111110;
assign LUT_1[24870] = 32'b00000000000000000011110011010011;
assign LUT_1[24871] = 32'b11111111111111111101000101001111;
assign LUT_1[24872] = 32'b11111111111111111111011001100000;
assign LUT_1[24873] = 32'b11111111111111111000101011011100;
assign LUT_1[24874] = 32'b11111111111111111011000111110001;
assign LUT_1[24875] = 32'b11111111111111110100011001101101;
assign LUT_1[24876] = 32'b00000000000000000111010010110111;
assign LUT_1[24877] = 32'b00000000000000000000100100110011;
assign LUT_1[24878] = 32'b00000000000000000011000001001000;
assign LUT_1[24879] = 32'b11111111111111111100010011000100;
assign LUT_1[24880] = 32'b00000000000000000010000111001101;
assign LUT_1[24881] = 32'b11111111111111111011011001001001;
assign LUT_1[24882] = 32'b11111111111111111101110101011110;
assign LUT_1[24883] = 32'b11111111111111110111000111011010;
assign LUT_1[24884] = 32'b00000000000000001010000000100100;
assign LUT_1[24885] = 32'b00000000000000000011010010100000;
assign LUT_1[24886] = 32'b00000000000000000101101110110101;
assign LUT_1[24887] = 32'b11111111111111111111000000110001;
assign LUT_1[24888] = 32'b00000000000000000001010101000010;
assign LUT_1[24889] = 32'b11111111111111111010100110111110;
assign LUT_1[24890] = 32'b11111111111111111101000011010011;
assign LUT_1[24891] = 32'b11111111111111110110010101001111;
assign LUT_1[24892] = 32'b00000000000000001001001110011001;
assign LUT_1[24893] = 32'b00000000000000000010100000010101;
assign LUT_1[24894] = 32'b00000000000000000100111100101010;
assign LUT_1[24895] = 32'b11111111111111111110001110100110;
assign LUT_1[24896] = 32'b00000000000000000001001110010100;
assign LUT_1[24897] = 32'b11111111111111111010100000010000;
assign LUT_1[24898] = 32'b11111111111111111100111100100101;
assign LUT_1[24899] = 32'b11111111111111110110001110100001;
assign LUT_1[24900] = 32'b00000000000000001001000111101011;
assign LUT_1[24901] = 32'b00000000000000000010011001100111;
assign LUT_1[24902] = 32'b00000000000000000100110101111100;
assign LUT_1[24903] = 32'b11111111111111111110000111111000;
assign LUT_1[24904] = 32'b00000000000000000000011100001001;
assign LUT_1[24905] = 32'b11111111111111111001101110000101;
assign LUT_1[24906] = 32'b11111111111111111100001010011010;
assign LUT_1[24907] = 32'b11111111111111110101011100010110;
assign LUT_1[24908] = 32'b00000000000000001000010101100000;
assign LUT_1[24909] = 32'b00000000000000000001100111011100;
assign LUT_1[24910] = 32'b00000000000000000100000011110001;
assign LUT_1[24911] = 32'b11111111111111111101010101101101;
assign LUT_1[24912] = 32'b00000000000000000011001001110110;
assign LUT_1[24913] = 32'b11111111111111111100011011110010;
assign LUT_1[24914] = 32'b11111111111111111110111000000111;
assign LUT_1[24915] = 32'b11111111111111111000001010000011;
assign LUT_1[24916] = 32'b00000000000000001011000011001101;
assign LUT_1[24917] = 32'b00000000000000000100010101001001;
assign LUT_1[24918] = 32'b00000000000000000110110001011110;
assign LUT_1[24919] = 32'b00000000000000000000000011011010;
assign LUT_1[24920] = 32'b00000000000000000010010111101011;
assign LUT_1[24921] = 32'b11111111111111111011101001100111;
assign LUT_1[24922] = 32'b11111111111111111110000101111100;
assign LUT_1[24923] = 32'b11111111111111110111010111111000;
assign LUT_1[24924] = 32'b00000000000000001010010001000010;
assign LUT_1[24925] = 32'b00000000000000000011100010111110;
assign LUT_1[24926] = 32'b00000000000000000101111111010011;
assign LUT_1[24927] = 32'b11111111111111111111010001001111;
assign LUT_1[24928] = 32'b00000000000000000010001001010011;
assign LUT_1[24929] = 32'b11111111111111111011011011001111;
assign LUT_1[24930] = 32'b11111111111111111101110111100100;
assign LUT_1[24931] = 32'b11111111111111110111001001100000;
assign LUT_1[24932] = 32'b00000000000000001010000010101010;
assign LUT_1[24933] = 32'b00000000000000000011010100100110;
assign LUT_1[24934] = 32'b00000000000000000101110000111011;
assign LUT_1[24935] = 32'b11111111111111111111000010110111;
assign LUT_1[24936] = 32'b00000000000000000001010111001000;
assign LUT_1[24937] = 32'b11111111111111111010101001000100;
assign LUT_1[24938] = 32'b11111111111111111101000101011001;
assign LUT_1[24939] = 32'b11111111111111110110010111010101;
assign LUT_1[24940] = 32'b00000000000000001001010000011111;
assign LUT_1[24941] = 32'b00000000000000000010100010011011;
assign LUT_1[24942] = 32'b00000000000000000100111110110000;
assign LUT_1[24943] = 32'b11111111111111111110010000101100;
assign LUT_1[24944] = 32'b00000000000000000100000100110101;
assign LUT_1[24945] = 32'b11111111111111111101010110110001;
assign LUT_1[24946] = 32'b11111111111111111111110011000110;
assign LUT_1[24947] = 32'b11111111111111111001000101000010;
assign LUT_1[24948] = 32'b00000000000000001011111110001100;
assign LUT_1[24949] = 32'b00000000000000000101010000001000;
assign LUT_1[24950] = 32'b00000000000000000111101100011101;
assign LUT_1[24951] = 32'b00000000000000000000111110011001;
assign LUT_1[24952] = 32'b00000000000000000011010010101010;
assign LUT_1[24953] = 32'b11111111111111111100100100100110;
assign LUT_1[24954] = 32'b11111111111111111111000000111011;
assign LUT_1[24955] = 32'b11111111111111111000010010110111;
assign LUT_1[24956] = 32'b00000000000000001011001100000001;
assign LUT_1[24957] = 32'b00000000000000000100011101111101;
assign LUT_1[24958] = 32'b00000000000000000110111010010010;
assign LUT_1[24959] = 32'b00000000000000000000001100001110;
assign LUT_1[24960] = 32'b00000000000000000010010000101111;
assign LUT_1[24961] = 32'b11111111111111111011100010101011;
assign LUT_1[24962] = 32'b11111111111111111101111111000000;
assign LUT_1[24963] = 32'b11111111111111110111010000111100;
assign LUT_1[24964] = 32'b00000000000000001010001010000110;
assign LUT_1[24965] = 32'b00000000000000000011011100000010;
assign LUT_1[24966] = 32'b00000000000000000101111000010111;
assign LUT_1[24967] = 32'b11111111111111111111001010010011;
assign LUT_1[24968] = 32'b00000000000000000001011110100100;
assign LUT_1[24969] = 32'b11111111111111111010110000100000;
assign LUT_1[24970] = 32'b11111111111111111101001100110101;
assign LUT_1[24971] = 32'b11111111111111110110011110110001;
assign LUT_1[24972] = 32'b00000000000000001001010111111011;
assign LUT_1[24973] = 32'b00000000000000000010101001110111;
assign LUT_1[24974] = 32'b00000000000000000101000110001100;
assign LUT_1[24975] = 32'b11111111111111111110011000001000;
assign LUT_1[24976] = 32'b00000000000000000100001100010001;
assign LUT_1[24977] = 32'b11111111111111111101011110001101;
assign LUT_1[24978] = 32'b11111111111111111111111010100010;
assign LUT_1[24979] = 32'b11111111111111111001001100011110;
assign LUT_1[24980] = 32'b00000000000000001100000101101000;
assign LUT_1[24981] = 32'b00000000000000000101010111100100;
assign LUT_1[24982] = 32'b00000000000000000111110011111001;
assign LUT_1[24983] = 32'b00000000000000000001000101110101;
assign LUT_1[24984] = 32'b00000000000000000011011010000110;
assign LUT_1[24985] = 32'b11111111111111111100101100000010;
assign LUT_1[24986] = 32'b11111111111111111111001000010111;
assign LUT_1[24987] = 32'b11111111111111111000011010010011;
assign LUT_1[24988] = 32'b00000000000000001011010011011101;
assign LUT_1[24989] = 32'b00000000000000000100100101011001;
assign LUT_1[24990] = 32'b00000000000000000111000001101110;
assign LUT_1[24991] = 32'b00000000000000000000010011101010;
assign LUT_1[24992] = 32'b00000000000000000011001011101110;
assign LUT_1[24993] = 32'b11111111111111111100011101101010;
assign LUT_1[24994] = 32'b11111111111111111110111001111111;
assign LUT_1[24995] = 32'b11111111111111111000001011111011;
assign LUT_1[24996] = 32'b00000000000000001011000101000101;
assign LUT_1[24997] = 32'b00000000000000000100010111000001;
assign LUT_1[24998] = 32'b00000000000000000110110011010110;
assign LUT_1[24999] = 32'b00000000000000000000000101010010;
assign LUT_1[25000] = 32'b00000000000000000010011001100011;
assign LUT_1[25001] = 32'b11111111111111111011101011011111;
assign LUT_1[25002] = 32'b11111111111111111110000111110100;
assign LUT_1[25003] = 32'b11111111111111110111011001110000;
assign LUT_1[25004] = 32'b00000000000000001010010010111010;
assign LUT_1[25005] = 32'b00000000000000000011100100110110;
assign LUT_1[25006] = 32'b00000000000000000110000001001011;
assign LUT_1[25007] = 32'b11111111111111111111010011000111;
assign LUT_1[25008] = 32'b00000000000000000101000111010000;
assign LUT_1[25009] = 32'b11111111111111111110011001001100;
assign LUT_1[25010] = 32'b00000000000000000000110101100001;
assign LUT_1[25011] = 32'b11111111111111111010000111011101;
assign LUT_1[25012] = 32'b00000000000000001101000000100111;
assign LUT_1[25013] = 32'b00000000000000000110010010100011;
assign LUT_1[25014] = 32'b00000000000000001000101110111000;
assign LUT_1[25015] = 32'b00000000000000000010000000110100;
assign LUT_1[25016] = 32'b00000000000000000100010101000101;
assign LUT_1[25017] = 32'b11111111111111111101100111000001;
assign LUT_1[25018] = 32'b00000000000000000000000011010110;
assign LUT_1[25019] = 32'b11111111111111111001010101010010;
assign LUT_1[25020] = 32'b00000000000000001100001110011100;
assign LUT_1[25021] = 32'b00000000000000000101100000011000;
assign LUT_1[25022] = 32'b00000000000000000111111100101101;
assign LUT_1[25023] = 32'b00000000000000000001001110101001;
assign LUT_1[25024] = 32'b00000000000000000100001110010111;
assign LUT_1[25025] = 32'b11111111111111111101100000010011;
assign LUT_1[25026] = 32'b11111111111111111111111100101000;
assign LUT_1[25027] = 32'b11111111111111111001001110100100;
assign LUT_1[25028] = 32'b00000000000000001100000111101110;
assign LUT_1[25029] = 32'b00000000000000000101011001101010;
assign LUT_1[25030] = 32'b00000000000000000111110101111111;
assign LUT_1[25031] = 32'b00000000000000000001000111111011;
assign LUT_1[25032] = 32'b00000000000000000011011100001100;
assign LUT_1[25033] = 32'b11111111111111111100101110001000;
assign LUT_1[25034] = 32'b11111111111111111111001010011101;
assign LUT_1[25035] = 32'b11111111111111111000011100011001;
assign LUT_1[25036] = 32'b00000000000000001011010101100011;
assign LUT_1[25037] = 32'b00000000000000000100100111011111;
assign LUT_1[25038] = 32'b00000000000000000111000011110100;
assign LUT_1[25039] = 32'b00000000000000000000010101110000;
assign LUT_1[25040] = 32'b00000000000000000110001001111001;
assign LUT_1[25041] = 32'b11111111111111111111011011110101;
assign LUT_1[25042] = 32'b00000000000000000001111000001010;
assign LUT_1[25043] = 32'b11111111111111111011001010000110;
assign LUT_1[25044] = 32'b00000000000000001110000011010000;
assign LUT_1[25045] = 32'b00000000000000000111010101001100;
assign LUT_1[25046] = 32'b00000000000000001001110001100001;
assign LUT_1[25047] = 32'b00000000000000000011000011011101;
assign LUT_1[25048] = 32'b00000000000000000101010111101110;
assign LUT_1[25049] = 32'b11111111111111111110101001101010;
assign LUT_1[25050] = 32'b00000000000000000001000101111111;
assign LUT_1[25051] = 32'b11111111111111111010010111111011;
assign LUT_1[25052] = 32'b00000000000000001101010001000101;
assign LUT_1[25053] = 32'b00000000000000000110100011000001;
assign LUT_1[25054] = 32'b00000000000000001000111111010110;
assign LUT_1[25055] = 32'b00000000000000000010010001010010;
assign LUT_1[25056] = 32'b00000000000000000101001001010110;
assign LUT_1[25057] = 32'b11111111111111111110011011010010;
assign LUT_1[25058] = 32'b00000000000000000000110111100111;
assign LUT_1[25059] = 32'b11111111111111111010001001100011;
assign LUT_1[25060] = 32'b00000000000000001101000010101101;
assign LUT_1[25061] = 32'b00000000000000000110010100101001;
assign LUT_1[25062] = 32'b00000000000000001000110000111110;
assign LUT_1[25063] = 32'b00000000000000000010000010111010;
assign LUT_1[25064] = 32'b00000000000000000100010111001011;
assign LUT_1[25065] = 32'b11111111111111111101101001000111;
assign LUT_1[25066] = 32'b00000000000000000000000101011100;
assign LUT_1[25067] = 32'b11111111111111111001010111011000;
assign LUT_1[25068] = 32'b00000000000000001100010000100010;
assign LUT_1[25069] = 32'b00000000000000000101100010011110;
assign LUT_1[25070] = 32'b00000000000000000111111110110011;
assign LUT_1[25071] = 32'b00000000000000000001010000101111;
assign LUT_1[25072] = 32'b00000000000000000111000100111000;
assign LUT_1[25073] = 32'b00000000000000000000010110110100;
assign LUT_1[25074] = 32'b00000000000000000010110011001001;
assign LUT_1[25075] = 32'b11111111111111111100000101000101;
assign LUT_1[25076] = 32'b00000000000000001110111110001111;
assign LUT_1[25077] = 32'b00000000000000001000010000001011;
assign LUT_1[25078] = 32'b00000000000000001010101100100000;
assign LUT_1[25079] = 32'b00000000000000000011111110011100;
assign LUT_1[25080] = 32'b00000000000000000110010010101101;
assign LUT_1[25081] = 32'b11111111111111111111100100101001;
assign LUT_1[25082] = 32'b00000000000000000010000000111110;
assign LUT_1[25083] = 32'b11111111111111111011010010111010;
assign LUT_1[25084] = 32'b00000000000000001110001100000100;
assign LUT_1[25085] = 32'b00000000000000000111011110000000;
assign LUT_1[25086] = 32'b00000000000000001001111010010101;
assign LUT_1[25087] = 32'b00000000000000000011001100010001;
assign LUT_1[25088] = 32'b11111111111111111011001010111101;
assign LUT_1[25089] = 32'b11111111111111110100011100111001;
assign LUT_1[25090] = 32'b11111111111111110110111001001110;
assign LUT_1[25091] = 32'b11111111111111110000001011001010;
assign LUT_1[25092] = 32'b00000000000000000011000100010100;
assign LUT_1[25093] = 32'b11111111111111111100010110010000;
assign LUT_1[25094] = 32'b11111111111111111110110010100101;
assign LUT_1[25095] = 32'b11111111111111111000000100100001;
assign LUT_1[25096] = 32'b11111111111111111010011000110010;
assign LUT_1[25097] = 32'b11111111111111110011101010101110;
assign LUT_1[25098] = 32'b11111111111111110110000111000011;
assign LUT_1[25099] = 32'b11111111111111101111011000111111;
assign LUT_1[25100] = 32'b00000000000000000010010010001001;
assign LUT_1[25101] = 32'b11111111111111111011100100000101;
assign LUT_1[25102] = 32'b11111111111111111110000000011010;
assign LUT_1[25103] = 32'b11111111111111110111010010010110;
assign LUT_1[25104] = 32'b11111111111111111101000110011111;
assign LUT_1[25105] = 32'b11111111111111110110011000011011;
assign LUT_1[25106] = 32'b11111111111111111000110100110000;
assign LUT_1[25107] = 32'b11111111111111110010000110101100;
assign LUT_1[25108] = 32'b00000000000000000100111111110110;
assign LUT_1[25109] = 32'b11111111111111111110010001110010;
assign LUT_1[25110] = 32'b00000000000000000000101110000111;
assign LUT_1[25111] = 32'b11111111111111111010000000000011;
assign LUT_1[25112] = 32'b11111111111111111100010100010100;
assign LUT_1[25113] = 32'b11111111111111110101100110010000;
assign LUT_1[25114] = 32'b11111111111111111000000010100101;
assign LUT_1[25115] = 32'b11111111111111110001010100100001;
assign LUT_1[25116] = 32'b00000000000000000100001101101011;
assign LUT_1[25117] = 32'b11111111111111111101011111100111;
assign LUT_1[25118] = 32'b11111111111111111111111011111100;
assign LUT_1[25119] = 32'b11111111111111111001001101111000;
assign LUT_1[25120] = 32'b11111111111111111100000101111100;
assign LUT_1[25121] = 32'b11111111111111110101010111111000;
assign LUT_1[25122] = 32'b11111111111111110111110100001101;
assign LUT_1[25123] = 32'b11111111111111110001000110001001;
assign LUT_1[25124] = 32'b00000000000000000011111111010011;
assign LUT_1[25125] = 32'b11111111111111111101010001001111;
assign LUT_1[25126] = 32'b11111111111111111111101101100100;
assign LUT_1[25127] = 32'b11111111111111111000111111100000;
assign LUT_1[25128] = 32'b11111111111111111011010011110001;
assign LUT_1[25129] = 32'b11111111111111110100100101101101;
assign LUT_1[25130] = 32'b11111111111111110111000010000010;
assign LUT_1[25131] = 32'b11111111111111110000010011111110;
assign LUT_1[25132] = 32'b00000000000000000011001101001000;
assign LUT_1[25133] = 32'b11111111111111111100011111000100;
assign LUT_1[25134] = 32'b11111111111111111110111011011001;
assign LUT_1[25135] = 32'b11111111111111111000001101010101;
assign LUT_1[25136] = 32'b11111111111111111110000001011110;
assign LUT_1[25137] = 32'b11111111111111110111010011011010;
assign LUT_1[25138] = 32'b11111111111111111001101111101111;
assign LUT_1[25139] = 32'b11111111111111110011000001101011;
assign LUT_1[25140] = 32'b00000000000000000101111010110101;
assign LUT_1[25141] = 32'b11111111111111111111001100110001;
assign LUT_1[25142] = 32'b00000000000000000001101001000110;
assign LUT_1[25143] = 32'b11111111111111111010111011000010;
assign LUT_1[25144] = 32'b11111111111111111101001111010011;
assign LUT_1[25145] = 32'b11111111111111110110100001001111;
assign LUT_1[25146] = 32'b11111111111111111000111101100100;
assign LUT_1[25147] = 32'b11111111111111110010001111100000;
assign LUT_1[25148] = 32'b00000000000000000101001000101010;
assign LUT_1[25149] = 32'b11111111111111111110011010100110;
assign LUT_1[25150] = 32'b00000000000000000000110110111011;
assign LUT_1[25151] = 32'b11111111111111111010001000110111;
assign LUT_1[25152] = 32'b11111111111111111101001000100101;
assign LUT_1[25153] = 32'b11111111111111110110011010100001;
assign LUT_1[25154] = 32'b11111111111111111000110110110110;
assign LUT_1[25155] = 32'b11111111111111110010001000110010;
assign LUT_1[25156] = 32'b00000000000000000101000001111100;
assign LUT_1[25157] = 32'b11111111111111111110010011111000;
assign LUT_1[25158] = 32'b00000000000000000000110000001101;
assign LUT_1[25159] = 32'b11111111111111111010000010001001;
assign LUT_1[25160] = 32'b11111111111111111100010110011010;
assign LUT_1[25161] = 32'b11111111111111110101101000010110;
assign LUT_1[25162] = 32'b11111111111111111000000100101011;
assign LUT_1[25163] = 32'b11111111111111110001010110100111;
assign LUT_1[25164] = 32'b00000000000000000100001111110001;
assign LUT_1[25165] = 32'b11111111111111111101100001101101;
assign LUT_1[25166] = 32'b11111111111111111111111110000010;
assign LUT_1[25167] = 32'b11111111111111111001001111111110;
assign LUT_1[25168] = 32'b11111111111111111111000100000111;
assign LUT_1[25169] = 32'b11111111111111111000010110000011;
assign LUT_1[25170] = 32'b11111111111111111010110010011000;
assign LUT_1[25171] = 32'b11111111111111110100000100010100;
assign LUT_1[25172] = 32'b00000000000000000110111101011110;
assign LUT_1[25173] = 32'b00000000000000000000001111011010;
assign LUT_1[25174] = 32'b00000000000000000010101011101111;
assign LUT_1[25175] = 32'b11111111111111111011111101101011;
assign LUT_1[25176] = 32'b11111111111111111110010001111100;
assign LUT_1[25177] = 32'b11111111111111110111100011111000;
assign LUT_1[25178] = 32'b11111111111111111010000000001101;
assign LUT_1[25179] = 32'b11111111111111110011010010001001;
assign LUT_1[25180] = 32'b00000000000000000110001011010011;
assign LUT_1[25181] = 32'b11111111111111111111011101001111;
assign LUT_1[25182] = 32'b00000000000000000001111001100100;
assign LUT_1[25183] = 32'b11111111111111111011001011100000;
assign LUT_1[25184] = 32'b11111111111111111110000011100100;
assign LUT_1[25185] = 32'b11111111111111110111010101100000;
assign LUT_1[25186] = 32'b11111111111111111001110001110101;
assign LUT_1[25187] = 32'b11111111111111110011000011110001;
assign LUT_1[25188] = 32'b00000000000000000101111100111011;
assign LUT_1[25189] = 32'b11111111111111111111001110110111;
assign LUT_1[25190] = 32'b00000000000000000001101011001100;
assign LUT_1[25191] = 32'b11111111111111111010111101001000;
assign LUT_1[25192] = 32'b11111111111111111101010001011001;
assign LUT_1[25193] = 32'b11111111111111110110100011010101;
assign LUT_1[25194] = 32'b11111111111111111000111111101010;
assign LUT_1[25195] = 32'b11111111111111110010010001100110;
assign LUT_1[25196] = 32'b00000000000000000101001010110000;
assign LUT_1[25197] = 32'b11111111111111111110011100101100;
assign LUT_1[25198] = 32'b00000000000000000000111001000001;
assign LUT_1[25199] = 32'b11111111111111111010001010111101;
assign LUT_1[25200] = 32'b11111111111111111111111111000110;
assign LUT_1[25201] = 32'b11111111111111111001010001000010;
assign LUT_1[25202] = 32'b11111111111111111011101101010111;
assign LUT_1[25203] = 32'b11111111111111110100111111010011;
assign LUT_1[25204] = 32'b00000000000000000111111000011101;
assign LUT_1[25205] = 32'b00000000000000000001001010011001;
assign LUT_1[25206] = 32'b00000000000000000011100110101110;
assign LUT_1[25207] = 32'b11111111111111111100111000101010;
assign LUT_1[25208] = 32'b11111111111111111111001100111011;
assign LUT_1[25209] = 32'b11111111111111111000011110110111;
assign LUT_1[25210] = 32'b11111111111111111010111011001100;
assign LUT_1[25211] = 32'b11111111111111110100001101001000;
assign LUT_1[25212] = 32'b00000000000000000111000110010010;
assign LUT_1[25213] = 32'b00000000000000000000011000001110;
assign LUT_1[25214] = 32'b00000000000000000010110100100011;
assign LUT_1[25215] = 32'b11111111111111111100000110011111;
assign LUT_1[25216] = 32'b11111111111111111110001011000000;
assign LUT_1[25217] = 32'b11111111111111110111011100111100;
assign LUT_1[25218] = 32'b11111111111111111001111001010001;
assign LUT_1[25219] = 32'b11111111111111110011001011001101;
assign LUT_1[25220] = 32'b00000000000000000110000100010111;
assign LUT_1[25221] = 32'b11111111111111111111010110010011;
assign LUT_1[25222] = 32'b00000000000000000001110010101000;
assign LUT_1[25223] = 32'b11111111111111111011000100100100;
assign LUT_1[25224] = 32'b11111111111111111101011000110101;
assign LUT_1[25225] = 32'b11111111111111110110101010110001;
assign LUT_1[25226] = 32'b11111111111111111001000111000110;
assign LUT_1[25227] = 32'b11111111111111110010011001000010;
assign LUT_1[25228] = 32'b00000000000000000101010010001100;
assign LUT_1[25229] = 32'b11111111111111111110100100001000;
assign LUT_1[25230] = 32'b00000000000000000001000000011101;
assign LUT_1[25231] = 32'b11111111111111111010010010011001;
assign LUT_1[25232] = 32'b00000000000000000000000110100010;
assign LUT_1[25233] = 32'b11111111111111111001011000011110;
assign LUT_1[25234] = 32'b11111111111111111011110100110011;
assign LUT_1[25235] = 32'b11111111111111110101000110101111;
assign LUT_1[25236] = 32'b00000000000000000111111111111001;
assign LUT_1[25237] = 32'b00000000000000000001010001110101;
assign LUT_1[25238] = 32'b00000000000000000011101110001010;
assign LUT_1[25239] = 32'b11111111111111111101000000000110;
assign LUT_1[25240] = 32'b11111111111111111111010100010111;
assign LUT_1[25241] = 32'b11111111111111111000100110010011;
assign LUT_1[25242] = 32'b11111111111111111011000010101000;
assign LUT_1[25243] = 32'b11111111111111110100010100100100;
assign LUT_1[25244] = 32'b00000000000000000111001101101110;
assign LUT_1[25245] = 32'b00000000000000000000011111101010;
assign LUT_1[25246] = 32'b00000000000000000010111011111111;
assign LUT_1[25247] = 32'b11111111111111111100001101111011;
assign LUT_1[25248] = 32'b11111111111111111111000101111111;
assign LUT_1[25249] = 32'b11111111111111111000010111111011;
assign LUT_1[25250] = 32'b11111111111111111010110100010000;
assign LUT_1[25251] = 32'b11111111111111110100000110001100;
assign LUT_1[25252] = 32'b00000000000000000110111111010110;
assign LUT_1[25253] = 32'b00000000000000000000010001010010;
assign LUT_1[25254] = 32'b00000000000000000010101101100111;
assign LUT_1[25255] = 32'b11111111111111111011111111100011;
assign LUT_1[25256] = 32'b11111111111111111110010011110100;
assign LUT_1[25257] = 32'b11111111111111110111100101110000;
assign LUT_1[25258] = 32'b11111111111111111010000010000101;
assign LUT_1[25259] = 32'b11111111111111110011010100000001;
assign LUT_1[25260] = 32'b00000000000000000110001101001011;
assign LUT_1[25261] = 32'b11111111111111111111011111000111;
assign LUT_1[25262] = 32'b00000000000000000001111011011100;
assign LUT_1[25263] = 32'b11111111111111111011001101011000;
assign LUT_1[25264] = 32'b00000000000000000001000001100001;
assign LUT_1[25265] = 32'b11111111111111111010010011011101;
assign LUT_1[25266] = 32'b11111111111111111100101111110010;
assign LUT_1[25267] = 32'b11111111111111110110000001101110;
assign LUT_1[25268] = 32'b00000000000000001000111010111000;
assign LUT_1[25269] = 32'b00000000000000000010001100110100;
assign LUT_1[25270] = 32'b00000000000000000100101001001001;
assign LUT_1[25271] = 32'b11111111111111111101111011000101;
assign LUT_1[25272] = 32'b00000000000000000000001111010110;
assign LUT_1[25273] = 32'b11111111111111111001100001010010;
assign LUT_1[25274] = 32'b11111111111111111011111101100111;
assign LUT_1[25275] = 32'b11111111111111110101001111100011;
assign LUT_1[25276] = 32'b00000000000000001000001000101101;
assign LUT_1[25277] = 32'b00000000000000000001011010101001;
assign LUT_1[25278] = 32'b00000000000000000011110110111110;
assign LUT_1[25279] = 32'b11111111111111111101001000111010;
assign LUT_1[25280] = 32'b00000000000000000000001000101000;
assign LUT_1[25281] = 32'b11111111111111111001011010100100;
assign LUT_1[25282] = 32'b11111111111111111011110110111001;
assign LUT_1[25283] = 32'b11111111111111110101001000110101;
assign LUT_1[25284] = 32'b00000000000000001000000001111111;
assign LUT_1[25285] = 32'b00000000000000000001010011111011;
assign LUT_1[25286] = 32'b00000000000000000011110000010000;
assign LUT_1[25287] = 32'b11111111111111111101000010001100;
assign LUT_1[25288] = 32'b11111111111111111111010110011101;
assign LUT_1[25289] = 32'b11111111111111111000101000011001;
assign LUT_1[25290] = 32'b11111111111111111011000100101110;
assign LUT_1[25291] = 32'b11111111111111110100010110101010;
assign LUT_1[25292] = 32'b00000000000000000111001111110100;
assign LUT_1[25293] = 32'b00000000000000000000100001110000;
assign LUT_1[25294] = 32'b00000000000000000010111110000101;
assign LUT_1[25295] = 32'b11111111111111111100010000000001;
assign LUT_1[25296] = 32'b00000000000000000010000100001010;
assign LUT_1[25297] = 32'b11111111111111111011010110000110;
assign LUT_1[25298] = 32'b11111111111111111101110010011011;
assign LUT_1[25299] = 32'b11111111111111110111000100010111;
assign LUT_1[25300] = 32'b00000000000000001001111101100001;
assign LUT_1[25301] = 32'b00000000000000000011001111011101;
assign LUT_1[25302] = 32'b00000000000000000101101011110010;
assign LUT_1[25303] = 32'b11111111111111111110111101101110;
assign LUT_1[25304] = 32'b00000000000000000001010001111111;
assign LUT_1[25305] = 32'b11111111111111111010100011111011;
assign LUT_1[25306] = 32'b11111111111111111101000000010000;
assign LUT_1[25307] = 32'b11111111111111110110010010001100;
assign LUT_1[25308] = 32'b00000000000000001001001011010110;
assign LUT_1[25309] = 32'b00000000000000000010011101010010;
assign LUT_1[25310] = 32'b00000000000000000100111001100111;
assign LUT_1[25311] = 32'b11111111111111111110001011100011;
assign LUT_1[25312] = 32'b00000000000000000001000011100111;
assign LUT_1[25313] = 32'b11111111111111111010010101100011;
assign LUT_1[25314] = 32'b11111111111111111100110001111000;
assign LUT_1[25315] = 32'b11111111111111110110000011110100;
assign LUT_1[25316] = 32'b00000000000000001000111100111110;
assign LUT_1[25317] = 32'b00000000000000000010001110111010;
assign LUT_1[25318] = 32'b00000000000000000100101011001111;
assign LUT_1[25319] = 32'b11111111111111111101111101001011;
assign LUT_1[25320] = 32'b00000000000000000000010001011100;
assign LUT_1[25321] = 32'b11111111111111111001100011011000;
assign LUT_1[25322] = 32'b11111111111111111011111111101101;
assign LUT_1[25323] = 32'b11111111111111110101010001101001;
assign LUT_1[25324] = 32'b00000000000000001000001010110011;
assign LUT_1[25325] = 32'b00000000000000000001011100101111;
assign LUT_1[25326] = 32'b00000000000000000011111001000100;
assign LUT_1[25327] = 32'b11111111111111111101001011000000;
assign LUT_1[25328] = 32'b00000000000000000010111111001001;
assign LUT_1[25329] = 32'b11111111111111111100010001000101;
assign LUT_1[25330] = 32'b11111111111111111110101101011010;
assign LUT_1[25331] = 32'b11111111111111110111111111010110;
assign LUT_1[25332] = 32'b00000000000000001010111000100000;
assign LUT_1[25333] = 32'b00000000000000000100001010011100;
assign LUT_1[25334] = 32'b00000000000000000110100110110001;
assign LUT_1[25335] = 32'b11111111111111111111111000101101;
assign LUT_1[25336] = 32'b00000000000000000010001100111110;
assign LUT_1[25337] = 32'b11111111111111111011011110111010;
assign LUT_1[25338] = 32'b11111111111111111101111011001111;
assign LUT_1[25339] = 32'b11111111111111110111001101001011;
assign LUT_1[25340] = 32'b00000000000000001010000110010101;
assign LUT_1[25341] = 32'b00000000000000000011011000010001;
assign LUT_1[25342] = 32'b00000000000000000101110100100110;
assign LUT_1[25343] = 32'b11111111111111111111000110100010;
assign LUT_1[25344] = 32'b11111111111111111000111111001001;
assign LUT_1[25345] = 32'b11111111111111110010010001000101;
assign LUT_1[25346] = 32'b11111111111111110100101101011010;
assign LUT_1[25347] = 32'b11111111111111101101111111010110;
assign LUT_1[25348] = 32'b00000000000000000000111000100000;
assign LUT_1[25349] = 32'b11111111111111111010001010011100;
assign LUT_1[25350] = 32'b11111111111111111100100110110001;
assign LUT_1[25351] = 32'b11111111111111110101111000101101;
assign LUT_1[25352] = 32'b11111111111111111000001100111110;
assign LUT_1[25353] = 32'b11111111111111110001011110111010;
assign LUT_1[25354] = 32'b11111111111111110011111011001111;
assign LUT_1[25355] = 32'b11111111111111101101001101001011;
assign LUT_1[25356] = 32'b00000000000000000000000110010101;
assign LUT_1[25357] = 32'b11111111111111111001011000010001;
assign LUT_1[25358] = 32'b11111111111111111011110100100110;
assign LUT_1[25359] = 32'b11111111111111110101000110100010;
assign LUT_1[25360] = 32'b11111111111111111010111010101011;
assign LUT_1[25361] = 32'b11111111111111110100001100100111;
assign LUT_1[25362] = 32'b11111111111111110110101000111100;
assign LUT_1[25363] = 32'b11111111111111101111111010111000;
assign LUT_1[25364] = 32'b00000000000000000010110100000010;
assign LUT_1[25365] = 32'b11111111111111111100000101111110;
assign LUT_1[25366] = 32'b11111111111111111110100010010011;
assign LUT_1[25367] = 32'b11111111111111110111110100001111;
assign LUT_1[25368] = 32'b11111111111111111010001000100000;
assign LUT_1[25369] = 32'b11111111111111110011011010011100;
assign LUT_1[25370] = 32'b11111111111111110101110110110001;
assign LUT_1[25371] = 32'b11111111111111101111001000101101;
assign LUT_1[25372] = 32'b00000000000000000010000001110111;
assign LUT_1[25373] = 32'b11111111111111111011010011110011;
assign LUT_1[25374] = 32'b11111111111111111101110000001000;
assign LUT_1[25375] = 32'b11111111111111110111000010000100;
assign LUT_1[25376] = 32'b11111111111111111001111010001000;
assign LUT_1[25377] = 32'b11111111111111110011001100000100;
assign LUT_1[25378] = 32'b11111111111111110101101000011001;
assign LUT_1[25379] = 32'b11111111111111101110111010010101;
assign LUT_1[25380] = 32'b00000000000000000001110011011111;
assign LUT_1[25381] = 32'b11111111111111111011000101011011;
assign LUT_1[25382] = 32'b11111111111111111101100001110000;
assign LUT_1[25383] = 32'b11111111111111110110110011101100;
assign LUT_1[25384] = 32'b11111111111111111001000111111101;
assign LUT_1[25385] = 32'b11111111111111110010011001111001;
assign LUT_1[25386] = 32'b11111111111111110100110110001110;
assign LUT_1[25387] = 32'b11111111111111101110001000001010;
assign LUT_1[25388] = 32'b00000000000000000001000001010100;
assign LUT_1[25389] = 32'b11111111111111111010010011010000;
assign LUT_1[25390] = 32'b11111111111111111100101111100101;
assign LUT_1[25391] = 32'b11111111111111110110000001100001;
assign LUT_1[25392] = 32'b11111111111111111011110101101010;
assign LUT_1[25393] = 32'b11111111111111110101000111100110;
assign LUT_1[25394] = 32'b11111111111111110111100011111011;
assign LUT_1[25395] = 32'b11111111111111110000110101110111;
assign LUT_1[25396] = 32'b00000000000000000011101111000001;
assign LUT_1[25397] = 32'b11111111111111111101000000111101;
assign LUT_1[25398] = 32'b11111111111111111111011101010010;
assign LUT_1[25399] = 32'b11111111111111111000101111001110;
assign LUT_1[25400] = 32'b11111111111111111011000011011111;
assign LUT_1[25401] = 32'b11111111111111110100010101011011;
assign LUT_1[25402] = 32'b11111111111111110110110001110000;
assign LUT_1[25403] = 32'b11111111111111110000000011101100;
assign LUT_1[25404] = 32'b00000000000000000010111100110110;
assign LUT_1[25405] = 32'b11111111111111111100001110110010;
assign LUT_1[25406] = 32'b11111111111111111110101011000111;
assign LUT_1[25407] = 32'b11111111111111110111111101000011;
assign LUT_1[25408] = 32'b11111111111111111010111100110001;
assign LUT_1[25409] = 32'b11111111111111110100001110101101;
assign LUT_1[25410] = 32'b11111111111111110110101011000010;
assign LUT_1[25411] = 32'b11111111111111101111111100111110;
assign LUT_1[25412] = 32'b00000000000000000010110110001000;
assign LUT_1[25413] = 32'b11111111111111111100001000000100;
assign LUT_1[25414] = 32'b11111111111111111110100100011001;
assign LUT_1[25415] = 32'b11111111111111110111110110010101;
assign LUT_1[25416] = 32'b11111111111111111010001010100110;
assign LUT_1[25417] = 32'b11111111111111110011011100100010;
assign LUT_1[25418] = 32'b11111111111111110101111000110111;
assign LUT_1[25419] = 32'b11111111111111101111001010110011;
assign LUT_1[25420] = 32'b00000000000000000010000011111101;
assign LUT_1[25421] = 32'b11111111111111111011010101111001;
assign LUT_1[25422] = 32'b11111111111111111101110010001110;
assign LUT_1[25423] = 32'b11111111111111110111000100001010;
assign LUT_1[25424] = 32'b11111111111111111100111000010011;
assign LUT_1[25425] = 32'b11111111111111110110001010001111;
assign LUT_1[25426] = 32'b11111111111111111000100110100100;
assign LUT_1[25427] = 32'b11111111111111110001111000100000;
assign LUT_1[25428] = 32'b00000000000000000100110001101010;
assign LUT_1[25429] = 32'b11111111111111111110000011100110;
assign LUT_1[25430] = 32'b00000000000000000000011111111011;
assign LUT_1[25431] = 32'b11111111111111111001110001110111;
assign LUT_1[25432] = 32'b11111111111111111100000110001000;
assign LUT_1[25433] = 32'b11111111111111110101011000000100;
assign LUT_1[25434] = 32'b11111111111111110111110100011001;
assign LUT_1[25435] = 32'b11111111111111110001000110010101;
assign LUT_1[25436] = 32'b00000000000000000011111111011111;
assign LUT_1[25437] = 32'b11111111111111111101010001011011;
assign LUT_1[25438] = 32'b11111111111111111111101101110000;
assign LUT_1[25439] = 32'b11111111111111111000111111101100;
assign LUT_1[25440] = 32'b11111111111111111011110111110000;
assign LUT_1[25441] = 32'b11111111111111110101001001101100;
assign LUT_1[25442] = 32'b11111111111111110111100110000001;
assign LUT_1[25443] = 32'b11111111111111110000110111111101;
assign LUT_1[25444] = 32'b00000000000000000011110001000111;
assign LUT_1[25445] = 32'b11111111111111111101000011000011;
assign LUT_1[25446] = 32'b11111111111111111111011111011000;
assign LUT_1[25447] = 32'b11111111111111111000110001010100;
assign LUT_1[25448] = 32'b11111111111111111011000101100101;
assign LUT_1[25449] = 32'b11111111111111110100010111100001;
assign LUT_1[25450] = 32'b11111111111111110110110011110110;
assign LUT_1[25451] = 32'b11111111111111110000000101110010;
assign LUT_1[25452] = 32'b00000000000000000010111110111100;
assign LUT_1[25453] = 32'b11111111111111111100010000111000;
assign LUT_1[25454] = 32'b11111111111111111110101101001101;
assign LUT_1[25455] = 32'b11111111111111110111111111001001;
assign LUT_1[25456] = 32'b11111111111111111101110011010010;
assign LUT_1[25457] = 32'b11111111111111110111000101001110;
assign LUT_1[25458] = 32'b11111111111111111001100001100011;
assign LUT_1[25459] = 32'b11111111111111110010110011011111;
assign LUT_1[25460] = 32'b00000000000000000101101100101001;
assign LUT_1[25461] = 32'b11111111111111111110111110100101;
assign LUT_1[25462] = 32'b00000000000000000001011010111010;
assign LUT_1[25463] = 32'b11111111111111111010101100110110;
assign LUT_1[25464] = 32'b11111111111111111101000001000111;
assign LUT_1[25465] = 32'b11111111111111110110010011000011;
assign LUT_1[25466] = 32'b11111111111111111000101111011000;
assign LUT_1[25467] = 32'b11111111111111110010000001010100;
assign LUT_1[25468] = 32'b00000000000000000100111010011110;
assign LUT_1[25469] = 32'b11111111111111111110001100011010;
assign LUT_1[25470] = 32'b00000000000000000000101000101111;
assign LUT_1[25471] = 32'b11111111111111111001111010101011;
assign LUT_1[25472] = 32'b11111111111111111011111111001100;
assign LUT_1[25473] = 32'b11111111111111110101010001001000;
assign LUT_1[25474] = 32'b11111111111111110111101101011101;
assign LUT_1[25475] = 32'b11111111111111110000111111011001;
assign LUT_1[25476] = 32'b00000000000000000011111000100011;
assign LUT_1[25477] = 32'b11111111111111111101001010011111;
assign LUT_1[25478] = 32'b11111111111111111111100110110100;
assign LUT_1[25479] = 32'b11111111111111111000111000110000;
assign LUT_1[25480] = 32'b11111111111111111011001101000001;
assign LUT_1[25481] = 32'b11111111111111110100011110111101;
assign LUT_1[25482] = 32'b11111111111111110110111011010010;
assign LUT_1[25483] = 32'b11111111111111110000001101001110;
assign LUT_1[25484] = 32'b00000000000000000011000110011000;
assign LUT_1[25485] = 32'b11111111111111111100011000010100;
assign LUT_1[25486] = 32'b11111111111111111110110100101001;
assign LUT_1[25487] = 32'b11111111111111111000000110100101;
assign LUT_1[25488] = 32'b11111111111111111101111010101110;
assign LUT_1[25489] = 32'b11111111111111110111001100101010;
assign LUT_1[25490] = 32'b11111111111111111001101000111111;
assign LUT_1[25491] = 32'b11111111111111110010111010111011;
assign LUT_1[25492] = 32'b00000000000000000101110100000101;
assign LUT_1[25493] = 32'b11111111111111111111000110000001;
assign LUT_1[25494] = 32'b00000000000000000001100010010110;
assign LUT_1[25495] = 32'b11111111111111111010110100010010;
assign LUT_1[25496] = 32'b11111111111111111101001000100011;
assign LUT_1[25497] = 32'b11111111111111110110011010011111;
assign LUT_1[25498] = 32'b11111111111111111000110110110100;
assign LUT_1[25499] = 32'b11111111111111110010001000110000;
assign LUT_1[25500] = 32'b00000000000000000101000001111010;
assign LUT_1[25501] = 32'b11111111111111111110010011110110;
assign LUT_1[25502] = 32'b00000000000000000000110000001011;
assign LUT_1[25503] = 32'b11111111111111111010000010000111;
assign LUT_1[25504] = 32'b11111111111111111100111010001011;
assign LUT_1[25505] = 32'b11111111111111110110001100000111;
assign LUT_1[25506] = 32'b11111111111111111000101000011100;
assign LUT_1[25507] = 32'b11111111111111110001111010011000;
assign LUT_1[25508] = 32'b00000000000000000100110011100010;
assign LUT_1[25509] = 32'b11111111111111111110000101011110;
assign LUT_1[25510] = 32'b00000000000000000000100001110011;
assign LUT_1[25511] = 32'b11111111111111111001110011101111;
assign LUT_1[25512] = 32'b11111111111111111100001000000000;
assign LUT_1[25513] = 32'b11111111111111110101011001111100;
assign LUT_1[25514] = 32'b11111111111111110111110110010001;
assign LUT_1[25515] = 32'b11111111111111110001001000001101;
assign LUT_1[25516] = 32'b00000000000000000100000001010111;
assign LUT_1[25517] = 32'b11111111111111111101010011010011;
assign LUT_1[25518] = 32'b11111111111111111111101111101000;
assign LUT_1[25519] = 32'b11111111111111111001000001100100;
assign LUT_1[25520] = 32'b11111111111111111110110101101101;
assign LUT_1[25521] = 32'b11111111111111111000000111101001;
assign LUT_1[25522] = 32'b11111111111111111010100011111110;
assign LUT_1[25523] = 32'b11111111111111110011110101111010;
assign LUT_1[25524] = 32'b00000000000000000110101111000100;
assign LUT_1[25525] = 32'b00000000000000000000000001000000;
assign LUT_1[25526] = 32'b00000000000000000010011101010101;
assign LUT_1[25527] = 32'b11111111111111111011101111010001;
assign LUT_1[25528] = 32'b11111111111111111110000011100010;
assign LUT_1[25529] = 32'b11111111111111110111010101011110;
assign LUT_1[25530] = 32'b11111111111111111001110001110011;
assign LUT_1[25531] = 32'b11111111111111110011000011101111;
assign LUT_1[25532] = 32'b00000000000000000101111100111001;
assign LUT_1[25533] = 32'b11111111111111111111001110110101;
assign LUT_1[25534] = 32'b00000000000000000001101011001010;
assign LUT_1[25535] = 32'b11111111111111111010111101000110;
assign LUT_1[25536] = 32'b11111111111111111101111100110100;
assign LUT_1[25537] = 32'b11111111111111110111001110110000;
assign LUT_1[25538] = 32'b11111111111111111001101011000101;
assign LUT_1[25539] = 32'b11111111111111110010111101000001;
assign LUT_1[25540] = 32'b00000000000000000101110110001011;
assign LUT_1[25541] = 32'b11111111111111111111001000000111;
assign LUT_1[25542] = 32'b00000000000000000001100100011100;
assign LUT_1[25543] = 32'b11111111111111111010110110011000;
assign LUT_1[25544] = 32'b11111111111111111101001010101001;
assign LUT_1[25545] = 32'b11111111111111110110011100100101;
assign LUT_1[25546] = 32'b11111111111111111000111000111010;
assign LUT_1[25547] = 32'b11111111111111110010001010110110;
assign LUT_1[25548] = 32'b00000000000000000101000100000000;
assign LUT_1[25549] = 32'b11111111111111111110010101111100;
assign LUT_1[25550] = 32'b00000000000000000000110010010001;
assign LUT_1[25551] = 32'b11111111111111111010000100001101;
assign LUT_1[25552] = 32'b11111111111111111111111000010110;
assign LUT_1[25553] = 32'b11111111111111111001001010010010;
assign LUT_1[25554] = 32'b11111111111111111011100110100111;
assign LUT_1[25555] = 32'b11111111111111110100111000100011;
assign LUT_1[25556] = 32'b00000000000000000111110001101101;
assign LUT_1[25557] = 32'b00000000000000000001000011101001;
assign LUT_1[25558] = 32'b00000000000000000011011111111110;
assign LUT_1[25559] = 32'b11111111111111111100110001111010;
assign LUT_1[25560] = 32'b11111111111111111111000110001011;
assign LUT_1[25561] = 32'b11111111111111111000011000000111;
assign LUT_1[25562] = 32'b11111111111111111010110100011100;
assign LUT_1[25563] = 32'b11111111111111110100000110011000;
assign LUT_1[25564] = 32'b00000000000000000110111111100010;
assign LUT_1[25565] = 32'b00000000000000000000010001011110;
assign LUT_1[25566] = 32'b00000000000000000010101101110011;
assign LUT_1[25567] = 32'b11111111111111111011111111101111;
assign LUT_1[25568] = 32'b11111111111111111110110111110011;
assign LUT_1[25569] = 32'b11111111111111111000001001101111;
assign LUT_1[25570] = 32'b11111111111111111010100110000100;
assign LUT_1[25571] = 32'b11111111111111110011111000000000;
assign LUT_1[25572] = 32'b00000000000000000110110001001010;
assign LUT_1[25573] = 32'b00000000000000000000000011000110;
assign LUT_1[25574] = 32'b00000000000000000010011111011011;
assign LUT_1[25575] = 32'b11111111111111111011110001010111;
assign LUT_1[25576] = 32'b11111111111111111110000101101000;
assign LUT_1[25577] = 32'b11111111111111110111010111100100;
assign LUT_1[25578] = 32'b11111111111111111001110011111001;
assign LUT_1[25579] = 32'b11111111111111110011000101110101;
assign LUT_1[25580] = 32'b00000000000000000101111110111111;
assign LUT_1[25581] = 32'b11111111111111111111010000111011;
assign LUT_1[25582] = 32'b00000000000000000001101101010000;
assign LUT_1[25583] = 32'b11111111111111111010111111001100;
assign LUT_1[25584] = 32'b00000000000000000000110011010101;
assign LUT_1[25585] = 32'b11111111111111111010000101010001;
assign LUT_1[25586] = 32'b11111111111111111100100001100110;
assign LUT_1[25587] = 32'b11111111111111110101110011100010;
assign LUT_1[25588] = 32'b00000000000000001000101100101100;
assign LUT_1[25589] = 32'b00000000000000000001111110101000;
assign LUT_1[25590] = 32'b00000000000000000100011010111101;
assign LUT_1[25591] = 32'b11111111111111111101101100111001;
assign LUT_1[25592] = 32'b00000000000000000000000001001010;
assign LUT_1[25593] = 32'b11111111111111111001010011000110;
assign LUT_1[25594] = 32'b11111111111111111011101111011011;
assign LUT_1[25595] = 32'b11111111111111110101000001010111;
assign LUT_1[25596] = 32'b00000000000000000111111010100001;
assign LUT_1[25597] = 32'b00000000000000000001001100011101;
assign LUT_1[25598] = 32'b00000000000000000011101000110010;
assign LUT_1[25599] = 32'b11111111111111111100111010101110;
assign LUT_1[25600] = 32'b00000000000000000111110011010000;
assign LUT_1[25601] = 32'b00000000000000000001000101001100;
assign LUT_1[25602] = 32'b00000000000000000011100001100001;
assign LUT_1[25603] = 32'b11111111111111111100110011011101;
assign LUT_1[25604] = 32'b00000000000000001111101100100111;
assign LUT_1[25605] = 32'b00000000000000001000111110100011;
assign LUT_1[25606] = 32'b00000000000000001011011010111000;
assign LUT_1[25607] = 32'b00000000000000000100101100110100;
assign LUT_1[25608] = 32'b00000000000000000111000001000101;
assign LUT_1[25609] = 32'b00000000000000000000010011000001;
assign LUT_1[25610] = 32'b00000000000000000010101111010110;
assign LUT_1[25611] = 32'b11111111111111111100000001010010;
assign LUT_1[25612] = 32'b00000000000000001110111010011100;
assign LUT_1[25613] = 32'b00000000000000001000001100011000;
assign LUT_1[25614] = 32'b00000000000000001010101000101101;
assign LUT_1[25615] = 32'b00000000000000000011111010101001;
assign LUT_1[25616] = 32'b00000000000000001001101110110010;
assign LUT_1[25617] = 32'b00000000000000000011000000101110;
assign LUT_1[25618] = 32'b00000000000000000101011101000011;
assign LUT_1[25619] = 32'b11111111111111111110101110111111;
assign LUT_1[25620] = 32'b00000000000000010001101000001001;
assign LUT_1[25621] = 32'b00000000000000001010111010000101;
assign LUT_1[25622] = 32'b00000000000000001101010110011010;
assign LUT_1[25623] = 32'b00000000000000000110101000010110;
assign LUT_1[25624] = 32'b00000000000000001000111100100111;
assign LUT_1[25625] = 32'b00000000000000000010001110100011;
assign LUT_1[25626] = 32'b00000000000000000100101010111000;
assign LUT_1[25627] = 32'b11111111111111111101111100110100;
assign LUT_1[25628] = 32'b00000000000000010000110101111110;
assign LUT_1[25629] = 32'b00000000000000001010000111111010;
assign LUT_1[25630] = 32'b00000000000000001100100100001111;
assign LUT_1[25631] = 32'b00000000000000000101110110001011;
assign LUT_1[25632] = 32'b00000000000000001000101110001111;
assign LUT_1[25633] = 32'b00000000000000000010000000001011;
assign LUT_1[25634] = 32'b00000000000000000100011100100000;
assign LUT_1[25635] = 32'b11111111111111111101101110011100;
assign LUT_1[25636] = 32'b00000000000000010000100111100110;
assign LUT_1[25637] = 32'b00000000000000001001111001100010;
assign LUT_1[25638] = 32'b00000000000000001100010101110111;
assign LUT_1[25639] = 32'b00000000000000000101100111110011;
assign LUT_1[25640] = 32'b00000000000000000111111100000100;
assign LUT_1[25641] = 32'b00000000000000000001001110000000;
assign LUT_1[25642] = 32'b00000000000000000011101010010101;
assign LUT_1[25643] = 32'b11111111111111111100111100010001;
assign LUT_1[25644] = 32'b00000000000000001111110101011011;
assign LUT_1[25645] = 32'b00000000000000001001000111010111;
assign LUT_1[25646] = 32'b00000000000000001011100011101100;
assign LUT_1[25647] = 32'b00000000000000000100110101101000;
assign LUT_1[25648] = 32'b00000000000000001010101001110001;
assign LUT_1[25649] = 32'b00000000000000000011111011101101;
assign LUT_1[25650] = 32'b00000000000000000110011000000010;
assign LUT_1[25651] = 32'b11111111111111111111101001111110;
assign LUT_1[25652] = 32'b00000000000000010010100011001000;
assign LUT_1[25653] = 32'b00000000000000001011110101000100;
assign LUT_1[25654] = 32'b00000000000000001110010001011001;
assign LUT_1[25655] = 32'b00000000000000000111100011010101;
assign LUT_1[25656] = 32'b00000000000000001001110111100110;
assign LUT_1[25657] = 32'b00000000000000000011001001100010;
assign LUT_1[25658] = 32'b00000000000000000101100101110111;
assign LUT_1[25659] = 32'b11111111111111111110110111110011;
assign LUT_1[25660] = 32'b00000000000000010001110000111101;
assign LUT_1[25661] = 32'b00000000000000001011000010111001;
assign LUT_1[25662] = 32'b00000000000000001101011111001110;
assign LUT_1[25663] = 32'b00000000000000000110110001001010;
assign LUT_1[25664] = 32'b00000000000000001001110000111000;
assign LUT_1[25665] = 32'b00000000000000000011000010110100;
assign LUT_1[25666] = 32'b00000000000000000101011111001001;
assign LUT_1[25667] = 32'b11111111111111111110110001000101;
assign LUT_1[25668] = 32'b00000000000000010001101010001111;
assign LUT_1[25669] = 32'b00000000000000001010111100001011;
assign LUT_1[25670] = 32'b00000000000000001101011000100000;
assign LUT_1[25671] = 32'b00000000000000000110101010011100;
assign LUT_1[25672] = 32'b00000000000000001000111110101101;
assign LUT_1[25673] = 32'b00000000000000000010010000101001;
assign LUT_1[25674] = 32'b00000000000000000100101100111110;
assign LUT_1[25675] = 32'b11111111111111111101111110111010;
assign LUT_1[25676] = 32'b00000000000000010000111000000100;
assign LUT_1[25677] = 32'b00000000000000001010001010000000;
assign LUT_1[25678] = 32'b00000000000000001100100110010101;
assign LUT_1[25679] = 32'b00000000000000000101111000010001;
assign LUT_1[25680] = 32'b00000000000000001011101100011010;
assign LUT_1[25681] = 32'b00000000000000000100111110010110;
assign LUT_1[25682] = 32'b00000000000000000111011010101011;
assign LUT_1[25683] = 32'b00000000000000000000101100100111;
assign LUT_1[25684] = 32'b00000000000000010011100101110001;
assign LUT_1[25685] = 32'b00000000000000001100110111101101;
assign LUT_1[25686] = 32'b00000000000000001111010100000010;
assign LUT_1[25687] = 32'b00000000000000001000100101111110;
assign LUT_1[25688] = 32'b00000000000000001010111010001111;
assign LUT_1[25689] = 32'b00000000000000000100001100001011;
assign LUT_1[25690] = 32'b00000000000000000110101000100000;
assign LUT_1[25691] = 32'b11111111111111111111111010011100;
assign LUT_1[25692] = 32'b00000000000000010010110011100110;
assign LUT_1[25693] = 32'b00000000000000001100000101100010;
assign LUT_1[25694] = 32'b00000000000000001110100001110111;
assign LUT_1[25695] = 32'b00000000000000000111110011110011;
assign LUT_1[25696] = 32'b00000000000000001010101011110111;
assign LUT_1[25697] = 32'b00000000000000000011111101110011;
assign LUT_1[25698] = 32'b00000000000000000110011010001000;
assign LUT_1[25699] = 32'b11111111111111111111101100000100;
assign LUT_1[25700] = 32'b00000000000000010010100101001110;
assign LUT_1[25701] = 32'b00000000000000001011110111001010;
assign LUT_1[25702] = 32'b00000000000000001110010011011111;
assign LUT_1[25703] = 32'b00000000000000000111100101011011;
assign LUT_1[25704] = 32'b00000000000000001001111001101100;
assign LUT_1[25705] = 32'b00000000000000000011001011101000;
assign LUT_1[25706] = 32'b00000000000000000101100111111101;
assign LUT_1[25707] = 32'b11111111111111111110111001111001;
assign LUT_1[25708] = 32'b00000000000000010001110011000011;
assign LUT_1[25709] = 32'b00000000000000001011000100111111;
assign LUT_1[25710] = 32'b00000000000000001101100001010100;
assign LUT_1[25711] = 32'b00000000000000000110110011010000;
assign LUT_1[25712] = 32'b00000000000000001100100111011001;
assign LUT_1[25713] = 32'b00000000000000000101111001010101;
assign LUT_1[25714] = 32'b00000000000000001000010101101010;
assign LUT_1[25715] = 32'b00000000000000000001100111100110;
assign LUT_1[25716] = 32'b00000000000000010100100000110000;
assign LUT_1[25717] = 32'b00000000000000001101110010101100;
assign LUT_1[25718] = 32'b00000000000000010000001111000001;
assign LUT_1[25719] = 32'b00000000000000001001100000111101;
assign LUT_1[25720] = 32'b00000000000000001011110101001110;
assign LUT_1[25721] = 32'b00000000000000000101000111001010;
assign LUT_1[25722] = 32'b00000000000000000111100011011111;
assign LUT_1[25723] = 32'b00000000000000000000110101011011;
assign LUT_1[25724] = 32'b00000000000000010011101110100101;
assign LUT_1[25725] = 32'b00000000000000001101000000100001;
assign LUT_1[25726] = 32'b00000000000000001111011100110110;
assign LUT_1[25727] = 32'b00000000000000001000101110110010;
assign LUT_1[25728] = 32'b00000000000000001010110011010011;
assign LUT_1[25729] = 32'b00000000000000000100000101001111;
assign LUT_1[25730] = 32'b00000000000000000110100001100100;
assign LUT_1[25731] = 32'b11111111111111111111110011100000;
assign LUT_1[25732] = 32'b00000000000000010010101100101010;
assign LUT_1[25733] = 32'b00000000000000001011111110100110;
assign LUT_1[25734] = 32'b00000000000000001110011010111011;
assign LUT_1[25735] = 32'b00000000000000000111101100110111;
assign LUT_1[25736] = 32'b00000000000000001010000001001000;
assign LUT_1[25737] = 32'b00000000000000000011010011000100;
assign LUT_1[25738] = 32'b00000000000000000101101111011001;
assign LUT_1[25739] = 32'b11111111111111111111000001010101;
assign LUT_1[25740] = 32'b00000000000000010001111010011111;
assign LUT_1[25741] = 32'b00000000000000001011001100011011;
assign LUT_1[25742] = 32'b00000000000000001101101000110000;
assign LUT_1[25743] = 32'b00000000000000000110111010101100;
assign LUT_1[25744] = 32'b00000000000000001100101110110101;
assign LUT_1[25745] = 32'b00000000000000000110000000110001;
assign LUT_1[25746] = 32'b00000000000000001000011101000110;
assign LUT_1[25747] = 32'b00000000000000000001101111000010;
assign LUT_1[25748] = 32'b00000000000000010100101000001100;
assign LUT_1[25749] = 32'b00000000000000001101111010001000;
assign LUT_1[25750] = 32'b00000000000000010000010110011101;
assign LUT_1[25751] = 32'b00000000000000001001101000011001;
assign LUT_1[25752] = 32'b00000000000000001011111100101010;
assign LUT_1[25753] = 32'b00000000000000000101001110100110;
assign LUT_1[25754] = 32'b00000000000000000111101010111011;
assign LUT_1[25755] = 32'b00000000000000000000111100110111;
assign LUT_1[25756] = 32'b00000000000000010011110110000001;
assign LUT_1[25757] = 32'b00000000000000001101000111111101;
assign LUT_1[25758] = 32'b00000000000000001111100100010010;
assign LUT_1[25759] = 32'b00000000000000001000110110001110;
assign LUT_1[25760] = 32'b00000000000000001011101110010010;
assign LUT_1[25761] = 32'b00000000000000000101000000001110;
assign LUT_1[25762] = 32'b00000000000000000111011100100011;
assign LUT_1[25763] = 32'b00000000000000000000101110011111;
assign LUT_1[25764] = 32'b00000000000000010011100111101001;
assign LUT_1[25765] = 32'b00000000000000001100111001100101;
assign LUT_1[25766] = 32'b00000000000000001111010101111010;
assign LUT_1[25767] = 32'b00000000000000001000100111110110;
assign LUT_1[25768] = 32'b00000000000000001010111100000111;
assign LUT_1[25769] = 32'b00000000000000000100001110000011;
assign LUT_1[25770] = 32'b00000000000000000110101010011000;
assign LUT_1[25771] = 32'b11111111111111111111111100010100;
assign LUT_1[25772] = 32'b00000000000000010010110101011110;
assign LUT_1[25773] = 32'b00000000000000001100000111011010;
assign LUT_1[25774] = 32'b00000000000000001110100011101111;
assign LUT_1[25775] = 32'b00000000000000000111110101101011;
assign LUT_1[25776] = 32'b00000000000000001101101001110100;
assign LUT_1[25777] = 32'b00000000000000000110111011110000;
assign LUT_1[25778] = 32'b00000000000000001001011000000101;
assign LUT_1[25779] = 32'b00000000000000000010101010000001;
assign LUT_1[25780] = 32'b00000000000000010101100011001011;
assign LUT_1[25781] = 32'b00000000000000001110110101000111;
assign LUT_1[25782] = 32'b00000000000000010001010001011100;
assign LUT_1[25783] = 32'b00000000000000001010100011011000;
assign LUT_1[25784] = 32'b00000000000000001100110111101001;
assign LUT_1[25785] = 32'b00000000000000000110001001100101;
assign LUT_1[25786] = 32'b00000000000000001000100101111010;
assign LUT_1[25787] = 32'b00000000000000000001110111110110;
assign LUT_1[25788] = 32'b00000000000000010100110001000000;
assign LUT_1[25789] = 32'b00000000000000001110000010111100;
assign LUT_1[25790] = 32'b00000000000000010000011111010001;
assign LUT_1[25791] = 32'b00000000000000001001110001001101;
assign LUT_1[25792] = 32'b00000000000000001100110000111011;
assign LUT_1[25793] = 32'b00000000000000000110000010110111;
assign LUT_1[25794] = 32'b00000000000000001000011111001100;
assign LUT_1[25795] = 32'b00000000000000000001110001001000;
assign LUT_1[25796] = 32'b00000000000000010100101010010010;
assign LUT_1[25797] = 32'b00000000000000001101111100001110;
assign LUT_1[25798] = 32'b00000000000000010000011000100011;
assign LUT_1[25799] = 32'b00000000000000001001101010011111;
assign LUT_1[25800] = 32'b00000000000000001011111110110000;
assign LUT_1[25801] = 32'b00000000000000000101010000101100;
assign LUT_1[25802] = 32'b00000000000000000111101101000001;
assign LUT_1[25803] = 32'b00000000000000000000111110111101;
assign LUT_1[25804] = 32'b00000000000000010011111000000111;
assign LUT_1[25805] = 32'b00000000000000001101001010000011;
assign LUT_1[25806] = 32'b00000000000000001111100110011000;
assign LUT_1[25807] = 32'b00000000000000001000111000010100;
assign LUT_1[25808] = 32'b00000000000000001110101100011101;
assign LUT_1[25809] = 32'b00000000000000000111111110011001;
assign LUT_1[25810] = 32'b00000000000000001010011010101110;
assign LUT_1[25811] = 32'b00000000000000000011101100101010;
assign LUT_1[25812] = 32'b00000000000000010110100101110100;
assign LUT_1[25813] = 32'b00000000000000001111110111110000;
assign LUT_1[25814] = 32'b00000000000000010010010100000101;
assign LUT_1[25815] = 32'b00000000000000001011100110000001;
assign LUT_1[25816] = 32'b00000000000000001101111010010010;
assign LUT_1[25817] = 32'b00000000000000000111001100001110;
assign LUT_1[25818] = 32'b00000000000000001001101000100011;
assign LUT_1[25819] = 32'b00000000000000000010111010011111;
assign LUT_1[25820] = 32'b00000000000000010101110011101001;
assign LUT_1[25821] = 32'b00000000000000001111000101100101;
assign LUT_1[25822] = 32'b00000000000000010001100001111010;
assign LUT_1[25823] = 32'b00000000000000001010110011110110;
assign LUT_1[25824] = 32'b00000000000000001101101011111010;
assign LUT_1[25825] = 32'b00000000000000000110111101110110;
assign LUT_1[25826] = 32'b00000000000000001001011010001011;
assign LUT_1[25827] = 32'b00000000000000000010101100000111;
assign LUT_1[25828] = 32'b00000000000000010101100101010001;
assign LUT_1[25829] = 32'b00000000000000001110110111001101;
assign LUT_1[25830] = 32'b00000000000000010001010011100010;
assign LUT_1[25831] = 32'b00000000000000001010100101011110;
assign LUT_1[25832] = 32'b00000000000000001100111001101111;
assign LUT_1[25833] = 32'b00000000000000000110001011101011;
assign LUT_1[25834] = 32'b00000000000000001000101000000000;
assign LUT_1[25835] = 32'b00000000000000000001111001111100;
assign LUT_1[25836] = 32'b00000000000000010100110011000110;
assign LUT_1[25837] = 32'b00000000000000001110000101000010;
assign LUT_1[25838] = 32'b00000000000000010000100001010111;
assign LUT_1[25839] = 32'b00000000000000001001110011010011;
assign LUT_1[25840] = 32'b00000000000000001111100111011100;
assign LUT_1[25841] = 32'b00000000000000001000111001011000;
assign LUT_1[25842] = 32'b00000000000000001011010101101101;
assign LUT_1[25843] = 32'b00000000000000000100100111101001;
assign LUT_1[25844] = 32'b00000000000000010111100000110011;
assign LUT_1[25845] = 32'b00000000000000010000110010101111;
assign LUT_1[25846] = 32'b00000000000000010011001111000100;
assign LUT_1[25847] = 32'b00000000000000001100100001000000;
assign LUT_1[25848] = 32'b00000000000000001110110101010001;
assign LUT_1[25849] = 32'b00000000000000001000000111001101;
assign LUT_1[25850] = 32'b00000000000000001010100011100010;
assign LUT_1[25851] = 32'b00000000000000000011110101011110;
assign LUT_1[25852] = 32'b00000000000000010110101110101000;
assign LUT_1[25853] = 32'b00000000000000010000000000100100;
assign LUT_1[25854] = 32'b00000000000000010010011100111001;
assign LUT_1[25855] = 32'b00000000000000001011101110110101;
assign LUT_1[25856] = 32'b00000000000000000101100111011100;
assign LUT_1[25857] = 32'b11111111111111111110111001011000;
assign LUT_1[25858] = 32'b00000000000000000001010101101101;
assign LUT_1[25859] = 32'b11111111111111111010100111101001;
assign LUT_1[25860] = 32'b00000000000000001101100000110011;
assign LUT_1[25861] = 32'b00000000000000000110110010101111;
assign LUT_1[25862] = 32'b00000000000000001001001111000100;
assign LUT_1[25863] = 32'b00000000000000000010100001000000;
assign LUT_1[25864] = 32'b00000000000000000100110101010001;
assign LUT_1[25865] = 32'b11111111111111111110000111001101;
assign LUT_1[25866] = 32'b00000000000000000000100011100010;
assign LUT_1[25867] = 32'b11111111111111111001110101011110;
assign LUT_1[25868] = 32'b00000000000000001100101110101000;
assign LUT_1[25869] = 32'b00000000000000000110000000100100;
assign LUT_1[25870] = 32'b00000000000000001000011100111001;
assign LUT_1[25871] = 32'b00000000000000000001101110110101;
assign LUT_1[25872] = 32'b00000000000000000111100010111110;
assign LUT_1[25873] = 32'b00000000000000000000110100111010;
assign LUT_1[25874] = 32'b00000000000000000011010001001111;
assign LUT_1[25875] = 32'b11111111111111111100100011001011;
assign LUT_1[25876] = 32'b00000000000000001111011100010101;
assign LUT_1[25877] = 32'b00000000000000001000101110010001;
assign LUT_1[25878] = 32'b00000000000000001011001010100110;
assign LUT_1[25879] = 32'b00000000000000000100011100100010;
assign LUT_1[25880] = 32'b00000000000000000110110000110011;
assign LUT_1[25881] = 32'b00000000000000000000000010101111;
assign LUT_1[25882] = 32'b00000000000000000010011111000100;
assign LUT_1[25883] = 32'b11111111111111111011110001000000;
assign LUT_1[25884] = 32'b00000000000000001110101010001010;
assign LUT_1[25885] = 32'b00000000000000000111111100000110;
assign LUT_1[25886] = 32'b00000000000000001010011000011011;
assign LUT_1[25887] = 32'b00000000000000000011101010010111;
assign LUT_1[25888] = 32'b00000000000000000110100010011011;
assign LUT_1[25889] = 32'b11111111111111111111110100010111;
assign LUT_1[25890] = 32'b00000000000000000010010000101100;
assign LUT_1[25891] = 32'b11111111111111111011100010101000;
assign LUT_1[25892] = 32'b00000000000000001110011011110010;
assign LUT_1[25893] = 32'b00000000000000000111101101101110;
assign LUT_1[25894] = 32'b00000000000000001010001010000011;
assign LUT_1[25895] = 32'b00000000000000000011011011111111;
assign LUT_1[25896] = 32'b00000000000000000101110000010000;
assign LUT_1[25897] = 32'b11111111111111111111000010001100;
assign LUT_1[25898] = 32'b00000000000000000001011110100001;
assign LUT_1[25899] = 32'b11111111111111111010110000011101;
assign LUT_1[25900] = 32'b00000000000000001101101001100111;
assign LUT_1[25901] = 32'b00000000000000000110111011100011;
assign LUT_1[25902] = 32'b00000000000000001001010111111000;
assign LUT_1[25903] = 32'b00000000000000000010101001110100;
assign LUT_1[25904] = 32'b00000000000000001000011101111101;
assign LUT_1[25905] = 32'b00000000000000000001101111111001;
assign LUT_1[25906] = 32'b00000000000000000100001100001110;
assign LUT_1[25907] = 32'b11111111111111111101011110001010;
assign LUT_1[25908] = 32'b00000000000000010000010111010100;
assign LUT_1[25909] = 32'b00000000000000001001101001010000;
assign LUT_1[25910] = 32'b00000000000000001100000101100101;
assign LUT_1[25911] = 32'b00000000000000000101010111100001;
assign LUT_1[25912] = 32'b00000000000000000111101011110010;
assign LUT_1[25913] = 32'b00000000000000000000111101101110;
assign LUT_1[25914] = 32'b00000000000000000011011010000011;
assign LUT_1[25915] = 32'b11111111111111111100101011111111;
assign LUT_1[25916] = 32'b00000000000000001111100101001001;
assign LUT_1[25917] = 32'b00000000000000001000110111000101;
assign LUT_1[25918] = 32'b00000000000000001011010011011010;
assign LUT_1[25919] = 32'b00000000000000000100100101010110;
assign LUT_1[25920] = 32'b00000000000000000111100101000100;
assign LUT_1[25921] = 32'b00000000000000000000110111000000;
assign LUT_1[25922] = 32'b00000000000000000011010011010101;
assign LUT_1[25923] = 32'b11111111111111111100100101010001;
assign LUT_1[25924] = 32'b00000000000000001111011110011011;
assign LUT_1[25925] = 32'b00000000000000001000110000010111;
assign LUT_1[25926] = 32'b00000000000000001011001100101100;
assign LUT_1[25927] = 32'b00000000000000000100011110101000;
assign LUT_1[25928] = 32'b00000000000000000110110010111001;
assign LUT_1[25929] = 32'b00000000000000000000000100110101;
assign LUT_1[25930] = 32'b00000000000000000010100001001010;
assign LUT_1[25931] = 32'b11111111111111111011110011000110;
assign LUT_1[25932] = 32'b00000000000000001110101100010000;
assign LUT_1[25933] = 32'b00000000000000000111111110001100;
assign LUT_1[25934] = 32'b00000000000000001010011010100001;
assign LUT_1[25935] = 32'b00000000000000000011101100011101;
assign LUT_1[25936] = 32'b00000000000000001001100000100110;
assign LUT_1[25937] = 32'b00000000000000000010110010100010;
assign LUT_1[25938] = 32'b00000000000000000101001110110111;
assign LUT_1[25939] = 32'b11111111111111111110100000110011;
assign LUT_1[25940] = 32'b00000000000000010001011001111101;
assign LUT_1[25941] = 32'b00000000000000001010101011111001;
assign LUT_1[25942] = 32'b00000000000000001101001000001110;
assign LUT_1[25943] = 32'b00000000000000000110011010001010;
assign LUT_1[25944] = 32'b00000000000000001000101110011011;
assign LUT_1[25945] = 32'b00000000000000000010000000010111;
assign LUT_1[25946] = 32'b00000000000000000100011100101100;
assign LUT_1[25947] = 32'b11111111111111111101101110101000;
assign LUT_1[25948] = 32'b00000000000000010000100111110010;
assign LUT_1[25949] = 32'b00000000000000001001111001101110;
assign LUT_1[25950] = 32'b00000000000000001100010110000011;
assign LUT_1[25951] = 32'b00000000000000000101100111111111;
assign LUT_1[25952] = 32'b00000000000000001000100000000011;
assign LUT_1[25953] = 32'b00000000000000000001110001111111;
assign LUT_1[25954] = 32'b00000000000000000100001110010100;
assign LUT_1[25955] = 32'b11111111111111111101100000010000;
assign LUT_1[25956] = 32'b00000000000000010000011001011010;
assign LUT_1[25957] = 32'b00000000000000001001101011010110;
assign LUT_1[25958] = 32'b00000000000000001100000111101011;
assign LUT_1[25959] = 32'b00000000000000000101011001100111;
assign LUT_1[25960] = 32'b00000000000000000111101101111000;
assign LUT_1[25961] = 32'b00000000000000000000111111110100;
assign LUT_1[25962] = 32'b00000000000000000011011100001001;
assign LUT_1[25963] = 32'b11111111111111111100101110000101;
assign LUT_1[25964] = 32'b00000000000000001111100111001111;
assign LUT_1[25965] = 32'b00000000000000001000111001001011;
assign LUT_1[25966] = 32'b00000000000000001011010101100000;
assign LUT_1[25967] = 32'b00000000000000000100100111011100;
assign LUT_1[25968] = 32'b00000000000000001010011011100101;
assign LUT_1[25969] = 32'b00000000000000000011101101100001;
assign LUT_1[25970] = 32'b00000000000000000110001001110110;
assign LUT_1[25971] = 32'b11111111111111111111011011110010;
assign LUT_1[25972] = 32'b00000000000000010010010100111100;
assign LUT_1[25973] = 32'b00000000000000001011100110111000;
assign LUT_1[25974] = 32'b00000000000000001110000011001101;
assign LUT_1[25975] = 32'b00000000000000000111010101001001;
assign LUT_1[25976] = 32'b00000000000000001001101001011010;
assign LUT_1[25977] = 32'b00000000000000000010111011010110;
assign LUT_1[25978] = 32'b00000000000000000101010111101011;
assign LUT_1[25979] = 32'b11111111111111111110101001100111;
assign LUT_1[25980] = 32'b00000000000000010001100010110001;
assign LUT_1[25981] = 32'b00000000000000001010110100101101;
assign LUT_1[25982] = 32'b00000000000000001101010001000010;
assign LUT_1[25983] = 32'b00000000000000000110100010111110;
assign LUT_1[25984] = 32'b00000000000000001000100111011111;
assign LUT_1[25985] = 32'b00000000000000000001111001011011;
assign LUT_1[25986] = 32'b00000000000000000100010101110000;
assign LUT_1[25987] = 32'b11111111111111111101100111101100;
assign LUT_1[25988] = 32'b00000000000000010000100000110110;
assign LUT_1[25989] = 32'b00000000000000001001110010110010;
assign LUT_1[25990] = 32'b00000000000000001100001111000111;
assign LUT_1[25991] = 32'b00000000000000000101100001000011;
assign LUT_1[25992] = 32'b00000000000000000111110101010100;
assign LUT_1[25993] = 32'b00000000000000000001000111010000;
assign LUT_1[25994] = 32'b00000000000000000011100011100101;
assign LUT_1[25995] = 32'b11111111111111111100110101100001;
assign LUT_1[25996] = 32'b00000000000000001111101110101011;
assign LUT_1[25997] = 32'b00000000000000001001000000100111;
assign LUT_1[25998] = 32'b00000000000000001011011100111100;
assign LUT_1[25999] = 32'b00000000000000000100101110111000;
assign LUT_1[26000] = 32'b00000000000000001010100011000001;
assign LUT_1[26001] = 32'b00000000000000000011110100111101;
assign LUT_1[26002] = 32'b00000000000000000110010001010010;
assign LUT_1[26003] = 32'b11111111111111111111100011001110;
assign LUT_1[26004] = 32'b00000000000000010010011100011000;
assign LUT_1[26005] = 32'b00000000000000001011101110010100;
assign LUT_1[26006] = 32'b00000000000000001110001010101001;
assign LUT_1[26007] = 32'b00000000000000000111011100100101;
assign LUT_1[26008] = 32'b00000000000000001001110000110110;
assign LUT_1[26009] = 32'b00000000000000000011000010110010;
assign LUT_1[26010] = 32'b00000000000000000101011111000111;
assign LUT_1[26011] = 32'b11111111111111111110110001000011;
assign LUT_1[26012] = 32'b00000000000000010001101010001101;
assign LUT_1[26013] = 32'b00000000000000001010111100001001;
assign LUT_1[26014] = 32'b00000000000000001101011000011110;
assign LUT_1[26015] = 32'b00000000000000000110101010011010;
assign LUT_1[26016] = 32'b00000000000000001001100010011110;
assign LUT_1[26017] = 32'b00000000000000000010110100011010;
assign LUT_1[26018] = 32'b00000000000000000101010000101111;
assign LUT_1[26019] = 32'b11111111111111111110100010101011;
assign LUT_1[26020] = 32'b00000000000000010001011011110101;
assign LUT_1[26021] = 32'b00000000000000001010101101110001;
assign LUT_1[26022] = 32'b00000000000000001101001010000110;
assign LUT_1[26023] = 32'b00000000000000000110011100000010;
assign LUT_1[26024] = 32'b00000000000000001000110000010011;
assign LUT_1[26025] = 32'b00000000000000000010000010001111;
assign LUT_1[26026] = 32'b00000000000000000100011110100100;
assign LUT_1[26027] = 32'b11111111111111111101110000100000;
assign LUT_1[26028] = 32'b00000000000000010000101001101010;
assign LUT_1[26029] = 32'b00000000000000001001111011100110;
assign LUT_1[26030] = 32'b00000000000000001100010111111011;
assign LUT_1[26031] = 32'b00000000000000000101101001110111;
assign LUT_1[26032] = 32'b00000000000000001011011110000000;
assign LUT_1[26033] = 32'b00000000000000000100101111111100;
assign LUT_1[26034] = 32'b00000000000000000111001100010001;
assign LUT_1[26035] = 32'b00000000000000000000011110001101;
assign LUT_1[26036] = 32'b00000000000000010011010111010111;
assign LUT_1[26037] = 32'b00000000000000001100101001010011;
assign LUT_1[26038] = 32'b00000000000000001111000101101000;
assign LUT_1[26039] = 32'b00000000000000001000010111100100;
assign LUT_1[26040] = 32'b00000000000000001010101011110101;
assign LUT_1[26041] = 32'b00000000000000000011111101110001;
assign LUT_1[26042] = 32'b00000000000000000110011010000110;
assign LUT_1[26043] = 32'b11111111111111111111101100000010;
assign LUT_1[26044] = 32'b00000000000000010010100101001100;
assign LUT_1[26045] = 32'b00000000000000001011110111001000;
assign LUT_1[26046] = 32'b00000000000000001110010011011101;
assign LUT_1[26047] = 32'b00000000000000000111100101011001;
assign LUT_1[26048] = 32'b00000000000000001010100101000111;
assign LUT_1[26049] = 32'b00000000000000000011110111000011;
assign LUT_1[26050] = 32'b00000000000000000110010011011000;
assign LUT_1[26051] = 32'b11111111111111111111100101010100;
assign LUT_1[26052] = 32'b00000000000000010010011110011110;
assign LUT_1[26053] = 32'b00000000000000001011110000011010;
assign LUT_1[26054] = 32'b00000000000000001110001100101111;
assign LUT_1[26055] = 32'b00000000000000000111011110101011;
assign LUT_1[26056] = 32'b00000000000000001001110010111100;
assign LUT_1[26057] = 32'b00000000000000000011000100111000;
assign LUT_1[26058] = 32'b00000000000000000101100001001101;
assign LUT_1[26059] = 32'b11111111111111111110110011001001;
assign LUT_1[26060] = 32'b00000000000000010001101100010011;
assign LUT_1[26061] = 32'b00000000000000001010111110001111;
assign LUT_1[26062] = 32'b00000000000000001101011010100100;
assign LUT_1[26063] = 32'b00000000000000000110101100100000;
assign LUT_1[26064] = 32'b00000000000000001100100000101001;
assign LUT_1[26065] = 32'b00000000000000000101110010100101;
assign LUT_1[26066] = 32'b00000000000000001000001110111010;
assign LUT_1[26067] = 32'b00000000000000000001100000110110;
assign LUT_1[26068] = 32'b00000000000000010100011010000000;
assign LUT_1[26069] = 32'b00000000000000001101101011111100;
assign LUT_1[26070] = 32'b00000000000000010000001000010001;
assign LUT_1[26071] = 32'b00000000000000001001011010001101;
assign LUT_1[26072] = 32'b00000000000000001011101110011110;
assign LUT_1[26073] = 32'b00000000000000000101000000011010;
assign LUT_1[26074] = 32'b00000000000000000111011100101111;
assign LUT_1[26075] = 32'b00000000000000000000101110101011;
assign LUT_1[26076] = 32'b00000000000000010011100111110101;
assign LUT_1[26077] = 32'b00000000000000001100111001110001;
assign LUT_1[26078] = 32'b00000000000000001111010110000110;
assign LUT_1[26079] = 32'b00000000000000001000101000000010;
assign LUT_1[26080] = 32'b00000000000000001011100000000110;
assign LUT_1[26081] = 32'b00000000000000000100110010000010;
assign LUT_1[26082] = 32'b00000000000000000111001110010111;
assign LUT_1[26083] = 32'b00000000000000000000100000010011;
assign LUT_1[26084] = 32'b00000000000000010011011001011101;
assign LUT_1[26085] = 32'b00000000000000001100101011011001;
assign LUT_1[26086] = 32'b00000000000000001111000111101110;
assign LUT_1[26087] = 32'b00000000000000001000011001101010;
assign LUT_1[26088] = 32'b00000000000000001010101101111011;
assign LUT_1[26089] = 32'b00000000000000000011111111110111;
assign LUT_1[26090] = 32'b00000000000000000110011100001100;
assign LUT_1[26091] = 32'b11111111111111111111101110001000;
assign LUT_1[26092] = 32'b00000000000000010010100111010010;
assign LUT_1[26093] = 32'b00000000000000001011111001001110;
assign LUT_1[26094] = 32'b00000000000000001110010101100011;
assign LUT_1[26095] = 32'b00000000000000000111100111011111;
assign LUT_1[26096] = 32'b00000000000000001101011011101000;
assign LUT_1[26097] = 32'b00000000000000000110101101100100;
assign LUT_1[26098] = 32'b00000000000000001001001001111001;
assign LUT_1[26099] = 32'b00000000000000000010011011110101;
assign LUT_1[26100] = 32'b00000000000000010101010100111111;
assign LUT_1[26101] = 32'b00000000000000001110100110111011;
assign LUT_1[26102] = 32'b00000000000000010001000011010000;
assign LUT_1[26103] = 32'b00000000000000001010010101001100;
assign LUT_1[26104] = 32'b00000000000000001100101001011101;
assign LUT_1[26105] = 32'b00000000000000000101111011011001;
assign LUT_1[26106] = 32'b00000000000000001000010111101110;
assign LUT_1[26107] = 32'b00000000000000000001101001101010;
assign LUT_1[26108] = 32'b00000000000000010100100010110100;
assign LUT_1[26109] = 32'b00000000000000001101110100110000;
assign LUT_1[26110] = 32'b00000000000000010000010001000101;
assign LUT_1[26111] = 32'b00000000000000001001100011000001;
assign LUT_1[26112] = 32'b00000000000000000001100001101101;
assign LUT_1[26113] = 32'b11111111111111111010110011101001;
assign LUT_1[26114] = 32'b11111111111111111101001111111110;
assign LUT_1[26115] = 32'b11111111111111110110100001111010;
assign LUT_1[26116] = 32'b00000000000000001001011011000100;
assign LUT_1[26117] = 32'b00000000000000000010101101000000;
assign LUT_1[26118] = 32'b00000000000000000101001001010101;
assign LUT_1[26119] = 32'b11111111111111111110011011010001;
assign LUT_1[26120] = 32'b00000000000000000000101111100010;
assign LUT_1[26121] = 32'b11111111111111111010000001011110;
assign LUT_1[26122] = 32'b11111111111111111100011101110011;
assign LUT_1[26123] = 32'b11111111111111110101101111101111;
assign LUT_1[26124] = 32'b00000000000000001000101000111001;
assign LUT_1[26125] = 32'b00000000000000000001111010110101;
assign LUT_1[26126] = 32'b00000000000000000100010111001010;
assign LUT_1[26127] = 32'b11111111111111111101101001000110;
assign LUT_1[26128] = 32'b00000000000000000011011101001111;
assign LUT_1[26129] = 32'b11111111111111111100101111001011;
assign LUT_1[26130] = 32'b11111111111111111111001011100000;
assign LUT_1[26131] = 32'b11111111111111111000011101011100;
assign LUT_1[26132] = 32'b00000000000000001011010110100110;
assign LUT_1[26133] = 32'b00000000000000000100101000100010;
assign LUT_1[26134] = 32'b00000000000000000111000100110111;
assign LUT_1[26135] = 32'b00000000000000000000010110110011;
assign LUT_1[26136] = 32'b00000000000000000010101011000100;
assign LUT_1[26137] = 32'b11111111111111111011111101000000;
assign LUT_1[26138] = 32'b11111111111111111110011001010101;
assign LUT_1[26139] = 32'b11111111111111110111101011010001;
assign LUT_1[26140] = 32'b00000000000000001010100100011011;
assign LUT_1[26141] = 32'b00000000000000000011110110010111;
assign LUT_1[26142] = 32'b00000000000000000110010010101100;
assign LUT_1[26143] = 32'b11111111111111111111100100101000;
assign LUT_1[26144] = 32'b00000000000000000010011100101100;
assign LUT_1[26145] = 32'b11111111111111111011101110101000;
assign LUT_1[26146] = 32'b11111111111111111110001010111101;
assign LUT_1[26147] = 32'b11111111111111110111011100111001;
assign LUT_1[26148] = 32'b00000000000000001010010110000011;
assign LUT_1[26149] = 32'b00000000000000000011100111111111;
assign LUT_1[26150] = 32'b00000000000000000110000100010100;
assign LUT_1[26151] = 32'b11111111111111111111010110010000;
assign LUT_1[26152] = 32'b00000000000000000001101010100001;
assign LUT_1[26153] = 32'b11111111111111111010111100011101;
assign LUT_1[26154] = 32'b11111111111111111101011000110010;
assign LUT_1[26155] = 32'b11111111111111110110101010101110;
assign LUT_1[26156] = 32'b00000000000000001001100011111000;
assign LUT_1[26157] = 32'b00000000000000000010110101110100;
assign LUT_1[26158] = 32'b00000000000000000101010010001001;
assign LUT_1[26159] = 32'b11111111111111111110100100000101;
assign LUT_1[26160] = 32'b00000000000000000100011000001110;
assign LUT_1[26161] = 32'b11111111111111111101101010001010;
assign LUT_1[26162] = 32'b00000000000000000000000110011111;
assign LUT_1[26163] = 32'b11111111111111111001011000011011;
assign LUT_1[26164] = 32'b00000000000000001100010001100101;
assign LUT_1[26165] = 32'b00000000000000000101100011100001;
assign LUT_1[26166] = 32'b00000000000000000111111111110110;
assign LUT_1[26167] = 32'b00000000000000000001010001110010;
assign LUT_1[26168] = 32'b00000000000000000011100110000011;
assign LUT_1[26169] = 32'b11111111111111111100110111111111;
assign LUT_1[26170] = 32'b11111111111111111111010100010100;
assign LUT_1[26171] = 32'b11111111111111111000100110010000;
assign LUT_1[26172] = 32'b00000000000000001011011111011010;
assign LUT_1[26173] = 32'b00000000000000000100110001010110;
assign LUT_1[26174] = 32'b00000000000000000111001101101011;
assign LUT_1[26175] = 32'b00000000000000000000011111100111;
assign LUT_1[26176] = 32'b00000000000000000011011111010101;
assign LUT_1[26177] = 32'b11111111111111111100110001010001;
assign LUT_1[26178] = 32'b11111111111111111111001101100110;
assign LUT_1[26179] = 32'b11111111111111111000011111100010;
assign LUT_1[26180] = 32'b00000000000000001011011000101100;
assign LUT_1[26181] = 32'b00000000000000000100101010101000;
assign LUT_1[26182] = 32'b00000000000000000111000110111101;
assign LUT_1[26183] = 32'b00000000000000000000011000111001;
assign LUT_1[26184] = 32'b00000000000000000010101101001010;
assign LUT_1[26185] = 32'b11111111111111111011111111000110;
assign LUT_1[26186] = 32'b11111111111111111110011011011011;
assign LUT_1[26187] = 32'b11111111111111110111101101010111;
assign LUT_1[26188] = 32'b00000000000000001010100110100001;
assign LUT_1[26189] = 32'b00000000000000000011111000011101;
assign LUT_1[26190] = 32'b00000000000000000110010100110010;
assign LUT_1[26191] = 32'b11111111111111111111100110101110;
assign LUT_1[26192] = 32'b00000000000000000101011010110111;
assign LUT_1[26193] = 32'b11111111111111111110101100110011;
assign LUT_1[26194] = 32'b00000000000000000001001001001000;
assign LUT_1[26195] = 32'b11111111111111111010011011000100;
assign LUT_1[26196] = 32'b00000000000000001101010100001110;
assign LUT_1[26197] = 32'b00000000000000000110100110001010;
assign LUT_1[26198] = 32'b00000000000000001001000010011111;
assign LUT_1[26199] = 32'b00000000000000000010010100011011;
assign LUT_1[26200] = 32'b00000000000000000100101000101100;
assign LUT_1[26201] = 32'b11111111111111111101111010101000;
assign LUT_1[26202] = 32'b00000000000000000000010110111101;
assign LUT_1[26203] = 32'b11111111111111111001101000111001;
assign LUT_1[26204] = 32'b00000000000000001100100010000011;
assign LUT_1[26205] = 32'b00000000000000000101110011111111;
assign LUT_1[26206] = 32'b00000000000000001000010000010100;
assign LUT_1[26207] = 32'b00000000000000000001100010010000;
assign LUT_1[26208] = 32'b00000000000000000100011010010100;
assign LUT_1[26209] = 32'b11111111111111111101101100010000;
assign LUT_1[26210] = 32'b00000000000000000000001000100101;
assign LUT_1[26211] = 32'b11111111111111111001011010100001;
assign LUT_1[26212] = 32'b00000000000000001100010011101011;
assign LUT_1[26213] = 32'b00000000000000000101100101100111;
assign LUT_1[26214] = 32'b00000000000000001000000001111100;
assign LUT_1[26215] = 32'b00000000000000000001010011111000;
assign LUT_1[26216] = 32'b00000000000000000011101000001001;
assign LUT_1[26217] = 32'b11111111111111111100111010000101;
assign LUT_1[26218] = 32'b11111111111111111111010110011010;
assign LUT_1[26219] = 32'b11111111111111111000101000010110;
assign LUT_1[26220] = 32'b00000000000000001011100001100000;
assign LUT_1[26221] = 32'b00000000000000000100110011011100;
assign LUT_1[26222] = 32'b00000000000000000111001111110001;
assign LUT_1[26223] = 32'b00000000000000000000100001101101;
assign LUT_1[26224] = 32'b00000000000000000110010101110110;
assign LUT_1[26225] = 32'b11111111111111111111100111110010;
assign LUT_1[26226] = 32'b00000000000000000010000100000111;
assign LUT_1[26227] = 32'b11111111111111111011010110000011;
assign LUT_1[26228] = 32'b00000000000000001110001111001101;
assign LUT_1[26229] = 32'b00000000000000000111100001001001;
assign LUT_1[26230] = 32'b00000000000000001001111101011110;
assign LUT_1[26231] = 32'b00000000000000000011001111011010;
assign LUT_1[26232] = 32'b00000000000000000101100011101011;
assign LUT_1[26233] = 32'b11111111111111111110110101100111;
assign LUT_1[26234] = 32'b00000000000000000001010001111100;
assign LUT_1[26235] = 32'b11111111111111111010100011111000;
assign LUT_1[26236] = 32'b00000000000000001101011101000010;
assign LUT_1[26237] = 32'b00000000000000000110101110111110;
assign LUT_1[26238] = 32'b00000000000000001001001011010011;
assign LUT_1[26239] = 32'b00000000000000000010011101001111;
assign LUT_1[26240] = 32'b00000000000000000100100001110000;
assign LUT_1[26241] = 32'b11111111111111111101110011101100;
assign LUT_1[26242] = 32'b00000000000000000000010000000001;
assign LUT_1[26243] = 32'b11111111111111111001100001111101;
assign LUT_1[26244] = 32'b00000000000000001100011011000111;
assign LUT_1[26245] = 32'b00000000000000000101101101000011;
assign LUT_1[26246] = 32'b00000000000000001000001001011000;
assign LUT_1[26247] = 32'b00000000000000000001011011010100;
assign LUT_1[26248] = 32'b00000000000000000011101111100101;
assign LUT_1[26249] = 32'b11111111111111111101000001100001;
assign LUT_1[26250] = 32'b11111111111111111111011101110110;
assign LUT_1[26251] = 32'b11111111111111111000101111110010;
assign LUT_1[26252] = 32'b00000000000000001011101000111100;
assign LUT_1[26253] = 32'b00000000000000000100111010111000;
assign LUT_1[26254] = 32'b00000000000000000111010111001101;
assign LUT_1[26255] = 32'b00000000000000000000101001001001;
assign LUT_1[26256] = 32'b00000000000000000110011101010010;
assign LUT_1[26257] = 32'b11111111111111111111101111001110;
assign LUT_1[26258] = 32'b00000000000000000010001011100011;
assign LUT_1[26259] = 32'b11111111111111111011011101011111;
assign LUT_1[26260] = 32'b00000000000000001110010110101001;
assign LUT_1[26261] = 32'b00000000000000000111101000100101;
assign LUT_1[26262] = 32'b00000000000000001010000100111010;
assign LUT_1[26263] = 32'b00000000000000000011010110110110;
assign LUT_1[26264] = 32'b00000000000000000101101011000111;
assign LUT_1[26265] = 32'b11111111111111111110111101000011;
assign LUT_1[26266] = 32'b00000000000000000001011001011000;
assign LUT_1[26267] = 32'b11111111111111111010101011010100;
assign LUT_1[26268] = 32'b00000000000000001101100100011110;
assign LUT_1[26269] = 32'b00000000000000000110110110011010;
assign LUT_1[26270] = 32'b00000000000000001001010010101111;
assign LUT_1[26271] = 32'b00000000000000000010100100101011;
assign LUT_1[26272] = 32'b00000000000000000101011100101111;
assign LUT_1[26273] = 32'b11111111111111111110101110101011;
assign LUT_1[26274] = 32'b00000000000000000001001011000000;
assign LUT_1[26275] = 32'b11111111111111111010011100111100;
assign LUT_1[26276] = 32'b00000000000000001101010110000110;
assign LUT_1[26277] = 32'b00000000000000000110101000000010;
assign LUT_1[26278] = 32'b00000000000000001001000100010111;
assign LUT_1[26279] = 32'b00000000000000000010010110010011;
assign LUT_1[26280] = 32'b00000000000000000100101010100100;
assign LUT_1[26281] = 32'b11111111111111111101111100100000;
assign LUT_1[26282] = 32'b00000000000000000000011000110101;
assign LUT_1[26283] = 32'b11111111111111111001101010110001;
assign LUT_1[26284] = 32'b00000000000000001100100011111011;
assign LUT_1[26285] = 32'b00000000000000000101110101110111;
assign LUT_1[26286] = 32'b00000000000000001000010010001100;
assign LUT_1[26287] = 32'b00000000000000000001100100001000;
assign LUT_1[26288] = 32'b00000000000000000111011000010001;
assign LUT_1[26289] = 32'b00000000000000000000101010001101;
assign LUT_1[26290] = 32'b00000000000000000011000110100010;
assign LUT_1[26291] = 32'b11111111111111111100011000011110;
assign LUT_1[26292] = 32'b00000000000000001111010001101000;
assign LUT_1[26293] = 32'b00000000000000001000100011100100;
assign LUT_1[26294] = 32'b00000000000000001010111111111001;
assign LUT_1[26295] = 32'b00000000000000000100010001110101;
assign LUT_1[26296] = 32'b00000000000000000110100110000110;
assign LUT_1[26297] = 32'b11111111111111111111111000000010;
assign LUT_1[26298] = 32'b00000000000000000010010100010111;
assign LUT_1[26299] = 32'b11111111111111111011100110010011;
assign LUT_1[26300] = 32'b00000000000000001110011111011101;
assign LUT_1[26301] = 32'b00000000000000000111110001011001;
assign LUT_1[26302] = 32'b00000000000000001010001101101110;
assign LUT_1[26303] = 32'b00000000000000000011011111101010;
assign LUT_1[26304] = 32'b00000000000000000110011111011000;
assign LUT_1[26305] = 32'b11111111111111111111110001010100;
assign LUT_1[26306] = 32'b00000000000000000010001101101001;
assign LUT_1[26307] = 32'b11111111111111111011011111100101;
assign LUT_1[26308] = 32'b00000000000000001110011000101111;
assign LUT_1[26309] = 32'b00000000000000000111101010101011;
assign LUT_1[26310] = 32'b00000000000000001010000111000000;
assign LUT_1[26311] = 32'b00000000000000000011011000111100;
assign LUT_1[26312] = 32'b00000000000000000101101101001101;
assign LUT_1[26313] = 32'b11111111111111111110111111001001;
assign LUT_1[26314] = 32'b00000000000000000001011011011110;
assign LUT_1[26315] = 32'b11111111111111111010101101011010;
assign LUT_1[26316] = 32'b00000000000000001101100110100100;
assign LUT_1[26317] = 32'b00000000000000000110111000100000;
assign LUT_1[26318] = 32'b00000000000000001001010100110101;
assign LUT_1[26319] = 32'b00000000000000000010100110110001;
assign LUT_1[26320] = 32'b00000000000000001000011010111010;
assign LUT_1[26321] = 32'b00000000000000000001101100110110;
assign LUT_1[26322] = 32'b00000000000000000100001001001011;
assign LUT_1[26323] = 32'b11111111111111111101011011000111;
assign LUT_1[26324] = 32'b00000000000000010000010100010001;
assign LUT_1[26325] = 32'b00000000000000001001100110001101;
assign LUT_1[26326] = 32'b00000000000000001100000010100010;
assign LUT_1[26327] = 32'b00000000000000000101010100011110;
assign LUT_1[26328] = 32'b00000000000000000111101000101111;
assign LUT_1[26329] = 32'b00000000000000000000111010101011;
assign LUT_1[26330] = 32'b00000000000000000011010111000000;
assign LUT_1[26331] = 32'b11111111111111111100101000111100;
assign LUT_1[26332] = 32'b00000000000000001111100010000110;
assign LUT_1[26333] = 32'b00000000000000001000110100000010;
assign LUT_1[26334] = 32'b00000000000000001011010000010111;
assign LUT_1[26335] = 32'b00000000000000000100100010010011;
assign LUT_1[26336] = 32'b00000000000000000111011010010111;
assign LUT_1[26337] = 32'b00000000000000000000101100010011;
assign LUT_1[26338] = 32'b00000000000000000011001000101000;
assign LUT_1[26339] = 32'b11111111111111111100011010100100;
assign LUT_1[26340] = 32'b00000000000000001111010011101110;
assign LUT_1[26341] = 32'b00000000000000001000100101101010;
assign LUT_1[26342] = 32'b00000000000000001011000001111111;
assign LUT_1[26343] = 32'b00000000000000000100010011111011;
assign LUT_1[26344] = 32'b00000000000000000110101000001100;
assign LUT_1[26345] = 32'b11111111111111111111111010001000;
assign LUT_1[26346] = 32'b00000000000000000010010110011101;
assign LUT_1[26347] = 32'b11111111111111111011101000011001;
assign LUT_1[26348] = 32'b00000000000000001110100001100011;
assign LUT_1[26349] = 32'b00000000000000000111110011011111;
assign LUT_1[26350] = 32'b00000000000000001010001111110100;
assign LUT_1[26351] = 32'b00000000000000000011100001110000;
assign LUT_1[26352] = 32'b00000000000000001001010101111001;
assign LUT_1[26353] = 32'b00000000000000000010100111110101;
assign LUT_1[26354] = 32'b00000000000000000101000100001010;
assign LUT_1[26355] = 32'b11111111111111111110010110000110;
assign LUT_1[26356] = 32'b00000000000000010001001111010000;
assign LUT_1[26357] = 32'b00000000000000001010100001001100;
assign LUT_1[26358] = 32'b00000000000000001100111101100001;
assign LUT_1[26359] = 32'b00000000000000000110001111011101;
assign LUT_1[26360] = 32'b00000000000000001000100011101110;
assign LUT_1[26361] = 32'b00000000000000000001110101101010;
assign LUT_1[26362] = 32'b00000000000000000100010001111111;
assign LUT_1[26363] = 32'b11111111111111111101100011111011;
assign LUT_1[26364] = 32'b00000000000000010000011101000101;
assign LUT_1[26365] = 32'b00000000000000001001101111000001;
assign LUT_1[26366] = 32'b00000000000000001100001011010110;
assign LUT_1[26367] = 32'b00000000000000000101011101010010;
assign LUT_1[26368] = 32'b11111111111111111111010101111001;
assign LUT_1[26369] = 32'b11111111111111111000100111110101;
assign LUT_1[26370] = 32'b11111111111111111011000100001010;
assign LUT_1[26371] = 32'b11111111111111110100010110000110;
assign LUT_1[26372] = 32'b00000000000000000111001111010000;
assign LUT_1[26373] = 32'b00000000000000000000100001001100;
assign LUT_1[26374] = 32'b00000000000000000010111101100001;
assign LUT_1[26375] = 32'b11111111111111111100001111011101;
assign LUT_1[26376] = 32'b11111111111111111110100011101110;
assign LUT_1[26377] = 32'b11111111111111110111110101101010;
assign LUT_1[26378] = 32'b11111111111111111010010001111111;
assign LUT_1[26379] = 32'b11111111111111110011100011111011;
assign LUT_1[26380] = 32'b00000000000000000110011101000101;
assign LUT_1[26381] = 32'b11111111111111111111101111000001;
assign LUT_1[26382] = 32'b00000000000000000010001011010110;
assign LUT_1[26383] = 32'b11111111111111111011011101010010;
assign LUT_1[26384] = 32'b00000000000000000001010001011011;
assign LUT_1[26385] = 32'b11111111111111111010100011010111;
assign LUT_1[26386] = 32'b11111111111111111100111111101100;
assign LUT_1[26387] = 32'b11111111111111110110010001101000;
assign LUT_1[26388] = 32'b00000000000000001001001010110010;
assign LUT_1[26389] = 32'b00000000000000000010011100101110;
assign LUT_1[26390] = 32'b00000000000000000100111001000011;
assign LUT_1[26391] = 32'b11111111111111111110001010111111;
assign LUT_1[26392] = 32'b00000000000000000000011111010000;
assign LUT_1[26393] = 32'b11111111111111111001110001001100;
assign LUT_1[26394] = 32'b11111111111111111100001101100001;
assign LUT_1[26395] = 32'b11111111111111110101011111011101;
assign LUT_1[26396] = 32'b00000000000000001000011000100111;
assign LUT_1[26397] = 32'b00000000000000000001101010100011;
assign LUT_1[26398] = 32'b00000000000000000100000110111000;
assign LUT_1[26399] = 32'b11111111111111111101011000110100;
assign LUT_1[26400] = 32'b00000000000000000000010000111000;
assign LUT_1[26401] = 32'b11111111111111111001100010110100;
assign LUT_1[26402] = 32'b11111111111111111011111111001001;
assign LUT_1[26403] = 32'b11111111111111110101010001000101;
assign LUT_1[26404] = 32'b00000000000000001000001010001111;
assign LUT_1[26405] = 32'b00000000000000000001011100001011;
assign LUT_1[26406] = 32'b00000000000000000011111000100000;
assign LUT_1[26407] = 32'b11111111111111111101001010011100;
assign LUT_1[26408] = 32'b11111111111111111111011110101101;
assign LUT_1[26409] = 32'b11111111111111111000110000101001;
assign LUT_1[26410] = 32'b11111111111111111011001100111110;
assign LUT_1[26411] = 32'b11111111111111110100011110111010;
assign LUT_1[26412] = 32'b00000000000000000111011000000100;
assign LUT_1[26413] = 32'b00000000000000000000101010000000;
assign LUT_1[26414] = 32'b00000000000000000011000110010101;
assign LUT_1[26415] = 32'b11111111111111111100011000010001;
assign LUT_1[26416] = 32'b00000000000000000010001100011010;
assign LUT_1[26417] = 32'b11111111111111111011011110010110;
assign LUT_1[26418] = 32'b11111111111111111101111010101011;
assign LUT_1[26419] = 32'b11111111111111110111001100100111;
assign LUT_1[26420] = 32'b00000000000000001010000101110001;
assign LUT_1[26421] = 32'b00000000000000000011010111101101;
assign LUT_1[26422] = 32'b00000000000000000101110100000010;
assign LUT_1[26423] = 32'b11111111111111111111000101111110;
assign LUT_1[26424] = 32'b00000000000000000001011010001111;
assign LUT_1[26425] = 32'b11111111111111111010101100001011;
assign LUT_1[26426] = 32'b11111111111111111101001000100000;
assign LUT_1[26427] = 32'b11111111111111110110011010011100;
assign LUT_1[26428] = 32'b00000000000000001001010011100110;
assign LUT_1[26429] = 32'b00000000000000000010100101100010;
assign LUT_1[26430] = 32'b00000000000000000101000001110111;
assign LUT_1[26431] = 32'b11111111111111111110010011110011;
assign LUT_1[26432] = 32'b00000000000000000001010011100001;
assign LUT_1[26433] = 32'b11111111111111111010100101011101;
assign LUT_1[26434] = 32'b11111111111111111101000001110010;
assign LUT_1[26435] = 32'b11111111111111110110010011101110;
assign LUT_1[26436] = 32'b00000000000000001001001100111000;
assign LUT_1[26437] = 32'b00000000000000000010011110110100;
assign LUT_1[26438] = 32'b00000000000000000100111011001001;
assign LUT_1[26439] = 32'b11111111111111111110001101000101;
assign LUT_1[26440] = 32'b00000000000000000000100001010110;
assign LUT_1[26441] = 32'b11111111111111111001110011010010;
assign LUT_1[26442] = 32'b11111111111111111100001111100111;
assign LUT_1[26443] = 32'b11111111111111110101100001100011;
assign LUT_1[26444] = 32'b00000000000000001000011010101101;
assign LUT_1[26445] = 32'b00000000000000000001101100101001;
assign LUT_1[26446] = 32'b00000000000000000100001000111110;
assign LUT_1[26447] = 32'b11111111111111111101011010111010;
assign LUT_1[26448] = 32'b00000000000000000011001111000011;
assign LUT_1[26449] = 32'b11111111111111111100100000111111;
assign LUT_1[26450] = 32'b11111111111111111110111101010100;
assign LUT_1[26451] = 32'b11111111111111111000001111010000;
assign LUT_1[26452] = 32'b00000000000000001011001000011010;
assign LUT_1[26453] = 32'b00000000000000000100011010010110;
assign LUT_1[26454] = 32'b00000000000000000110110110101011;
assign LUT_1[26455] = 32'b00000000000000000000001000100111;
assign LUT_1[26456] = 32'b00000000000000000010011100111000;
assign LUT_1[26457] = 32'b11111111111111111011101110110100;
assign LUT_1[26458] = 32'b11111111111111111110001011001001;
assign LUT_1[26459] = 32'b11111111111111110111011101000101;
assign LUT_1[26460] = 32'b00000000000000001010010110001111;
assign LUT_1[26461] = 32'b00000000000000000011101000001011;
assign LUT_1[26462] = 32'b00000000000000000110000100100000;
assign LUT_1[26463] = 32'b11111111111111111111010110011100;
assign LUT_1[26464] = 32'b00000000000000000010001110100000;
assign LUT_1[26465] = 32'b11111111111111111011100000011100;
assign LUT_1[26466] = 32'b11111111111111111101111100110001;
assign LUT_1[26467] = 32'b11111111111111110111001110101101;
assign LUT_1[26468] = 32'b00000000000000001010000111110111;
assign LUT_1[26469] = 32'b00000000000000000011011001110011;
assign LUT_1[26470] = 32'b00000000000000000101110110001000;
assign LUT_1[26471] = 32'b11111111111111111111001000000100;
assign LUT_1[26472] = 32'b00000000000000000001011100010101;
assign LUT_1[26473] = 32'b11111111111111111010101110010001;
assign LUT_1[26474] = 32'b11111111111111111101001010100110;
assign LUT_1[26475] = 32'b11111111111111110110011100100010;
assign LUT_1[26476] = 32'b00000000000000001001010101101100;
assign LUT_1[26477] = 32'b00000000000000000010100111101000;
assign LUT_1[26478] = 32'b00000000000000000101000011111101;
assign LUT_1[26479] = 32'b11111111111111111110010101111001;
assign LUT_1[26480] = 32'b00000000000000000100001010000010;
assign LUT_1[26481] = 32'b11111111111111111101011011111110;
assign LUT_1[26482] = 32'b11111111111111111111111000010011;
assign LUT_1[26483] = 32'b11111111111111111001001010001111;
assign LUT_1[26484] = 32'b00000000000000001100000011011001;
assign LUT_1[26485] = 32'b00000000000000000101010101010101;
assign LUT_1[26486] = 32'b00000000000000000111110001101010;
assign LUT_1[26487] = 32'b00000000000000000001000011100110;
assign LUT_1[26488] = 32'b00000000000000000011010111110111;
assign LUT_1[26489] = 32'b11111111111111111100101001110011;
assign LUT_1[26490] = 32'b11111111111111111111000110001000;
assign LUT_1[26491] = 32'b11111111111111111000011000000100;
assign LUT_1[26492] = 32'b00000000000000001011010001001110;
assign LUT_1[26493] = 32'b00000000000000000100100011001010;
assign LUT_1[26494] = 32'b00000000000000000110111111011111;
assign LUT_1[26495] = 32'b00000000000000000000010001011011;
assign LUT_1[26496] = 32'b00000000000000000010010101111100;
assign LUT_1[26497] = 32'b11111111111111111011100111111000;
assign LUT_1[26498] = 32'b11111111111111111110000100001101;
assign LUT_1[26499] = 32'b11111111111111110111010110001001;
assign LUT_1[26500] = 32'b00000000000000001010001111010011;
assign LUT_1[26501] = 32'b00000000000000000011100001001111;
assign LUT_1[26502] = 32'b00000000000000000101111101100100;
assign LUT_1[26503] = 32'b11111111111111111111001111100000;
assign LUT_1[26504] = 32'b00000000000000000001100011110001;
assign LUT_1[26505] = 32'b11111111111111111010110101101101;
assign LUT_1[26506] = 32'b11111111111111111101010010000010;
assign LUT_1[26507] = 32'b11111111111111110110100011111110;
assign LUT_1[26508] = 32'b00000000000000001001011101001000;
assign LUT_1[26509] = 32'b00000000000000000010101111000100;
assign LUT_1[26510] = 32'b00000000000000000101001011011001;
assign LUT_1[26511] = 32'b11111111111111111110011101010101;
assign LUT_1[26512] = 32'b00000000000000000100010001011110;
assign LUT_1[26513] = 32'b11111111111111111101100011011010;
assign LUT_1[26514] = 32'b11111111111111111111111111101111;
assign LUT_1[26515] = 32'b11111111111111111001010001101011;
assign LUT_1[26516] = 32'b00000000000000001100001010110101;
assign LUT_1[26517] = 32'b00000000000000000101011100110001;
assign LUT_1[26518] = 32'b00000000000000000111111001000110;
assign LUT_1[26519] = 32'b00000000000000000001001011000010;
assign LUT_1[26520] = 32'b00000000000000000011011111010011;
assign LUT_1[26521] = 32'b11111111111111111100110001001111;
assign LUT_1[26522] = 32'b11111111111111111111001101100100;
assign LUT_1[26523] = 32'b11111111111111111000011111100000;
assign LUT_1[26524] = 32'b00000000000000001011011000101010;
assign LUT_1[26525] = 32'b00000000000000000100101010100110;
assign LUT_1[26526] = 32'b00000000000000000111000110111011;
assign LUT_1[26527] = 32'b00000000000000000000011000110111;
assign LUT_1[26528] = 32'b00000000000000000011010000111011;
assign LUT_1[26529] = 32'b11111111111111111100100010110111;
assign LUT_1[26530] = 32'b11111111111111111110111111001100;
assign LUT_1[26531] = 32'b11111111111111111000010001001000;
assign LUT_1[26532] = 32'b00000000000000001011001010010010;
assign LUT_1[26533] = 32'b00000000000000000100011100001110;
assign LUT_1[26534] = 32'b00000000000000000110111000100011;
assign LUT_1[26535] = 32'b00000000000000000000001010011111;
assign LUT_1[26536] = 32'b00000000000000000010011110110000;
assign LUT_1[26537] = 32'b11111111111111111011110000101100;
assign LUT_1[26538] = 32'b11111111111111111110001101000001;
assign LUT_1[26539] = 32'b11111111111111110111011110111101;
assign LUT_1[26540] = 32'b00000000000000001010011000000111;
assign LUT_1[26541] = 32'b00000000000000000011101010000011;
assign LUT_1[26542] = 32'b00000000000000000110000110011000;
assign LUT_1[26543] = 32'b11111111111111111111011000010100;
assign LUT_1[26544] = 32'b00000000000000000101001100011101;
assign LUT_1[26545] = 32'b11111111111111111110011110011001;
assign LUT_1[26546] = 32'b00000000000000000000111010101110;
assign LUT_1[26547] = 32'b11111111111111111010001100101010;
assign LUT_1[26548] = 32'b00000000000000001101000101110100;
assign LUT_1[26549] = 32'b00000000000000000110010111110000;
assign LUT_1[26550] = 32'b00000000000000001000110100000101;
assign LUT_1[26551] = 32'b00000000000000000010000110000001;
assign LUT_1[26552] = 32'b00000000000000000100011010010010;
assign LUT_1[26553] = 32'b11111111111111111101101100001110;
assign LUT_1[26554] = 32'b00000000000000000000001000100011;
assign LUT_1[26555] = 32'b11111111111111111001011010011111;
assign LUT_1[26556] = 32'b00000000000000001100010011101001;
assign LUT_1[26557] = 32'b00000000000000000101100101100101;
assign LUT_1[26558] = 32'b00000000000000001000000001111010;
assign LUT_1[26559] = 32'b00000000000000000001010011110110;
assign LUT_1[26560] = 32'b00000000000000000100010011100100;
assign LUT_1[26561] = 32'b11111111111111111101100101100000;
assign LUT_1[26562] = 32'b00000000000000000000000001110101;
assign LUT_1[26563] = 32'b11111111111111111001010011110001;
assign LUT_1[26564] = 32'b00000000000000001100001100111011;
assign LUT_1[26565] = 32'b00000000000000000101011110110111;
assign LUT_1[26566] = 32'b00000000000000000111111011001100;
assign LUT_1[26567] = 32'b00000000000000000001001101001000;
assign LUT_1[26568] = 32'b00000000000000000011100001011001;
assign LUT_1[26569] = 32'b11111111111111111100110011010101;
assign LUT_1[26570] = 32'b11111111111111111111001111101010;
assign LUT_1[26571] = 32'b11111111111111111000100001100110;
assign LUT_1[26572] = 32'b00000000000000001011011010110000;
assign LUT_1[26573] = 32'b00000000000000000100101100101100;
assign LUT_1[26574] = 32'b00000000000000000111001001000001;
assign LUT_1[26575] = 32'b00000000000000000000011010111101;
assign LUT_1[26576] = 32'b00000000000000000110001111000110;
assign LUT_1[26577] = 32'b11111111111111111111100001000010;
assign LUT_1[26578] = 32'b00000000000000000001111101010111;
assign LUT_1[26579] = 32'b11111111111111111011001111010011;
assign LUT_1[26580] = 32'b00000000000000001110001000011101;
assign LUT_1[26581] = 32'b00000000000000000111011010011001;
assign LUT_1[26582] = 32'b00000000000000001001110110101110;
assign LUT_1[26583] = 32'b00000000000000000011001000101010;
assign LUT_1[26584] = 32'b00000000000000000101011100111011;
assign LUT_1[26585] = 32'b11111111111111111110101110110111;
assign LUT_1[26586] = 32'b00000000000000000001001011001100;
assign LUT_1[26587] = 32'b11111111111111111010011101001000;
assign LUT_1[26588] = 32'b00000000000000001101010110010010;
assign LUT_1[26589] = 32'b00000000000000000110101000001110;
assign LUT_1[26590] = 32'b00000000000000001001000100100011;
assign LUT_1[26591] = 32'b00000000000000000010010110011111;
assign LUT_1[26592] = 32'b00000000000000000101001110100011;
assign LUT_1[26593] = 32'b11111111111111111110100000011111;
assign LUT_1[26594] = 32'b00000000000000000000111100110100;
assign LUT_1[26595] = 32'b11111111111111111010001110110000;
assign LUT_1[26596] = 32'b00000000000000001101000111111010;
assign LUT_1[26597] = 32'b00000000000000000110011001110110;
assign LUT_1[26598] = 32'b00000000000000001000110110001011;
assign LUT_1[26599] = 32'b00000000000000000010001000000111;
assign LUT_1[26600] = 32'b00000000000000000100011100011000;
assign LUT_1[26601] = 32'b11111111111111111101101110010100;
assign LUT_1[26602] = 32'b00000000000000000000001010101001;
assign LUT_1[26603] = 32'b11111111111111111001011100100101;
assign LUT_1[26604] = 32'b00000000000000001100010101101111;
assign LUT_1[26605] = 32'b00000000000000000101100111101011;
assign LUT_1[26606] = 32'b00000000000000001000000100000000;
assign LUT_1[26607] = 32'b00000000000000000001010101111100;
assign LUT_1[26608] = 32'b00000000000000000111001010000101;
assign LUT_1[26609] = 32'b00000000000000000000011100000001;
assign LUT_1[26610] = 32'b00000000000000000010111000010110;
assign LUT_1[26611] = 32'b11111111111111111100001010010010;
assign LUT_1[26612] = 32'b00000000000000001111000011011100;
assign LUT_1[26613] = 32'b00000000000000001000010101011000;
assign LUT_1[26614] = 32'b00000000000000001010110001101101;
assign LUT_1[26615] = 32'b00000000000000000100000011101001;
assign LUT_1[26616] = 32'b00000000000000000110010111111010;
assign LUT_1[26617] = 32'b11111111111111111111101001110110;
assign LUT_1[26618] = 32'b00000000000000000010000110001011;
assign LUT_1[26619] = 32'b11111111111111111011011000000111;
assign LUT_1[26620] = 32'b00000000000000001110010001010001;
assign LUT_1[26621] = 32'b00000000000000000111100011001101;
assign LUT_1[26622] = 32'b00000000000000001001111111100010;
assign LUT_1[26623] = 32'b00000000000000000011010001011110;
assign LUT_1[26624] = 32'b00000000000000000010011110011011;
assign LUT_1[26625] = 32'b11111111111111111011110000010111;
assign LUT_1[26626] = 32'b11111111111111111110001100101100;
assign LUT_1[26627] = 32'b11111111111111110111011110101000;
assign LUT_1[26628] = 32'b00000000000000001010010111110010;
assign LUT_1[26629] = 32'b00000000000000000011101001101110;
assign LUT_1[26630] = 32'b00000000000000000110000110000011;
assign LUT_1[26631] = 32'b11111111111111111111010111111111;
assign LUT_1[26632] = 32'b00000000000000000001101100010000;
assign LUT_1[26633] = 32'b11111111111111111010111110001100;
assign LUT_1[26634] = 32'b11111111111111111101011010100001;
assign LUT_1[26635] = 32'b11111111111111110110101100011101;
assign LUT_1[26636] = 32'b00000000000000001001100101100111;
assign LUT_1[26637] = 32'b00000000000000000010110111100011;
assign LUT_1[26638] = 32'b00000000000000000101010011111000;
assign LUT_1[26639] = 32'b11111111111111111110100101110100;
assign LUT_1[26640] = 32'b00000000000000000100011001111101;
assign LUT_1[26641] = 32'b11111111111111111101101011111001;
assign LUT_1[26642] = 32'b00000000000000000000001000001110;
assign LUT_1[26643] = 32'b11111111111111111001011010001010;
assign LUT_1[26644] = 32'b00000000000000001100010011010100;
assign LUT_1[26645] = 32'b00000000000000000101100101010000;
assign LUT_1[26646] = 32'b00000000000000001000000001100101;
assign LUT_1[26647] = 32'b00000000000000000001010011100001;
assign LUT_1[26648] = 32'b00000000000000000011100111110010;
assign LUT_1[26649] = 32'b11111111111111111100111001101110;
assign LUT_1[26650] = 32'b11111111111111111111010110000011;
assign LUT_1[26651] = 32'b11111111111111111000100111111111;
assign LUT_1[26652] = 32'b00000000000000001011100001001001;
assign LUT_1[26653] = 32'b00000000000000000100110011000101;
assign LUT_1[26654] = 32'b00000000000000000111001111011010;
assign LUT_1[26655] = 32'b00000000000000000000100001010110;
assign LUT_1[26656] = 32'b00000000000000000011011001011010;
assign LUT_1[26657] = 32'b11111111111111111100101011010110;
assign LUT_1[26658] = 32'b11111111111111111111000111101011;
assign LUT_1[26659] = 32'b11111111111111111000011001100111;
assign LUT_1[26660] = 32'b00000000000000001011010010110001;
assign LUT_1[26661] = 32'b00000000000000000100100100101101;
assign LUT_1[26662] = 32'b00000000000000000111000001000010;
assign LUT_1[26663] = 32'b00000000000000000000010010111110;
assign LUT_1[26664] = 32'b00000000000000000010100111001111;
assign LUT_1[26665] = 32'b11111111111111111011111001001011;
assign LUT_1[26666] = 32'b11111111111111111110010101100000;
assign LUT_1[26667] = 32'b11111111111111110111100111011100;
assign LUT_1[26668] = 32'b00000000000000001010100000100110;
assign LUT_1[26669] = 32'b00000000000000000011110010100010;
assign LUT_1[26670] = 32'b00000000000000000110001110110111;
assign LUT_1[26671] = 32'b11111111111111111111100000110011;
assign LUT_1[26672] = 32'b00000000000000000101010100111100;
assign LUT_1[26673] = 32'b11111111111111111110100110111000;
assign LUT_1[26674] = 32'b00000000000000000001000011001101;
assign LUT_1[26675] = 32'b11111111111111111010010101001001;
assign LUT_1[26676] = 32'b00000000000000001101001110010011;
assign LUT_1[26677] = 32'b00000000000000000110100000001111;
assign LUT_1[26678] = 32'b00000000000000001000111100100100;
assign LUT_1[26679] = 32'b00000000000000000010001110100000;
assign LUT_1[26680] = 32'b00000000000000000100100010110001;
assign LUT_1[26681] = 32'b11111111111111111101110100101101;
assign LUT_1[26682] = 32'b00000000000000000000010001000010;
assign LUT_1[26683] = 32'b11111111111111111001100010111110;
assign LUT_1[26684] = 32'b00000000000000001100011100001000;
assign LUT_1[26685] = 32'b00000000000000000101101110000100;
assign LUT_1[26686] = 32'b00000000000000001000001010011001;
assign LUT_1[26687] = 32'b00000000000000000001011100010101;
assign LUT_1[26688] = 32'b00000000000000000100011100000011;
assign LUT_1[26689] = 32'b11111111111111111101101101111111;
assign LUT_1[26690] = 32'b00000000000000000000001010010100;
assign LUT_1[26691] = 32'b11111111111111111001011100010000;
assign LUT_1[26692] = 32'b00000000000000001100010101011010;
assign LUT_1[26693] = 32'b00000000000000000101100111010110;
assign LUT_1[26694] = 32'b00000000000000001000000011101011;
assign LUT_1[26695] = 32'b00000000000000000001010101100111;
assign LUT_1[26696] = 32'b00000000000000000011101001111000;
assign LUT_1[26697] = 32'b11111111111111111100111011110100;
assign LUT_1[26698] = 32'b11111111111111111111011000001001;
assign LUT_1[26699] = 32'b11111111111111111000101010000101;
assign LUT_1[26700] = 32'b00000000000000001011100011001111;
assign LUT_1[26701] = 32'b00000000000000000100110101001011;
assign LUT_1[26702] = 32'b00000000000000000111010001100000;
assign LUT_1[26703] = 32'b00000000000000000000100011011100;
assign LUT_1[26704] = 32'b00000000000000000110010111100101;
assign LUT_1[26705] = 32'b11111111111111111111101001100001;
assign LUT_1[26706] = 32'b00000000000000000010000101110110;
assign LUT_1[26707] = 32'b11111111111111111011010111110010;
assign LUT_1[26708] = 32'b00000000000000001110010000111100;
assign LUT_1[26709] = 32'b00000000000000000111100010111000;
assign LUT_1[26710] = 32'b00000000000000001001111111001101;
assign LUT_1[26711] = 32'b00000000000000000011010001001001;
assign LUT_1[26712] = 32'b00000000000000000101100101011010;
assign LUT_1[26713] = 32'b11111111111111111110110111010110;
assign LUT_1[26714] = 32'b00000000000000000001010011101011;
assign LUT_1[26715] = 32'b11111111111111111010100101100111;
assign LUT_1[26716] = 32'b00000000000000001101011110110001;
assign LUT_1[26717] = 32'b00000000000000000110110000101101;
assign LUT_1[26718] = 32'b00000000000000001001001101000010;
assign LUT_1[26719] = 32'b00000000000000000010011110111110;
assign LUT_1[26720] = 32'b00000000000000000101010111000010;
assign LUT_1[26721] = 32'b11111111111111111110101000111110;
assign LUT_1[26722] = 32'b00000000000000000001000101010011;
assign LUT_1[26723] = 32'b11111111111111111010010111001111;
assign LUT_1[26724] = 32'b00000000000000001101010000011001;
assign LUT_1[26725] = 32'b00000000000000000110100010010101;
assign LUT_1[26726] = 32'b00000000000000001000111110101010;
assign LUT_1[26727] = 32'b00000000000000000010010000100110;
assign LUT_1[26728] = 32'b00000000000000000100100100110111;
assign LUT_1[26729] = 32'b11111111111111111101110110110011;
assign LUT_1[26730] = 32'b00000000000000000000010011001000;
assign LUT_1[26731] = 32'b11111111111111111001100101000100;
assign LUT_1[26732] = 32'b00000000000000001100011110001110;
assign LUT_1[26733] = 32'b00000000000000000101110000001010;
assign LUT_1[26734] = 32'b00000000000000001000001100011111;
assign LUT_1[26735] = 32'b00000000000000000001011110011011;
assign LUT_1[26736] = 32'b00000000000000000111010010100100;
assign LUT_1[26737] = 32'b00000000000000000000100100100000;
assign LUT_1[26738] = 32'b00000000000000000011000000110101;
assign LUT_1[26739] = 32'b11111111111111111100010010110001;
assign LUT_1[26740] = 32'b00000000000000001111001011111011;
assign LUT_1[26741] = 32'b00000000000000001000011101110111;
assign LUT_1[26742] = 32'b00000000000000001010111010001100;
assign LUT_1[26743] = 32'b00000000000000000100001100001000;
assign LUT_1[26744] = 32'b00000000000000000110100000011001;
assign LUT_1[26745] = 32'b11111111111111111111110010010101;
assign LUT_1[26746] = 32'b00000000000000000010001110101010;
assign LUT_1[26747] = 32'b11111111111111111011100000100110;
assign LUT_1[26748] = 32'b00000000000000001110011001110000;
assign LUT_1[26749] = 32'b00000000000000000111101011101100;
assign LUT_1[26750] = 32'b00000000000000001010001000000001;
assign LUT_1[26751] = 32'b00000000000000000011011001111101;
assign LUT_1[26752] = 32'b00000000000000000101011110011110;
assign LUT_1[26753] = 32'b11111111111111111110110000011010;
assign LUT_1[26754] = 32'b00000000000000000001001100101111;
assign LUT_1[26755] = 32'b11111111111111111010011110101011;
assign LUT_1[26756] = 32'b00000000000000001101010111110101;
assign LUT_1[26757] = 32'b00000000000000000110101001110001;
assign LUT_1[26758] = 32'b00000000000000001001000110000110;
assign LUT_1[26759] = 32'b00000000000000000010011000000010;
assign LUT_1[26760] = 32'b00000000000000000100101100010011;
assign LUT_1[26761] = 32'b11111111111111111101111110001111;
assign LUT_1[26762] = 32'b00000000000000000000011010100100;
assign LUT_1[26763] = 32'b11111111111111111001101100100000;
assign LUT_1[26764] = 32'b00000000000000001100100101101010;
assign LUT_1[26765] = 32'b00000000000000000101110111100110;
assign LUT_1[26766] = 32'b00000000000000001000010011111011;
assign LUT_1[26767] = 32'b00000000000000000001100101110111;
assign LUT_1[26768] = 32'b00000000000000000111011010000000;
assign LUT_1[26769] = 32'b00000000000000000000101011111100;
assign LUT_1[26770] = 32'b00000000000000000011001000010001;
assign LUT_1[26771] = 32'b11111111111111111100011010001101;
assign LUT_1[26772] = 32'b00000000000000001111010011010111;
assign LUT_1[26773] = 32'b00000000000000001000100101010011;
assign LUT_1[26774] = 32'b00000000000000001011000001101000;
assign LUT_1[26775] = 32'b00000000000000000100010011100100;
assign LUT_1[26776] = 32'b00000000000000000110100111110101;
assign LUT_1[26777] = 32'b11111111111111111111111001110001;
assign LUT_1[26778] = 32'b00000000000000000010010110000110;
assign LUT_1[26779] = 32'b11111111111111111011101000000010;
assign LUT_1[26780] = 32'b00000000000000001110100001001100;
assign LUT_1[26781] = 32'b00000000000000000111110011001000;
assign LUT_1[26782] = 32'b00000000000000001010001111011101;
assign LUT_1[26783] = 32'b00000000000000000011100001011001;
assign LUT_1[26784] = 32'b00000000000000000110011001011101;
assign LUT_1[26785] = 32'b11111111111111111111101011011001;
assign LUT_1[26786] = 32'b00000000000000000010000111101110;
assign LUT_1[26787] = 32'b11111111111111111011011001101010;
assign LUT_1[26788] = 32'b00000000000000001110010010110100;
assign LUT_1[26789] = 32'b00000000000000000111100100110000;
assign LUT_1[26790] = 32'b00000000000000001010000001000101;
assign LUT_1[26791] = 32'b00000000000000000011010011000001;
assign LUT_1[26792] = 32'b00000000000000000101100111010010;
assign LUT_1[26793] = 32'b11111111111111111110111001001110;
assign LUT_1[26794] = 32'b00000000000000000001010101100011;
assign LUT_1[26795] = 32'b11111111111111111010100111011111;
assign LUT_1[26796] = 32'b00000000000000001101100000101001;
assign LUT_1[26797] = 32'b00000000000000000110110010100101;
assign LUT_1[26798] = 32'b00000000000000001001001110111010;
assign LUT_1[26799] = 32'b00000000000000000010100000110110;
assign LUT_1[26800] = 32'b00000000000000001000010100111111;
assign LUT_1[26801] = 32'b00000000000000000001100110111011;
assign LUT_1[26802] = 32'b00000000000000000100000011010000;
assign LUT_1[26803] = 32'b11111111111111111101010101001100;
assign LUT_1[26804] = 32'b00000000000000010000001110010110;
assign LUT_1[26805] = 32'b00000000000000001001100000010010;
assign LUT_1[26806] = 32'b00000000000000001011111100100111;
assign LUT_1[26807] = 32'b00000000000000000101001110100011;
assign LUT_1[26808] = 32'b00000000000000000111100010110100;
assign LUT_1[26809] = 32'b00000000000000000000110100110000;
assign LUT_1[26810] = 32'b00000000000000000011010001000101;
assign LUT_1[26811] = 32'b11111111111111111100100011000001;
assign LUT_1[26812] = 32'b00000000000000001111011100001011;
assign LUT_1[26813] = 32'b00000000000000001000101110000111;
assign LUT_1[26814] = 32'b00000000000000001011001010011100;
assign LUT_1[26815] = 32'b00000000000000000100011100011000;
assign LUT_1[26816] = 32'b00000000000000000111011100000110;
assign LUT_1[26817] = 32'b00000000000000000000101110000010;
assign LUT_1[26818] = 32'b00000000000000000011001010010111;
assign LUT_1[26819] = 32'b11111111111111111100011100010011;
assign LUT_1[26820] = 32'b00000000000000001111010101011101;
assign LUT_1[26821] = 32'b00000000000000001000100111011001;
assign LUT_1[26822] = 32'b00000000000000001011000011101110;
assign LUT_1[26823] = 32'b00000000000000000100010101101010;
assign LUT_1[26824] = 32'b00000000000000000110101001111011;
assign LUT_1[26825] = 32'b11111111111111111111111011110111;
assign LUT_1[26826] = 32'b00000000000000000010011000001100;
assign LUT_1[26827] = 32'b11111111111111111011101010001000;
assign LUT_1[26828] = 32'b00000000000000001110100011010010;
assign LUT_1[26829] = 32'b00000000000000000111110101001110;
assign LUT_1[26830] = 32'b00000000000000001010010001100011;
assign LUT_1[26831] = 32'b00000000000000000011100011011111;
assign LUT_1[26832] = 32'b00000000000000001001010111101000;
assign LUT_1[26833] = 32'b00000000000000000010101001100100;
assign LUT_1[26834] = 32'b00000000000000000101000101111001;
assign LUT_1[26835] = 32'b11111111111111111110010111110101;
assign LUT_1[26836] = 32'b00000000000000010001010000111111;
assign LUT_1[26837] = 32'b00000000000000001010100010111011;
assign LUT_1[26838] = 32'b00000000000000001100111111010000;
assign LUT_1[26839] = 32'b00000000000000000110010001001100;
assign LUT_1[26840] = 32'b00000000000000001000100101011101;
assign LUT_1[26841] = 32'b00000000000000000001110111011001;
assign LUT_1[26842] = 32'b00000000000000000100010011101110;
assign LUT_1[26843] = 32'b11111111111111111101100101101010;
assign LUT_1[26844] = 32'b00000000000000010000011110110100;
assign LUT_1[26845] = 32'b00000000000000001001110000110000;
assign LUT_1[26846] = 32'b00000000000000001100001101000101;
assign LUT_1[26847] = 32'b00000000000000000101011111000001;
assign LUT_1[26848] = 32'b00000000000000001000010111000101;
assign LUT_1[26849] = 32'b00000000000000000001101001000001;
assign LUT_1[26850] = 32'b00000000000000000100000101010110;
assign LUT_1[26851] = 32'b11111111111111111101010111010010;
assign LUT_1[26852] = 32'b00000000000000010000010000011100;
assign LUT_1[26853] = 32'b00000000000000001001100010011000;
assign LUT_1[26854] = 32'b00000000000000001011111110101101;
assign LUT_1[26855] = 32'b00000000000000000101010000101001;
assign LUT_1[26856] = 32'b00000000000000000111100100111010;
assign LUT_1[26857] = 32'b00000000000000000000110110110110;
assign LUT_1[26858] = 32'b00000000000000000011010011001011;
assign LUT_1[26859] = 32'b11111111111111111100100101000111;
assign LUT_1[26860] = 32'b00000000000000001111011110010001;
assign LUT_1[26861] = 32'b00000000000000001000110000001101;
assign LUT_1[26862] = 32'b00000000000000001011001100100010;
assign LUT_1[26863] = 32'b00000000000000000100011110011110;
assign LUT_1[26864] = 32'b00000000000000001010010010100111;
assign LUT_1[26865] = 32'b00000000000000000011100100100011;
assign LUT_1[26866] = 32'b00000000000000000110000000111000;
assign LUT_1[26867] = 32'b11111111111111111111010010110100;
assign LUT_1[26868] = 32'b00000000000000010010001011111110;
assign LUT_1[26869] = 32'b00000000000000001011011101111010;
assign LUT_1[26870] = 32'b00000000000000001101111010001111;
assign LUT_1[26871] = 32'b00000000000000000111001100001011;
assign LUT_1[26872] = 32'b00000000000000001001100000011100;
assign LUT_1[26873] = 32'b00000000000000000010110010011000;
assign LUT_1[26874] = 32'b00000000000000000101001110101101;
assign LUT_1[26875] = 32'b11111111111111111110100000101001;
assign LUT_1[26876] = 32'b00000000000000010001011001110011;
assign LUT_1[26877] = 32'b00000000000000001010101011101111;
assign LUT_1[26878] = 32'b00000000000000001101001000000100;
assign LUT_1[26879] = 32'b00000000000000000110011010000000;
assign LUT_1[26880] = 32'b00000000000000000000010010100111;
assign LUT_1[26881] = 32'b11111111111111111001100100100011;
assign LUT_1[26882] = 32'b11111111111111111100000000111000;
assign LUT_1[26883] = 32'b11111111111111110101010010110100;
assign LUT_1[26884] = 32'b00000000000000001000001011111110;
assign LUT_1[26885] = 32'b00000000000000000001011101111010;
assign LUT_1[26886] = 32'b00000000000000000011111010001111;
assign LUT_1[26887] = 32'b11111111111111111101001100001011;
assign LUT_1[26888] = 32'b11111111111111111111100000011100;
assign LUT_1[26889] = 32'b11111111111111111000110010011000;
assign LUT_1[26890] = 32'b11111111111111111011001110101101;
assign LUT_1[26891] = 32'b11111111111111110100100000101001;
assign LUT_1[26892] = 32'b00000000000000000111011001110011;
assign LUT_1[26893] = 32'b00000000000000000000101011101111;
assign LUT_1[26894] = 32'b00000000000000000011001000000100;
assign LUT_1[26895] = 32'b11111111111111111100011010000000;
assign LUT_1[26896] = 32'b00000000000000000010001110001001;
assign LUT_1[26897] = 32'b11111111111111111011100000000101;
assign LUT_1[26898] = 32'b11111111111111111101111100011010;
assign LUT_1[26899] = 32'b11111111111111110111001110010110;
assign LUT_1[26900] = 32'b00000000000000001010000111100000;
assign LUT_1[26901] = 32'b00000000000000000011011001011100;
assign LUT_1[26902] = 32'b00000000000000000101110101110001;
assign LUT_1[26903] = 32'b11111111111111111111000111101101;
assign LUT_1[26904] = 32'b00000000000000000001011011111110;
assign LUT_1[26905] = 32'b11111111111111111010101101111010;
assign LUT_1[26906] = 32'b11111111111111111101001010001111;
assign LUT_1[26907] = 32'b11111111111111110110011100001011;
assign LUT_1[26908] = 32'b00000000000000001001010101010101;
assign LUT_1[26909] = 32'b00000000000000000010100111010001;
assign LUT_1[26910] = 32'b00000000000000000101000011100110;
assign LUT_1[26911] = 32'b11111111111111111110010101100010;
assign LUT_1[26912] = 32'b00000000000000000001001101100110;
assign LUT_1[26913] = 32'b11111111111111111010011111100010;
assign LUT_1[26914] = 32'b11111111111111111100111011110111;
assign LUT_1[26915] = 32'b11111111111111110110001101110011;
assign LUT_1[26916] = 32'b00000000000000001001000110111101;
assign LUT_1[26917] = 32'b00000000000000000010011000111001;
assign LUT_1[26918] = 32'b00000000000000000100110101001110;
assign LUT_1[26919] = 32'b11111111111111111110000111001010;
assign LUT_1[26920] = 32'b00000000000000000000011011011011;
assign LUT_1[26921] = 32'b11111111111111111001101101010111;
assign LUT_1[26922] = 32'b11111111111111111100001001101100;
assign LUT_1[26923] = 32'b11111111111111110101011011101000;
assign LUT_1[26924] = 32'b00000000000000001000010100110010;
assign LUT_1[26925] = 32'b00000000000000000001100110101110;
assign LUT_1[26926] = 32'b00000000000000000100000011000011;
assign LUT_1[26927] = 32'b11111111111111111101010100111111;
assign LUT_1[26928] = 32'b00000000000000000011001001001000;
assign LUT_1[26929] = 32'b11111111111111111100011011000100;
assign LUT_1[26930] = 32'b11111111111111111110110111011001;
assign LUT_1[26931] = 32'b11111111111111111000001001010101;
assign LUT_1[26932] = 32'b00000000000000001011000010011111;
assign LUT_1[26933] = 32'b00000000000000000100010100011011;
assign LUT_1[26934] = 32'b00000000000000000110110000110000;
assign LUT_1[26935] = 32'b00000000000000000000000010101100;
assign LUT_1[26936] = 32'b00000000000000000010010110111101;
assign LUT_1[26937] = 32'b11111111111111111011101000111001;
assign LUT_1[26938] = 32'b11111111111111111110000101001110;
assign LUT_1[26939] = 32'b11111111111111110111010111001010;
assign LUT_1[26940] = 32'b00000000000000001010010000010100;
assign LUT_1[26941] = 32'b00000000000000000011100010010000;
assign LUT_1[26942] = 32'b00000000000000000101111110100101;
assign LUT_1[26943] = 32'b11111111111111111111010000100001;
assign LUT_1[26944] = 32'b00000000000000000010010000001111;
assign LUT_1[26945] = 32'b11111111111111111011100010001011;
assign LUT_1[26946] = 32'b11111111111111111101111110100000;
assign LUT_1[26947] = 32'b11111111111111110111010000011100;
assign LUT_1[26948] = 32'b00000000000000001010001001100110;
assign LUT_1[26949] = 32'b00000000000000000011011011100010;
assign LUT_1[26950] = 32'b00000000000000000101110111110111;
assign LUT_1[26951] = 32'b11111111111111111111001001110011;
assign LUT_1[26952] = 32'b00000000000000000001011110000100;
assign LUT_1[26953] = 32'b11111111111111111010110000000000;
assign LUT_1[26954] = 32'b11111111111111111101001100010101;
assign LUT_1[26955] = 32'b11111111111111110110011110010001;
assign LUT_1[26956] = 32'b00000000000000001001010111011011;
assign LUT_1[26957] = 32'b00000000000000000010101001010111;
assign LUT_1[26958] = 32'b00000000000000000101000101101100;
assign LUT_1[26959] = 32'b11111111111111111110010111101000;
assign LUT_1[26960] = 32'b00000000000000000100001011110001;
assign LUT_1[26961] = 32'b11111111111111111101011101101101;
assign LUT_1[26962] = 32'b11111111111111111111111010000010;
assign LUT_1[26963] = 32'b11111111111111111001001011111110;
assign LUT_1[26964] = 32'b00000000000000001100000101001000;
assign LUT_1[26965] = 32'b00000000000000000101010111000100;
assign LUT_1[26966] = 32'b00000000000000000111110011011001;
assign LUT_1[26967] = 32'b00000000000000000001000101010101;
assign LUT_1[26968] = 32'b00000000000000000011011001100110;
assign LUT_1[26969] = 32'b11111111111111111100101011100010;
assign LUT_1[26970] = 32'b11111111111111111111000111110111;
assign LUT_1[26971] = 32'b11111111111111111000011001110011;
assign LUT_1[26972] = 32'b00000000000000001011010010111101;
assign LUT_1[26973] = 32'b00000000000000000100100100111001;
assign LUT_1[26974] = 32'b00000000000000000111000001001110;
assign LUT_1[26975] = 32'b00000000000000000000010011001010;
assign LUT_1[26976] = 32'b00000000000000000011001011001110;
assign LUT_1[26977] = 32'b11111111111111111100011101001010;
assign LUT_1[26978] = 32'b11111111111111111110111001011111;
assign LUT_1[26979] = 32'b11111111111111111000001011011011;
assign LUT_1[26980] = 32'b00000000000000001011000100100101;
assign LUT_1[26981] = 32'b00000000000000000100010110100001;
assign LUT_1[26982] = 32'b00000000000000000110110010110110;
assign LUT_1[26983] = 32'b00000000000000000000000100110010;
assign LUT_1[26984] = 32'b00000000000000000010011001000011;
assign LUT_1[26985] = 32'b11111111111111111011101010111111;
assign LUT_1[26986] = 32'b11111111111111111110000111010100;
assign LUT_1[26987] = 32'b11111111111111110111011001010000;
assign LUT_1[26988] = 32'b00000000000000001010010010011010;
assign LUT_1[26989] = 32'b00000000000000000011100100010110;
assign LUT_1[26990] = 32'b00000000000000000110000000101011;
assign LUT_1[26991] = 32'b11111111111111111111010010100111;
assign LUT_1[26992] = 32'b00000000000000000101000110110000;
assign LUT_1[26993] = 32'b11111111111111111110011000101100;
assign LUT_1[26994] = 32'b00000000000000000000110101000001;
assign LUT_1[26995] = 32'b11111111111111111010000110111101;
assign LUT_1[26996] = 32'b00000000000000001101000000000111;
assign LUT_1[26997] = 32'b00000000000000000110010010000011;
assign LUT_1[26998] = 32'b00000000000000001000101110011000;
assign LUT_1[26999] = 32'b00000000000000000010000000010100;
assign LUT_1[27000] = 32'b00000000000000000100010100100101;
assign LUT_1[27001] = 32'b11111111111111111101100110100001;
assign LUT_1[27002] = 32'b00000000000000000000000010110110;
assign LUT_1[27003] = 32'b11111111111111111001010100110010;
assign LUT_1[27004] = 32'b00000000000000001100001101111100;
assign LUT_1[27005] = 32'b00000000000000000101011111111000;
assign LUT_1[27006] = 32'b00000000000000000111111100001101;
assign LUT_1[27007] = 32'b00000000000000000001001110001001;
assign LUT_1[27008] = 32'b00000000000000000011010010101010;
assign LUT_1[27009] = 32'b11111111111111111100100100100110;
assign LUT_1[27010] = 32'b11111111111111111111000000111011;
assign LUT_1[27011] = 32'b11111111111111111000010010110111;
assign LUT_1[27012] = 32'b00000000000000001011001100000001;
assign LUT_1[27013] = 32'b00000000000000000100011101111101;
assign LUT_1[27014] = 32'b00000000000000000110111010010010;
assign LUT_1[27015] = 32'b00000000000000000000001100001110;
assign LUT_1[27016] = 32'b00000000000000000010100000011111;
assign LUT_1[27017] = 32'b11111111111111111011110010011011;
assign LUT_1[27018] = 32'b11111111111111111110001110110000;
assign LUT_1[27019] = 32'b11111111111111110111100000101100;
assign LUT_1[27020] = 32'b00000000000000001010011001110110;
assign LUT_1[27021] = 32'b00000000000000000011101011110010;
assign LUT_1[27022] = 32'b00000000000000000110001000000111;
assign LUT_1[27023] = 32'b11111111111111111111011010000011;
assign LUT_1[27024] = 32'b00000000000000000101001110001100;
assign LUT_1[27025] = 32'b11111111111111111110100000001000;
assign LUT_1[27026] = 32'b00000000000000000000111100011101;
assign LUT_1[27027] = 32'b11111111111111111010001110011001;
assign LUT_1[27028] = 32'b00000000000000001101000111100011;
assign LUT_1[27029] = 32'b00000000000000000110011001011111;
assign LUT_1[27030] = 32'b00000000000000001000110101110100;
assign LUT_1[27031] = 32'b00000000000000000010000111110000;
assign LUT_1[27032] = 32'b00000000000000000100011100000001;
assign LUT_1[27033] = 32'b11111111111111111101101101111101;
assign LUT_1[27034] = 32'b00000000000000000000001010010010;
assign LUT_1[27035] = 32'b11111111111111111001011100001110;
assign LUT_1[27036] = 32'b00000000000000001100010101011000;
assign LUT_1[27037] = 32'b00000000000000000101100111010100;
assign LUT_1[27038] = 32'b00000000000000001000000011101001;
assign LUT_1[27039] = 32'b00000000000000000001010101100101;
assign LUT_1[27040] = 32'b00000000000000000100001101101001;
assign LUT_1[27041] = 32'b11111111111111111101011111100101;
assign LUT_1[27042] = 32'b11111111111111111111111011111010;
assign LUT_1[27043] = 32'b11111111111111111001001101110110;
assign LUT_1[27044] = 32'b00000000000000001100000111000000;
assign LUT_1[27045] = 32'b00000000000000000101011000111100;
assign LUT_1[27046] = 32'b00000000000000000111110101010001;
assign LUT_1[27047] = 32'b00000000000000000001000111001101;
assign LUT_1[27048] = 32'b00000000000000000011011011011110;
assign LUT_1[27049] = 32'b11111111111111111100101101011010;
assign LUT_1[27050] = 32'b11111111111111111111001001101111;
assign LUT_1[27051] = 32'b11111111111111111000011011101011;
assign LUT_1[27052] = 32'b00000000000000001011010100110101;
assign LUT_1[27053] = 32'b00000000000000000100100110110001;
assign LUT_1[27054] = 32'b00000000000000000111000011000110;
assign LUT_1[27055] = 32'b00000000000000000000010101000010;
assign LUT_1[27056] = 32'b00000000000000000110001001001011;
assign LUT_1[27057] = 32'b11111111111111111111011011000111;
assign LUT_1[27058] = 32'b00000000000000000001110111011100;
assign LUT_1[27059] = 32'b11111111111111111011001001011000;
assign LUT_1[27060] = 32'b00000000000000001110000010100010;
assign LUT_1[27061] = 32'b00000000000000000111010100011110;
assign LUT_1[27062] = 32'b00000000000000001001110000110011;
assign LUT_1[27063] = 32'b00000000000000000011000010101111;
assign LUT_1[27064] = 32'b00000000000000000101010111000000;
assign LUT_1[27065] = 32'b11111111111111111110101000111100;
assign LUT_1[27066] = 32'b00000000000000000001000101010001;
assign LUT_1[27067] = 32'b11111111111111111010010111001101;
assign LUT_1[27068] = 32'b00000000000000001101010000010111;
assign LUT_1[27069] = 32'b00000000000000000110100010010011;
assign LUT_1[27070] = 32'b00000000000000001000111110101000;
assign LUT_1[27071] = 32'b00000000000000000010010000100100;
assign LUT_1[27072] = 32'b00000000000000000101010000010010;
assign LUT_1[27073] = 32'b11111111111111111110100010001110;
assign LUT_1[27074] = 32'b00000000000000000000111110100011;
assign LUT_1[27075] = 32'b11111111111111111010010000011111;
assign LUT_1[27076] = 32'b00000000000000001101001001101001;
assign LUT_1[27077] = 32'b00000000000000000110011011100101;
assign LUT_1[27078] = 32'b00000000000000001000110111111010;
assign LUT_1[27079] = 32'b00000000000000000010001001110110;
assign LUT_1[27080] = 32'b00000000000000000100011110000111;
assign LUT_1[27081] = 32'b11111111111111111101110000000011;
assign LUT_1[27082] = 32'b00000000000000000000001100011000;
assign LUT_1[27083] = 32'b11111111111111111001011110010100;
assign LUT_1[27084] = 32'b00000000000000001100010111011110;
assign LUT_1[27085] = 32'b00000000000000000101101001011010;
assign LUT_1[27086] = 32'b00000000000000001000000101101111;
assign LUT_1[27087] = 32'b00000000000000000001010111101011;
assign LUT_1[27088] = 32'b00000000000000000111001011110100;
assign LUT_1[27089] = 32'b00000000000000000000011101110000;
assign LUT_1[27090] = 32'b00000000000000000010111010000101;
assign LUT_1[27091] = 32'b11111111111111111100001100000001;
assign LUT_1[27092] = 32'b00000000000000001111000101001011;
assign LUT_1[27093] = 32'b00000000000000001000010111000111;
assign LUT_1[27094] = 32'b00000000000000001010110011011100;
assign LUT_1[27095] = 32'b00000000000000000100000101011000;
assign LUT_1[27096] = 32'b00000000000000000110011001101001;
assign LUT_1[27097] = 32'b11111111111111111111101011100101;
assign LUT_1[27098] = 32'b00000000000000000010000111111010;
assign LUT_1[27099] = 32'b11111111111111111011011001110110;
assign LUT_1[27100] = 32'b00000000000000001110010011000000;
assign LUT_1[27101] = 32'b00000000000000000111100100111100;
assign LUT_1[27102] = 32'b00000000000000001010000001010001;
assign LUT_1[27103] = 32'b00000000000000000011010011001101;
assign LUT_1[27104] = 32'b00000000000000000110001011010001;
assign LUT_1[27105] = 32'b11111111111111111111011101001101;
assign LUT_1[27106] = 32'b00000000000000000001111001100010;
assign LUT_1[27107] = 32'b11111111111111111011001011011110;
assign LUT_1[27108] = 32'b00000000000000001110000100101000;
assign LUT_1[27109] = 32'b00000000000000000111010110100100;
assign LUT_1[27110] = 32'b00000000000000001001110010111001;
assign LUT_1[27111] = 32'b00000000000000000011000100110101;
assign LUT_1[27112] = 32'b00000000000000000101011001000110;
assign LUT_1[27113] = 32'b11111111111111111110101011000010;
assign LUT_1[27114] = 32'b00000000000000000001000111010111;
assign LUT_1[27115] = 32'b11111111111111111010011001010011;
assign LUT_1[27116] = 32'b00000000000000001101010010011101;
assign LUT_1[27117] = 32'b00000000000000000110100100011001;
assign LUT_1[27118] = 32'b00000000000000001001000000101110;
assign LUT_1[27119] = 32'b00000000000000000010010010101010;
assign LUT_1[27120] = 32'b00000000000000001000000110110011;
assign LUT_1[27121] = 32'b00000000000000000001011000101111;
assign LUT_1[27122] = 32'b00000000000000000011110101000100;
assign LUT_1[27123] = 32'b11111111111111111101000111000000;
assign LUT_1[27124] = 32'b00000000000000010000000000001010;
assign LUT_1[27125] = 32'b00000000000000001001010010000110;
assign LUT_1[27126] = 32'b00000000000000001011101110011011;
assign LUT_1[27127] = 32'b00000000000000000101000000010111;
assign LUT_1[27128] = 32'b00000000000000000111010100101000;
assign LUT_1[27129] = 32'b00000000000000000000100110100100;
assign LUT_1[27130] = 32'b00000000000000000011000010111001;
assign LUT_1[27131] = 32'b11111111111111111100010100110101;
assign LUT_1[27132] = 32'b00000000000000001111001101111111;
assign LUT_1[27133] = 32'b00000000000000001000011111111011;
assign LUT_1[27134] = 32'b00000000000000001010111100010000;
assign LUT_1[27135] = 32'b00000000000000000100001110001100;
assign LUT_1[27136] = 32'b11111111111111111100001100111000;
assign LUT_1[27137] = 32'b11111111111111110101011110110100;
assign LUT_1[27138] = 32'b11111111111111110111111011001001;
assign LUT_1[27139] = 32'b11111111111111110001001101000101;
assign LUT_1[27140] = 32'b00000000000000000100000110001111;
assign LUT_1[27141] = 32'b11111111111111111101011000001011;
assign LUT_1[27142] = 32'b11111111111111111111110100100000;
assign LUT_1[27143] = 32'b11111111111111111001000110011100;
assign LUT_1[27144] = 32'b11111111111111111011011010101101;
assign LUT_1[27145] = 32'b11111111111111110100101100101001;
assign LUT_1[27146] = 32'b11111111111111110111001000111110;
assign LUT_1[27147] = 32'b11111111111111110000011010111010;
assign LUT_1[27148] = 32'b00000000000000000011010100000100;
assign LUT_1[27149] = 32'b11111111111111111100100110000000;
assign LUT_1[27150] = 32'b11111111111111111111000010010101;
assign LUT_1[27151] = 32'b11111111111111111000010100010001;
assign LUT_1[27152] = 32'b11111111111111111110001000011010;
assign LUT_1[27153] = 32'b11111111111111110111011010010110;
assign LUT_1[27154] = 32'b11111111111111111001110110101011;
assign LUT_1[27155] = 32'b11111111111111110011001000100111;
assign LUT_1[27156] = 32'b00000000000000000110000001110001;
assign LUT_1[27157] = 32'b11111111111111111111010011101101;
assign LUT_1[27158] = 32'b00000000000000000001110000000010;
assign LUT_1[27159] = 32'b11111111111111111011000001111110;
assign LUT_1[27160] = 32'b11111111111111111101010110001111;
assign LUT_1[27161] = 32'b11111111111111110110101000001011;
assign LUT_1[27162] = 32'b11111111111111111001000100100000;
assign LUT_1[27163] = 32'b11111111111111110010010110011100;
assign LUT_1[27164] = 32'b00000000000000000101001111100110;
assign LUT_1[27165] = 32'b11111111111111111110100001100010;
assign LUT_1[27166] = 32'b00000000000000000000111101110111;
assign LUT_1[27167] = 32'b11111111111111111010001111110011;
assign LUT_1[27168] = 32'b11111111111111111101000111110111;
assign LUT_1[27169] = 32'b11111111111111110110011001110011;
assign LUT_1[27170] = 32'b11111111111111111000110110001000;
assign LUT_1[27171] = 32'b11111111111111110010001000000100;
assign LUT_1[27172] = 32'b00000000000000000101000001001110;
assign LUT_1[27173] = 32'b11111111111111111110010011001010;
assign LUT_1[27174] = 32'b00000000000000000000101111011111;
assign LUT_1[27175] = 32'b11111111111111111010000001011011;
assign LUT_1[27176] = 32'b11111111111111111100010101101100;
assign LUT_1[27177] = 32'b11111111111111110101100111101000;
assign LUT_1[27178] = 32'b11111111111111111000000011111101;
assign LUT_1[27179] = 32'b11111111111111110001010101111001;
assign LUT_1[27180] = 32'b00000000000000000100001111000011;
assign LUT_1[27181] = 32'b11111111111111111101100000111111;
assign LUT_1[27182] = 32'b11111111111111111111111101010100;
assign LUT_1[27183] = 32'b11111111111111111001001111010000;
assign LUT_1[27184] = 32'b11111111111111111111000011011001;
assign LUT_1[27185] = 32'b11111111111111111000010101010101;
assign LUT_1[27186] = 32'b11111111111111111010110001101010;
assign LUT_1[27187] = 32'b11111111111111110100000011100110;
assign LUT_1[27188] = 32'b00000000000000000110111100110000;
assign LUT_1[27189] = 32'b00000000000000000000001110101100;
assign LUT_1[27190] = 32'b00000000000000000010101011000001;
assign LUT_1[27191] = 32'b11111111111111111011111100111101;
assign LUT_1[27192] = 32'b11111111111111111110010001001110;
assign LUT_1[27193] = 32'b11111111111111110111100011001010;
assign LUT_1[27194] = 32'b11111111111111111001111111011111;
assign LUT_1[27195] = 32'b11111111111111110011010001011011;
assign LUT_1[27196] = 32'b00000000000000000110001010100101;
assign LUT_1[27197] = 32'b11111111111111111111011100100001;
assign LUT_1[27198] = 32'b00000000000000000001111000110110;
assign LUT_1[27199] = 32'b11111111111111111011001010110010;
assign LUT_1[27200] = 32'b11111111111111111110001010100000;
assign LUT_1[27201] = 32'b11111111111111110111011100011100;
assign LUT_1[27202] = 32'b11111111111111111001111000110001;
assign LUT_1[27203] = 32'b11111111111111110011001010101101;
assign LUT_1[27204] = 32'b00000000000000000110000011110111;
assign LUT_1[27205] = 32'b11111111111111111111010101110011;
assign LUT_1[27206] = 32'b00000000000000000001110010001000;
assign LUT_1[27207] = 32'b11111111111111111011000100000100;
assign LUT_1[27208] = 32'b11111111111111111101011000010101;
assign LUT_1[27209] = 32'b11111111111111110110101010010001;
assign LUT_1[27210] = 32'b11111111111111111001000110100110;
assign LUT_1[27211] = 32'b11111111111111110010011000100010;
assign LUT_1[27212] = 32'b00000000000000000101010001101100;
assign LUT_1[27213] = 32'b11111111111111111110100011101000;
assign LUT_1[27214] = 32'b00000000000000000000111111111101;
assign LUT_1[27215] = 32'b11111111111111111010010001111001;
assign LUT_1[27216] = 32'b00000000000000000000000110000010;
assign LUT_1[27217] = 32'b11111111111111111001010111111110;
assign LUT_1[27218] = 32'b11111111111111111011110100010011;
assign LUT_1[27219] = 32'b11111111111111110101000110001111;
assign LUT_1[27220] = 32'b00000000000000000111111111011001;
assign LUT_1[27221] = 32'b00000000000000000001010001010101;
assign LUT_1[27222] = 32'b00000000000000000011101101101010;
assign LUT_1[27223] = 32'b11111111111111111100111111100110;
assign LUT_1[27224] = 32'b11111111111111111111010011110111;
assign LUT_1[27225] = 32'b11111111111111111000100101110011;
assign LUT_1[27226] = 32'b11111111111111111011000010001000;
assign LUT_1[27227] = 32'b11111111111111110100010100000100;
assign LUT_1[27228] = 32'b00000000000000000111001101001110;
assign LUT_1[27229] = 32'b00000000000000000000011111001010;
assign LUT_1[27230] = 32'b00000000000000000010111011011111;
assign LUT_1[27231] = 32'b11111111111111111100001101011011;
assign LUT_1[27232] = 32'b11111111111111111111000101011111;
assign LUT_1[27233] = 32'b11111111111111111000010111011011;
assign LUT_1[27234] = 32'b11111111111111111010110011110000;
assign LUT_1[27235] = 32'b11111111111111110100000101101100;
assign LUT_1[27236] = 32'b00000000000000000110111110110110;
assign LUT_1[27237] = 32'b00000000000000000000010000110010;
assign LUT_1[27238] = 32'b00000000000000000010101101000111;
assign LUT_1[27239] = 32'b11111111111111111011111111000011;
assign LUT_1[27240] = 32'b11111111111111111110010011010100;
assign LUT_1[27241] = 32'b11111111111111110111100101010000;
assign LUT_1[27242] = 32'b11111111111111111010000001100101;
assign LUT_1[27243] = 32'b11111111111111110011010011100001;
assign LUT_1[27244] = 32'b00000000000000000110001100101011;
assign LUT_1[27245] = 32'b11111111111111111111011110100111;
assign LUT_1[27246] = 32'b00000000000000000001111010111100;
assign LUT_1[27247] = 32'b11111111111111111011001100111000;
assign LUT_1[27248] = 32'b00000000000000000001000001000001;
assign LUT_1[27249] = 32'b11111111111111111010010010111101;
assign LUT_1[27250] = 32'b11111111111111111100101111010010;
assign LUT_1[27251] = 32'b11111111111111110110000001001110;
assign LUT_1[27252] = 32'b00000000000000001000111010011000;
assign LUT_1[27253] = 32'b00000000000000000010001100010100;
assign LUT_1[27254] = 32'b00000000000000000100101000101001;
assign LUT_1[27255] = 32'b11111111111111111101111010100101;
assign LUT_1[27256] = 32'b00000000000000000000001110110110;
assign LUT_1[27257] = 32'b11111111111111111001100000110010;
assign LUT_1[27258] = 32'b11111111111111111011111101000111;
assign LUT_1[27259] = 32'b11111111111111110101001111000011;
assign LUT_1[27260] = 32'b00000000000000001000001000001101;
assign LUT_1[27261] = 32'b00000000000000000001011010001001;
assign LUT_1[27262] = 32'b00000000000000000011110110011110;
assign LUT_1[27263] = 32'b11111111111111111101001000011010;
assign LUT_1[27264] = 32'b11111111111111111111001100111011;
assign LUT_1[27265] = 32'b11111111111111111000011110110111;
assign LUT_1[27266] = 32'b11111111111111111010111011001100;
assign LUT_1[27267] = 32'b11111111111111110100001101001000;
assign LUT_1[27268] = 32'b00000000000000000111000110010010;
assign LUT_1[27269] = 32'b00000000000000000000011000001110;
assign LUT_1[27270] = 32'b00000000000000000010110100100011;
assign LUT_1[27271] = 32'b11111111111111111100000110011111;
assign LUT_1[27272] = 32'b11111111111111111110011010110000;
assign LUT_1[27273] = 32'b11111111111111110111101100101100;
assign LUT_1[27274] = 32'b11111111111111111010001001000001;
assign LUT_1[27275] = 32'b11111111111111110011011010111101;
assign LUT_1[27276] = 32'b00000000000000000110010100000111;
assign LUT_1[27277] = 32'b11111111111111111111100110000011;
assign LUT_1[27278] = 32'b00000000000000000010000010011000;
assign LUT_1[27279] = 32'b11111111111111111011010100010100;
assign LUT_1[27280] = 32'b00000000000000000001001000011101;
assign LUT_1[27281] = 32'b11111111111111111010011010011001;
assign LUT_1[27282] = 32'b11111111111111111100110110101110;
assign LUT_1[27283] = 32'b11111111111111110110001000101010;
assign LUT_1[27284] = 32'b00000000000000001001000001110100;
assign LUT_1[27285] = 32'b00000000000000000010010011110000;
assign LUT_1[27286] = 32'b00000000000000000100110000000101;
assign LUT_1[27287] = 32'b11111111111111111110000010000001;
assign LUT_1[27288] = 32'b00000000000000000000010110010010;
assign LUT_1[27289] = 32'b11111111111111111001101000001110;
assign LUT_1[27290] = 32'b11111111111111111100000100100011;
assign LUT_1[27291] = 32'b11111111111111110101010110011111;
assign LUT_1[27292] = 32'b00000000000000001000001111101001;
assign LUT_1[27293] = 32'b00000000000000000001100001100101;
assign LUT_1[27294] = 32'b00000000000000000011111101111010;
assign LUT_1[27295] = 32'b11111111111111111101001111110110;
assign LUT_1[27296] = 32'b00000000000000000000000111111010;
assign LUT_1[27297] = 32'b11111111111111111001011001110110;
assign LUT_1[27298] = 32'b11111111111111111011110110001011;
assign LUT_1[27299] = 32'b11111111111111110101001000000111;
assign LUT_1[27300] = 32'b00000000000000001000000001010001;
assign LUT_1[27301] = 32'b00000000000000000001010011001101;
assign LUT_1[27302] = 32'b00000000000000000011101111100010;
assign LUT_1[27303] = 32'b11111111111111111101000001011110;
assign LUT_1[27304] = 32'b11111111111111111111010101101111;
assign LUT_1[27305] = 32'b11111111111111111000100111101011;
assign LUT_1[27306] = 32'b11111111111111111011000100000000;
assign LUT_1[27307] = 32'b11111111111111110100010101111100;
assign LUT_1[27308] = 32'b00000000000000000111001111000110;
assign LUT_1[27309] = 32'b00000000000000000000100001000010;
assign LUT_1[27310] = 32'b00000000000000000010111101010111;
assign LUT_1[27311] = 32'b11111111111111111100001111010011;
assign LUT_1[27312] = 32'b00000000000000000010000011011100;
assign LUT_1[27313] = 32'b11111111111111111011010101011000;
assign LUT_1[27314] = 32'b11111111111111111101110001101101;
assign LUT_1[27315] = 32'b11111111111111110111000011101001;
assign LUT_1[27316] = 32'b00000000000000001001111100110011;
assign LUT_1[27317] = 32'b00000000000000000011001110101111;
assign LUT_1[27318] = 32'b00000000000000000101101011000100;
assign LUT_1[27319] = 32'b11111111111111111110111101000000;
assign LUT_1[27320] = 32'b00000000000000000001010001010001;
assign LUT_1[27321] = 32'b11111111111111111010100011001101;
assign LUT_1[27322] = 32'b11111111111111111100111111100010;
assign LUT_1[27323] = 32'b11111111111111110110010001011110;
assign LUT_1[27324] = 32'b00000000000000001001001010101000;
assign LUT_1[27325] = 32'b00000000000000000010011100100100;
assign LUT_1[27326] = 32'b00000000000000000100111000111001;
assign LUT_1[27327] = 32'b11111111111111111110001010110101;
assign LUT_1[27328] = 32'b00000000000000000001001010100011;
assign LUT_1[27329] = 32'b11111111111111111010011100011111;
assign LUT_1[27330] = 32'b11111111111111111100111000110100;
assign LUT_1[27331] = 32'b11111111111111110110001010110000;
assign LUT_1[27332] = 32'b00000000000000001001000011111010;
assign LUT_1[27333] = 32'b00000000000000000010010101110110;
assign LUT_1[27334] = 32'b00000000000000000100110010001011;
assign LUT_1[27335] = 32'b11111111111111111110000100000111;
assign LUT_1[27336] = 32'b00000000000000000000011000011000;
assign LUT_1[27337] = 32'b11111111111111111001101010010100;
assign LUT_1[27338] = 32'b11111111111111111100000110101001;
assign LUT_1[27339] = 32'b11111111111111110101011000100101;
assign LUT_1[27340] = 32'b00000000000000001000010001101111;
assign LUT_1[27341] = 32'b00000000000000000001100011101011;
assign LUT_1[27342] = 32'b00000000000000000100000000000000;
assign LUT_1[27343] = 32'b11111111111111111101010001111100;
assign LUT_1[27344] = 32'b00000000000000000011000110000101;
assign LUT_1[27345] = 32'b11111111111111111100011000000001;
assign LUT_1[27346] = 32'b11111111111111111110110100010110;
assign LUT_1[27347] = 32'b11111111111111111000000110010010;
assign LUT_1[27348] = 32'b00000000000000001010111111011100;
assign LUT_1[27349] = 32'b00000000000000000100010001011000;
assign LUT_1[27350] = 32'b00000000000000000110101101101101;
assign LUT_1[27351] = 32'b11111111111111111111111111101001;
assign LUT_1[27352] = 32'b00000000000000000010010011111010;
assign LUT_1[27353] = 32'b11111111111111111011100101110110;
assign LUT_1[27354] = 32'b11111111111111111110000010001011;
assign LUT_1[27355] = 32'b11111111111111110111010100000111;
assign LUT_1[27356] = 32'b00000000000000001010001101010001;
assign LUT_1[27357] = 32'b00000000000000000011011111001101;
assign LUT_1[27358] = 32'b00000000000000000101111011100010;
assign LUT_1[27359] = 32'b11111111111111111111001101011110;
assign LUT_1[27360] = 32'b00000000000000000010000101100010;
assign LUT_1[27361] = 32'b11111111111111111011010111011110;
assign LUT_1[27362] = 32'b11111111111111111101110011110011;
assign LUT_1[27363] = 32'b11111111111111110111000101101111;
assign LUT_1[27364] = 32'b00000000000000001001111110111001;
assign LUT_1[27365] = 32'b00000000000000000011010000110101;
assign LUT_1[27366] = 32'b00000000000000000101101101001010;
assign LUT_1[27367] = 32'b11111111111111111110111111000110;
assign LUT_1[27368] = 32'b00000000000000000001010011010111;
assign LUT_1[27369] = 32'b11111111111111111010100101010011;
assign LUT_1[27370] = 32'b11111111111111111101000001101000;
assign LUT_1[27371] = 32'b11111111111111110110010011100100;
assign LUT_1[27372] = 32'b00000000000000001001001100101110;
assign LUT_1[27373] = 32'b00000000000000000010011110101010;
assign LUT_1[27374] = 32'b00000000000000000100111010111111;
assign LUT_1[27375] = 32'b11111111111111111110001100111011;
assign LUT_1[27376] = 32'b00000000000000000100000001000100;
assign LUT_1[27377] = 32'b11111111111111111101010011000000;
assign LUT_1[27378] = 32'b11111111111111111111101111010101;
assign LUT_1[27379] = 32'b11111111111111111001000001010001;
assign LUT_1[27380] = 32'b00000000000000001011111010011011;
assign LUT_1[27381] = 32'b00000000000000000101001100010111;
assign LUT_1[27382] = 32'b00000000000000000111101000101100;
assign LUT_1[27383] = 32'b00000000000000000000111010101000;
assign LUT_1[27384] = 32'b00000000000000000011001110111001;
assign LUT_1[27385] = 32'b11111111111111111100100000110101;
assign LUT_1[27386] = 32'b11111111111111111110111101001010;
assign LUT_1[27387] = 32'b11111111111111111000001111000110;
assign LUT_1[27388] = 32'b00000000000000001011001000010000;
assign LUT_1[27389] = 32'b00000000000000000100011010001100;
assign LUT_1[27390] = 32'b00000000000000000110110110100001;
assign LUT_1[27391] = 32'b00000000000000000000001000011101;
assign LUT_1[27392] = 32'b11111111111111111010000001000100;
assign LUT_1[27393] = 32'b11111111111111110011010011000000;
assign LUT_1[27394] = 32'b11111111111111110101101111010101;
assign LUT_1[27395] = 32'b11111111111111101111000001010001;
assign LUT_1[27396] = 32'b00000000000000000001111010011011;
assign LUT_1[27397] = 32'b11111111111111111011001100010111;
assign LUT_1[27398] = 32'b11111111111111111101101000101100;
assign LUT_1[27399] = 32'b11111111111111110110111010101000;
assign LUT_1[27400] = 32'b11111111111111111001001110111001;
assign LUT_1[27401] = 32'b11111111111111110010100000110101;
assign LUT_1[27402] = 32'b11111111111111110100111101001010;
assign LUT_1[27403] = 32'b11111111111111101110001111000110;
assign LUT_1[27404] = 32'b00000000000000000001001000010000;
assign LUT_1[27405] = 32'b11111111111111111010011010001100;
assign LUT_1[27406] = 32'b11111111111111111100110110100001;
assign LUT_1[27407] = 32'b11111111111111110110001000011101;
assign LUT_1[27408] = 32'b11111111111111111011111100100110;
assign LUT_1[27409] = 32'b11111111111111110101001110100010;
assign LUT_1[27410] = 32'b11111111111111110111101010110111;
assign LUT_1[27411] = 32'b11111111111111110000111100110011;
assign LUT_1[27412] = 32'b00000000000000000011110101111101;
assign LUT_1[27413] = 32'b11111111111111111101000111111001;
assign LUT_1[27414] = 32'b11111111111111111111100100001110;
assign LUT_1[27415] = 32'b11111111111111111000110110001010;
assign LUT_1[27416] = 32'b11111111111111111011001010011011;
assign LUT_1[27417] = 32'b11111111111111110100011100010111;
assign LUT_1[27418] = 32'b11111111111111110110111000101100;
assign LUT_1[27419] = 32'b11111111111111110000001010101000;
assign LUT_1[27420] = 32'b00000000000000000011000011110010;
assign LUT_1[27421] = 32'b11111111111111111100010101101110;
assign LUT_1[27422] = 32'b11111111111111111110110010000011;
assign LUT_1[27423] = 32'b11111111111111111000000011111111;
assign LUT_1[27424] = 32'b11111111111111111010111100000011;
assign LUT_1[27425] = 32'b11111111111111110100001101111111;
assign LUT_1[27426] = 32'b11111111111111110110101010010100;
assign LUT_1[27427] = 32'b11111111111111101111111100010000;
assign LUT_1[27428] = 32'b00000000000000000010110101011010;
assign LUT_1[27429] = 32'b11111111111111111100000111010110;
assign LUT_1[27430] = 32'b11111111111111111110100011101011;
assign LUT_1[27431] = 32'b11111111111111110111110101100111;
assign LUT_1[27432] = 32'b11111111111111111010001001111000;
assign LUT_1[27433] = 32'b11111111111111110011011011110100;
assign LUT_1[27434] = 32'b11111111111111110101111000001001;
assign LUT_1[27435] = 32'b11111111111111101111001010000101;
assign LUT_1[27436] = 32'b00000000000000000010000011001111;
assign LUT_1[27437] = 32'b11111111111111111011010101001011;
assign LUT_1[27438] = 32'b11111111111111111101110001100000;
assign LUT_1[27439] = 32'b11111111111111110111000011011100;
assign LUT_1[27440] = 32'b11111111111111111100110111100101;
assign LUT_1[27441] = 32'b11111111111111110110001001100001;
assign LUT_1[27442] = 32'b11111111111111111000100101110110;
assign LUT_1[27443] = 32'b11111111111111110001110111110010;
assign LUT_1[27444] = 32'b00000000000000000100110000111100;
assign LUT_1[27445] = 32'b11111111111111111110000010111000;
assign LUT_1[27446] = 32'b00000000000000000000011111001101;
assign LUT_1[27447] = 32'b11111111111111111001110001001001;
assign LUT_1[27448] = 32'b11111111111111111100000101011010;
assign LUT_1[27449] = 32'b11111111111111110101010111010110;
assign LUT_1[27450] = 32'b11111111111111110111110011101011;
assign LUT_1[27451] = 32'b11111111111111110001000101100111;
assign LUT_1[27452] = 32'b00000000000000000011111110110001;
assign LUT_1[27453] = 32'b11111111111111111101010000101101;
assign LUT_1[27454] = 32'b11111111111111111111101101000010;
assign LUT_1[27455] = 32'b11111111111111111000111110111110;
assign LUT_1[27456] = 32'b11111111111111111011111110101100;
assign LUT_1[27457] = 32'b11111111111111110101010000101000;
assign LUT_1[27458] = 32'b11111111111111110111101100111101;
assign LUT_1[27459] = 32'b11111111111111110000111110111001;
assign LUT_1[27460] = 32'b00000000000000000011111000000011;
assign LUT_1[27461] = 32'b11111111111111111101001001111111;
assign LUT_1[27462] = 32'b11111111111111111111100110010100;
assign LUT_1[27463] = 32'b11111111111111111000111000010000;
assign LUT_1[27464] = 32'b11111111111111111011001100100001;
assign LUT_1[27465] = 32'b11111111111111110100011110011101;
assign LUT_1[27466] = 32'b11111111111111110110111010110010;
assign LUT_1[27467] = 32'b11111111111111110000001100101110;
assign LUT_1[27468] = 32'b00000000000000000011000101111000;
assign LUT_1[27469] = 32'b11111111111111111100010111110100;
assign LUT_1[27470] = 32'b11111111111111111110110100001001;
assign LUT_1[27471] = 32'b11111111111111111000000110000101;
assign LUT_1[27472] = 32'b11111111111111111101111010001110;
assign LUT_1[27473] = 32'b11111111111111110111001100001010;
assign LUT_1[27474] = 32'b11111111111111111001101000011111;
assign LUT_1[27475] = 32'b11111111111111110010111010011011;
assign LUT_1[27476] = 32'b00000000000000000101110011100101;
assign LUT_1[27477] = 32'b11111111111111111111000101100001;
assign LUT_1[27478] = 32'b00000000000000000001100001110110;
assign LUT_1[27479] = 32'b11111111111111111010110011110010;
assign LUT_1[27480] = 32'b11111111111111111101001000000011;
assign LUT_1[27481] = 32'b11111111111111110110011001111111;
assign LUT_1[27482] = 32'b11111111111111111000110110010100;
assign LUT_1[27483] = 32'b11111111111111110010001000010000;
assign LUT_1[27484] = 32'b00000000000000000101000001011010;
assign LUT_1[27485] = 32'b11111111111111111110010011010110;
assign LUT_1[27486] = 32'b00000000000000000000101111101011;
assign LUT_1[27487] = 32'b11111111111111111010000001100111;
assign LUT_1[27488] = 32'b11111111111111111100111001101011;
assign LUT_1[27489] = 32'b11111111111111110110001011100111;
assign LUT_1[27490] = 32'b11111111111111111000100111111100;
assign LUT_1[27491] = 32'b11111111111111110001111001111000;
assign LUT_1[27492] = 32'b00000000000000000100110011000010;
assign LUT_1[27493] = 32'b11111111111111111110000100111110;
assign LUT_1[27494] = 32'b00000000000000000000100001010011;
assign LUT_1[27495] = 32'b11111111111111111001110011001111;
assign LUT_1[27496] = 32'b11111111111111111100000111100000;
assign LUT_1[27497] = 32'b11111111111111110101011001011100;
assign LUT_1[27498] = 32'b11111111111111110111110101110001;
assign LUT_1[27499] = 32'b11111111111111110001000111101101;
assign LUT_1[27500] = 32'b00000000000000000100000000110111;
assign LUT_1[27501] = 32'b11111111111111111101010010110011;
assign LUT_1[27502] = 32'b11111111111111111111101111001000;
assign LUT_1[27503] = 32'b11111111111111111001000001000100;
assign LUT_1[27504] = 32'b11111111111111111110110101001101;
assign LUT_1[27505] = 32'b11111111111111111000000111001001;
assign LUT_1[27506] = 32'b11111111111111111010100011011110;
assign LUT_1[27507] = 32'b11111111111111110011110101011010;
assign LUT_1[27508] = 32'b00000000000000000110101110100100;
assign LUT_1[27509] = 32'b00000000000000000000000000100000;
assign LUT_1[27510] = 32'b00000000000000000010011100110101;
assign LUT_1[27511] = 32'b11111111111111111011101110110001;
assign LUT_1[27512] = 32'b11111111111111111110000011000010;
assign LUT_1[27513] = 32'b11111111111111110111010100111110;
assign LUT_1[27514] = 32'b11111111111111111001110001010011;
assign LUT_1[27515] = 32'b11111111111111110011000011001111;
assign LUT_1[27516] = 32'b00000000000000000101111100011001;
assign LUT_1[27517] = 32'b11111111111111111111001110010101;
assign LUT_1[27518] = 32'b00000000000000000001101010101010;
assign LUT_1[27519] = 32'b11111111111111111010111100100110;
assign LUT_1[27520] = 32'b11111111111111111101000001000111;
assign LUT_1[27521] = 32'b11111111111111110110010011000011;
assign LUT_1[27522] = 32'b11111111111111111000101111011000;
assign LUT_1[27523] = 32'b11111111111111110010000001010100;
assign LUT_1[27524] = 32'b00000000000000000100111010011110;
assign LUT_1[27525] = 32'b11111111111111111110001100011010;
assign LUT_1[27526] = 32'b00000000000000000000101000101111;
assign LUT_1[27527] = 32'b11111111111111111001111010101011;
assign LUT_1[27528] = 32'b11111111111111111100001110111100;
assign LUT_1[27529] = 32'b11111111111111110101100000111000;
assign LUT_1[27530] = 32'b11111111111111110111111101001101;
assign LUT_1[27531] = 32'b11111111111111110001001111001001;
assign LUT_1[27532] = 32'b00000000000000000100001000010011;
assign LUT_1[27533] = 32'b11111111111111111101011010001111;
assign LUT_1[27534] = 32'b11111111111111111111110110100100;
assign LUT_1[27535] = 32'b11111111111111111001001000100000;
assign LUT_1[27536] = 32'b11111111111111111110111100101001;
assign LUT_1[27537] = 32'b11111111111111111000001110100101;
assign LUT_1[27538] = 32'b11111111111111111010101010111010;
assign LUT_1[27539] = 32'b11111111111111110011111100110110;
assign LUT_1[27540] = 32'b00000000000000000110110110000000;
assign LUT_1[27541] = 32'b00000000000000000000000111111100;
assign LUT_1[27542] = 32'b00000000000000000010100100010001;
assign LUT_1[27543] = 32'b11111111111111111011110110001101;
assign LUT_1[27544] = 32'b11111111111111111110001010011110;
assign LUT_1[27545] = 32'b11111111111111110111011100011010;
assign LUT_1[27546] = 32'b11111111111111111001111000101111;
assign LUT_1[27547] = 32'b11111111111111110011001010101011;
assign LUT_1[27548] = 32'b00000000000000000110000011110101;
assign LUT_1[27549] = 32'b11111111111111111111010101110001;
assign LUT_1[27550] = 32'b00000000000000000001110010000110;
assign LUT_1[27551] = 32'b11111111111111111011000100000010;
assign LUT_1[27552] = 32'b11111111111111111101111100000110;
assign LUT_1[27553] = 32'b11111111111111110111001110000010;
assign LUT_1[27554] = 32'b11111111111111111001101010010111;
assign LUT_1[27555] = 32'b11111111111111110010111100010011;
assign LUT_1[27556] = 32'b00000000000000000101110101011101;
assign LUT_1[27557] = 32'b11111111111111111111000111011001;
assign LUT_1[27558] = 32'b00000000000000000001100011101110;
assign LUT_1[27559] = 32'b11111111111111111010110101101010;
assign LUT_1[27560] = 32'b11111111111111111101001001111011;
assign LUT_1[27561] = 32'b11111111111111110110011011110111;
assign LUT_1[27562] = 32'b11111111111111111000111000001100;
assign LUT_1[27563] = 32'b11111111111111110010001010001000;
assign LUT_1[27564] = 32'b00000000000000000101000011010010;
assign LUT_1[27565] = 32'b11111111111111111110010101001110;
assign LUT_1[27566] = 32'b00000000000000000000110001100011;
assign LUT_1[27567] = 32'b11111111111111111010000011011111;
assign LUT_1[27568] = 32'b11111111111111111111110111101000;
assign LUT_1[27569] = 32'b11111111111111111001001001100100;
assign LUT_1[27570] = 32'b11111111111111111011100101111001;
assign LUT_1[27571] = 32'b11111111111111110100110111110101;
assign LUT_1[27572] = 32'b00000000000000000111110000111111;
assign LUT_1[27573] = 32'b00000000000000000001000010111011;
assign LUT_1[27574] = 32'b00000000000000000011011111010000;
assign LUT_1[27575] = 32'b11111111111111111100110001001100;
assign LUT_1[27576] = 32'b11111111111111111111000101011101;
assign LUT_1[27577] = 32'b11111111111111111000010111011001;
assign LUT_1[27578] = 32'b11111111111111111010110011101110;
assign LUT_1[27579] = 32'b11111111111111110100000101101010;
assign LUT_1[27580] = 32'b00000000000000000110111110110100;
assign LUT_1[27581] = 32'b00000000000000000000010000110000;
assign LUT_1[27582] = 32'b00000000000000000010101101000101;
assign LUT_1[27583] = 32'b11111111111111111011111111000001;
assign LUT_1[27584] = 32'b11111111111111111110111110101111;
assign LUT_1[27585] = 32'b11111111111111111000010000101011;
assign LUT_1[27586] = 32'b11111111111111111010101101000000;
assign LUT_1[27587] = 32'b11111111111111110011111110111100;
assign LUT_1[27588] = 32'b00000000000000000110111000000110;
assign LUT_1[27589] = 32'b00000000000000000000001010000010;
assign LUT_1[27590] = 32'b00000000000000000010100110010111;
assign LUT_1[27591] = 32'b11111111111111111011111000010011;
assign LUT_1[27592] = 32'b11111111111111111110001100100100;
assign LUT_1[27593] = 32'b11111111111111110111011110100000;
assign LUT_1[27594] = 32'b11111111111111111001111010110101;
assign LUT_1[27595] = 32'b11111111111111110011001100110001;
assign LUT_1[27596] = 32'b00000000000000000110000101111011;
assign LUT_1[27597] = 32'b11111111111111111111010111110111;
assign LUT_1[27598] = 32'b00000000000000000001110100001100;
assign LUT_1[27599] = 32'b11111111111111111011000110001000;
assign LUT_1[27600] = 32'b00000000000000000000111010010001;
assign LUT_1[27601] = 32'b11111111111111111010001100001101;
assign LUT_1[27602] = 32'b11111111111111111100101000100010;
assign LUT_1[27603] = 32'b11111111111111110101111010011110;
assign LUT_1[27604] = 32'b00000000000000001000110011101000;
assign LUT_1[27605] = 32'b00000000000000000010000101100100;
assign LUT_1[27606] = 32'b00000000000000000100100001111001;
assign LUT_1[27607] = 32'b11111111111111111101110011110101;
assign LUT_1[27608] = 32'b00000000000000000000001000000110;
assign LUT_1[27609] = 32'b11111111111111111001011010000010;
assign LUT_1[27610] = 32'b11111111111111111011110110010111;
assign LUT_1[27611] = 32'b11111111111111110101001000010011;
assign LUT_1[27612] = 32'b00000000000000001000000001011101;
assign LUT_1[27613] = 32'b00000000000000000001010011011001;
assign LUT_1[27614] = 32'b00000000000000000011101111101110;
assign LUT_1[27615] = 32'b11111111111111111101000001101010;
assign LUT_1[27616] = 32'b11111111111111111111111001101110;
assign LUT_1[27617] = 32'b11111111111111111001001011101010;
assign LUT_1[27618] = 32'b11111111111111111011100111111111;
assign LUT_1[27619] = 32'b11111111111111110100111001111011;
assign LUT_1[27620] = 32'b00000000000000000111110011000101;
assign LUT_1[27621] = 32'b00000000000000000001000101000001;
assign LUT_1[27622] = 32'b00000000000000000011100001010110;
assign LUT_1[27623] = 32'b11111111111111111100110011010010;
assign LUT_1[27624] = 32'b11111111111111111111000111100011;
assign LUT_1[27625] = 32'b11111111111111111000011001011111;
assign LUT_1[27626] = 32'b11111111111111111010110101110100;
assign LUT_1[27627] = 32'b11111111111111110100000111110000;
assign LUT_1[27628] = 32'b00000000000000000111000000111010;
assign LUT_1[27629] = 32'b00000000000000000000010010110110;
assign LUT_1[27630] = 32'b00000000000000000010101111001011;
assign LUT_1[27631] = 32'b11111111111111111100000001000111;
assign LUT_1[27632] = 32'b00000000000000000001110101010000;
assign LUT_1[27633] = 32'b11111111111111111011000111001100;
assign LUT_1[27634] = 32'b11111111111111111101100011100001;
assign LUT_1[27635] = 32'b11111111111111110110110101011101;
assign LUT_1[27636] = 32'b00000000000000001001101110100111;
assign LUT_1[27637] = 32'b00000000000000000011000000100011;
assign LUT_1[27638] = 32'b00000000000000000101011100111000;
assign LUT_1[27639] = 32'b11111111111111111110101110110100;
assign LUT_1[27640] = 32'b00000000000000000001000011000101;
assign LUT_1[27641] = 32'b11111111111111111010010101000001;
assign LUT_1[27642] = 32'b11111111111111111100110001010110;
assign LUT_1[27643] = 32'b11111111111111110110000011010010;
assign LUT_1[27644] = 32'b00000000000000001000111100011100;
assign LUT_1[27645] = 32'b00000000000000000010001110011000;
assign LUT_1[27646] = 32'b00000000000000000100101010101101;
assign LUT_1[27647] = 32'b11111111111111111101111100101001;
assign LUT_1[27648] = 32'b00000000000000001000110101001011;
assign LUT_1[27649] = 32'b00000000000000000010000111000111;
assign LUT_1[27650] = 32'b00000000000000000100100011011100;
assign LUT_1[27651] = 32'b11111111111111111101110101011000;
assign LUT_1[27652] = 32'b00000000000000010000101110100010;
assign LUT_1[27653] = 32'b00000000000000001010000000011110;
assign LUT_1[27654] = 32'b00000000000000001100011100110011;
assign LUT_1[27655] = 32'b00000000000000000101101110101111;
assign LUT_1[27656] = 32'b00000000000000001000000011000000;
assign LUT_1[27657] = 32'b00000000000000000001010100111100;
assign LUT_1[27658] = 32'b00000000000000000011110001010001;
assign LUT_1[27659] = 32'b11111111111111111101000011001101;
assign LUT_1[27660] = 32'b00000000000000001111111100010111;
assign LUT_1[27661] = 32'b00000000000000001001001110010011;
assign LUT_1[27662] = 32'b00000000000000001011101010101000;
assign LUT_1[27663] = 32'b00000000000000000100111100100100;
assign LUT_1[27664] = 32'b00000000000000001010110000101101;
assign LUT_1[27665] = 32'b00000000000000000100000010101001;
assign LUT_1[27666] = 32'b00000000000000000110011110111110;
assign LUT_1[27667] = 32'b11111111111111111111110000111010;
assign LUT_1[27668] = 32'b00000000000000010010101010000100;
assign LUT_1[27669] = 32'b00000000000000001011111100000000;
assign LUT_1[27670] = 32'b00000000000000001110011000010101;
assign LUT_1[27671] = 32'b00000000000000000111101010010001;
assign LUT_1[27672] = 32'b00000000000000001001111110100010;
assign LUT_1[27673] = 32'b00000000000000000011010000011110;
assign LUT_1[27674] = 32'b00000000000000000101101100110011;
assign LUT_1[27675] = 32'b11111111111111111110111110101111;
assign LUT_1[27676] = 32'b00000000000000010001110111111001;
assign LUT_1[27677] = 32'b00000000000000001011001001110101;
assign LUT_1[27678] = 32'b00000000000000001101100110001010;
assign LUT_1[27679] = 32'b00000000000000000110111000000110;
assign LUT_1[27680] = 32'b00000000000000001001110000001010;
assign LUT_1[27681] = 32'b00000000000000000011000010000110;
assign LUT_1[27682] = 32'b00000000000000000101011110011011;
assign LUT_1[27683] = 32'b11111111111111111110110000010111;
assign LUT_1[27684] = 32'b00000000000000010001101001100001;
assign LUT_1[27685] = 32'b00000000000000001010111011011101;
assign LUT_1[27686] = 32'b00000000000000001101010111110010;
assign LUT_1[27687] = 32'b00000000000000000110101001101110;
assign LUT_1[27688] = 32'b00000000000000001000111101111111;
assign LUT_1[27689] = 32'b00000000000000000010001111111011;
assign LUT_1[27690] = 32'b00000000000000000100101100010000;
assign LUT_1[27691] = 32'b11111111111111111101111110001100;
assign LUT_1[27692] = 32'b00000000000000010000110111010110;
assign LUT_1[27693] = 32'b00000000000000001010001001010010;
assign LUT_1[27694] = 32'b00000000000000001100100101100111;
assign LUT_1[27695] = 32'b00000000000000000101110111100011;
assign LUT_1[27696] = 32'b00000000000000001011101011101100;
assign LUT_1[27697] = 32'b00000000000000000100111101101000;
assign LUT_1[27698] = 32'b00000000000000000111011001111101;
assign LUT_1[27699] = 32'b00000000000000000000101011111001;
assign LUT_1[27700] = 32'b00000000000000010011100101000011;
assign LUT_1[27701] = 32'b00000000000000001100110110111111;
assign LUT_1[27702] = 32'b00000000000000001111010011010100;
assign LUT_1[27703] = 32'b00000000000000001000100101010000;
assign LUT_1[27704] = 32'b00000000000000001010111001100001;
assign LUT_1[27705] = 32'b00000000000000000100001011011101;
assign LUT_1[27706] = 32'b00000000000000000110100111110010;
assign LUT_1[27707] = 32'b11111111111111111111111001101110;
assign LUT_1[27708] = 32'b00000000000000010010110010111000;
assign LUT_1[27709] = 32'b00000000000000001100000100110100;
assign LUT_1[27710] = 32'b00000000000000001110100001001001;
assign LUT_1[27711] = 32'b00000000000000000111110011000101;
assign LUT_1[27712] = 32'b00000000000000001010110010110011;
assign LUT_1[27713] = 32'b00000000000000000100000100101111;
assign LUT_1[27714] = 32'b00000000000000000110100001000100;
assign LUT_1[27715] = 32'b11111111111111111111110011000000;
assign LUT_1[27716] = 32'b00000000000000010010101100001010;
assign LUT_1[27717] = 32'b00000000000000001011111110000110;
assign LUT_1[27718] = 32'b00000000000000001110011010011011;
assign LUT_1[27719] = 32'b00000000000000000111101100010111;
assign LUT_1[27720] = 32'b00000000000000001010000000101000;
assign LUT_1[27721] = 32'b00000000000000000011010010100100;
assign LUT_1[27722] = 32'b00000000000000000101101110111001;
assign LUT_1[27723] = 32'b11111111111111111111000000110101;
assign LUT_1[27724] = 32'b00000000000000010001111001111111;
assign LUT_1[27725] = 32'b00000000000000001011001011111011;
assign LUT_1[27726] = 32'b00000000000000001101101000010000;
assign LUT_1[27727] = 32'b00000000000000000110111010001100;
assign LUT_1[27728] = 32'b00000000000000001100101110010101;
assign LUT_1[27729] = 32'b00000000000000000110000000010001;
assign LUT_1[27730] = 32'b00000000000000001000011100100110;
assign LUT_1[27731] = 32'b00000000000000000001101110100010;
assign LUT_1[27732] = 32'b00000000000000010100100111101100;
assign LUT_1[27733] = 32'b00000000000000001101111001101000;
assign LUT_1[27734] = 32'b00000000000000010000010101111101;
assign LUT_1[27735] = 32'b00000000000000001001100111111001;
assign LUT_1[27736] = 32'b00000000000000001011111100001010;
assign LUT_1[27737] = 32'b00000000000000000101001110000110;
assign LUT_1[27738] = 32'b00000000000000000111101010011011;
assign LUT_1[27739] = 32'b00000000000000000000111100010111;
assign LUT_1[27740] = 32'b00000000000000010011110101100001;
assign LUT_1[27741] = 32'b00000000000000001101000111011101;
assign LUT_1[27742] = 32'b00000000000000001111100011110010;
assign LUT_1[27743] = 32'b00000000000000001000110101101110;
assign LUT_1[27744] = 32'b00000000000000001011101101110010;
assign LUT_1[27745] = 32'b00000000000000000100111111101110;
assign LUT_1[27746] = 32'b00000000000000000111011100000011;
assign LUT_1[27747] = 32'b00000000000000000000101101111111;
assign LUT_1[27748] = 32'b00000000000000010011100111001001;
assign LUT_1[27749] = 32'b00000000000000001100111001000101;
assign LUT_1[27750] = 32'b00000000000000001111010101011010;
assign LUT_1[27751] = 32'b00000000000000001000100111010110;
assign LUT_1[27752] = 32'b00000000000000001010111011100111;
assign LUT_1[27753] = 32'b00000000000000000100001101100011;
assign LUT_1[27754] = 32'b00000000000000000110101001111000;
assign LUT_1[27755] = 32'b11111111111111111111111011110100;
assign LUT_1[27756] = 32'b00000000000000010010110100111110;
assign LUT_1[27757] = 32'b00000000000000001100000110111010;
assign LUT_1[27758] = 32'b00000000000000001110100011001111;
assign LUT_1[27759] = 32'b00000000000000000111110101001011;
assign LUT_1[27760] = 32'b00000000000000001101101001010100;
assign LUT_1[27761] = 32'b00000000000000000110111011010000;
assign LUT_1[27762] = 32'b00000000000000001001010111100101;
assign LUT_1[27763] = 32'b00000000000000000010101001100001;
assign LUT_1[27764] = 32'b00000000000000010101100010101011;
assign LUT_1[27765] = 32'b00000000000000001110110100100111;
assign LUT_1[27766] = 32'b00000000000000010001010000111100;
assign LUT_1[27767] = 32'b00000000000000001010100010111000;
assign LUT_1[27768] = 32'b00000000000000001100110111001001;
assign LUT_1[27769] = 32'b00000000000000000110001001000101;
assign LUT_1[27770] = 32'b00000000000000001000100101011010;
assign LUT_1[27771] = 32'b00000000000000000001110111010110;
assign LUT_1[27772] = 32'b00000000000000010100110000100000;
assign LUT_1[27773] = 32'b00000000000000001110000010011100;
assign LUT_1[27774] = 32'b00000000000000010000011110110001;
assign LUT_1[27775] = 32'b00000000000000001001110000101101;
assign LUT_1[27776] = 32'b00000000000000001011110101001110;
assign LUT_1[27777] = 32'b00000000000000000101000111001010;
assign LUT_1[27778] = 32'b00000000000000000111100011011111;
assign LUT_1[27779] = 32'b00000000000000000000110101011011;
assign LUT_1[27780] = 32'b00000000000000010011101110100101;
assign LUT_1[27781] = 32'b00000000000000001101000000100001;
assign LUT_1[27782] = 32'b00000000000000001111011100110110;
assign LUT_1[27783] = 32'b00000000000000001000101110110010;
assign LUT_1[27784] = 32'b00000000000000001011000011000011;
assign LUT_1[27785] = 32'b00000000000000000100010100111111;
assign LUT_1[27786] = 32'b00000000000000000110110001010100;
assign LUT_1[27787] = 32'b00000000000000000000000011010000;
assign LUT_1[27788] = 32'b00000000000000010010111100011010;
assign LUT_1[27789] = 32'b00000000000000001100001110010110;
assign LUT_1[27790] = 32'b00000000000000001110101010101011;
assign LUT_1[27791] = 32'b00000000000000000111111100100111;
assign LUT_1[27792] = 32'b00000000000000001101110000110000;
assign LUT_1[27793] = 32'b00000000000000000111000010101100;
assign LUT_1[27794] = 32'b00000000000000001001011111000001;
assign LUT_1[27795] = 32'b00000000000000000010110000111101;
assign LUT_1[27796] = 32'b00000000000000010101101010000111;
assign LUT_1[27797] = 32'b00000000000000001110111100000011;
assign LUT_1[27798] = 32'b00000000000000010001011000011000;
assign LUT_1[27799] = 32'b00000000000000001010101010010100;
assign LUT_1[27800] = 32'b00000000000000001100111110100101;
assign LUT_1[27801] = 32'b00000000000000000110010000100001;
assign LUT_1[27802] = 32'b00000000000000001000101100110110;
assign LUT_1[27803] = 32'b00000000000000000001111110110010;
assign LUT_1[27804] = 32'b00000000000000010100110111111100;
assign LUT_1[27805] = 32'b00000000000000001110001001111000;
assign LUT_1[27806] = 32'b00000000000000010000100110001101;
assign LUT_1[27807] = 32'b00000000000000001001111000001001;
assign LUT_1[27808] = 32'b00000000000000001100110000001101;
assign LUT_1[27809] = 32'b00000000000000000110000010001001;
assign LUT_1[27810] = 32'b00000000000000001000011110011110;
assign LUT_1[27811] = 32'b00000000000000000001110000011010;
assign LUT_1[27812] = 32'b00000000000000010100101001100100;
assign LUT_1[27813] = 32'b00000000000000001101111011100000;
assign LUT_1[27814] = 32'b00000000000000010000010111110101;
assign LUT_1[27815] = 32'b00000000000000001001101001110001;
assign LUT_1[27816] = 32'b00000000000000001011111110000010;
assign LUT_1[27817] = 32'b00000000000000000101001111111110;
assign LUT_1[27818] = 32'b00000000000000000111101100010011;
assign LUT_1[27819] = 32'b00000000000000000000111110001111;
assign LUT_1[27820] = 32'b00000000000000010011110111011001;
assign LUT_1[27821] = 32'b00000000000000001101001001010101;
assign LUT_1[27822] = 32'b00000000000000001111100101101010;
assign LUT_1[27823] = 32'b00000000000000001000110111100110;
assign LUT_1[27824] = 32'b00000000000000001110101011101111;
assign LUT_1[27825] = 32'b00000000000000000111111101101011;
assign LUT_1[27826] = 32'b00000000000000001010011010000000;
assign LUT_1[27827] = 32'b00000000000000000011101011111100;
assign LUT_1[27828] = 32'b00000000000000010110100101000110;
assign LUT_1[27829] = 32'b00000000000000001111110111000010;
assign LUT_1[27830] = 32'b00000000000000010010010011010111;
assign LUT_1[27831] = 32'b00000000000000001011100101010011;
assign LUT_1[27832] = 32'b00000000000000001101111001100100;
assign LUT_1[27833] = 32'b00000000000000000111001011100000;
assign LUT_1[27834] = 32'b00000000000000001001100111110101;
assign LUT_1[27835] = 32'b00000000000000000010111001110001;
assign LUT_1[27836] = 32'b00000000000000010101110010111011;
assign LUT_1[27837] = 32'b00000000000000001111000100110111;
assign LUT_1[27838] = 32'b00000000000000010001100001001100;
assign LUT_1[27839] = 32'b00000000000000001010110011001000;
assign LUT_1[27840] = 32'b00000000000000001101110010110110;
assign LUT_1[27841] = 32'b00000000000000000111000100110010;
assign LUT_1[27842] = 32'b00000000000000001001100001000111;
assign LUT_1[27843] = 32'b00000000000000000010110011000011;
assign LUT_1[27844] = 32'b00000000000000010101101100001101;
assign LUT_1[27845] = 32'b00000000000000001110111110001001;
assign LUT_1[27846] = 32'b00000000000000010001011010011110;
assign LUT_1[27847] = 32'b00000000000000001010101100011010;
assign LUT_1[27848] = 32'b00000000000000001101000000101011;
assign LUT_1[27849] = 32'b00000000000000000110010010100111;
assign LUT_1[27850] = 32'b00000000000000001000101110111100;
assign LUT_1[27851] = 32'b00000000000000000010000000111000;
assign LUT_1[27852] = 32'b00000000000000010100111010000010;
assign LUT_1[27853] = 32'b00000000000000001110001011111110;
assign LUT_1[27854] = 32'b00000000000000010000101000010011;
assign LUT_1[27855] = 32'b00000000000000001001111010001111;
assign LUT_1[27856] = 32'b00000000000000001111101110011000;
assign LUT_1[27857] = 32'b00000000000000001001000000010100;
assign LUT_1[27858] = 32'b00000000000000001011011100101001;
assign LUT_1[27859] = 32'b00000000000000000100101110100101;
assign LUT_1[27860] = 32'b00000000000000010111100111101111;
assign LUT_1[27861] = 32'b00000000000000010000111001101011;
assign LUT_1[27862] = 32'b00000000000000010011010110000000;
assign LUT_1[27863] = 32'b00000000000000001100100111111100;
assign LUT_1[27864] = 32'b00000000000000001110111100001101;
assign LUT_1[27865] = 32'b00000000000000001000001110001001;
assign LUT_1[27866] = 32'b00000000000000001010101010011110;
assign LUT_1[27867] = 32'b00000000000000000011111100011010;
assign LUT_1[27868] = 32'b00000000000000010110110101100100;
assign LUT_1[27869] = 32'b00000000000000010000000111100000;
assign LUT_1[27870] = 32'b00000000000000010010100011110101;
assign LUT_1[27871] = 32'b00000000000000001011110101110001;
assign LUT_1[27872] = 32'b00000000000000001110101101110101;
assign LUT_1[27873] = 32'b00000000000000000111111111110001;
assign LUT_1[27874] = 32'b00000000000000001010011100000110;
assign LUT_1[27875] = 32'b00000000000000000011101110000010;
assign LUT_1[27876] = 32'b00000000000000010110100111001100;
assign LUT_1[27877] = 32'b00000000000000001111111001001000;
assign LUT_1[27878] = 32'b00000000000000010010010101011101;
assign LUT_1[27879] = 32'b00000000000000001011100111011001;
assign LUT_1[27880] = 32'b00000000000000001101111011101010;
assign LUT_1[27881] = 32'b00000000000000000111001101100110;
assign LUT_1[27882] = 32'b00000000000000001001101001111011;
assign LUT_1[27883] = 32'b00000000000000000010111011110111;
assign LUT_1[27884] = 32'b00000000000000010101110101000001;
assign LUT_1[27885] = 32'b00000000000000001111000110111101;
assign LUT_1[27886] = 32'b00000000000000010001100011010010;
assign LUT_1[27887] = 32'b00000000000000001010110101001110;
assign LUT_1[27888] = 32'b00000000000000010000101001010111;
assign LUT_1[27889] = 32'b00000000000000001001111011010011;
assign LUT_1[27890] = 32'b00000000000000001100010111101000;
assign LUT_1[27891] = 32'b00000000000000000101101001100100;
assign LUT_1[27892] = 32'b00000000000000011000100010101110;
assign LUT_1[27893] = 32'b00000000000000010001110100101010;
assign LUT_1[27894] = 32'b00000000000000010100010000111111;
assign LUT_1[27895] = 32'b00000000000000001101100010111011;
assign LUT_1[27896] = 32'b00000000000000001111110111001100;
assign LUT_1[27897] = 32'b00000000000000001001001001001000;
assign LUT_1[27898] = 32'b00000000000000001011100101011101;
assign LUT_1[27899] = 32'b00000000000000000100110111011001;
assign LUT_1[27900] = 32'b00000000000000010111110000100011;
assign LUT_1[27901] = 32'b00000000000000010001000010011111;
assign LUT_1[27902] = 32'b00000000000000010011011110110100;
assign LUT_1[27903] = 32'b00000000000000001100110000110000;
assign LUT_1[27904] = 32'b00000000000000000110101001010111;
assign LUT_1[27905] = 32'b11111111111111111111111011010011;
assign LUT_1[27906] = 32'b00000000000000000010010111101000;
assign LUT_1[27907] = 32'b11111111111111111011101001100100;
assign LUT_1[27908] = 32'b00000000000000001110100010101110;
assign LUT_1[27909] = 32'b00000000000000000111110100101010;
assign LUT_1[27910] = 32'b00000000000000001010010000111111;
assign LUT_1[27911] = 32'b00000000000000000011100010111011;
assign LUT_1[27912] = 32'b00000000000000000101110111001100;
assign LUT_1[27913] = 32'b11111111111111111111001001001000;
assign LUT_1[27914] = 32'b00000000000000000001100101011101;
assign LUT_1[27915] = 32'b11111111111111111010110111011001;
assign LUT_1[27916] = 32'b00000000000000001101110000100011;
assign LUT_1[27917] = 32'b00000000000000000111000010011111;
assign LUT_1[27918] = 32'b00000000000000001001011110110100;
assign LUT_1[27919] = 32'b00000000000000000010110000110000;
assign LUT_1[27920] = 32'b00000000000000001000100100111001;
assign LUT_1[27921] = 32'b00000000000000000001110110110101;
assign LUT_1[27922] = 32'b00000000000000000100010011001010;
assign LUT_1[27923] = 32'b11111111111111111101100101000110;
assign LUT_1[27924] = 32'b00000000000000010000011110010000;
assign LUT_1[27925] = 32'b00000000000000001001110000001100;
assign LUT_1[27926] = 32'b00000000000000001100001100100001;
assign LUT_1[27927] = 32'b00000000000000000101011110011101;
assign LUT_1[27928] = 32'b00000000000000000111110010101110;
assign LUT_1[27929] = 32'b00000000000000000001000100101010;
assign LUT_1[27930] = 32'b00000000000000000011100000111111;
assign LUT_1[27931] = 32'b11111111111111111100110010111011;
assign LUT_1[27932] = 32'b00000000000000001111101100000101;
assign LUT_1[27933] = 32'b00000000000000001000111110000001;
assign LUT_1[27934] = 32'b00000000000000001011011010010110;
assign LUT_1[27935] = 32'b00000000000000000100101100010010;
assign LUT_1[27936] = 32'b00000000000000000111100100010110;
assign LUT_1[27937] = 32'b00000000000000000000110110010010;
assign LUT_1[27938] = 32'b00000000000000000011010010100111;
assign LUT_1[27939] = 32'b11111111111111111100100100100011;
assign LUT_1[27940] = 32'b00000000000000001111011101101101;
assign LUT_1[27941] = 32'b00000000000000001000101111101001;
assign LUT_1[27942] = 32'b00000000000000001011001011111110;
assign LUT_1[27943] = 32'b00000000000000000100011101111010;
assign LUT_1[27944] = 32'b00000000000000000110110010001011;
assign LUT_1[27945] = 32'b00000000000000000000000100000111;
assign LUT_1[27946] = 32'b00000000000000000010100000011100;
assign LUT_1[27947] = 32'b11111111111111111011110010011000;
assign LUT_1[27948] = 32'b00000000000000001110101011100010;
assign LUT_1[27949] = 32'b00000000000000000111111101011110;
assign LUT_1[27950] = 32'b00000000000000001010011001110011;
assign LUT_1[27951] = 32'b00000000000000000011101011101111;
assign LUT_1[27952] = 32'b00000000000000001001011111111000;
assign LUT_1[27953] = 32'b00000000000000000010110001110100;
assign LUT_1[27954] = 32'b00000000000000000101001110001001;
assign LUT_1[27955] = 32'b11111111111111111110100000000101;
assign LUT_1[27956] = 32'b00000000000000010001011001001111;
assign LUT_1[27957] = 32'b00000000000000001010101011001011;
assign LUT_1[27958] = 32'b00000000000000001101000111100000;
assign LUT_1[27959] = 32'b00000000000000000110011001011100;
assign LUT_1[27960] = 32'b00000000000000001000101101101101;
assign LUT_1[27961] = 32'b00000000000000000001111111101001;
assign LUT_1[27962] = 32'b00000000000000000100011011111110;
assign LUT_1[27963] = 32'b11111111111111111101101101111010;
assign LUT_1[27964] = 32'b00000000000000010000100111000100;
assign LUT_1[27965] = 32'b00000000000000001001111001000000;
assign LUT_1[27966] = 32'b00000000000000001100010101010101;
assign LUT_1[27967] = 32'b00000000000000000101100111010001;
assign LUT_1[27968] = 32'b00000000000000001000100110111111;
assign LUT_1[27969] = 32'b00000000000000000001111000111011;
assign LUT_1[27970] = 32'b00000000000000000100010101010000;
assign LUT_1[27971] = 32'b11111111111111111101100111001100;
assign LUT_1[27972] = 32'b00000000000000010000100000010110;
assign LUT_1[27973] = 32'b00000000000000001001110010010010;
assign LUT_1[27974] = 32'b00000000000000001100001110100111;
assign LUT_1[27975] = 32'b00000000000000000101100000100011;
assign LUT_1[27976] = 32'b00000000000000000111110100110100;
assign LUT_1[27977] = 32'b00000000000000000001000110110000;
assign LUT_1[27978] = 32'b00000000000000000011100011000101;
assign LUT_1[27979] = 32'b11111111111111111100110101000001;
assign LUT_1[27980] = 32'b00000000000000001111101110001011;
assign LUT_1[27981] = 32'b00000000000000001001000000000111;
assign LUT_1[27982] = 32'b00000000000000001011011100011100;
assign LUT_1[27983] = 32'b00000000000000000100101110011000;
assign LUT_1[27984] = 32'b00000000000000001010100010100001;
assign LUT_1[27985] = 32'b00000000000000000011110100011101;
assign LUT_1[27986] = 32'b00000000000000000110010000110010;
assign LUT_1[27987] = 32'b11111111111111111111100010101110;
assign LUT_1[27988] = 32'b00000000000000010010011011111000;
assign LUT_1[27989] = 32'b00000000000000001011101101110100;
assign LUT_1[27990] = 32'b00000000000000001110001010001001;
assign LUT_1[27991] = 32'b00000000000000000111011100000101;
assign LUT_1[27992] = 32'b00000000000000001001110000010110;
assign LUT_1[27993] = 32'b00000000000000000011000010010010;
assign LUT_1[27994] = 32'b00000000000000000101011110100111;
assign LUT_1[27995] = 32'b11111111111111111110110000100011;
assign LUT_1[27996] = 32'b00000000000000010001101001101101;
assign LUT_1[27997] = 32'b00000000000000001010111011101001;
assign LUT_1[27998] = 32'b00000000000000001101010111111110;
assign LUT_1[27999] = 32'b00000000000000000110101001111010;
assign LUT_1[28000] = 32'b00000000000000001001100001111110;
assign LUT_1[28001] = 32'b00000000000000000010110011111010;
assign LUT_1[28002] = 32'b00000000000000000101010000001111;
assign LUT_1[28003] = 32'b11111111111111111110100010001011;
assign LUT_1[28004] = 32'b00000000000000010001011011010101;
assign LUT_1[28005] = 32'b00000000000000001010101101010001;
assign LUT_1[28006] = 32'b00000000000000001101001001100110;
assign LUT_1[28007] = 32'b00000000000000000110011011100010;
assign LUT_1[28008] = 32'b00000000000000001000101111110011;
assign LUT_1[28009] = 32'b00000000000000000010000001101111;
assign LUT_1[28010] = 32'b00000000000000000100011110000100;
assign LUT_1[28011] = 32'b11111111111111111101110000000000;
assign LUT_1[28012] = 32'b00000000000000010000101001001010;
assign LUT_1[28013] = 32'b00000000000000001001111011000110;
assign LUT_1[28014] = 32'b00000000000000001100010111011011;
assign LUT_1[28015] = 32'b00000000000000000101101001010111;
assign LUT_1[28016] = 32'b00000000000000001011011101100000;
assign LUT_1[28017] = 32'b00000000000000000100101111011100;
assign LUT_1[28018] = 32'b00000000000000000111001011110001;
assign LUT_1[28019] = 32'b00000000000000000000011101101101;
assign LUT_1[28020] = 32'b00000000000000010011010110110111;
assign LUT_1[28021] = 32'b00000000000000001100101000110011;
assign LUT_1[28022] = 32'b00000000000000001111000101001000;
assign LUT_1[28023] = 32'b00000000000000001000010111000100;
assign LUT_1[28024] = 32'b00000000000000001010101011010101;
assign LUT_1[28025] = 32'b00000000000000000011111101010001;
assign LUT_1[28026] = 32'b00000000000000000110011001100110;
assign LUT_1[28027] = 32'b11111111111111111111101011100010;
assign LUT_1[28028] = 32'b00000000000000010010100100101100;
assign LUT_1[28029] = 32'b00000000000000001011110110101000;
assign LUT_1[28030] = 32'b00000000000000001110010010111101;
assign LUT_1[28031] = 32'b00000000000000000111100100111001;
assign LUT_1[28032] = 32'b00000000000000001001101001011010;
assign LUT_1[28033] = 32'b00000000000000000010111011010110;
assign LUT_1[28034] = 32'b00000000000000000101010111101011;
assign LUT_1[28035] = 32'b11111111111111111110101001100111;
assign LUT_1[28036] = 32'b00000000000000010001100010110001;
assign LUT_1[28037] = 32'b00000000000000001010110100101101;
assign LUT_1[28038] = 32'b00000000000000001101010001000010;
assign LUT_1[28039] = 32'b00000000000000000110100010111110;
assign LUT_1[28040] = 32'b00000000000000001000110111001111;
assign LUT_1[28041] = 32'b00000000000000000010001001001011;
assign LUT_1[28042] = 32'b00000000000000000100100101100000;
assign LUT_1[28043] = 32'b11111111111111111101110111011100;
assign LUT_1[28044] = 32'b00000000000000010000110000100110;
assign LUT_1[28045] = 32'b00000000000000001010000010100010;
assign LUT_1[28046] = 32'b00000000000000001100011110110111;
assign LUT_1[28047] = 32'b00000000000000000101110000110011;
assign LUT_1[28048] = 32'b00000000000000001011100100111100;
assign LUT_1[28049] = 32'b00000000000000000100110110111000;
assign LUT_1[28050] = 32'b00000000000000000111010011001101;
assign LUT_1[28051] = 32'b00000000000000000000100101001001;
assign LUT_1[28052] = 32'b00000000000000010011011110010011;
assign LUT_1[28053] = 32'b00000000000000001100110000001111;
assign LUT_1[28054] = 32'b00000000000000001111001100100100;
assign LUT_1[28055] = 32'b00000000000000001000011110100000;
assign LUT_1[28056] = 32'b00000000000000001010110010110001;
assign LUT_1[28057] = 32'b00000000000000000100000100101101;
assign LUT_1[28058] = 32'b00000000000000000110100001000010;
assign LUT_1[28059] = 32'b11111111111111111111110010111110;
assign LUT_1[28060] = 32'b00000000000000010010101100001000;
assign LUT_1[28061] = 32'b00000000000000001011111110000100;
assign LUT_1[28062] = 32'b00000000000000001110011010011001;
assign LUT_1[28063] = 32'b00000000000000000111101100010101;
assign LUT_1[28064] = 32'b00000000000000001010100100011001;
assign LUT_1[28065] = 32'b00000000000000000011110110010101;
assign LUT_1[28066] = 32'b00000000000000000110010010101010;
assign LUT_1[28067] = 32'b11111111111111111111100100100110;
assign LUT_1[28068] = 32'b00000000000000010010011101110000;
assign LUT_1[28069] = 32'b00000000000000001011101111101100;
assign LUT_1[28070] = 32'b00000000000000001110001100000001;
assign LUT_1[28071] = 32'b00000000000000000111011101111101;
assign LUT_1[28072] = 32'b00000000000000001001110010001110;
assign LUT_1[28073] = 32'b00000000000000000011000100001010;
assign LUT_1[28074] = 32'b00000000000000000101100000011111;
assign LUT_1[28075] = 32'b11111111111111111110110010011011;
assign LUT_1[28076] = 32'b00000000000000010001101011100101;
assign LUT_1[28077] = 32'b00000000000000001010111101100001;
assign LUT_1[28078] = 32'b00000000000000001101011001110110;
assign LUT_1[28079] = 32'b00000000000000000110101011110010;
assign LUT_1[28080] = 32'b00000000000000001100011111111011;
assign LUT_1[28081] = 32'b00000000000000000101110001110111;
assign LUT_1[28082] = 32'b00000000000000001000001110001100;
assign LUT_1[28083] = 32'b00000000000000000001100000001000;
assign LUT_1[28084] = 32'b00000000000000010100011001010010;
assign LUT_1[28085] = 32'b00000000000000001101101011001110;
assign LUT_1[28086] = 32'b00000000000000010000000111100011;
assign LUT_1[28087] = 32'b00000000000000001001011001011111;
assign LUT_1[28088] = 32'b00000000000000001011101101110000;
assign LUT_1[28089] = 32'b00000000000000000100111111101100;
assign LUT_1[28090] = 32'b00000000000000000111011100000001;
assign LUT_1[28091] = 32'b00000000000000000000101101111101;
assign LUT_1[28092] = 32'b00000000000000010011100111000111;
assign LUT_1[28093] = 32'b00000000000000001100111001000011;
assign LUT_1[28094] = 32'b00000000000000001111010101011000;
assign LUT_1[28095] = 32'b00000000000000001000100111010100;
assign LUT_1[28096] = 32'b00000000000000001011100111000010;
assign LUT_1[28097] = 32'b00000000000000000100111000111110;
assign LUT_1[28098] = 32'b00000000000000000111010101010011;
assign LUT_1[28099] = 32'b00000000000000000000100111001111;
assign LUT_1[28100] = 32'b00000000000000010011100000011001;
assign LUT_1[28101] = 32'b00000000000000001100110010010101;
assign LUT_1[28102] = 32'b00000000000000001111001110101010;
assign LUT_1[28103] = 32'b00000000000000001000100000100110;
assign LUT_1[28104] = 32'b00000000000000001010110100110111;
assign LUT_1[28105] = 32'b00000000000000000100000110110011;
assign LUT_1[28106] = 32'b00000000000000000110100011001000;
assign LUT_1[28107] = 32'b11111111111111111111110101000100;
assign LUT_1[28108] = 32'b00000000000000010010101110001110;
assign LUT_1[28109] = 32'b00000000000000001100000000001010;
assign LUT_1[28110] = 32'b00000000000000001110011100011111;
assign LUT_1[28111] = 32'b00000000000000000111101110011011;
assign LUT_1[28112] = 32'b00000000000000001101100010100100;
assign LUT_1[28113] = 32'b00000000000000000110110100100000;
assign LUT_1[28114] = 32'b00000000000000001001010000110101;
assign LUT_1[28115] = 32'b00000000000000000010100010110001;
assign LUT_1[28116] = 32'b00000000000000010101011011111011;
assign LUT_1[28117] = 32'b00000000000000001110101101110111;
assign LUT_1[28118] = 32'b00000000000000010001001010001100;
assign LUT_1[28119] = 32'b00000000000000001010011100001000;
assign LUT_1[28120] = 32'b00000000000000001100110000011001;
assign LUT_1[28121] = 32'b00000000000000000110000010010101;
assign LUT_1[28122] = 32'b00000000000000001000011110101010;
assign LUT_1[28123] = 32'b00000000000000000001110000100110;
assign LUT_1[28124] = 32'b00000000000000010100101001110000;
assign LUT_1[28125] = 32'b00000000000000001101111011101100;
assign LUT_1[28126] = 32'b00000000000000010000011000000001;
assign LUT_1[28127] = 32'b00000000000000001001101001111101;
assign LUT_1[28128] = 32'b00000000000000001100100010000001;
assign LUT_1[28129] = 32'b00000000000000000101110011111101;
assign LUT_1[28130] = 32'b00000000000000001000010000010010;
assign LUT_1[28131] = 32'b00000000000000000001100010001110;
assign LUT_1[28132] = 32'b00000000000000010100011011011000;
assign LUT_1[28133] = 32'b00000000000000001101101101010100;
assign LUT_1[28134] = 32'b00000000000000010000001001101001;
assign LUT_1[28135] = 32'b00000000000000001001011011100101;
assign LUT_1[28136] = 32'b00000000000000001011101111110110;
assign LUT_1[28137] = 32'b00000000000000000101000001110010;
assign LUT_1[28138] = 32'b00000000000000000111011110000111;
assign LUT_1[28139] = 32'b00000000000000000000110000000011;
assign LUT_1[28140] = 32'b00000000000000010011101001001101;
assign LUT_1[28141] = 32'b00000000000000001100111011001001;
assign LUT_1[28142] = 32'b00000000000000001111010111011110;
assign LUT_1[28143] = 32'b00000000000000001000101001011010;
assign LUT_1[28144] = 32'b00000000000000001110011101100011;
assign LUT_1[28145] = 32'b00000000000000000111101111011111;
assign LUT_1[28146] = 32'b00000000000000001010001011110100;
assign LUT_1[28147] = 32'b00000000000000000011011101110000;
assign LUT_1[28148] = 32'b00000000000000010110010110111010;
assign LUT_1[28149] = 32'b00000000000000001111101000110110;
assign LUT_1[28150] = 32'b00000000000000010010000101001011;
assign LUT_1[28151] = 32'b00000000000000001011010111000111;
assign LUT_1[28152] = 32'b00000000000000001101101011011000;
assign LUT_1[28153] = 32'b00000000000000000110111101010100;
assign LUT_1[28154] = 32'b00000000000000001001011001101001;
assign LUT_1[28155] = 32'b00000000000000000010101011100101;
assign LUT_1[28156] = 32'b00000000000000010101100100101111;
assign LUT_1[28157] = 32'b00000000000000001110110110101011;
assign LUT_1[28158] = 32'b00000000000000010001010011000000;
assign LUT_1[28159] = 32'b00000000000000001010100100111100;
assign LUT_1[28160] = 32'b00000000000000000010100011101000;
assign LUT_1[28161] = 32'b11111111111111111011110101100100;
assign LUT_1[28162] = 32'b11111111111111111110010001111001;
assign LUT_1[28163] = 32'b11111111111111110111100011110101;
assign LUT_1[28164] = 32'b00000000000000001010011100111111;
assign LUT_1[28165] = 32'b00000000000000000011101110111011;
assign LUT_1[28166] = 32'b00000000000000000110001011010000;
assign LUT_1[28167] = 32'b11111111111111111111011101001100;
assign LUT_1[28168] = 32'b00000000000000000001110001011101;
assign LUT_1[28169] = 32'b11111111111111111011000011011001;
assign LUT_1[28170] = 32'b11111111111111111101011111101110;
assign LUT_1[28171] = 32'b11111111111111110110110001101010;
assign LUT_1[28172] = 32'b00000000000000001001101010110100;
assign LUT_1[28173] = 32'b00000000000000000010111100110000;
assign LUT_1[28174] = 32'b00000000000000000101011001000101;
assign LUT_1[28175] = 32'b11111111111111111110101011000001;
assign LUT_1[28176] = 32'b00000000000000000100011111001010;
assign LUT_1[28177] = 32'b11111111111111111101110001000110;
assign LUT_1[28178] = 32'b00000000000000000000001101011011;
assign LUT_1[28179] = 32'b11111111111111111001011111010111;
assign LUT_1[28180] = 32'b00000000000000001100011000100001;
assign LUT_1[28181] = 32'b00000000000000000101101010011101;
assign LUT_1[28182] = 32'b00000000000000001000000110110010;
assign LUT_1[28183] = 32'b00000000000000000001011000101110;
assign LUT_1[28184] = 32'b00000000000000000011101100111111;
assign LUT_1[28185] = 32'b11111111111111111100111110111011;
assign LUT_1[28186] = 32'b11111111111111111111011011010000;
assign LUT_1[28187] = 32'b11111111111111111000101101001100;
assign LUT_1[28188] = 32'b00000000000000001011100110010110;
assign LUT_1[28189] = 32'b00000000000000000100111000010010;
assign LUT_1[28190] = 32'b00000000000000000111010100100111;
assign LUT_1[28191] = 32'b00000000000000000000100110100011;
assign LUT_1[28192] = 32'b00000000000000000011011110100111;
assign LUT_1[28193] = 32'b11111111111111111100110000100011;
assign LUT_1[28194] = 32'b11111111111111111111001100111000;
assign LUT_1[28195] = 32'b11111111111111111000011110110100;
assign LUT_1[28196] = 32'b00000000000000001011010111111110;
assign LUT_1[28197] = 32'b00000000000000000100101001111010;
assign LUT_1[28198] = 32'b00000000000000000111000110001111;
assign LUT_1[28199] = 32'b00000000000000000000011000001011;
assign LUT_1[28200] = 32'b00000000000000000010101100011100;
assign LUT_1[28201] = 32'b11111111111111111011111110011000;
assign LUT_1[28202] = 32'b11111111111111111110011010101101;
assign LUT_1[28203] = 32'b11111111111111110111101100101001;
assign LUT_1[28204] = 32'b00000000000000001010100101110011;
assign LUT_1[28205] = 32'b00000000000000000011110111101111;
assign LUT_1[28206] = 32'b00000000000000000110010100000100;
assign LUT_1[28207] = 32'b11111111111111111111100110000000;
assign LUT_1[28208] = 32'b00000000000000000101011010001001;
assign LUT_1[28209] = 32'b11111111111111111110101100000101;
assign LUT_1[28210] = 32'b00000000000000000001001000011010;
assign LUT_1[28211] = 32'b11111111111111111010011010010110;
assign LUT_1[28212] = 32'b00000000000000001101010011100000;
assign LUT_1[28213] = 32'b00000000000000000110100101011100;
assign LUT_1[28214] = 32'b00000000000000001001000001110001;
assign LUT_1[28215] = 32'b00000000000000000010010011101101;
assign LUT_1[28216] = 32'b00000000000000000100100111111110;
assign LUT_1[28217] = 32'b11111111111111111101111001111010;
assign LUT_1[28218] = 32'b00000000000000000000010110001111;
assign LUT_1[28219] = 32'b11111111111111111001101000001011;
assign LUT_1[28220] = 32'b00000000000000001100100001010101;
assign LUT_1[28221] = 32'b00000000000000000101110011010001;
assign LUT_1[28222] = 32'b00000000000000001000001111100110;
assign LUT_1[28223] = 32'b00000000000000000001100001100010;
assign LUT_1[28224] = 32'b00000000000000000100100001010000;
assign LUT_1[28225] = 32'b11111111111111111101110011001100;
assign LUT_1[28226] = 32'b00000000000000000000001111100001;
assign LUT_1[28227] = 32'b11111111111111111001100001011101;
assign LUT_1[28228] = 32'b00000000000000001100011010100111;
assign LUT_1[28229] = 32'b00000000000000000101101100100011;
assign LUT_1[28230] = 32'b00000000000000001000001000111000;
assign LUT_1[28231] = 32'b00000000000000000001011010110100;
assign LUT_1[28232] = 32'b00000000000000000011101111000101;
assign LUT_1[28233] = 32'b11111111111111111101000001000001;
assign LUT_1[28234] = 32'b11111111111111111111011101010110;
assign LUT_1[28235] = 32'b11111111111111111000101111010010;
assign LUT_1[28236] = 32'b00000000000000001011101000011100;
assign LUT_1[28237] = 32'b00000000000000000100111010011000;
assign LUT_1[28238] = 32'b00000000000000000111010110101101;
assign LUT_1[28239] = 32'b00000000000000000000101000101001;
assign LUT_1[28240] = 32'b00000000000000000110011100110010;
assign LUT_1[28241] = 32'b11111111111111111111101110101110;
assign LUT_1[28242] = 32'b00000000000000000010001011000011;
assign LUT_1[28243] = 32'b11111111111111111011011100111111;
assign LUT_1[28244] = 32'b00000000000000001110010110001001;
assign LUT_1[28245] = 32'b00000000000000000111101000000101;
assign LUT_1[28246] = 32'b00000000000000001010000100011010;
assign LUT_1[28247] = 32'b00000000000000000011010110010110;
assign LUT_1[28248] = 32'b00000000000000000101101010100111;
assign LUT_1[28249] = 32'b11111111111111111110111100100011;
assign LUT_1[28250] = 32'b00000000000000000001011000111000;
assign LUT_1[28251] = 32'b11111111111111111010101010110100;
assign LUT_1[28252] = 32'b00000000000000001101100011111110;
assign LUT_1[28253] = 32'b00000000000000000110110101111010;
assign LUT_1[28254] = 32'b00000000000000001001010010001111;
assign LUT_1[28255] = 32'b00000000000000000010100100001011;
assign LUT_1[28256] = 32'b00000000000000000101011100001111;
assign LUT_1[28257] = 32'b11111111111111111110101110001011;
assign LUT_1[28258] = 32'b00000000000000000001001010100000;
assign LUT_1[28259] = 32'b11111111111111111010011100011100;
assign LUT_1[28260] = 32'b00000000000000001101010101100110;
assign LUT_1[28261] = 32'b00000000000000000110100111100010;
assign LUT_1[28262] = 32'b00000000000000001001000011110111;
assign LUT_1[28263] = 32'b00000000000000000010010101110011;
assign LUT_1[28264] = 32'b00000000000000000100101010000100;
assign LUT_1[28265] = 32'b11111111111111111101111100000000;
assign LUT_1[28266] = 32'b00000000000000000000011000010101;
assign LUT_1[28267] = 32'b11111111111111111001101010010001;
assign LUT_1[28268] = 32'b00000000000000001100100011011011;
assign LUT_1[28269] = 32'b00000000000000000101110101010111;
assign LUT_1[28270] = 32'b00000000000000001000010001101100;
assign LUT_1[28271] = 32'b00000000000000000001100011101000;
assign LUT_1[28272] = 32'b00000000000000000111010111110001;
assign LUT_1[28273] = 32'b00000000000000000000101001101101;
assign LUT_1[28274] = 32'b00000000000000000011000110000010;
assign LUT_1[28275] = 32'b11111111111111111100010111111110;
assign LUT_1[28276] = 32'b00000000000000001111010001001000;
assign LUT_1[28277] = 32'b00000000000000001000100011000100;
assign LUT_1[28278] = 32'b00000000000000001010111111011001;
assign LUT_1[28279] = 32'b00000000000000000100010001010101;
assign LUT_1[28280] = 32'b00000000000000000110100101100110;
assign LUT_1[28281] = 32'b11111111111111111111110111100010;
assign LUT_1[28282] = 32'b00000000000000000010010011110111;
assign LUT_1[28283] = 32'b11111111111111111011100101110011;
assign LUT_1[28284] = 32'b00000000000000001110011110111101;
assign LUT_1[28285] = 32'b00000000000000000111110000111001;
assign LUT_1[28286] = 32'b00000000000000001010001101001110;
assign LUT_1[28287] = 32'b00000000000000000011011111001010;
assign LUT_1[28288] = 32'b00000000000000000101100011101011;
assign LUT_1[28289] = 32'b11111111111111111110110101100111;
assign LUT_1[28290] = 32'b00000000000000000001010001111100;
assign LUT_1[28291] = 32'b11111111111111111010100011111000;
assign LUT_1[28292] = 32'b00000000000000001101011101000010;
assign LUT_1[28293] = 32'b00000000000000000110101110111110;
assign LUT_1[28294] = 32'b00000000000000001001001011010011;
assign LUT_1[28295] = 32'b00000000000000000010011101001111;
assign LUT_1[28296] = 32'b00000000000000000100110001100000;
assign LUT_1[28297] = 32'b11111111111111111110000011011100;
assign LUT_1[28298] = 32'b00000000000000000000011111110001;
assign LUT_1[28299] = 32'b11111111111111111001110001101101;
assign LUT_1[28300] = 32'b00000000000000001100101010110111;
assign LUT_1[28301] = 32'b00000000000000000101111100110011;
assign LUT_1[28302] = 32'b00000000000000001000011001001000;
assign LUT_1[28303] = 32'b00000000000000000001101011000100;
assign LUT_1[28304] = 32'b00000000000000000111011111001101;
assign LUT_1[28305] = 32'b00000000000000000000110001001001;
assign LUT_1[28306] = 32'b00000000000000000011001101011110;
assign LUT_1[28307] = 32'b11111111111111111100011111011010;
assign LUT_1[28308] = 32'b00000000000000001111011000100100;
assign LUT_1[28309] = 32'b00000000000000001000101010100000;
assign LUT_1[28310] = 32'b00000000000000001011000110110101;
assign LUT_1[28311] = 32'b00000000000000000100011000110001;
assign LUT_1[28312] = 32'b00000000000000000110101101000010;
assign LUT_1[28313] = 32'b11111111111111111111111110111110;
assign LUT_1[28314] = 32'b00000000000000000010011011010011;
assign LUT_1[28315] = 32'b11111111111111111011101101001111;
assign LUT_1[28316] = 32'b00000000000000001110100110011001;
assign LUT_1[28317] = 32'b00000000000000000111111000010101;
assign LUT_1[28318] = 32'b00000000000000001010010100101010;
assign LUT_1[28319] = 32'b00000000000000000011100110100110;
assign LUT_1[28320] = 32'b00000000000000000110011110101010;
assign LUT_1[28321] = 32'b11111111111111111111110000100110;
assign LUT_1[28322] = 32'b00000000000000000010001100111011;
assign LUT_1[28323] = 32'b11111111111111111011011110110111;
assign LUT_1[28324] = 32'b00000000000000001110011000000001;
assign LUT_1[28325] = 32'b00000000000000000111101001111101;
assign LUT_1[28326] = 32'b00000000000000001010000110010010;
assign LUT_1[28327] = 32'b00000000000000000011011000001110;
assign LUT_1[28328] = 32'b00000000000000000101101100011111;
assign LUT_1[28329] = 32'b11111111111111111110111110011011;
assign LUT_1[28330] = 32'b00000000000000000001011010110000;
assign LUT_1[28331] = 32'b11111111111111111010101100101100;
assign LUT_1[28332] = 32'b00000000000000001101100101110110;
assign LUT_1[28333] = 32'b00000000000000000110110111110010;
assign LUT_1[28334] = 32'b00000000000000001001010100000111;
assign LUT_1[28335] = 32'b00000000000000000010100110000011;
assign LUT_1[28336] = 32'b00000000000000001000011010001100;
assign LUT_1[28337] = 32'b00000000000000000001101100001000;
assign LUT_1[28338] = 32'b00000000000000000100001000011101;
assign LUT_1[28339] = 32'b11111111111111111101011010011001;
assign LUT_1[28340] = 32'b00000000000000010000010011100011;
assign LUT_1[28341] = 32'b00000000000000001001100101011111;
assign LUT_1[28342] = 32'b00000000000000001100000001110100;
assign LUT_1[28343] = 32'b00000000000000000101010011110000;
assign LUT_1[28344] = 32'b00000000000000000111101000000001;
assign LUT_1[28345] = 32'b00000000000000000000111001111101;
assign LUT_1[28346] = 32'b00000000000000000011010110010010;
assign LUT_1[28347] = 32'b11111111111111111100101000001110;
assign LUT_1[28348] = 32'b00000000000000001111100001011000;
assign LUT_1[28349] = 32'b00000000000000001000110011010100;
assign LUT_1[28350] = 32'b00000000000000001011001111101001;
assign LUT_1[28351] = 32'b00000000000000000100100001100101;
assign LUT_1[28352] = 32'b00000000000000000111100001010011;
assign LUT_1[28353] = 32'b00000000000000000000110011001111;
assign LUT_1[28354] = 32'b00000000000000000011001111100100;
assign LUT_1[28355] = 32'b11111111111111111100100001100000;
assign LUT_1[28356] = 32'b00000000000000001111011010101010;
assign LUT_1[28357] = 32'b00000000000000001000101100100110;
assign LUT_1[28358] = 32'b00000000000000001011001000111011;
assign LUT_1[28359] = 32'b00000000000000000100011010110111;
assign LUT_1[28360] = 32'b00000000000000000110101111001000;
assign LUT_1[28361] = 32'b00000000000000000000000001000100;
assign LUT_1[28362] = 32'b00000000000000000010011101011001;
assign LUT_1[28363] = 32'b11111111111111111011101111010101;
assign LUT_1[28364] = 32'b00000000000000001110101000011111;
assign LUT_1[28365] = 32'b00000000000000000111111010011011;
assign LUT_1[28366] = 32'b00000000000000001010010110110000;
assign LUT_1[28367] = 32'b00000000000000000011101000101100;
assign LUT_1[28368] = 32'b00000000000000001001011100110101;
assign LUT_1[28369] = 32'b00000000000000000010101110110001;
assign LUT_1[28370] = 32'b00000000000000000101001011000110;
assign LUT_1[28371] = 32'b11111111111111111110011101000010;
assign LUT_1[28372] = 32'b00000000000000010001010110001100;
assign LUT_1[28373] = 32'b00000000000000001010101000001000;
assign LUT_1[28374] = 32'b00000000000000001101000100011101;
assign LUT_1[28375] = 32'b00000000000000000110010110011001;
assign LUT_1[28376] = 32'b00000000000000001000101010101010;
assign LUT_1[28377] = 32'b00000000000000000001111100100110;
assign LUT_1[28378] = 32'b00000000000000000100011000111011;
assign LUT_1[28379] = 32'b11111111111111111101101010110111;
assign LUT_1[28380] = 32'b00000000000000010000100100000001;
assign LUT_1[28381] = 32'b00000000000000001001110101111101;
assign LUT_1[28382] = 32'b00000000000000001100010010010010;
assign LUT_1[28383] = 32'b00000000000000000101100100001110;
assign LUT_1[28384] = 32'b00000000000000001000011100010010;
assign LUT_1[28385] = 32'b00000000000000000001101110001110;
assign LUT_1[28386] = 32'b00000000000000000100001010100011;
assign LUT_1[28387] = 32'b11111111111111111101011100011111;
assign LUT_1[28388] = 32'b00000000000000010000010101101001;
assign LUT_1[28389] = 32'b00000000000000001001100111100101;
assign LUT_1[28390] = 32'b00000000000000001100000011111010;
assign LUT_1[28391] = 32'b00000000000000000101010101110110;
assign LUT_1[28392] = 32'b00000000000000000111101010000111;
assign LUT_1[28393] = 32'b00000000000000000000111100000011;
assign LUT_1[28394] = 32'b00000000000000000011011000011000;
assign LUT_1[28395] = 32'b11111111111111111100101010010100;
assign LUT_1[28396] = 32'b00000000000000001111100011011110;
assign LUT_1[28397] = 32'b00000000000000001000110101011010;
assign LUT_1[28398] = 32'b00000000000000001011010001101111;
assign LUT_1[28399] = 32'b00000000000000000100100011101011;
assign LUT_1[28400] = 32'b00000000000000001010010111110100;
assign LUT_1[28401] = 32'b00000000000000000011101001110000;
assign LUT_1[28402] = 32'b00000000000000000110000110000101;
assign LUT_1[28403] = 32'b11111111111111111111011000000001;
assign LUT_1[28404] = 32'b00000000000000010010010001001011;
assign LUT_1[28405] = 32'b00000000000000001011100011000111;
assign LUT_1[28406] = 32'b00000000000000001101111111011100;
assign LUT_1[28407] = 32'b00000000000000000111010001011000;
assign LUT_1[28408] = 32'b00000000000000001001100101101001;
assign LUT_1[28409] = 32'b00000000000000000010110111100101;
assign LUT_1[28410] = 32'b00000000000000000101010011111010;
assign LUT_1[28411] = 32'b11111111111111111110100101110110;
assign LUT_1[28412] = 32'b00000000000000010001011111000000;
assign LUT_1[28413] = 32'b00000000000000001010110000111100;
assign LUT_1[28414] = 32'b00000000000000001101001101010001;
assign LUT_1[28415] = 32'b00000000000000000110011111001101;
assign LUT_1[28416] = 32'b00000000000000000000010111110100;
assign LUT_1[28417] = 32'b11111111111111111001101001110000;
assign LUT_1[28418] = 32'b11111111111111111100000110000101;
assign LUT_1[28419] = 32'b11111111111111110101011000000001;
assign LUT_1[28420] = 32'b00000000000000001000010001001011;
assign LUT_1[28421] = 32'b00000000000000000001100011000111;
assign LUT_1[28422] = 32'b00000000000000000011111111011100;
assign LUT_1[28423] = 32'b11111111111111111101010001011000;
assign LUT_1[28424] = 32'b11111111111111111111100101101001;
assign LUT_1[28425] = 32'b11111111111111111000110111100101;
assign LUT_1[28426] = 32'b11111111111111111011010011111010;
assign LUT_1[28427] = 32'b11111111111111110100100101110110;
assign LUT_1[28428] = 32'b00000000000000000111011111000000;
assign LUT_1[28429] = 32'b00000000000000000000110000111100;
assign LUT_1[28430] = 32'b00000000000000000011001101010001;
assign LUT_1[28431] = 32'b11111111111111111100011111001101;
assign LUT_1[28432] = 32'b00000000000000000010010011010110;
assign LUT_1[28433] = 32'b11111111111111111011100101010010;
assign LUT_1[28434] = 32'b11111111111111111110000001100111;
assign LUT_1[28435] = 32'b11111111111111110111010011100011;
assign LUT_1[28436] = 32'b00000000000000001010001100101101;
assign LUT_1[28437] = 32'b00000000000000000011011110101001;
assign LUT_1[28438] = 32'b00000000000000000101111010111110;
assign LUT_1[28439] = 32'b11111111111111111111001100111010;
assign LUT_1[28440] = 32'b00000000000000000001100001001011;
assign LUT_1[28441] = 32'b11111111111111111010110011000111;
assign LUT_1[28442] = 32'b11111111111111111101001111011100;
assign LUT_1[28443] = 32'b11111111111111110110100001011000;
assign LUT_1[28444] = 32'b00000000000000001001011010100010;
assign LUT_1[28445] = 32'b00000000000000000010101100011110;
assign LUT_1[28446] = 32'b00000000000000000101001000110011;
assign LUT_1[28447] = 32'b11111111111111111110011010101111;
assign LUT_1[28448] = 32'b00000000000000000001010010110011;
assign LUT_1[28449] = 32'b11111111111111111010100100101111;
assign LUT_1[28450] = 32'b11111111111111111101000001000100;
assign LUT_1[28451] = 32'b11111111111111110110010011000000;
assign LUT_1[28452] = 32'b00000000000000001001001100001010;
assign LUT_1[28453] = 32'b00000000000000000010011110000110;
assign LUT_1[28454] = 32'b00000000000000000100111010011011;
assign LUT_1[28455] = 32'b11111111111111111110001100010111;
assign LUT_1[28456] = 32'b00000000000000000000100000101000;
assign LUT_1[28457] = 32'b11111111111111111001110010100100;
assign LUT_1[28458] = 32'b11111111111111111100001110111001;
assign LUT_1[28459] = 32'b11111111111111110101100000110101;
assign LUT_1[28460] = 32'b00000000000000001000011001111111;
assign LUT_1[28461] = 32'b00000000000000000001101011111011;
assign LUT_1[28462] = 32'b00000000000000000100001000010000;
assign LUT_1[28463] = 32'b11111111111111111101011010001100;
assign LUT_1[28464] = 32'b00000000000000000011001110010101;
assign LUT_1[28465] = 32'b11111111111111111100100000010001;
assign LUT_1[28466] = 32'b11111111111111111110111100100110;
assign LUT_1[28467] = 32'b11111111111111111000001110100010;
assign LUT_1[28468] = 32'b00000000000000001011000111101100;
assign LUT_1[28469] = 32'b00000000000000000100011001101000;
assign LUT_1[28470] = 32'b00000000000000000110110101111101;
assign LUT_1[28471] = 32'b00000000000000000000000111111001;
assign LUT_1[28472] = 32'b00000000000000000010011100001010;
assign LUT_1[28473] = 32'b11111111111111111011101110000110;
assign LUT_1[28474] = 32'b11111111111111111110001010011011;
assign LUT_1[28475] = 32'b11111111111111110111011100010111;
assign LUT_1[28476] = 32'b00000000000000001010010101100001;
assign LUT_1[28477] = 32'b00000000000000000011100111011101;
assign LUT_1[28478] = 32'b00000000000000000110000011110010;
assign LUT_1[28479] = 32'b11111111111111111111010101101110;
assign LUT_1[28480] = 32'b00000000000000000010010101011100;
assign LUT_1[28481] = 32'b11111111111111111011100111011000;
assign LUT_1[28482] = 32'b11111111111111111110000011101101;
assign LUT_1[28483] = 32'b11111111111111110111010101101001;
assign LUT_1[28484] = 32'b00000000000000001010001110110011;
assign LUT_1[28485] = 32'b00000000000000000011100000101111;
assign LUT_1[28486] = 32'b00000000000000000101111101000100;
assign LUT_1[28487] = 32'b11111111111111111111001111000000;
assign LUT_1[28488] = 32'b00000000000000000001100011010001;
assign LUT_1[28489] = 32'b11111111111111111010110101001101;
assign LUT_1[28490] = 32'b11111111111111111101010001100010;
assign LUT_1[28491] = 32'b11111111111111110110100011011110;
assign LUT_1[28492] = 32'b00000000000000001001011100101000;
assign LUT_1[28493] = 32'b00000000000000000010101110100100;
assign LUT_1[28494] = 32'b00000000000000000101001010111001;
assign LUT_1[28495] = 32'b11111111111111111110011100110101;
assign LUT_1[28496] = 32'b00000000000000000100010000111110;
assign LUT_1[28497] = 32'b11111111111111111101100010111010;
assign LUT_1[28498] = 32'b11111111111111111111111111001111;
assign LUT_1[28499] = 32'b11111111111111111001010001001011;
assign LUT_1[28500] = 32'b00000000000000001100001010010101;
assign LUT_1[28501] = 32'b00000000000000000101011100010001;
assign LUT_1[28502] = 32'b00000000000000000111111000100110;
assign LUT_1[28503] = 32'b00000000000000000001001010100010;
assign LUT_1[28504] = 32'b00000000000000000011011110110011;
assign LUT_1[28505] = 32'b11111111111111111100110000101111;
assign LUT_1[28506] = 32'b11111111111111111111001101000100;
assign LUT_1[28507] = 32'b11111111111111111000011111000000;
assign LUT_1[28508] = 32'b00000000000000001011011000001010;
assign LUT_1[28509] = 32'b00000000000000000100101010000110;
assign LUT_1[28510] = 32'b00000000000000000111000110011011;
assign LUT_1[28511] = 32'b00000000000000000000011000010111;
assign LUT_1[28512] = 32'b00000000000000000011010000011011;
assign LUT_1[28513] = 32'b11111111111111111100100010010111;
assign LUT_1[28514] = 32'b11111111111111111110111110101100;
assign LUT_1[28515] = 32'b11111111111111111000010000101000;
assign LUT_1[28516] = 32'b00000000000000001011001001110010;
assign LUT_1[28517] = 32'b00000000000000000100011011101110;
assign LUT_1[28518] = 32'b00000000000000000110111000000011;
assign LUT_1[28519] = 32'b00000000000000000000001001111111;
assign LUT_1[28520] = 32'b00000000000000000010011110010000;
assign LUT_1[28521] = 32'b11111111111111111011110000001100;
assign LUT_1[28522] = 32'b11111111111111111110001100100001;
assign LUT_1[28523] = 32'b11111111111111110111011110011101;
assign LUT_1[28524] = 32'b00000000000000001010010111100111;
assign LUT_1[28525] = 32'b00000000000000000011101001100011;
assign LUT_1[28526] = 32'b00000000000000000110000101111000;
assign LUT_1[28527] = 32'b11111111111111111111010111110100;
assign LUT_1[28528] = 32'b00000000000000000101001011111101;
assign LUT_1[28529] = 32'b11111111111111111110011101111001;
assign LUT_1[28530] = 32'b00000000000000000000111010001110;
assign LUT_1[28531] = 32'b11111111111111111010001100001010;
assign LUT_1[28532] = 32'b00000000000000001101000101010100;
assign LUT_1[28533] = 32'b00000000000000000110010111010000;
assign LUT_1[28534] = 32'b00000000000000001000110011100101;
assign LUT_1[28535] = 32'b00000000000000000010000101100001;
assign LUT_1[28536] = 32'b00000000000000000100011001110010;
assign LUT_1[28537] = 32'b11111111111111111101101011101110;
assign LUT_1[28538] = 32'b00000000000000000000001000000011;
assign LUT_1[28539] = 32'b11111111111111111001011001111111;
assign LUT_1[28540] = 32'b00000000000000001100010011001001;
assign LUT_1[28541] = 32'b00000000000000000101100101000101;
assign LUT_1[28542] = 32'b00000000000000001000000001011010;
assign LUT_1[28543] = 32'b00000000000000000001010011010110;
assign LUT_1[28544] = 32'b00000000000000000011010111110111;
assign LUT_1[28545] = 32'b11111111111111111100101001110011;
assign LUT_1[28546] = 32'b11111111111111111111000110001000;
assign LUT_1[28547] = 32'b11111111111111111000011000000100;
assign LUT_1[28548] = 32'b00000000000000001011010001001110;
assign LUT_1[28549] = 32'b00000000000000000100100011001010;
assign LUT_1[28550] = 32'b00000000000000000110111111011111;
assign LUT_1[28551] = 32'b00000000000000000000010001011011;
assign LUT_1[28552] = 32'b00000000000000000010100101101100;
assign LUT_1[28553] = 32'b11111111111111111011110111101000;
assign LUT_1[28554] = 32'b11111111111111111110010011111101;
assign LUT_1[28555] = 32'b11111111111111110111100101111001;
assign LUT_1[28556] = 32'b00000000000000001010011111000011;
assign LUT_1[28557] = 32'b00000000000000000011110000111111;
assign LUT_1[28558] = 32'b00000000000000000110001101010100;
assign LUT_1[28559] = 32'b11111111111111111111011111010000;
assign LUT_1[28560] = 32'b00000000000000000101010011011001;
assign LUT_1[28561] = 32'b11111111111111111110100101010101;
assign LUT_1[28562] = 32'b00000000000000000001000001101010;
assign LUT_1[28563] = 32'b11111111111111111010010011100110;
assign LUT_1[28564] = 32'b00000000000000001101001100110000;
assign LUT_1[28565] = 32'b00000000000000000110011110101100;
assign LUT_1[28566] = 32'b00000000000000001000111011000001;
assign LUT_1[28567] = 32'b00000000000000000010001100111101;
assign LUT_1[28568] = 32'b00000000000000000100100001001110;
assign LUT_1[28569] = 32'b11111111111111111101110011001010;
assign LUT_1[28570] = 32'b00000000000000000000001111011111;
assign LUT_1[28571] = 32'b11111111111111111001100001011011;
assign LUT_1[28572] = 32'b00000000000000001100011010100101;
assign LUT_1[28573] = 32'b00000000000000000101101100100001;
assign LUT_1[28574] = 32'b00000000000000001000001000110110;
assign LUT_1[28575] = 32'b00000000000000000001011010110010;
assign LUT_1[28576] = 32'b00000000000000000100010010110110;
assign LUT_1[28577] = 32'b11111111111111111101100100110010;
assign LUT_1[28578] = 32'b00000000000000000000000001000111;
assign LUT_1[28579] = 32'b11111111111111111001010011000011;
assign LUT_1[28580] = 32'b00000000000000001100001100001101;
assign LUT_1[28581] = 32'b00000000000000000101011110001001;
assign LUT_1[28582] = 32'b00000000000000000111111010011110;
assign LUT_1[28583] = 32'b00000000000000000001001100011010;
assign LUT_1[28584] = 32'b00000000000000000011100000101011;
assign LUT_1[28585] = 32'b11111111111111111100110010100111;
assign LUT_1[28586] = 32'b11111111111111111111001110111100;
assign LUT_1[28587] = 32'b11111111111111111000100000111000;
assign LUT_1[28588] = 32'b00000000000000001011011010000010;
assign LUT_1[28589] = 32'b00000000000000000100101011111110;
assign LUT_1[28590] = 32'b00000000000000000111001000010011;
assign LUT_1[28591] = 32'b00000000000000000000011010001111;
assign LUT_1[28592] = 32'b00000000000000000110001110011000;
assign LUT_1[28593] = 32'b11111111111111111111100000010100;
assign LUT_1[28594] = 32'b00000000000000000001111100101001;
assign LUT_1[28595] = 32'b11111111111111111011001110100101;
assign LUT_1[28596] = 32'b00000000000000001110000111101111;
assign LUT_1[28597] = 32'b00000000000000000111011001101011;
assign LUT_1[28598] = 32'b00000000000000001001110110000000;
assign LUT_1[28599] = 32'b00000000000000000011000111111100;
assign LUT_1[28600] = 32'b00000000000000000101011100001101;
assign LUT_1[28601] = 32'b11111111111111111110101110001001;
assign LUT_1[28602] = 32'b00000000000000000001001010011110;
assign LUT_1[28603] = 32'b11111111111111111010011100011010;
assign LUT_1[28604] = 32'b00000000000000001101010101100100;
assign LUT_1[28605] = 32'b00000000000000000110100111100000;
assign LUT_1[28606] = 32'b00000000000000001001000011110101;
assign LUT_1[28607] = 32'b00000000000000000010010101110001;
assign LUT_1[28608] = 32'b00000000000000000101010101011111;
assign LUT_1[28609] = 32'b11111111111111111110100111011011;
assign LUT_1[28610] = 32'b00000000000000000001000011110000;
assign LUT_1[28611] = 32'b11111111111111111010010101101100;
assign LUT_1[28612] = 32'b00000000000000001101001110110110;
assign LUT_1[28613] = 32'b00000000000000000110100000110010;
assign LUT_1[28614] = 32'b00000000000000001000111101000111;
assign LUT_1[28615] = 32'b00000000000000000010001111000011;
assign LUT_1[28616] = 32'b00000000000000000100100011010100;
assign LUT_1[28617] = 32'b11111111111111111101110101010000;
assign LUT_1[28618] = 32'b00000000000000000000010001100101;
assign LUT_1[28619] = 32'b11111111111111111001100011100001;
assign LUT_1[28620] = 32'b00000000000000001100011100101011;
assign LUT_1[28621] = 32'b00000000000000000101101110100111;
assign LUT_1[28622] = 32'b00000000000000001000001010111100;
assign LUT_1[28623] = 32'b00000000000000000001011100111000;
assign LUT_1[28624] = 32'b00000000000000000111010001000001;
assign LUT_1[28625] = 32'b00000000000000000000100010111101;
assign LUT_1[28626] = 32'b00000000000000000010111111010010;
assign LUT_1[28627] = 32'b11111111111111111100010001001110;
assign LUT_1[28628] = 32'b00000000000000001111001010011000;
assign LUT_1[28629] = 32'b00000000000000001000011100010100;
assign LUT_1[28630] = 32'b00000000000000001010111000101001;
assign LUT_1[28631] = 32'b00000000000000000100001010100101;
assign LUT_1[28632] = 32'b00000000000000000110011110110110;
assign LUT_1[28633] = 32'b11111111111111111111110000110010;
assign LUT_1[28634] = 32'b00000000000000000010001101000111;
assign LUT_1[28635] = 32'b11111111111111111011011111000011;
assign LUT_1[28636] = 32'b00000000000000001110011000001101;
assign LUT_1[28637] = 32'b00000000000000000111101010001001;
assign LUT_1[28638] = 32'b00000000000000001010000110011110;
assign LUT_1[28639] = 32'b00000000000000000011011000011010;
assign LUT_1[28640] = 32'b00000000000000000110010000011110;
assign LUT_1[28641] = 32'b11111111111111111111100010011010;
assign LUT_1[28642] = 32'b00000000000000000001111110101111;
assign LUT_1[28643] = 32'b11111111111111111011010000101011;
assign LUT_1[28644] = 32'b00000000000000001110001001110101;
assign LUT_1[28645] = 32'b00000000000000000111011011110001;
assign LUT_1[28646] = 32'b00000000000000001001111000000110;
assign LUT_1[28647] = 32'b00000000000000000011001010000010;
assign LUT_1[28648] = 32'b00000000000000000101011110010011;
assign LUT_1[28649] = 32'b11111111111111111110110000001111;
assign LUT_1[28650] = 32'b00000000000000000001001100100100;
assign LUT_1[28651] = 32'b11111111111111111010011110100000;
assign LUT_1[28652] = 32'b00000000000000001101010111101010;
assign LUT_1[28653] = 32'b00000000000000000110101001100110;
assign LUT_1[28654] = 32'b00000000000000001001000101111011;
assign LUT_1[28655] = 32'b00000000000000000010010111110111;
assign LUT_1[28656] = 32'b00000000000000001000001100000000;
assign LUT_1[28657] = 32'b00000000000000000001011101111100;
assign LUT_1[28658] = 32'b00000000000000000011111010010001;
assign LUT_1[28659] = 32'b11111111111111111101001100001101;
assign LUT_1[28660] = 32'b00000000000000010000000101010111;
assign LUT_1[28661] = 32'b00000000000000001001010111010011;
assign LUT_1[28662] = 32'b00000000000000001011110011101000;
assign LUT_1[28663] = 32'b00000000000000000101000101100100;
assign LUT_1[28664] = 32'b00000000000000000111011001110101;
assign LUT_1[28665] = 32'b00000000000000000000101011110001;
assign LUT_1[28666] = 32'b00000000000000000011001000000110;
assign LUT_1[28667] = 32'b11111111111111111100011010000010;
assign LUT_1[28668] = 32'b00000000000000001111010011001100;
assign LUT_1[28669] = 32'b00000000000000001000100101001000;
assign LUT_1[28670] = 32'b00000000000000001011000001011101;
assign LUT_1[28671] = 32'b00000000000000000100010011011001;
assign LUT_1[28672] = 32'b00000000000000000001010001100110;
assign LUT_1[28673] = 32'b11111111111111111010100011100010;
assign LUT_1[28674] = 32'b11111111111111111100111111110111;
assign LUT_1[28675] = 32'b11111111111111110110010001110011;
assign LUT_1[28676] = 32'b00000000000000001001001010111101;
assign LUT_1[28677] = 32'b00000000000000000010011100111001;
assign LUT_1[28678] = 32'b00000000000000000100111001001110;
assign LUT_1[28679] = 32'b11111111111111111110001011001010;
assign LUT_1[28680] = 32'b00000000000000000000011111011011;
assign LUT_1[28681] = 32'b11111111111111111001110001010111;
assign LUT_1[28682] = 32'b11111111111111111100001101101100;
assign LUT_1[28683] = 32'b11111111111111110101011111101000;
assign LUT_1[28684] = 32'b00000000000000001000011000110010;
assign LUT_1[28685] = 32'b00000000000000000001101010101110;
assign LUT_1[28686] = 32'b00000000000000000100000111000011;
assign LUT_1[28687] = 32'b11111111111111111101011000111111;
assign LUT_1[28688] = 32'b00000000000000000011001101001000;
assign LUT_1[28689] = 32'b11111111111111111100011111000100;
assign LUT_1[28690] = 32'b11111111111111111110111011011001;
assign LUT_1[28691] = 32'b11111111111111111000001101010101;
assign LUT_1[28692] = 32'b00000000000000001011000110011111;
assign LUT_1[28693] = 32'b00000000000000000100011000011011;
assign LUT_1[28694] = 32'b00000000000000000110110100110000;
assign LUT_1[28695] = 32'b00000000000000000000000110101100;
assign LUT_1[28696] = 32'b00000000000000000010011010111101;
assign LUT_1[28697] = 32'b11111111111111111011101100111001;
assign LUT_1[28698] = 32'b11111111111111111110001001001110;
assign LUT_1[28699] = 32'b11111111111111110111011011001010;
assign LUT_1[28700] = 32'b00000000000000001010010100010100;
assign LUT_1[28701] = 32'b00000000000000000011100110010000;
assign LUT_1[28702] = 32'b00000000000000000110000010100101;
assign LUT_1[28703] = 32'b11111111111111111111010100100001;
assign LUT_1[28704] = 32'b00000000000000000010001100100101;
assign LUT_1[28705] = 32'b11111111111111111011011110100001;
assign LUT_1[28706] = 32'b11111111111111111101111010110110;
assign LUT_1[28707] = 32'b11111111111111110111001100110010;
assign LUT_1[28708] = 32'b00000000000000001010000101111100;
assign LUT_1[28709] = 32'b00000000000000000011010111111000;
assign LUT_1[28710] = 32'b00000000000000000101110100001101;
assign LUT_1[28711] = 32'b11111111111111111111000110001001;
assign LUT_1[28712] = 32'b00000000000000000001011010011010;
assign LUT_1[28713] = 32'b11111111111111111010101100010110;
assign LUT_1[28714] = 32'b11111111111111111101001000101011;
assign LUT_1[28715] = 32'b11111111111111110110011010100111;
assign LUT_1[28716] = 32'b00000000000000001001010011110001;
assign LUT_1[28717] = 32'b00000000000000000010100101101101;
assign LUT_1[28718] = 32'b00000000000000000101000010000010;
assign LUT_1[28719] = 32'b11111111111111111110010011111110;
assign LUT_1[28720] = 32'b00000000000000000100001000000111;
assign LUT_1[28721] = 32'b11111111111111111101011010000011;
assign LUT_1[28722] = 32'b11111111111111111111110110011000;
assign LUT_1[28723] = 32'b11111111111111111001001000010100;
assign LUT_1[28724] = 32'b00000000000000001100000001011110;
assign LUT_1[28725] = 32'b00000000000000000101010011011010;
assign LUT_1[28726] = 32'b00000000000000000111101111101111;
assign LUT_1[28727] = 32'b00000000000000000001000001101011;
assign LUT_1[28728] = 32'b00000000000000000011010101111100;
assign LUT_1[28729] = 32'b11111111111111111100100111111000;
assign LUT_1[28730] = 32'b11111111111111111111000100001101;
assign LUT_1[28731] = 32'b11111111111111111000010110001001;
assign LUT_1[28732] = 32'b00000000000000001011001111010011;
assign LUT_1[28733] = 32'b00000000000000000100100001001111;
assign LUT_1[28734] = 32'b00000000000000000110111101100100;
assign LUT_1[28735] = 32'b00000000000000000000001111100000;
assign LUT_1[28736] = 32'b00000000000000000011001111001110;
assign LUT_1[28737] = 32'b11111111111111111100100001001010;
assign LUT_1[28738] = 32'b11111111111111111110111101011111;
assign LUT_1[28739] = 32'b11111111111111111000001111011011;
assign LUT_1[28740] = 32'b00000000000000001011001000100101;
assign LUT_1[28741] = 32'b00000000000000000100011010100001;
assign LUT_1[28742] = 32'b00000000000000000110110110110110;
assign LUT_1[28743] = 32'b00000000000000000000001000110010;
assign LUT_1[28744] = 32'b00000000000000000010011101000011;
assign LUT_1[28745] = 32'b11111111111111111011101110111111;
assign LUT_1[28746] = 32'b11111111111111111110001011010100;
assign LUT_1[28747] = 32'b11111111111111110111011101010000;
assign LUT_1[28748] = 32'b00000000000000001010010110011010;
assign LUT_1[28749] = 32'b00000000000000000011101000010110;
assign LUT_1[28750] = 32'b00000000000000000110000100101011;
assign LUT_1[28751] = 32'b11111111111111111111010110100111;
assign LUT_1[28752] = 32'b00000000000000000101001010110000;
assign LUT_1[28753] = 32'b11111111111111111110011100101100;
assign LUT_1[28754] = 32'b00000000000000000000111001000001;
assign LUT_1[28755] = 32'b11111111111111111010001010111101;
assign LUT_1[28756] = 32'b00000000000000001101000100000111;
assign LUT_1[28757] = 32'b00000000000000000110010110000011;
assign LUT_1[28758] = 32'b00000000000000001000110010011000;
assign LUT_1[28759] = 32'b00000000000000000010000100010100;
assign LUT_1[28760] = 32'b00000000000000000100011000100101;
assign LUT_1[28761] = 32'b11111111111111111101101010100001;
assign LUT_1[28762] = 32'b00000000000000000000000110110110;
assign LUT_1[28763] = 32'b11111111111111111001011000110010;
assign LUT_1[28764] = 32'b00000000000000001100010001111100;
assign LUT_1[28765] = 32'b00000000000000000101100011111000;
assign LUT_1[28766] = 32'b00000000000000001000000000001101;
assign LUT_1[28767] = 32'b00000000000000000001010010001001;
assign LUT_1[28768] = 32'b00000000000000000100001010001101;
assign LUT_1[28769] = 32'b11111111111111111101011100001001;
assign LUT_1[28770] = 32'b11111111111111111111111000011110;
assign LUT_1[28771] = 32'b11111111111111111001001010011010;
assign LUT_1[28772] = 32'b00000000000000001100000011100100;
assign LUT_1[28773] = 32'b00000000000000000101010101100000;
assign LUT_1[28774] = 32'b00000000000000000111110001110101;
assign LUT_1[28775] = 32'b00000000000000000001000011110001;
assign LUT_1[28776] = 32'b00000000000000000011011000000010;
assign LUT_1[28777] = 32'b11111111111111111100101001111110;
assign LUT_1[28778] = 32'b11111111111111111111000110010011;
assign LUT_1[28779] = 32'b11111111111111111000011000001111;
assign LUT_1[28780] = 32'b00000000000000001011010001011001;
assign LUT_1[28781] = 32'b00000000000000000100100011010101;
assign LUT_1[28782] = 32'b00000000000000000110111111101010;
assign LUT_1[28783] = 32'b00000000000000000000010001100110;
assign LUT_1[28784] = 32'b00000000000000000110000101101111;
assign LUT_1[28785] = 32'b11111111111111111111010111101011;
assign LUT_1[28786] = 32'b00000000000000000001110100000000;
assign LUT_1[28787] = 32'b11111111111111111011000101111100;
assign LUT_1[28788] = 32'b00000000000000001101111111000110;
assign LUT_1[28789] = 32'b00000000000000000111010001000010;
assign LUT_1[28790] = 32'b00000000000000001001101101010111;
assign LUT_1[28791] = 32'b00000000000000000010111111010011;
assign LUT_1[28792] = 32'b00000000000000000101010011100100;
assign LUT_1[28793] = 32'b11111111111111111110100101100000;
assign LUT_1[28794] = 32'b00000000000000000001000001110101;
assign LUT_1[28795] = 32'b11111111111111111010010011110001;
assign LUT_1[28796] = 32'b00000000000000001101001100111011;
assign LUT_1[28797] = 32'b00000000000000000110011110110111;
assign LUT_1[28798] = 32'b00000000000000001000111011001100;
assign LUT_1[28799] = 32'b00000000000000000010001101001000;
assign LUT_1[28800] = 32'b00000000000000000100010001101001;
assign LUT_1[28801] = 32'b11111111111111111101100011100101;
assign LUT_1[28802] = 32'b11111111111111111111111111111010;
assign LUT_1[28803] = 32'b11111111111111111001010001110110;
assign LUT_1[28804] = 32'b00000000000000001100001011000000;
assign LUT_1[28805] = 32'b00000000000000000101011100111100;
assign LUT_1[28806] = 32'b00000000000000000111111001010001;
assign LUT_1[28807] = 32'b00000000000000000001001011001101;
assign LUT_1[28808] = 32'b00000000000000000011011111011110;
assign LUT_1[28809] = 32'b11111111111111111100110001011010;
assign LUT_1[28810] = 32'b11111111111111111111001101101111;
assign LUT_1[28811] = 32'b11111111111111111000011111101011;
assign LUT_1[28812] = 32'b00000000000000001011011000110101;
assign LUT_1[28813] = 32'b00000000000000000100101010110001;
assign LUT_1[28814] = 32'b00000000000000000111000111000110;
assign LUT_1[28815] = 32'b00000000000000000000011001000010;
assign LUT_1[28816] = 32'b00000000000000000110001101001011;
assign LUT_1[28817] = 32'b11111111111111111111011111000111;
assign LUT_1[28818] = 32'b00000000000000000001111011011100;
assign LUT_1[28819] = 32'b11111111111111111011001101011000;
assign LUT_1[28820] = 32'b00000000000000001110000110100010;
assign LUT_1[28821] = 32'b00000000000000000111011000011110;
assign LUT_1[28822] = 32'b00000000000000001001110100110011;
assign LUT_1[28823] = 32'b00000000000000000011000110101111;
assign LUT_1[28824] = 32'b00000000000000000101011011000000;
assign LUT_1[28825] = 32'b11111111111111111110101100111100;
assign LUT_1[28826] = 32'b00000000000000000001001001010001;
assign LUT_1[28827] = 32'b11111111111111111010011011001101;
assign LUT_1[28828] = 32'b00000000000000001101010100010111;
assign LUT_1[28829] = 32'b00000000000000000110100110010011;
assign LUT_1[28830] = 32'b00000000000000001001000010101000;
assign LUT_1[28831] = 32'b00000000000000000010010100100100;
assign LUT_1[28832] = 32'b00000000000000000101001100101000;
assign LUT_1[28833] = 32'b11111111111111111110011110100100;
assign LUT_1[28834] = 32'b00000000000000000000111010111001;
assign LUT_1[28835] = 32'b11111111111111111010001100110101;
assign LUT_1[28836] = 32'b00000000000000001101000101111111;
assign LUT_1[28837] = 32'b00000000000000000110010111111011;
assign LUT_1[28838] = 32'b00000000000000001000110100010000;
assign LUT_1[28839] = 32'b00000000000000000010000110001100;
assign LUT_1[28840] = 32'b00000000000000000100011010011101;
assign LUT_1[28841] = 32'b11111111111111111101101100011001;
assign LUT_1[28842] = 32'b00000000000000000000001000101110;
assign LUT_1[28843] = 32'b11111111111111111001011010101010;
assign LUT_1[28844] = 32'b00000000000000001100010011110100;
assign LUT_1[28845] = 32'b00000000000000000101100101110000;
assign LUT_1[28846] = 32'b00000000000000001000000010000101;
assign LUT_1[28847] = 32'b00000000000000000001010100000001;
assign LUT_1[28848] = 32'b00000000000000000111001000001010;
assign LUT_1[28849] = 32'b00000000000000000000011010000110;
assign LUT_1[28850] = 32'b00000000000000000010110110011011;
assign LUT_1[28851] = 32'b11111111111111111100001000010111;
assign LUT_1[28852] = 32'b00000000000000001111000001100001;
assign LUT_1[28853] = 32'b00000000000000001000010011011101;
assign LUT_1[28854] = 32'b00000000000000001010101111110010;
assign LUT_1[28855] = 32'b00000000000000000100000001101110;
assign LUT_1[28856] = 32'b00000000000000000110010101111111;
assign LUT_1[28857] = 32'b11111111111111111111100111111011;
assign LUT_1[28858] = 32'b00000000000000000010000100010000;
assign LUT_1[28859] = 32'b11111111111111111011010110001100;
assign LUT_1[28860] = 32'b00000000000000001110001111010110;
assign LUT_1[28861] = 32'b00000000000000000111100001010010;
assign LUT_1[28862] = 32'b00000000000000001001111101100111;
assign LUT_1[28863] = 32'b00000000000000000011001111100011;
assign LUT_1[28864] = 32'b00000000000000000110001111010001;
assign LUT_1[28865] = 32'b11111111111111111111100001001101;
assign LUT_1[28866] = 32'b00000000000000000001111101100010;
assign LUT_1[28867] = 32'b11111111111111111011001111011110;
assign LUT_1[28868] = 32'b00000000000000001110001000101000;
assign LUT_1[28869] = 32'b00000000000000000111011010100100;
assign LUT_1[28870] = 32'b00000000000000001001110110111001;
assign LUT_1[28871] = 32'b00000000000000000011001000110101;
assign LUT_1[28872] = 32'b00000000000000000101011101000110;
assign LUT_1[28873] = 32'b11111111111111111110101111000010;
assign LUT_1[28874] = 32'b00000000000000000001001011010111;
assign LUT_1[28875] = 32'b11111111111111111010011101010011;
assign LUT_1[28876] = 32'b00000000000000001101010110011101;
assign LUT_1[28877] = 32'b00000000000000000110101000011001;
assign LUT_1[28878] = 32'b00000000000000001001000100101110;
assign LUT_1[28879] = 32'b00000000000000000010010110101010;
assign LUT_1[28880] = 32'b00000000000000001000001010110011;
assign LUT_1[28881] = 32'b00000000000000000001011100101111;
assign LUT_1[28882] = 32'b00000000000000000011111001000100;
assign LUT_1[28883] = 32'b11111111111111111101001011000000;
assign LUT_1[28884] = 32'b00000000000000010000000100001010;
assign LUT_1[28885] = 32'b00000000000000001001010110000110;
assign LUT_1[28886] = 32'b00000000000000001011110010011011;
assign LUT_1[28887] = 32'b00000000000000000101000100010111;
assign LUT_1[28888] = 32'b00000000000000000111011000101000;
assign LUT_1[28889] = 32'b00000000000000000000101010100100;
assign LUT_1[28890] = 32'b00000000000000000011000110111001;
assign LUT_1[28891] = 32'b11111111111111111100011000110101;
assign LUT_1[28892] = 32'b00000000000000001111010001111111;
assign LUT_1[28893] = 32'b00000000000000001000100011111011;
assign LUT_1[28894] = 32'b00000000000000001011000000010000;
assign LUT_1[28895] = 32'b00000000000000000100010010001100;
assign LUT_1[28896] = 32'b00000000000000000111001010010000;
assign LUT_1[28897] = 32'b00000000000000000000011100001100;
assign LUT_1[28898] = 32'b00000000000000000010111000100001;
assign LUT_1[28899] = 32'b11111111111111111100001010011101;
assign LUT_1[28900] = 32'b00000000000000001111000011100111;
assign LUT_1[28901] = 32'b00000000000000001000010101100011;
assign LUT_1[28902] = 32'b00000000000000001010110001111000;
assign LUT_1[28903] = 32'b00000000000000000100000011110100;
assign LUT_1[28904] = 32'b00000000000000000110011000000101;
assign LUT_1[28905] = 32'b11111111111111111111101010000001;
assign LUT_1[28906] = 32'b00000000000000000010000110010110;
assign LUT_1[28907] = 32'b11111111111111111011011000010010;
assign LUT_1[28908] = 32'b00000000000000001110010001011100;
assign LUT_1[28909] = 32'b00000000000000000111100011011000;
assign LUT_1[28910] = 32'b00000000000000001001111111101101;
assign LUT_1[28911] = 32'b00000000000000000011010001101001;
assign LUT_1[28912] = 32'b00000000000000001001000101110010;
assign LUT_1[28913] = 32'b00000000000000000010010111101110;
assign LUT_1[28914] = 32'b00000000000000000100110100000011;
assign LUT_1[28915] = 32'b11111111111111111110000101111111;
assign LUT_1[28916] = 32'b00000000000000010000111111001001;
assign LUT_1[28917] = 32'b00000000000000001010010001000101;
assign LUT_1[28918] = 32'b00000000000000001100101101011010;
assign LUT_1[28919] = 32'b00000000000000000101111111010110;
assign LUT_1[28920] = 32'b00000000000000001000010011100111;
assign LUT_1[28921] = 32'b00000000000000000001100101100011;
assign LUT_1[28922] = 32'b00000000000000000100000001111000;
assign LUT_1[28923] = 32'b11111111111111111101010011110100;
assign LUT_1[28924] = 32'b00000000000000010000001100111110;
assign LUT_1[28925] = 32'b00000000000000001001011110111010;
assign LUT_1[28926] = 32'b00000000000000001011111011001111;
assign LUT_1[28927] = 32'b00000000000000000101001101001011;
assign LUT_1[28928] = 32'b11111111111111111111000101110010;
assign LUT_1[28929] = 32'b11111111111111111000010111101110;
assign LUT_1[28930] = 32'b11111111111111111010110100000011;
assign LUT_1[28931] = 32'b11111111111111110100000101111111;
assign LUT_1[28932] = 32'b00000000000000000110111111001001;
assign LUT_1[28933] = 32'b00000000000000000000010001000101;
assign LUT_1[28934] = 32'b00000000000000000010101101011010;
assign LUT_1[28935] = 32'b11111111111111111011111111010110;
assign LUT_1[28936] = 32'b11111111111111111110010011100111;
assign LUT_1[28937] = 32'b11111111111111110111100101100011;
assign LUT_1[28938] = 32'b11111111111111111010000001111000;
assign LUT_1[28939] = 32'b11111111111111110011010011110100;
assign LUT_1[28940] = 32'b00000000000000000110001100111110;
assign LUT_1[28941] = 32'b11111111111111111111011110111010;
assign LUT_1[28942] = 32'b00000000000000000001111011001111;
assign LUT_1[28943] = 32'b11111111111111111011001101001011;
assign LUT_1[28944] = 32'b00000000000000000001000001010100;
assign LUT_1[28945] = 32'b11111111111111111010010011010000;
assign LUT_1[28946] = 32'b11111111111111111100101111100101;
assign LUT_1[28947] = 32'b11111111111111110110000001100001;
assign LUT_1[28948] = 32'b00000000000000001000111010101011;
assign LUT_1[28949] = 32'b00000000000000000010001100100111;
assign LUT_1[28950] = 32'b00000000000000000100101000111100;
assign LUT_1[28951] = 32'b11111111111111111101111010111000;
assign LUT_1[28952] = 32'b00000000000000000000001111001001;
assign LUT_1[28953] = 32'b11111111111111111001100001000101;
assign LUT_1[28954] = 32'b11111111111111111011111101011010;
assign LUT_1[28955] = 32'b11111111111111110101001111010110;
assign LUT_1[28956] = 32'b00000000000000001000001000100000;
assign LUT_1[28957] = 32'b00000000000000000001011010011100;
assign LUT_1[28958] = 32'b00000000000000000011110110110001;
assign LUT_1[28959] = 32'b11111111111111111101001000101101;
assign LUT_1[28960] = 32'b00000000000000000000000000110001;
assign LUT_1[28961] = 32'b11111111111111111001010010101101;
assign LUT_1[28962] = 32'b11111111111111111011101111000010;
assign LUT_1[28963] = 32'b11111111111111110101000000111110;
assign LUT_1[28964] = 32'b00000000000000000111111010001000;
assign LUT_1[28965] = 32'b00000000000000000001001100000100;
assign LUT_1[28966] = 32'b00000000000000000011101000011001;
assign LUT_1[28967] = 32'b11111111111111111100111010010101;
assign LUT_1[28968] = 32'b11111111111111111111001110100110;
assign LUT_1[28969] = 32'b11111111111111111000100000100010;
assign LUT_1[28970] = 32'b11111111111111111010111100110111;
assign LUT_1[28971] = 32'b11111111111111110100001110110011;
assign LUT_1[28972] = 32'b00000000000000000111000111111101;
assign LUT_1[28973] = 32'b00000000000000000000011001111001;
assign LUT_1[28974] = 32'b00000000000000000010110110001110;
assign LUT_1[28975] = 32'b11111111111111111100001000001010;
assign LUT_1[28976] = 32'b00000000000000000001111100010011;
assign LUT_1[28977] = 32'b11111111111111111011001110001111;
assign LUT_1[28978] = 32'b11111111111111111101101010100100;
assign LUT_1[28979] = 32'b11111111111111110110111100100000;
assign LUT_1[28980] = 32'b00000000000000001001110101101010;
assign LUT_1[28981] = 32'b00000000000000000011000111100110;
assign LUT_1[28982] = 32'b00000000000000000101100011111011;
assign LUT_1[28983] = 32'b11111111111111111110110101110111;
assign LUT_1[28984] = 32'b00000000000000000001001010001000;
assign LUT_1[28985] = 32'b11111111111111111010011100000100;
assign LUT_1[28986] = 32'b11111111111111111100111000011001;
assign LUT_1[28987] = 32'b11111111111111110110001010010101;
assign LUT_1[28988] = 32'b00000000000000001001000011011111;
assign LUT_1[28989] = 32'b00000000000000000010010101011011;
assign LUT_1[28990] = 32'b00000000000000000100110001110000;
assign LUT_1[28991] = 32'b11111111111111111110000011101100;
assign LUT_1[28992] = 32'b00000000000000000001000011011010;
assign LUT_1[28993] = 32'b11111111111111111010010101010110;
assign LUT_1[28994] = 32'b11111111111111111100110001101011;
assign LUT_1[28995] = 32'b11111111111111110110000011100111;
assign LUT_1[28996] = 32'b00000000000000001000111100110001;
assign LUT_1[28997] = 32'b00000000000000000010001110101101;
assign LUT_1[28998] = 32'b00000000000000000100101011000010;
assign LUT_1[28999] = 32'b11111111111111111101111100111110;
assign LUT_1[29000] = 32'b00000000000000000000010001001111;
assign LUT_1[29001] = 32'b11111111111111111001100011001011;
assign LUT_1[29002] = 32'b11111111111111111011111111100000;
assign LUT_1[29003] = 32'b11111111111111110101010001011100;
assign LUT_1[29004] = 32'b00000000000000001000001010100110;
assign LUT_1[29005] = 32'b00000000000000000001011100100010;
assign LUT_1[29006] = 32'b00000000000000000011111000110111;
assign LUT_1[29007] = 32'b11111111111111111101001010110011;
assign LUT_1[29008] = 32'b00000000000000000010111110111100;
assign LUT_1[29009] = 32'b11111111111111111100010000111000;
assign LUT_1[29010] = 32'b11111111111111111110101101001101;
assign LUT_1[29011] = 32'b11111111111111110111111111001001;
assign LUT_1[29012] = 32'b00000000000000001010111000010011;
assign LUT_1[29013] = 32'b00000000000000000100001010001111;
assign LUT_1[29014] = 32'b00000000000000000110100110100100;
assign LUT_1[29015] = 32'b11111111111111111111111000100000;
assign LUT_1[29016] = 32'b00000000000000000010001100110001;
assign LUT_1[29017] = 32'b11111111111111111011011110101101;
assign LUT_1[29018] = 32'b11111111111111111101111011000010;
assign LUT_1[29019] = 32'b11111111111111110111001100111110;
assign LUT_1[29020] = 32'b00000000000000001010000110001000;
assign LUT_1[29021] = 32'b00000000000000000011011000000100;
assign LUT_1[29022] = 32'b00000000000000000101110100011001;
assign LUT_1[29023] = 32'b11111111111111111111000110010101;
assign LUT_1[29024] = 32'b00000000000000000001111110011001;
assign LUT_1[29025] = 32'b11111111111111111011010000010101;
assign LUT_1[29026] = 32'b11111111111111111101101100101010;
assign LUT_1[29027] = 32'b11111111111111110110111110100110;
assign LUT_1[29028] = 32'b00000000000000001001110111110000;
assign LUT_1[29029] = 32'b00000000000000000011001001101100;
assign LUT_1[29030] = 32'b00000000000000000101100110000001;
assign LUT_1[29031] = 32'b11111111111111111110110111111101;
assign LUT_1[29032] = 32'b00000000000000000001001100001110;
assign LUT_1[29033] = 32'b11111111111111111010011110001010;
assign LUT_1[29034] = 32'b11111111111111111100111010011111;
assign LUT_1[29035] = 32'b11111111111111110110001100011011;
assign LUT_1[29036] = 32'b00000000000000001001000101100101;
assign LUT_1[29037] = 32'b00000000000000000010010111100001;
assign LUT_1[29038] = 32'b00000000000000000100110011110110;
assign LUT_1[29039] = 32'b11111111111111111110000101110010;
assign LUT_1[29040] = 32'b00000000000000000011111001111011;
assign LUT_1[29041] = 32'b11111111111111111101001011110111;
assign LUT_1[29042] = 32'b11111111111111111111101000001100;
assign LUT_1[29043] = 32'b11111111111111111000111010001000;
assign LUT_1[29044] = 32'b00000000000000001011110011010010;
assign LUT_1[29045] = 32'b00000000000000000101000101001110;
assign LUT_1[29046] = 32'b00000000000000000111100001100011;
assign LUT_1[29047] = 32'b00000000000000000000110011011111;
assign LUT_1[29048] = 32'b00000000000000000011000111110000;
assign LUT_1[29049] = 32'b11111111111111111100011001101100;
assign LUT_1[29050] = 32'b11111111111111111110110110000001;
assign LUT_1[29051] = 32'b11111111111111111000000111111101;
assign LUT_1[29052] = 32'b00000000000000001011000001000111;
assign LUT_1[29053] = 32'b00000000000000000100010011000011;
assign LUT_1[29054] = 32'b00000000000000000110101111011000;
assign LUT_1[29055] = 32'b00000000000000000000000001010100;
assign LUT_1[29056] = 32'b00000000000000000010000101110101;
assign LUT_1[29057] = 32'b11111111111111111011010111110001;
assign LUT_1[29058] = 32'b11111111111111111101110100000110;
assign LUT_1[29059] = 32'b11111111111111110111000110000010;
assign LUT_1[29060] = 32'b00000000000000001001111111001100;
assign LUT_1[29061] = 32'b00000000000000000011010001001000;
assign LUT_1[29062] = 32'b00000000000000000101101101011101;
assign LUT_1[29063] = 32'b11111111111111111110111111011001;
assign LUT_1[29064] = 32'b00000000000000000001010011101010;
assign LUT_1[29065] = 32'b11111111111111111010100101100110;
assign LUT_1[29066] = 32'b11111111111111111101000001111011;
assign LUT_1[29067] = 32'b11111111111111110110010011110111;
assign LUT_1[29068] = 32'b00000000000000001001001101000001;
assign LUT_1[29069] = 32'b00000000000000000010011110111101;
assign LUT_1[29070] = 32'b00000000000000000100111011010010;
assign LUT_1[29071] = 32'b11111111111111111110001101001110;
assign LUT_1[29072] = 32'b00000000000000000100000001010111;
assign LUT_1[29073] = 32'b11111111111111111101010011010011;
assign LUT_1[29074] = 32'b11111111111111111111101111101000;
assign LUT_1[29075] = 32'b11111111111111111001000001100100;
assign LUT_1[29076] = 32'b00000000000000001011111010101110;
assign LUT_1[29077] = 32'b00000000000000000101001100101010;
assign LUT_1[29078] = 32'b00000000000000000111101000111111;
assign LUT_1[29079] = 32'b00000000000000000000111010111011;
assign LUT_1[29080] = 32'b00000000000000000011001111001100;
assign LUT_1[29081] = 32'b11111111111111111100100001001000;
assign LUT_1[29082] = 32'b11111111111111111110111101011101;
assign LUT_1[29083] = 32'b11111111111111111000001111011001;
assign LUT_1[29084] = 32'b00000000000000001011001000100011;
assign LUT_1[29085] = 32'b00000000000000000100011010011111;
assign LUT_1[29086] = 32'b00000000000000000110110110110100;
assign LUT_1[29087] = 32'b00000000000000000000001000110000;
assign LUT_1[29088] = 32'b00000000000000000011000000110100;
assign LUT_1[29089] = 32'b11111111111111111100010010110000;
assign LUT_1[29090] = 32'b11111111111111111110101111000101;
assign LUT_1[29091] = 32'b11111111111111111000000001000001;
assign LUT_1[29092] = 32'b00000000000000001010111010001011;
assign LUT_1[29093] = 32'b00000000000000000100001100000111;
assign LUT_1[29094] = 32'b00000000000000000110101000011100;
assign LUT_1[29095] = 32'b11111111111111111111111010011000;
assign LUT_1[29096] = 32'b00000000000000000010001110101001;
assign LUT_1[29097] = 32'b11111111111111111011100000100101;
assign LUT_1[29098] = 32'b11111111111111111101111100111010;
assign LUT_1[29099] = 32'b11111111111111110111001110110110;
assign LUT_1[29100] = 32'b00000000000000001010001000000000;
assign LUT_1[29101] = 32'b00000000000000000011011001111100;
assign LUT_1[29102] = 32'b00000000000000000101110110010001;
assign LUT_1[29103] = 32'b11111111111111111111001000001101;
assign LUT_1[29104] = 32'b00000000000000000100111100010110;
assign LUT_1[29105] = 32'b11111111111111111110001110010010;
assign LUT_1[29106] = 32'b00000000000000000000101010100111;
assign LUT_1[29107] = 32'b11111111111111111001111100100011;
assign LUT_1[29108] = 32'b00000000000000001100110101101101;
assign LUT_1[29109] = 32'b00000000000000000110000111101001;
assign LUT_1[29110] = 32'b00000000000000001000100011111110;
assign LUT_1[29111] = 32'b00000000000000000001110101111010;
assign LUT_1[29112] = 32'b00000000000000000100001010001011;
assign LUT_1[29113] = 32'b11111111111111111101011100000111;
assign LUT_1[29114] = 32'b11111111111111111111111000011100;
assign LUT_1[29115] = 32'b11111111111111111001001010011000;
assign LUT_1[29116] = 32'b00000000000000001100000011100010;
assign LUT_1[29117] = 32'b00000000000000000101010101011110;
assign LUT_1[29118] = 32'b00000000000000000111110001110011;
assign LUT_1[29119] = 32'b00000000000000000001000011101111;
assign LUT_1[29120] = 32'b00000000000000000100000011011101;
assign LUT_1[29121] = 32'b11111111111111111101010101011001;
assign LUT_1[29122] = 32'b11111111111111111111110001101110;
assign LUT_1[29123] = 32'b11111111111111111001000011101010;
assign LUT_1[29124] = 32'b00000000000000001011111100110100;
assign LUT_1[29125] = 32'b00000000000000000101001110110000;
assign LUT_1[29126] = 32'b00000000000000000111101011000101;
assign LUT_1[29127] = 32'b00000000000000000000111101000001;
assign LUT_1[29128] = 32'b00000000000000000011010001010010;
assign LUT_1[29129] = 32'b11111111111111111100100011001110;
assign LUT_1[29130] = 32'b11111111111111111110111111100011;
assign LUT_1[29131] = 32'b11111111111111111000010001011111;
assign LUT_1[29132] = 32'b00000000000000001011001010101001;
assign LUT_1[29133] = 32'b00000000000000000100011100100101;
assign LUT_1[29134] = 32'b00000000000000000110111000111010;
assign LUT_1[29135] = 32'b00000000000000000000001010110110;
assign LUT_1[29136] = 32'b00000000000000000101111110111111;
assign LUT_1[29137] = 32'b11111111111111111111010000111011;
assign LUT_1[29138] = 32'b00000000000000000001101101010000;
assign LUT_1[29139] = 32'b11111111111111111010111111001100;
assign LUT_1[29140] = 32'b00000000000000001101111000010110;
assign LUT_1[29141] = 32'b00000000000000000111001010010010;
assign LUT_1[29142] = 32'b00000000000000001001100110100111;
assign LUT_1[29143] = 32'b00000000000000000010111000100011;
assign LUT_1[29144] = 32'b00000000000000000101001100110100;
assign LUT_1[29145] = 32'b11111111111111111110011110110000;
assign LUT_1[29146] = 32'b00000000000000000000111011000101;
assign LUT_1[29147] = 32'b11111111111111111010001101000001;
assign LUT_1[29148] = 32'b00000000000000001101000110001011;
assign LUT_1[29149] = 32'b00000000000000000110011000000111;
assign LUT_1[29150] = 32'b00000000000000001000110100011100;
assign LUT_1[29151] = 32'b00000000000000000010000110011000;
assign LUT_1[29152] = 32'b00000000000000000100111110011100;
assign LUT_1[29153] = 32'b11111111111111111110010000011000;
assign LUT_1[29154] = 32'b00000000000000000000101100101101;
assign LUT_1[29155] = 32'b11111111111111111001111110101001;
assign LUT_1[29156] = 32'b00000000000000001100110111110011;
assign LUT_1[29157] = 32'b00000000000000000110001001101111;
assign LUT_1[29158] = 32'b00000000000000001000100110000100;
assign LUT_1[29159] = 32'b00000000000000000001111000000000;
assign LUT_1[29160] = 32'b00000000000000000100001100010001;
assign LUT_1[29161] = 32'b11111111111111111101011110001101;
assign LUT_1[29162] = 32'b11111111111111111111111010100010;
assign LUT_1[29163] = 32'b11111111111111111001001100011110;
assign LUT_1[29164] = 32'b00000000000000001100000101101000;
assign LUT_1[29165] = 32'b00000000000000000101010111100100;
assign LUT_1[29166] = 32'b00000000000000000111110011111001;
assign LUT_1[29167] = 32'b00000000000000000001000101110101;
assign LUT_1[29168] = 32'b00000000000000000110111001111110;
assign LUT_1[29169] = 32'b00000000000000000000001011111010;
assign LUT_1[29170] = 32'b00000000000000000010101000001111;
assign LUT_1[29171] = 32'b11111111111111111011111010001011;
assign LUT_1[29172] = 32'b00000000000000001110110011010101;
assign LUT_1[29173] = 32'b00000000000000001000000101010001;
assign LUT_1[29174] = 32'b00000000000000001010100001100110;
assign LUT_1[29175] = 32'b00000000000000000011110011100010;
assign LUT_1[29176] = 32'b00000000000000000110000111110011;
assign LUT_1[29177] = 32'b11111111111111111111011001101111;
assign LUT_1[29178] = 32'b00000000000000000001110110000100;
assign LUT_1[29179] = 32'b11111111111111111011001000000000;
assign LUT_1[29180] = 32'b00000000000000001110000001001010;
assign LUT_1[29181] = 32'b00000000000000000111010011000110;
assign LUT_1[29182] = 32'b00000000000000001001101111011011;
assign LUT_1[29183] = 32'b00000000000000000011000001010111;
assign LUT_1[29184] = 32'b11111111111111111011000000000011;
assign LUT_1[29185] = 32'b11111111111111110100010001111111;
assign LUT_1[29186] = 32'b11111111111111110110101110010100;
assign LUT_1[29187] = 32'b11111111111111110000000000010000;
assign LUT_1[29188] = 32'b00000000000000000010111001011010;
assign LUT_1[29189] = 32'b11111111111111111100001011010110;
assign LUT_1[29190] = 32'b11111111111111111110100111101011;
assign LUT_1[29191] = 32'b11111111111111110111111001100111;
assign LUT_1[29192] = 32'b11111111111111111010001101111000;
assign LUT_1[29193] = 32'b11111111111111110011011111110100;
assign LUT_1[29194] = 32'b11111111111111110101111100001001;
assign LUT_1[29195] = 32'b11111111111111101111001110000101;
assign LUT_1[29196] = 32'b00000000000000000010000111001111;
assign LUT_1[29197] = 32'b11111111111111111011011001001011;
assign LUT_1[29198] = 32'b11111111111111111101110101100000;
assign LUT_1[29199] = 32'b11111111111111110111000111011100;
assign LUT_1[29200] = 32'b11111111111111111100111011100101;
assign LUT_1[29201] = 32'b11111111111111110110001101100001;
assign LUT_1[29202] = 32'b11111111111111111000101001110110;
assign LUT_1[29203] = 32'b11111111111111110001111011110010;
assign LUT_1[29204] = 32'b00000000000000000100110100111100;
assign LUT_1[29205] = 32'b11111111111111111110000110111000;
assign LUT_1[29206] = 32'b00000000000000000000100011001101;
assign LUT_1[29207] = 32'b11111111111111111001110101001001;
assign LUT_1[29208] = 32'b11111111111111111100001001011010;
assign LUT_1[29209] = 32'b11111111111111110101011011010110;
assign LUT_1[29210] = 32'b11111111111111110111110111101011;
assign LUT_1[29211] = 32'b11111111111111110001001001100111;
assign LUT_1[29212] = 32'b00000000000000000100000010110001;
assign LUT_1[29213] = 32'b11111111111111111101010100101101;
assign LUT_1[29214] = 32'b11111111111111111111110001000010;
assign LUT_1[29215] = 32'b11111111111111111001000010111110;
assign LUT_1[29216] = 32'b11111111111111111011111011000010;
assign LUT_1[29217] = 32'b11111111111111110101001100111110;
assign LUT_1[29218] = 32'b11111111111111110111101001010011;
assign LUT_1[29219] = 32'b11111111111111110000111011001111;
assign LUT_1[29220] = 32'b00000000000000000011110100011001;
assign LUT_1[29221] = 32'b11111111111111111101000110010101;
assign LUT_1[29222] = 32'b11111111111111111111100010101010;
assign LUT_1[29223] = 32'b11111111111111111000110100100110;
assign LUT_1[29224] = 32'b11111111111111111011001000110111;
assign LUT_1[29225] = 32'b11111111111111110100011010110011;
assign LUT_1[29226] = 32'b11111111111111110110110111001000;
assign LUT_1[29227] = 32'b11111111111111110000001001000100;
assign LUT_1[29228] = 32'b00000000000000000011000010001110;
assign LUT_1[29229] = 32'b11111111111111111100010100001010;
assign LUT_1[29230] = 32'b11111111111111111110110000011111;
assign LUT_1[29231] = 32'b11111111111111111000000010011011;
assign LUT_1[29232] = 32'b11111111111111111101110110100100;
assign LUT_1[29233] = 32'b11111111111111110111001000100000;
assign LUT_1[29234] = 32'b11111111111111111001100100110101;
assign LUT_1[29235] = 32'b11111111111111110010110110110001;
assign LUT_1[29236] = 32'b00000000000000000101101111111011;
assign LUT_1[29237] = 32'b11111111111111111111000001110111;
assign LUT_1[29238] = 32'b00000000000000000001011110001100;
assign LUT_1[29239] = 32'b11111111111111111010110000001000;
assign LUT_1[29240] = 32'b11111111111111111101000100011001;
assign LUT_1[29241] = 32'b11111111111111110110010110010101;
assign LUT_1[29242] = 32'b11111111111111111000110010101010;
assign LUT_1[29243] = 32'b11111111111111110010000100100110;
assign LUT_1[29244] = 32'b00000000000000000100111101110000;
assign LUT_1[29245] = 32'b11111111111111111110001111101100;
assign LUT_1[29246] = 32'b00000000000000000000101100000001;
assign LUT_1[29247] = 32'b11111111111111111001111101111101;
assign LUT_1[29248] = 32'b11111111111111111100111101101011;
assign LUT_1[29249] = 32'b11111111111111110110001111100111;
assign LUT_1[29250] = 32'b11111111111111111000101011111100;
assign LUT_1[29251] = 32'b11111111111111110001111101111000;
assign LUT_1[29252] = 32'b00000000000000000100110111000010;
assign LUT_1[29253] = 32'b11111111111111111110001000111110;
assign LUT_1[29254] = 32'b00000000000000000000100101010011;
assign LUT_1[29255] = 32'b11111111111111111001110111001111;
assign LUT_1[29256] = 32'b11111111111111111100001011100000;
assign LUT_1[29257] = 32'b11111111111111110101011101011100;
assign LUT_1[29258] = 32'b11111111111111110111111001110001;
assign LUT_1[29259] = 32'b11111111111111110001001011101101;
assign LUT_1[29260] = 32'b00000000000000000100000100110111;
assign LUT_1[29261] = 32'b11111111111111111101010110110011;
assign LUT_1[29262] = 32'b11111111111111111111110011001000;
assign LUT_1[29263] = 32'b11111111111111111001000101000100;
assign LUT_1[29264] = 32'b11111111111111111110111001001101;
assign LUT_1[29265] = 32'b11111111111111111000001011001001;
assign LUT_1[29266] = 32'b11111111111111111010100111011110;
assign LUT_1[29267] = 32'b11111111111111110011111001011010;
assign LUT_1[29268] = 32'b00000000000000000110110010100100;
assign LUT_1[29269] = 32'b00000000000000000000000100100000;
assign LUT_1[29270] = 32'b00000000000000000010100000110101;
assign LUT_1[29271] = 32'b11111111111111111011110010110001;
assign LUT_1[29272] = 32'b11111111111111111110000111000010;
assign LUT_1[29273] = 32'b11111111111111110111011000111110;
assign LUT_1[29274] = 32'b11111111111111111001110101010011;
assign LUT_1[29275] = 32'b11111111111111110011000111001111;
assign LUT_1[29276] = 32'b00000000000000000110000000011001;
assign LUT_1[29277] = 32'b11111111111111111111010010010101;
assign LUT_1[29278] = 32'b00000000000000000001101110101010;
assign LUT_1[29279] = 32'b11111111111111111011000000100110;
assign LUT_1[29280] = 32'b11111111111111111101111000101010;
assign LUT_1[29281] = 32'b11111111111111110111001010100110;
assign LUT_1[29282] = 32'b11111111111111111001100110111011;
assign LUT_1[29283] = 32'b11111111111111110010111000110111;
assign LUT_1[29284] = 32'b00000000000000000101110010000001;
assign LUT_1[29285] = 32'b11111111111111111111000011111101;
assign LUT_1[29286] = 32'b00000000000000000001100000010010;
assign LUT_1[29287] = 32'b11111111111111111010110010001110;
assign LUT_1[29288] = 32'b11111111111111111101000110011111;
assign LUT_1[29289] = 32'b11111111111111110110011000011011;
assign LUT_1[29290] = 32'b11111111111111111000110100110000;
assign LUT_1[29291] = 32'b11111111111111110010000110101100;
assign LUT_1[29292] = 32'b00000000000000000100111111110110;
assign LUT_1[29293] = 32'b11111111111111111110010001110010;
assign LUT_1[29294] = 32'b00000000000000000000101110000111;
assign LUT_1[29295] = 32'b11111111111111111010000000000011;
assign LUT_1[29296] = 32'b11111111111111111111110100001100;
assign LUT_1[29297] = 32'b11111111111111111001000110001000;
assign LUT_1[29298] = 32'b11111111111111111011100010011101;
assign LUT_1[29299] = 32'b11111111111111110100110100011001;
assign LUT_1[29300] = 32'b00000000000000000111101101100011;
assign LUT_1[29301] = 32'b00000000000000000000111111011111;
assign LUT_1[29302] = 32'b00000000000000000011011011110100;
assign LUT_1[29303] = 32'b11111111111111111100101101110000;
assign LUT_1[29304] = 32'b11111111111111111111000010000001;
assign LUT_1[29305] = 32'b11111111111111111000010011111101;
assign LUT_1[29306] = 32'b11111111111111111010110000010010;
assign LUT_1[29307] = 32'b11111111111111110100000010001110;
assign LUT_1[29308] = 32'b00000000000000000110111011011000;
assign LUT_1[29309] = 32'b00000000000000000000001101010100;
assign LUT_1[29310] = 32'b00000000000000000010101001101001;
assign LUT_1[29311] = 32'b11111111111111111011111011100101;
assign LUT_1[29312] = 32'b11111111111111111110000000000110;
assign LUT_1[29313] = 32'b11111111111111110111010010000010;
assign LUT_1[29314] = 32'b11111111111111111001101110010111;
assign LUT_1[29315] = 32'b11111111111111110011000000010011;
assign LUT_1[29316] = 32'b00000000000000000101111001011101;
assign LUT_1[29317] = 32'b11111111111111111111001011011001;
assign LUT_1[29318] = 32'b00000000000000000001100111101110;
assign LUT_1[29319] = 32'b11111111111111111010111001101010;
assign LUT_1[29320] = 32'b11111111111111111101001101111011;
assign LUT_1[29321] = 32'b11111111111111110110011111110111;
assign LUT_1[29322] = 32'b11111111111111111000111100001100;
assign LUT_1[29323] = 32'b11111111111111110010001110001000;
assign LUT_1[29324] = 32'b00000000000000000101000111010010;
assign LUT_1[29325] = 32'b11111111111111111110011001001110;
assign LUT_1[29326] = 32'b00000000000000000000110101100011;
assign LUT_1[29327] = 32'b11111111111111111010000111011111;
assign LUT_1[29328] = 32'b11111111111111111111111011101000;
assign LUT_1[29329] = 32'b11111111111111111001001101100100;
assign LUT_1[29330] = 32'b11111111111111111011101001111001;
assign LUT_1[29331] = 32'b11111111111111110100111011110101;
assign LUT_1[29332] = 32'b00000000000000000111110100111111;
assign LUT_1[29333] = 32'b00000000000000000001000110111011;
assign LUT_1[29334] = 32'b00000000000000000011100011010000;
assign LUT_1[29335] = 32'b11111111111111111100110101001100;
assign LUT_1[29336] = 32'b11111111111111111111001001011101;
assign LUT_1[29337] = 32'b11111111111111111000011011011001;
assign LUT_1[29338] = 32'b11111111111111111010110111101110;
assign LUT_1[29339] = 32'b11111111111111110100001001101010;
assign LUT_1[29340] = 32'b00000000000000000111000010110100;
assign LUT_1[29341] = 32'b00000000000000000000010100110000;
assign LUT_1[29342] = 32'b00000000000000000010110001000101;
assign LUT_1[29343] = 32'b11111111111111111100000011000001;
assign LUT_1[29344] = 32'b11111111111111111110111011000101;
assign LUT_1[29345] = 32'b11111111111111111000001101000001;
assign LUT_1[29346] = 32'b11111111111111111010101001010110;
assign LUT_1[29347] = 32'b11111111111111110011111011010010;
assign LUT_1[29348] = 32'b00000000000000000110110100011100;
assign LUT_1[29349] = 32'b00000000000000000000000110011000;
assign LUT_1[29350] = 32'b00000000000000000010100010101101;
assign LUT_1[29351] = 32'b11111111111111111011110100101001;
assign LUT_1[29352] = 32'b11111111111111111110001000111010;
assign LUT_1[29353] = 32'b11111111111111110111011010110110;
assign LUT_1[29354] = 32'b11111111111111111001110111001011;
assign LUT_1[29355] = 32'b11111111111111110011001001000111;
assign LUT_1[29356] = 32'b00000000000000000110000010010001;
assign LUT_1[29357] = 32'b11111111111111111111010100001101;
assign LUT_1[29358] = 32'b00000000000000000001110000100010;
assign LUT_1[29359] = 32'b11111111111111111011000010011110;
assign LUT_1[29360] = 32'b00000000000000000000110110100111;
assign LUT_1[29361] = 32'b11111111111111111010001000100011;
assign LUT_1[29362] = 32'b11111111111111111100100100111000;
assign LUT_1[29363] = 32'b11111111111111110101110110110100;
assign LUT_1[29364] = 32'b00000000000000001000101111111110;
assign LUT_1[29365] = 32'b00000000000000000010000001111010;
assign LUT_1[29366] = 32'b00000000000000000100011110001111;
assign LUT_1[29367] = 32'b11111111111111111101110000001011;
assign LUT_1[29368] = 32'b00000000000000000000000100011100;
assign LUT_1[29369] = 32'b11111111111111111001010110011000;
assign LUT_1[29370] = 32'b11111111111111111011110010101101;
assign LUT_1[29371] = 32'b11111111111111110101000100101001;
assign LUT_1[29372] = 32'b00000000000000000111111101110011;
assign LUT_1[29373] = 32'b00000000000000000001001111101111;
assign LUT_1[29374] = 32'b00000000000000000011101100000100;
assign LUT_1[29375] = 32'b11111111111111111100111110000000;
assign LUT_1[29376] = 32'b11111111111111111111111101101110;
assign LUT_1[29377] = 32'b11111111111111111001001111101010;
assign LUT_1[29378] = 32'b11111111111111111011101011111111;
assign LUT_1[29379] = 32'b11111111111111110100111101111011;
assign LUT_1[29380] = 32'b00000000000000000111110111000101;
assign LUT_1[29381] = 32'b00000000000000000001001001000001;
assign LUT_1[29382] = 32'b00000000000000000011100101010110;
assign LUT_1[29383] = 32'b11111111111111111100110111010010;
assign LUT_1[29384] = 32'b11111111111111111111001011100011;
assign LUT_1[29385] = 32'b11111111111111111000011101011111;
assign LUT_1[29386] = 32'b11111111111111111010111001110100;
assign LUT_1[29387] = 32'b11111111111111110100001011110000;
assign LUT_1[29388] = 32'b00000000000000000111000100111010;
assign LUT_1[29389] = 32'b00000000000000000000010110110110;
assign LUT_1[29390] = 32'b00000000000000000010110011001011;
assign LUT_1[29391] = 32'b11111111111111111100000101000111;
assign LUT_1[29392] = 32'b00000000000000000001111001010000;
assign LUT_1[29393] = 32'b11111111111111111011001011001100;
assign LUT_1[29394] = 32'b11111111111111111101100111100001;
assign LUT_1[29395] = 32'b11111111111111110110111001011101;
assign LUT_1[29396] = 32'b00000000000000001001110010100111;
assign LUT_1[29397] = 32'b00000000000000000011000100100011;
assign LUT_1[29398] = 32'b00000000000000000101100000111000;
assign LUT_1[29399] = 32'b11111111111111111110110010110100;
assign LUT_1[29400] = 32'b00000000000000000001000111000101;
assign LUT_1[29401] = 32'b11111111111111111010011001000001;
assign LUT_1[29402] = 32'b11111111111111111100110101010110;
assign LUT_1[29403] = 32'b11111111111111110110000111010010;
assign LUT_1[29404] = 32'b00000000000000001001000000011100;
assign LUT_1[29405] = 32'b00000000000000000010010010011000;
assign LUT_1[29406] = 32'b00000000000000000100101110101101;
assign LUT_1[29407] = 32'b11111111111111111110000000101001;
assign LUT_1[29408] = 32'b00000000000000000000111000101101;
assign LUT_1[29409] = 32'b11111111111111111010001010101001;
assign LUT_1[29410] = 32'b11111111111111111100100110111110;
assign LUT_1[29411] = 32'b11111111111111110101111000111010;
assign LUT_1[29412] = 32'b00000000000000001000110010000100;
assign LUT_1[29413] = 32'b00000000000000000010000100000000;
assign LUT_1[29414] = 32'b00000000000000000100100000010101;
assign LUT_1[29415] = 32'b11111111111111111101110010010001;
assign LUT_1[29416] = 32'b00000000000000000000000110100010;
assign LUT_1[29417] = 32'b11111111111111111001011000011110;
assign LUT_1[29418] = 32'b11111111111111111011110100110011;
assign LUT_1[29419] = 32'b11111111111111110101000110101111;
assign LUT_1[29420] = 32'b00000000000000000111111111111001;
assign LUT_1[29421] = 32'b00000000000000000001010001110101;
assign LUT_1[29422] = 32'b00000000000000000011101110001010;
assign LUT_1[29423] = 32'b11111111111111111101000000000110;
assign LUT_1[29424] = 32'b00000000000000000010110100001111;
assign LUT_1[29425] = 32'b11111111111111111100000110001011;
assign LUT_1[29426] = 32'b11111111111111111110100010100000;
assign LUT_1[29427] = 32'b11111111111111110111110100011100;
assign LUT_1[29428] = 32'b00000000000000001010101101100110;
assign LUT_1[29429] = 32'b00000000000000000011111111100010;
assign LUT_1[29430] = 32'b00000000000000000110011011110111;
assign LUT_1[29431] = 32'b11111111111111111111101101110011;
assign LUT_1[29432] = 32'b00000000000000000010000010000100;
assign LUT_1[29433] = 32'b11111111111111111011010100000000;
assign LUT_1[29434] = 32'b11111111111111111101110000010101;
assign LUT_1[29435] = 32'b11111111111111110111000010010001;
assign LUT_1[29436] = 32'b00000000000000001001111011011011;
assign LUT_1[29437] = 32'b00000000000000000011001101010111;
assign LUT_1[29438] = 32'b00000000000000000101101001101100;
assign LUT_1[29439] = 32'b11111111111111111110111011101000;
assign LUT_1[29440] = 32'b11111111111111111000110100001111;
assign LUT_1[29441] = 32'b11111111111111110010000110001011;
assign LUT_1[29442] = 32'b11111111111111110100100010100000;
assign LUT_1[29443] = 32'b11111111111111101101110100011100;
assign LUT_1[29444] = 32'b00000000000000000000101101100110;
assign LUT_1[29445] = 32'b11111111111111111001111111100010;
assign LUT_1[29446] = 32'b11111111111111111100011011110111;
assign LUT_1[29447] = 32'b11111111111111110101101101110011;
assign LUT_1[29448] = 32'b11111111111111111000000010000100;
assign LUT_1[29449] = 32'b11111111111111110001010100000000;
assign LUT_1[29450] = 32'b11111111111111110011110000010101;
assign LUT_1[29451] = 32'b11111111111111101101000010010001;
assign LUT_1[29452] = 32'b11111111111111111111111011011011;
assign LUT_1[29453] = 32'b11111111111111111001001101010111;
assign LUT_1[29454] = 32'b11111111111111111011101001101100;
assign LUT_1[29455] = 32'b11111111111111110100111011101000;
assign LUT_1[29456] = 32'b11111111111111111010101111110001;
assign LUT_1[29457] = 32'b11111111111111110100000001101101;
assign LUT_1[29458] = 32'b11111111111111110110011110000010;
assign LUT_1[29459] = 32'b11111111111111101111101111111110;
assign LUT_1[29460] = 32'b00000000000000000010101001001000;
assign LUT_1[29461] = 32'b11111111111111111011111011000100;
assign LUT_1[29462] = 32'b11111111111111111110010111011001;
assign LUT_1[29463] = 32'b11111111111111110111101001010101;
assign LUT_1[29464] = 32'b11111111111111111001111101100110;
assign LUT_1[29465] = 32'b11111111111111110011001111100010;
assign LUT_1[29466] = 32'b11111111111111110101101011110111;
assign LUT_1[29467] = 32'b11111111111111101110111101110011;
assign LUT_1[29468] = 32'b00000000000000000001110110111101;
assign LUT_1[29469] = 32'b11111111111111111011001000111001;
assign LUT_1[29470] = 32'b11111111111111111101100101001110;
assign LUT_1[29471] = 32'b11111111111111110110110111001010;
assign LUT_1[29472] = 32'b11111111111111111001101111001110;
assign LUT_1[29473] = 32'b11111111111111110011000001001010;
assign LUT_1[29474] = 32'b11111111111111110101011101011111;
assign LUT_1[29475] = 32'b11111111111111101110101111011011;
assign LUT_1[29476] = 32'b00000000000000000001101000100101;
assign LUT_1[29477] = 32'b11111111111111111010111010100001;
assign LUT_1[29478] = 32'b11111111111111111101010110110110;
assign LUT_1[29479] = 32'b11111111111111110110101000110010;
assign LUT_1[29480] = 32'b11111111111111111000111101000011;
assign LUT_1[29481] = 32'b11111111111111110010001110111111;
assign LUT_1[29482] = 32'b11111111111111110100101011010100;
assign LUT_1[29483] = 32'b11111111111111101101111101010000;
assign LUT_1[29484] = 32'b00000000000000000000110110011010;
assign LUT_1[29485] = 32'b11111111111111111010001000010110;
assign LUT_1[29486] = 32'b11111111111111111100100100101011;
assign LUT_1[29487] = 32'b11111111111111110101110110100111;
assign LUT_1[29488] = 32'b11111111111111111011101010110000;
assign LUT_1[29489] = 32'b11111111111111110100111100101100;
assign LUT_1[29490] = 32'b11111111111111110111011001000001;
assign LUT_1[29491] = 32'b11111111111111110000101010111101;
assign LUT_1[29492] = 32'b00000000000000000011100100000111;
assign LUT_1[29493] = 32'b11111111111111111100110110000011;
assign LUT_1[29494] = 32'b11111111111111111111010010011000;
assign LUT_1[29495] = 32'b11111111111111111000100100010100;
assign LUT_1[29496] = 32'b11111111111111111010111000100101;
assign LUT_1[29497] = 32'b11111111111111110100001010100001;
assign LUT_1[29498] = 32'b11111111111111110110100110110110;
assign LUT_1[29499] = 32'b11111111111111101111111000110010;
assign LUT_1[29500] = 32'b00000000000000000010110001111100;
assign LUT_1[29501] = 32'b11111111111111111100000011111000;
assign LUT_1[29502] = 32'b11111111111111111110100000001101;
assign LUT_1[29503] = 32'b11111111111111110111110010001001;
assign LUT_1[29504] = 32'b11111111111111111010110001110111;
assign LUT_1[29505] = 32'b11111111111111110100000011110011;
assign LUT_1[29506] = 32'b11111111111111110110100000001000;
assign LUT_1[29507] = 32'b11111111111111101111110010000100;
assign LUT_1[29508] = 32'b00000000000000000010101011001110;
assign LUT_1[29509] = 32'b11111111111111111011111101001010;
assign LUT_1[29510] = 32'b11111111111111111110011001011111;
assign LUT_1[29511] = 32'b11111111111111110111101011011011;
assign LUT_1[29512] = 32'b11111111111111111001111111101100;
assign LUT_1[29513] = 32'b11111111111111110011010001101000;
assign LUT_1[29514] = 32'b11111111111111110101101101111101;
assign LUT_1[29515] = 32'b11111111111111101110111111111001;
assign LUT_1[29516] = 32'b00000000000000000001111001000011;
assign LUT_1[29517] = 32'b11111111111111111011001010111111;
assign LUT_1[29518] = 32'b11111111111111111101100111010100;
assign LUT_1[29519] = 32'b11111111111111110110111001010000;
assign LUT_1[29520] = 32'b11111111111111111100101101011001;
assign LUT_1[29521] = 32'b11111111111111110101111111010101;
assign LUT_1[29522] = 32'b11111111111111111000011011101010;
assign LUT_1[29523] = 32'b11111111111111110001101101100110;
assign LUT_1[29524] = 32'b00000000000000000100100110110000;
assign LUT_1[29525] = 32'b11111111111111111101111000101100;
assign LUT_1[29526] = 32'b00000000000000000000010101000001;
assign LUT_1[29527] = 32'b11111111111111111001100110111101;
assign LUT_1[29528] = 32'b11111111111111111011111011001110;
assign LUT_1[29529] = 32'b11111111111111110101001101001010;
assign LUT_1[29530] = 32'b11111111111111110111101001011111;
assign LUT_1[29531] = 32'b11111111111111110000111011011011;
assign LUT_1[29532] = 32'b00000000000000000011110100100101;
assign LUT_1[29533] = 32'b11111111111111111101000110100001;
assign LUT_1[29534] = 32'b11111111111111111111100010110110;
assign LUT_1[29535] = 32'b11111111111111111000110100110010;
assign LUT_1[29536] = 32'b11111111111111111011101100110110;
assign LUT_1[29537] = 32'b11111111111111110100111110110010;
assign LUT_1[29538] = 32'b11111111111111110111011011000111;
assign LUT_1[29539] = 32'b11111111111111110000101101000011;
assign LUT_1[29540] = 32'b00000000000000000011100110001101;
assign LUT_1[29541] = 32'b11111111111111111100111000001001;
assign LUT_1[29542] = 32'b11111111111111111111010100011110;
assign LUT_1[29543] = 32'b11111111111111111000100110011010;
assign LUT_1[29544] = 32'b11111111111111111010111010101011;
assign LUT_1[29545] = 32'b11111111111111110100001100100111;
assign LUT_1[29546] = 32'b11111111111111110110101000111100;
assign LUT_1[29547] = 32'b11111111111111101111111010111000;
assign LUT_1[29548] = 32'b00000000000000000010110100000010;
assign LUT_1[29549] = 32'b11111111111111111100000101111110;
assign LUT_1[29550] = 32'b11111111111111111110100010010011;
assign LUT_1[29551] = 32'b11111111111111110111110100001111;
assign LUT_1[29552] = 32'b11111111111111111101101000011000;
assign LUT_1[29553] = 32'b11111111111111110110111010010100;
assign LUT_1[29554] = 32'b11111111111111111001010110101001;
assign LUT_1[29555] = 32'b11111111111111110010101000100101;
assign LUT_1[29556] = 32'b00000000000000000101100001101111;
assign LUT_1[29557] = 32'b11111111111111111110110011101011;
assign LUT_1[29558] = 32'b00000000000000000001010000000000;
assign LUT_1[29559] = 32'b11111111111111111010100001111100;
assign LUT_1[29560] = 32'b11111111111111111100110110001101;
assign LUT_1[29561] = 32'b11111111111111110110001000001001;
assign LUT_1[29562] = 32'b11111111111111111000100100011110;
assign LUT_1[29563] = 32'b11111111111111110001110110011010;
assign LUT_1[29564] = 32'b00000000000000000100101111100100;
assign LUT_1[29565] = 32'b11111111111111111110000001100000;
assign LUT_1[29566] = 32'b00000000000000000000011101110101;
assign LUT_1[29567] = 32'b11111111111111111001101111110001;
assign LUT_1[29568] = 32'b11111111111111111011110100010010;
assign LUT_1[29569] = 32'b11111111111111110101000110001110;
assign LUT_1[29570] = 32'b11111111111111110111100010100011;
assign LUT_1[29571] = 32'b11111111111111110000110100011111;
assign LUT_1[29572] = 32'b00000000000000000011101101101001;
assign LUT_1[29573] = 32'b11111111111111111100111111100101;
assign LUT_1[29574] = 32'b11111111111111111111011011111010;
assign LUT_1[29575] = 32'b11111111111111111000101101110110;
assign LUT_1[29576] = 32'b11111111111111111011000010000111;
assign LUT_1[29577] = 32'b11111111111111110100010100000011;
assign LUT_1[29578] = 32'b11111111111111110110110000011000;
assign LUT_1[29579] = 32'b11111111111111110000000010010100;
assign LUT_1[29580] = 32'b00000000000000000010111011011110;
assign LUT_1[29581] = 32'b11111111111111111100001101011010;
assign LUT_1[29582] = 32'b11111111111111111110101001101111;
assign LUT_1[29583] = 32'b11111111111111110111111011101011;
assign LUT_1[29584] = 32'b11111111111111111101101111110100;
assign LUT_1[29585] = 32'b11111111111111110111000001110000;
assign LUT_1[29586] = 32'b11111111111111111001011110000101;
assign LUT_1[29587] = 32'b11111111111111110010110000000001;
assign LUT_1[29588] = 32'b00000000000000000101101001001011;
assign LUT_1[29589] = 32'b11111111111111111110111011000111;
assign LUT_1[29590] = 32'b00000000000000000001010111011100;
assign LUT_1[29591] = 32'b11111111111111111010101001011000;
assign LUT_1[29592] = 32'b11111111111111111100111101101001;
assign LUT_1[29593] = 32'b11111111111111110110001111100101;
assign LUT_1[29594] = 32'b11111111111111111000101011111010;
assign LUT_1[29595] = 32'b11111111111111110001111101110110;
assign LUT_1[29596] = 32'b00000000000000000100110111000000;
assign LUT_1[29597] = 32'b11111111111111111110001000111100;
assign LUT_1[29598] = 32'b00000000000000000000100101010001;
assign LUT_1[29599] = 32'b11111111111111111001110111001101;
assign LUT_1[29600] = 32'b11111111111111111100101111010001;
assign LUT_1[29601] = 32'b11111111111111110110000001001101;
assign LUT_1[29602] = 32'b11111111111111111000011101100010;
assign LUT_1[29603] = 32'b11111111111111110001101111011110;
assign LUT_1[29604] = 32'b00000000000000000100101000101000;
assign LUT_1[29605] = 32'b11111111111111111101111010100100;
assign LUT_1[29606] = 32'b00000000000000000000010110111001;
assign LUT_1[29607] = 32'b11111111111111111001101000110101;
assign LUT_1[29608] = 32'b11111111111111111011111101000110;
assign LUT_1[29609] = 32'b11111111111111110101001111000010;
assign LUT_1[29610] = 32'b11111111111111110111101011010111;
assign LUT_1[29611] = 32'b11111111111111110000111101010011;
assign LUT_1[29612] = 32'b00000000000000000011110110011101;
assign LUT_1[29613] = 32'b11111111111111111101001000011001;
assign LUT_1[29614] = 32'b11111111111111111111100100101110;
assign LUT_1[29615] = 32'b11111111111111111000110110101010;
assign LUT_1[29616] = 32'b11111111111111111110101010110011;
assign LUT_1[29617] = 32'b11111111111111110111111100101111;
assign LUT_1[29618] = 32'b11111111111111111010011001000100;
assign LUT_1[29619] = 32'b11111111111111110011101011000000;
assign LUT_1[29620] = 32'b00000000000000000110100100001010;
assign LUT_1[29621] = 32'b11111111111111111111110110000110;
assign LUT_1[29622] = 32'b00000000000000000010010010011011;
assign LUT_1[29623] = 32'b11111111111111111011100100010111;
assign LUT_1[29624] = 32'b11111111111111111101111000101000;
assign LUT_1[29625] = 32'b11111111111111110111001010100100;
assign LUT_1[29626] = 32'b11111111111111111001100110111001;
assign LUT_1[29627] = 32'b11111111111111110010111000110101;
assign LUT_1[29628] = 32'b00000000000000000101110001111111;
assign LUT_1[29629] = 32'b11111111111111111111000011111011;
assign LUT_1[29630] = 32'b00000000000000000001100000010000;
assign LUT_1[29631] = 32'b11111111111111111010110010001100;
assign LUT_1[29632] = 32'b11111111111111111101110001111010;
assign LUT_1[29633] = 32'b11111111111111110111000011110110;
assign LUT_1[29634] = 32'b11111111111111111001100000001011;
assign LUT_1[29635] = 32'b11111111111111110010110010000111;
assign LUT_1[29636] = 32'b00000000000000000101101011010001;
assign LUT_1[29637] = 32'b11111111111111111110111101001101;
assign LUT_1[29638] = 32'b00000000000000000001011001100010;
assign LUT_1[29639] = 32'b11111111111111111010101011011110;
assign LUT_1[29640] = 32'b11111111111111111100111111101111;
assign LUT_1[29641] = 32'b11111111111111110110010001101011;
assign LUT_1[29642] = 32'b11111111111111111000101110000000;
assign LUT_1[29643] = 32'b11111111111111110001111111111100;
assign LUT_1[29644] = 32'b00000000000000000100111001000110;
assign LUT_1[29645] = 32'b11111111111111111110001011000010;
assign LUT_1[29646] = 32'b00000000000000000000100111010111;
assign LUT_1[29647] = 32'b11111111111111111001111001010011;
assign LUT_1[29648] = 32'b11111111111111111111101101011100;
assign LUT_1[29649] = 32'b11111111111111111000111111011000;
assign LUT_1[29650] = 32'b11111111111111111011011011101101;
assign LUT_1[29651] = 32'b11111111111111110100101101101001;
assign LUT_1[29652] = 32'b00000000000000000111100110110011;
assign LUT_1[29653] = 32'b00000000000000000000111000101111;
assign LUT_1[29654] = 32'b00000000000000000011010101000100;
assign LUT_1[29655] = 32'b11111111111111111100100111000000;
assign LUT_1[29656] = 32'b11111111111111111110111011010001;
assign LUT_1[29657] = 32'b11111111111111111000001101001101;
assign LUT_1[29658] = 32'b11111111111111111010101001100010;
assign LUT_1[29659] = 32'b11111111111111110011111011011110;
assign LUT_1[29660] = 32'b00000000000000000110110100101000;
assign LUT_1[29661] = 32'b00000000000000000000000110100100;
assign LUT_1[29662] = 32'b00000000000000000010100010111001;
assign LUT_1[29663] = 32'b11111111111111111011110100110101;
assign LUT_1[29664] = 32'b11111111111111111110101100111001;
assign LUT_1[29665] = 32'b11111111111111110111111110110101;
assign LUT_1[29666] = 32'b11111111111111111010011011001010;
assign LUT_1[29667] = 32'b11111111111111110011101101000110;
assign LUT_1[29668] = 32'b00000000000000000110100110010000;
assign LUT_1[29669] = 32'b11111111111111111111111000001100;
assign LUT_1[29670] = 32'b00000000000000000010010100100001;
assign LUT_1[29671] = 32'b11111111111111111011100110011101;
assign LUT_1[29672] = 32'b11111111111111111101111010101110;
assign LUT_1[29673] = 32'b11111111111111110111001100101010;
assign LUT_1[29674] = 32'b11111111111111111001101000111111;
assign LUT_1[29675] = 32'b11111111111111110010111010111011;
assign LUT_1[29676] = 32'b00000000000000000101110100000101;
assign LUT_1[29677] = 32'b11111111111111111111000110000001;
assign LUT_1[29678] = 32'b00000000000000000001100010010110;
assign LUT_1[29679] = 32'b11111111111111111010110100010010;
assign LUT_1[29680] = 32'b00000000000000000000101000011011;
assign LUT_1[29681] = 32'b11111111111111111001111010010111;
assign LUT_1[29682] = 32'b11111111111111111100010110101100;
assign LUT_1[29683] = 32'b11111111111111110101101000101000;
assign LUT_1[29684] = 32'b00000000000000001000100001110010;
assign LUT_1[29685] = 32'b00000000000000000001110011101110;
assign LUT_1[29686] = 32'b00000000000000000100010000000011;
assign LUT_1[29687] = 32'b11111111111111111101100001111111;
assign LUT_1[29688] = 32'b11111111111111111111110110010000;
assign LUT_1[29689] = 32'b11111111111111111001001000001100;
assign LUT_1[29690] = 32'b11111111111111111011100100100001;
assign LUT_1[29691] = 32'b11111111111111110100110110011101;
assign LUT_1[29692] = 32'b00000000000000000111101111100111;
assign LUT_1[29693] = 32'b00000000000000000001000001100011;
assign LUT_1[29694] = 32'b00000000000000000011011101111000;
assign LUT_1[29695] = 32'b11111111111111111100101111110100;
assign LUT_1[29696] = 32'b00000000000000000111101000010110;
assign LUT_1[29697] = 32'b00000000000000000000111010010010;
assign LUT_1[29698] = 32'b00000000000000000011010110100111;
assign LUT_1[29699] = 32'b11111111111111111100101000100011;
assign LUT_1[29700] = 32'b00000000000000001111100001101101;
assign LUT_1[29701] = 32'b00000000000000001000110011101001;
assign LUT_1[29702] = 32'b00000000000000001011001111111110;
assign LUT_1[29703] = 32'b00000000000000000100100001111010;
assign LUT_1[29704] = 32'b00000000000000000110110110001011;
assign LUT_1[29705] = 32'b00000000000000000000001000000111;
assign LUT_1[29706] = 32'b00000000000000000010100100011100;
assign LUT_1[29707] = 32'b11111111111111111011110110011000;
assign LUT_1[29708] = 32'b00000000000000001110101111100010;
assign LUT_1[29709] = 32'b00000000000000001000000001011110;
assign LUT_1[29710] = 32'b00000000000000001010011101110011;
assign LUT_1[29711] = 32'b00000000000000000011101111101111;
assign LUT_1[29712] = 32'b00000000000000001001100011111000;
assign LUT_1[29713] = 32'b00000000000000000010110101110100;
assign LUT_1[29714] = 32'b00000000000000000101010010001001;
assign LUT_1[29715] = 32'b11111111111111111110100100000101;
assign LUT_1[29716] = 32'b00000000000000010001011101001111;
assign LUT_1[29717] = 32'b00000000000000001010101111001011;
assign LUT_1[29718] = 32'b00000000000000001101001011100000;
assign LUT_1[29719] = 32'b00000000000000000110011101011100;
assign LUT_1[29720] = 32'b00000000000000001000110001101101;
assign LUT_1[29721] = 32'b00000000000000000010000011101001;
assign LUT_1[29722] = 32'b00000000000000000100011111111110;
assign LUT_1[29723] = 32'b11111111111111111101110001111010;
assign LUT_1[29724] = 32'b00000000000000010000101011000100;
assign LUT_1[29725] = 32'b00000000000000001001111101000000;
assign LUT_1[29726] = 32'b00000000000000001100011001010101;
assign LUT_1[29727] = 32'b00000000000000000101101011010001;
assign LUT_1[29728] = 32'b00000000000000001000100011010101;
assign LUT_1[29729] = 32'b00000000000000000001110101010001;
assign LUT_1[29730] = 32'b00000000000000000100010001100110;
assign LUT_1[29731] = 32'b11111111111111111101100011100010;
assign LUT_1[29732] = 32'b00000000000000010000011100101100;
assign LUT_1[29733] = 32'b00000000000000001001101110101000;
assign LUT_1[29734] = 32'b00000000000000001100001010111101;
assign LUT_1[29735] = 32'b00000000000000000101011100111001;
assign LUT_1[29736] = 32'b00000000000000000111110001001010;
assign LUT_1[29737] = 32'b00000000000000000001000011000110;
assign LUT_1[29738] = 32'b00000000000000000011011111011011;
assign LUT_1[29739] = 32'b11111111111111111100110001010111;
assign LUT_1[29740] = 32'b00000000000000001111101010100001;
assign LUT_1[29741] = 32'b00000000000000001000111100011101;
assign LUT_1[29742] = 32'b00000000000000001011011000110010;
assign LUT_1[29743] = 32'b00000000000000000100101010101110;
assign LUT_1[29744] = 32'b00000000000000001010011110110111;
assign LUT_1[29745] = 32'b00000000000000000011110000110011;
assign LUT_1[29746] = 32'b00000000000000000110001101001000;
assign LUT_1[29747] = 32'b11111111111111111111011111000100;
assign LUT_1[29748] = 32'b00000000000000010010011000001110;
assign LUT_1[29749] = 32'b00000000000000001011101010001010;
assign LUT_1[29750] = 32'b00000000000000001110000110011111;
assign LUT_1[29751] = 32'b00000000000000000111011000011011;
assign LUT_1[29752] = 32'b00000000000000001001101100101100;
assign LUT_1[29753] = 32'b00000000000000000010111110101000;
assign LUT_1[29754] = 32'b00000000000000000101011010111101;
assign LUT_1[29755] = 32'b11111111111111111110101100111001;
assign LUT_1[29756] = 32'b00000000000000010001100110000011;
assign LUT_1[29757] = 32'b00000000000000001010110111111111;
assign LUT_1[29758] = 32'b00000000000000001101010100010100;
assign LUT_1[29759] = 32'b00000000000000000110100110010000;
assign LUT_1[29760] = 32'b00000000000000001001100101111110;
assign LUT_1[29761] = 32'b00000000000000000010110111111010;
assign LUT_1[29762] = 32'b00000000000000000101010100001111;
assign LUT_1[29763] = 32'b11111111111111111110100110001011;
assign LUT_1[29764] = 32'b00000000000000010001011111010101;
assign LUT_1[29765] = 32'b00000000000000001010110001010001;
assign LUT_1[29766] = 32'b00000000000000001101001101100110;
assign LUT_1[29767] = 32'b00000000000000000110011111100010;
assign LUT_1[29768] = 32'b00000000000000001000110011110011;
assign LUT_1[29769] = 32'b00000000000000000010000101101111;
assign LUT_1[29770] = 32'b00000000000000000100100010000100;
assign LUT_1[29771] = 32'b11111111111111111101110100000000;
assign LUT_1[29772] = 32'b00000000000000010000101101001010;
assign LUT_1[29773] = 32'b00000000000000001001111111000110;
assign LUT_1[29774] = 32'b00000000000000001100011011011011;
assign LUT_1[29775] = 32'b00000000000000000101101101010111;
assign LUT_1[29776] = 32'b00000000000000001011100001100000;
assign LUT_1[29777] = 32'b00000000000000000100110011011100;
assign LUT_1[29778] = 32'b00000000000000000111001111110001;
assign LUT_1[29779] = 32'b00000000000000000000100001101101;
assign LUT_1[29780] = 32'b00000000000000010011011010110111;
assign LUT_1[29781] = 32'b00000000000000001100101100110011;
assign LUT_1[29782] = 32'b00000000000000001111001001001000;
assign LUT_1[29783] = 32'b00000000000000001000011011000100;
assign LUT_1[29784] = 32'b00000000000000001010101111010101;
assign LUT_1[29785] = 32'b00000000000000000100000001010001;
assign LUT_1[29786] = 32'b00000000000000000110011101100110;
assign LUT_1[29787] = 32'b11111111111111111111101111100010;
assign LUT_1[29788] = 32'b00000000000000010010101000101100;
assign LUT_1[29789] = 32'b00000000000000001011111010101000;
assign LUT_1[29790] = 32'b00000000000000001110010110111101;
assign LUT_1[29791] = 32'b00000000000000000111101000111001;
assign LUT_1[29792] = 32'b00000000000000001010100000111101;
assign LUT_1[29793] = 32'b00000000000000000011110010111001;
assign LUT_1[29794] = 32'b00000000000000000110001111001110;
assign LUT_1[29795] = 32'b11111111111111111111100001001010;
assign LUT_1[29796] = 32'b00000000000000010010011010010100;
assign LUT_1[29797] = 32'b00000000000000001011101100010000;
assign LUT_1[29798] = 32'b00000000000000001110001000100101;
assign LUT_1[29799] = 32'b00000000000000000111011010100001;
assign LUT_1[29800] = 32'b00000000000000001001101110110010;
assign LUT_1[29801] = 32'b00000000000000000011000000101110;
assign LUT_1[29802] = 32'b00000000000000000101011101000011;
assign LUT_1[29803] = 32'b11111111111111111110101110111111;
assign LUT_1[29804] = 32'b00000000000000010001101000001001;
assign LUT_1[29805] = 32'b00000000000000001010111010000101;
assign LUT_1[29806] = 32'b00000000000000001101010110011010;
assign LUT_1[29807] = 32'b00000000000000000110101000010110;
assign LUT_1[29808] = 32'b00000000000000001100011100011111;
assign LUT_1[29809] = 32'b00000000000000000101101110011011;
assign LUT_1[29810] = 32'b00000000000000001000001010110000;
assign LUT_1[29811] = 32'b00000000000000000001011100101100;
assign LUT_1[29812] = 32'b00000000000000010100010101110110;
assign LUT_1[29813] = 32'b00000000000000001101100111110010;
assign LUT_1[29814] = 32'b00000000000000010000000100000111;
assign LUT_1[29815] = 32'b00000000000000001001010110000011;
assign LUT_1[29816] = 32'b00000000000000001011101010010100;
assign LUT_1[29817] = 32'b00000000000000000100111100010000;
assign LUT_1[29818] = 32'b00000000000000000111011000100101;
assign LUT_1[29819] = 32'b00000000000000000000101010100001;
assign LUT_1[29820] = 32'b00000000000000010011100011101011;
assign LUT_1[29821] = 32'b00000000000000001100110101100111;
assign LUT_1[29822] = 32'b00000000000000001111010001111100;
assign LUT_1[29823] = 32'b00000000000000001000100011111000;
assign LUT_1[29824] = 32'b00000000000000001010101000011001;
assign LUT_1[29825] = 32'b00000000000000000011111010010101;
assign LUT_1[29826] = 32'b00000000000000000110010110101010;
assign LUT_1[29827] = 32'b11111111111111111111101000100110;
assign LUT_1[29828] = 32'b00000000000000010010100001110000;
assign LUT_1[29829] = 32'b00000000000000001011110011101100;
assign LUT_1[29830] = 32'b00000000000000001110010000000001;
assign LUT_1[29831] = 32'b00000000000000000111100001111101;
assign LUT_1[29832] = 32'b00000000000000001001110110001110;
assign LUT_1[29833] = 32'b00000000000000000011001000001010;
assign LUT_1[29834] = 32'b00000000000000000101100100011111;
assign LUT_1[29835] = 32'b11111111111111111110110110011011;
assign LUT_1[29836] = 32'b00000000000000010001101111100101;
assign LUT_1[29837] = 32'b00000000000000001011000001100001;
assign LUT_1[29838] = 32'b00000000000000001101011101110110;
assign LUT_1[29839] = 32'b00000000000000000110101111110010;
assign LUT_1[29840] = 32'b00000000000000001100100011111011;
assign LUT_1[29841] = 32'b00000000000000000101110101110111;
assign LUT_1[29842] = 32'b00000000000000001000010010001100;
assign LUT_1[29843] = 32'b00000000000000000001100100001000;
assign LUT_1[29844] = 32'b00000000000000010100011101010010;
assign LUT_1[29845] = 32'b00000000000000001101101111001110;
assign LUT_1[29846] = 32'b00000000000000010000001011100011;
assign LUT_1[29847] = 32'b00000000000000001001011101011111;
assign LUT_1[29848] = 32'b00000000000000001011110001110000;
assign LUT_1[29849] = 32'b00000000000000000101000011101100;
assign LUT_1[29850] = 32'b00000000000000000111100000000001;
assign LUT_1[29851] = 32'b00000000000000000000110001111101;
assign LUT_1[29852] = 32'b00000000000000010011101011000111;
assign LUT_1[29853] = 32'b00000000000000001100111101000011;
assign LUT_1[29854] = 32'b00000000000000001111011001011000;
assign LUT_1[29855] = 32'b00000000000000001000101011010100;
assign LUT_1[29856] = 32'b00000000000000001011100011011000;
assign LUT_1[29857] = 32'b00000000000000000100110101010100;
assign LUT_1[29858] = 32'b00000000000000000111010001101001;
assign LUT_1[29859] = 32'b00000000000000000000100011100101;
assign LUT_1[29860] = 32'b00000000000000010011011100101111;
assign LUT_1[29861] = 32'b00000000000000001100101110101011;
assign LUT_1[29862] = 32'b00000000000000001111001011000000;
assign LUT_1[29863] = 32'b00000000000000001000011100111100;
assign LUT_1[29864] = 32'b00000000000000001010110001001101;
assign LUT_1[29865] = 32'b00000000000000000100000011001001;
assign LUT_1[29866] = 32'b00000000000000000110011111011110;
assign LUT_1[29867] = 32'b11111111111111111111110001011010;
assign LUT_1[29868] = 32'b00000000000000010010101010100100;
assign LUT_1[29869] = 32'b00000000000000001011111100100000;
assign LUT_1[29870] = 32'b00000000000000001110011000110101;
assign LUT_1[29871] = 32'b00000000000000000111101010110001;
assign LUT_1[29872] = 32'b00000000000000001101011110111010;
assign LUT_1[29873] = 32'b00000000000000000110110000110110;
assign LUT_1[29874] = 32'b00000000000000001001001101001011;
assign LUT_1[29875] = 32'b00000000000000000010011111000111;
assign LUT_1[29876] = 32'b00000000000000010101011000010001;
assign LUT_1[29877] = 32'b00000000000000001110101010001101;
assign LUT_1[29878] = 32'b00000000000000010001000110100010;
assign LUT_1[29879] = 32'b00000000000000001010011000011110;
assign LUT_1[29880] = 32'b00000000000000001100101100101111;
assign LUT_1[29881] = 32'b00000000000000000101111110101011;
assign LUT_1[29882] = 32'b00000000000000001000011011000000;
assign LUT_1[29883] = 32'b00000000000000000001101100111100;
assign LUT_1[29884] = 32'b00000000000000010100100110000110;
assign LUT_1[29885] = 32'b00000000000000001101111000000010;
assign LUT_1[29886] = 32'b00000000000000010000010100010111;
assign LUT_1[29887] = 32'b00000000000000001001100110010011;
assign LUT_1[29888] = 32'b00000000000000001100100110000001;
assign LUT_1[29889] = 32'b00000000000000000101110111111101;
assign LUT_1[29890] = 32'b00000000000000001000010100010010;
assign LUT_1[29891] = 32'b00000000000000000001100110001110;
assign LUT_1[29892] = 32'b00000000000000010100011111011000;
assign LUT_1[29893] = 32'b00000000000000001101110001010100;
assign LUT_1[29894] = 32'b00000000000000010000001101101001;
assign LUT_1[29895] = 32'b00000000000000001001011111100101;
assign LUT_1[29896] = 32'b00000000000000001011110011110110;
assign LUT_1[29897] = 32'b00000000000000000101000101110010;
assign LUT_1[29898] = 32'b00000000000000000111100010000111;
assign LUT_1[29899] = 32'b00000000000000000000110100000011;
assign LUT_1[29900] = 32'b00000000000000010011101101001101;
assign LUT_1[29901] = 32'b00000000000000001100111111001001;
assign LUT_1[29902] = 32'b00000000000000001111011011011110;
assign LUT_1[29903] = 32'b00000000000000001000101101011010;
assign LUT_1[29904] = 32'b00000000000000001110100001100011;
assign LUT_1[29905] = 32'b00000000000000000111110011011111;
assign LUT_1[29906] = 32'b00000000000000001010001111110100;
assign LUT_1[29907] = 32'b00000000000000000011100001110000;
assign LUT_1[29908] = 32'b00000000000000010110011010111010;
assign LUT_1[29909] = 32'b00000000000000001111101100110110;
assign LUT_1[29910] = 32'b00000000000000010010001001001011;
assign LUT_1[29911] = 32'b00000000000000001011011011000111;
assign LUT_1[29912] = 32'b00000000000000001101101111011000;
assign LUT_1[29913] = 32'b00000000000000000111000001010100;
assign LUT_1[29914] = 32'b00000000000000001001011101101001;
assign LUT_1[29915] = 32'b00000000000000000010101111100101;
assign LUT_1[29916] = 32'b00000000000000010101101000101111;
assign LUT_1[29917] = 32'b00000000000000001110111010101011;
assign LUT_1[29918] = 32'b00000000000000010001010111000000;
assign LUT_1[29919] = 32'b00000000000000001010101000111100;
assign LUT_1[29920] = 32'b00000000000000001101100001000000;
assign LUT_1[29921] = 32'b00000000000000000110110010111100;
assign LUT_1[29922] = 32'b00000000000000001001001111010001;
assign LUT_1[29923] = 32'b00000000000000000010100001001101;
assign LUT_1[29924] = 32'b00000000000000010101011010010111;
assign LUT_1[29925] = 32'b00000000000000001110101100010011;
assign LUT_1[29926] = 32'b00000000000000010001001000101000;
assign LUT_1[29927] = 32'b00000000000000001010011010100100;
assign LUT_1[29928] = 32'b00000000000000001100101110110101;
assign LUT_1[29929] = 32'b00000000000000000110000000110001;
assign LUT_1[29930] = 32'b00000000000000001000011101000110;
assign LUT_1[29931] = 32'b00000000000000000001101111000010;
assign LUT_1[29932] = 32'b00000000000000010100101000001100;
assign LUT_1[29933] = 32'b00000000000000001101111010001000;
assign LUT_1[29934] = 32'b00000000000000010000010110011101;
assign LUT_1[29935] = 32'b00000000000000001001101000011001;
assign LUT_1[29936] = 32'b00000000000000001111011100100010;
assign LUT_1[29937] = 32'b00000000000000001000101110011110;
assign LUT_1[29938] = 32'b00000000000000001011001010110011;
assign LUT_1[29939] = 32'b00000000000000000100011100101111;
assign LUT_1[29940] = 32'b00000000000000010111010101111001;
assign LUT_1[29941] = 32'b00000000000000010000100111110101;
assign LUT_1[29942] = 32'b00000000000000010011000100001010;
assign LUT_1[29943] = 32'b00000000000000001100010110000110;
assign LUT_1[29944] = 32'b00000000000000001110101010010111;
assign LUT_1[29945] = 32'b00000000000000000111111100010011;
assign LUT_1[29946] = 32'b00000000000000001010011000101000;
assign LUT_1[29947] = 32'b00000000000000000011101010100100;
assign LUT_1[29948] = 32'b00000000000000010110100011101110;
assign LUT_1[29949] = 32'b00000000000000001111110101101010;
assign LUT_1[29950] = 32'b00000000000000010010010001111111;
assign LUT_1[29951] = 32'b00000000000000001011100011111011;
assign LUT_1[29952] = 32'b00000000000000000101011100100010;
assign LUT_1[29953] = 32'b11111111111111111110101110011110;
assign LUT_1[29954] = 32'b00000000000000000001001010110011;
assign LUT_1[29955] = 32'b11111111111111111010011100101111;
assign LUT_1[29956] = 32'b00000000000000001101010101111001;
assign LUT_1[29957] = 32'b00000000000000000110100111110101;
assign LUT_1[29958] = 32'b00000000000000001001000100001010;
assign LUT_1[29959] = 32'b00000000000000000010010110000110;
assign LUT_1[29960] = 32'b00000000000000000100101010010111;
assign LUT_1[29961] = 32'b11111111111111111101111100010011;
assign LUT_1[29962] = 32'b00000000000000000000011000101000;
assign LUT_1[29963] = 32'b11111111111111111001101010100100;
assign LUT_1[29964] = 32'b00000000000000001100100011101110;
assign LUT_1[29965] = 32'b00000000000000000101110101101010;
assign LUT_1[29966] = 32'b00000000000000001000010001111111;
assign LUT_1[29967] = 32'b00000000000000000001100011111011;
assign LUT_1[29968] = 32'b00000000000000000111011000000100;
assign LUT_1[29969] = 32'b00000000000000000000101010000000;
assign LUT_1[29970] = 32'b00000000000000000011000110010101;
assign LUT_1[29971] = 32'b11111111111111111100011000010001;
assign LUT_1[29972] = 32'b00000000000000001111010001011011;
assign LUT_1[29973] = 32'b00000000000000001000100011010111;
assign LUT_1[29974] = 32'b00000000000000001010111111101100;
assign LUT_1[29975] = 32'b00000000000000000100010001101000;
assign LUT_1[29976] = 32'b00000000000000000110100101111001;
assign LUT_1[29977] = 32'b11111111111111111111110111110101;
assign LUT_1[29978] = 32'b00000000000000000010010100001010;
assign LUT_1[29979] = 32'b11111111111111111011100110000110;
assign LUT_1[29980] = 32'b00000000000000001110011111010000;
assign LUT_1[29981] = 32'b00000000000000000111110001001100;
assign LUT_1[29982] = 32'b00000000000000001010001101100001;
assign LUT_1[29983] = 32'b00000000000000000011011111011101;
assign LUT_1[29984] = 32'b00000000000000000110010111100001;
assign LUT_1[29985] = 32'b11111111111111111111101001011101;
assign LUT_1[29986] = 32'b00000000000000000010000101110010;
assign LUT_1[29987] = 32'b11111111111111111011010111101110;
assign LUT_1[29988] = 32'b00000000000000001110010000111000;
assign LUT_1[29989] = 32'b00000000000000000111100010110100;
assign LUT_1[29990] = 32'b00000000000000001001111111001001;
assign LUT_1[29991] = 32'b00000000000000000011010001000101;
assign LUT_1[29992] = 32'b00000000000000000101100101010110;
assign LUT_1[29993] = 32'b11111111111111111110110111010010;
assign LUT_1[29994] = 32'b00000000000000000001010011100111;
assign LUT_1[29995] = 32'b11111111111111111010100101100011;
assign LUT_1[29996] = 32'b00000000000000001101011110101101;
assign LUT_1[29997] = 32'b00000000000000000110110000101001;
assign LUT_1[29998] = 32'b00000000000000001001001100111110;
assign LUT_1[29999] = 32'b00000000000000000010011110111010;
assign LUT_1[30000] = 32'b00000000000000001000010011000011;
assign LUT_1[30001] = 32'b00000000000000000001100100111111;
assign LUT_1[30002] = 32'b00000000000000000100000001010100;
assign LUT_1[30003] = 32'b11111111111111111101010011010000;
assign LUT_1[30004] = 32'b00000000000000010000001100011010;
assign LUT_1[30005] = 32'b00000000000000001001011110010110;
assign LUT_1[30006] = 32'b00000000000000001011111010101011;
assign LUT_1[30007] = 32'b00000000000000000101001100100111;
assign LUT_1[30008] = 32'b00000000000000000111100000111000;
assign LUT_1[30009] = 32'b00000000000000000000110010110100;
assign LUT_1[30010] = 32'b00000000000000000011001111001001;
assign LUT_1[30011] = 32'b11111111111111111100100001000101;
assign LUT_1[30012] = 32'b00000000000000001111011010001111;
assign LUT_1[30013] = 32'b00000000000000001000101100001011;
assign LUT_1[30014] = 32'b00000000000000001011001000100000;
assign LUT_1[30015] = 32'b00000000000000000100011010011100;
assign LUT_1[30016] = 32'b00000000000000000111011010001010;
assign LUT_1[30017] = 32'b00000000000000000000101100000110;
assign LUT_1[30018] = 32'b00000000000000000011001000011011;
assign LUT_1[30019] = 32'b11111111111111111100011010010111;
assign LUT_1[30020] = 32'b00000000000000001111010011100001;
assign LUT_1[30021] = 32'b00000000000000001000100101011101;
assign LUT_1[30022] = 32'b00000000000000001011000001110010;
assign LUT_1[30023] = 32'b00000000000000000100010011101110;
assign LUT_1[30024] = 32'b00000000000000000110100111111111;
assign LUT_1[30025] = 32'b11111111111111111111111001111011;
assign LUT_1[30026] = 32'b00000000000000000010010110010000;
assign LUT_1[30027] = 32'b11111111111111111011101000001100;
assign LUT_1[30028] = 32'b00000000000000001110100001010110;
assign LUT_1[30029] = 32'b00000000000000000111110011010010;
assign LUT_1[30030] = 32'b00000000000000001010001111100111;
assign LUT_1[30031] = 32'b00000000000000000011100001100011;
assign LUT_1[30032] = 32'b00000000000000001001010101101100;
assign LUT_1[30033] = 32'b00000000000000000010100111101000;
assign LUT_1[30034] = 32'b00000000000000000101000011111101;
assign LUT_1[30035] = 32'b11111111111111111110010101111001;
assign LUT_1[30036] = 32'b00000000000000010001001111000011;
assign LUT_1[30037] = 32'b00000000000000001010100000111111;
assign LUT_1[30038] = 32'b00000000000000001100111101010100;
assign LUT_1[30039] = 32'b00000000000000000110001111010000;
assign LUT_1[30040] = 32'b00000000000000001000100011100001;
assign LUT_1[30041] = 32'b00000000000000000001110101011101;
assign LUT_1[30042] = 32'b00000000000000000100010001110010;
assign LUT_1[30043] = 32'b11111111111111111101100011101110;
assign LUT_1[30044] = 32'b00000000000000010000011100111000;
assign LUT_1[30045] = 32'b00000000000000001001101110110100;
assign LUT_1[30046] = 32'b00000000000000001100001011001001;
assign LUT_1[30047] = 32'b00000000000000000101011101000101;
assign LUT_1[30048] = 32'b00000000000000001000010101001001;
assign LUT_1[30049] = 32'b00000000000000000001100111000101;
assign LUT_1[30050] = 32'b00000000000000000100000011011010;
assign LUT_1[30051] = 32'b11111111111111111101010101010110;
assign LUT_1[30052] = 32'b00000000000000010000001110100000;
assign LUT_1[30053] = 32'b00000000000000001001100000011100;
assign LUT_1[30054] = 32'b00000000000000001011111100110001;
assign LUT_1[30055] = 32'b00000000000000000101001110101101;
assign LUT_1[30056] = 32'b00000000000000000111100010111110;
assign LUT_1[30057] = 32'b00000000000000000000110100111010;
assign LUT_1[30058] = 32'b00000000000000000011010001001111;
assign LUT_1[30059] = 32'b11111111111111111100100011001011;
assign LUT_1[30060] = 32'b00000000000000001111011100010101;
assign LUT_1[30061] = 32'b00000000000000001000101110010001;
assign LUT_1[30062] = 32'b00000000000000001011001010100110;
assign LUT_1[30063] = 32'b00000000000000000100011100100010;
assign LUT_1[30064] = 32'b00000000000000001010010000101011;
assign LUT_1[30065] = 32'b00000000000000000011100010100111;
assign LUT_1[30066] = 32'b00000000000000000101111110111100;
assign LUT_1[30067] = 32'b11111111111111111111010000111000;
assign LUT_1[30068] = 32'b00000000000000010010001010000010;
assign LUT_1[30069] = 32'b00000000000000001011011011111110;
assign LUT_1[30070] = 32'b00000000000000001101111000010011;
assign LUT_1[30071] = 32'b00000000000000000111001010001111;
assign LUT_1[30072] = 32'b00000000000000001001011110100000;
assign LUT_1[30073] = 32'b00000000000000000010110000011100;
assign LUT_1[30074] = 32'b00000000000000000101001100110001;
assign LUT_1[30075] = 32'b11111111111111111110011110101101;
assign LUT_1[30076] = 32'b00000000000000010001010111110111;
assign LUT_1[30077] = 32'b00000000000000001010101001110011;
assign LUT_1[30078] = 32'b00000000000000001101000110001000;
assign LUT_1[30079] = 32'b00000000000000000110011000000100;
assign LUT_1[30080] = 32'b00000000000000001000011100100101;
assign LUT_1[30081] = 32'b00000000000000000001101110100001;
assign LUT_1[30082] = 32'b00000000000000000100001010110110;
assign LUT_1[30083] = 32'b11111111111111111101011100110010;
assign LUT_1[30084] = 32'b00000000000000010000010101111100;
assign LUT_1[30085] = 32'b00000000000000001001100111111000;
assign LUT_1[30086] = 32'b00000000000000001100000100001101;
assign LUT_1[30087] = 32'b00000000000000000101010110001001;
assign LUT_1[30088] = 32'b00000000000000000111101010011010;
assign LUT_1[30089] = 32'b00000000000000000000111100010110;
assign LUT_1[30090] = 32'b00000000000000000011011000101011;
assign LUT_1[30091] = 32'b11111111111111111100101010100111;
assign LUT_1[30092] = 32'b00000000000000001111100011110001;
assign LUT_1[30093] = 32'b00000000000000001000110101101101;
assign LUT_1[30094] = 32'b00000000000000001011010010000010;
assign LUT_1[30095] = 32'b00000000000000000100100011111110;
assign LUT_1[30096] = 32'b00000000000000001010011000000111;
assign LUT_1[30097] = 32'b00000000000000000011101010000011;
assign LUT_1[30098] = 32'b00000000000000000110000110011000;
assign LUT_1[30099] = 32'b11111111111111111111011000010100;
assign LUT_1[30100] = 32'b00000000000000010010010001011110;
assign LUT_1[30101] = 32'b00000000000000001011100011011010;
assign LUT_1[30102] = 32'b00000000000000001101111111101111;
assign LUT_1[30103] = 32'b00000000000000000111010001101011;
assign LUT_1[30104] = 32'b00000000000000001001100101111100;
assign LUT_1[30105] = 32'b00000000000000000010110111111000;
assign LUT_1[30106] = 32'b00000000000000000101010100001101;
assign LUT_1[30107] = 32'b11111111111111111110100110001001;
assign LUT_1[30108] = 32'b00000000000000010001011111010011;
assign LUT_1[30109] = 32'b00000000000000001010110001001111;
assign LUT_1[30110] = 32'b00000000000000001101001101100100;
assign LUT_1[30111] = 32'b00000000000000000110011111100000;
assign LUT_1[30112] = 32'b00000000000000001001010111100100;
assign LUT_1[30113] = 32'b00000000000000000010101001100000;
assign LUT_1[30114] = 32'b00000000000000000101000101110101;
assign LUT_1[30115] = 32'b11111111111111111110010111110001;
assign LUT_1[30116] = 32'b00000000000000010001010000111011;
assign LUT_1[30117] = 32'b00000000000000001010100010110111;
assign LUT_1[30118] = 32'b00000000000000001100111111001100;
assign LUT_1[30119] = 32'b00000000000000000110010001001000;
assign LUT_1[30120] = 32'b00000000000000001000100101011001;
assign LUT_1[30121] = 32'b00000000000000000001110111010101;
assign LUT_1[30122] = 32'b00000000000000000100010011101010;
assign LUT_1[30123] = 32'b11111111111111111101100101100110;
assign LUT_1[30124] = 32'b00000000000000010000011110110000;
assign LUT_1[30125] = 32'b00000000000000001001110000101100;
assign LUT_1[30126] = 32'b00000000000000001100001101000001;
assign LUT_1[30127] = 32'b00000000000000000101011110111101;
assign LUT_1[30128] = 32'b00000000000000001011010011000110;
assign LUT_1[30129] = 32'b00000000000000000100100101000010;
assign LUT_1[30130] = 32'b00000000000000000111000001010111;
assign LUT_1[30131] = 32'b00000000000000000000010011010011;
assign LUT_1[30132] = 32'b00000000000000010011001100011101;
assign LUT_1[30133] = 32'b00000000000000001100011110011001;
assign LUT_1[30134] = 32'b00000000000000001110111010101110;
assign LUT_1[30135] = 32'b00000000000000001000001100101010;
assign LUT_1[30136] = 32'b00000000000000001010100000111011;
assign LUT_1[30137] = 32'b00000000000000000011110010110111;
assign LUT_1[30138] = 32'b00000000000000000110001111001100;
assign LUT_1[30139] = 32'b11111111111111111111100001001000;
assign LUT_1[30140] = 32'b00000000000000010010011010010010;
assign LUT_1[30141] = 32'b00000000000000001011101100001110;
assign LUT_1[30142] = 32'b00000000000000001110001000100011;
assign LUT_1[30143] = 32'b00000000000000000111011010011111;
assign LUT_1[30144] = 32'b00000000000000001010011010001101;
assign LUT_1[30145] = 32'b00000000000000000011101100001001;
assign LUT_1[30146] = 32'b00000000000000000110001000011110;
assign LUT_1[30147] = 32'b11111111111111111111011010011010;
assign LUT_1[30148] = 32'b00000000000000010010010011100100;
assign LUT_1[30149] = 32'b00000000000000001011100101100000;
assign LUT_1[30150] = 32'b00000000000000001110000001110101;
assign LUT_1[30151] = 32'b00000000000000000111010011110001;
assign LUT_1[30152] = 32'b00000000000000001001101000000010;
assign LUT_1[30153] = 32'b00000000000000000010111001111110;
assign LUT_1[30154] = 32'b00000000000000000101010110010011;
assign LUT_1[30155] = 32'b11111111111111111110101000001111;
assign LUT_1[30156] = 32'b00000000000000010001100001011001;
assign LUT_1[30157] = 32'b00000000000000001010110011010101;
assign LUT_1[30158] = 32'b00000000000000001101001111101010;
assign LUT_1[30159] = 32'b00000000000000000110100001100110;
assign LUT_1[30160] = 32'b00000000000000001100010101101111;
assign LUT_1[30161] = 32'b00000000000000000101100111101011;
assign LUT_1[30162] = 32'b00000000000000001000000100000000;
assign LUT_1[30163] = 32'b00000000000000000001010101111100;
assign LUT_1[30164] = 32'b00000000000000010100001111000110;
assign LUT_1[30165] = 32'b00000000000000001101100001000010;
assign LUT_1[30166] = 32'b00000000000000001111111101010111;
assign LUT_1[30167] = 32'b00000000000000001001001111010011;
assign LUT_1[30168] = 32'b00000000000000001011100011100100;
assign LUT_1[30169] = 32'b00000000000000000100110101100000;
assign LUT_1[30170] = 32'b00000000000000000111010001110101;
assign LUT_1[30171] = 32'b00000000000000000000100011110001;
assign LUT_1[30172] = 32'b00000000000000010011011100111011;
assign LUT_1[30173] = 32'b00000000000000001100101110110111;
assign LUT_1[30174] = 32'b00000000000000001111001011001100;
assign LUT_1[30175] = 32'b00000000000000001000011101001000;
assign LUT_1[30176] = 32'b00000000000000001011010101001100;
assign LUT_1[30177] = 32'b00000000000000000100100111001000;
assign LUT_1[30178] = 32'b00000000000000000111000011011101;
assign LUT_1[30179] = 32'b00000000000000000000010101011001;
assign LUT_1[30180] = 32'b00000000000000010011001110100011;
assign LUT_1[30181] = 32'b00000000000000001100100000011111;
assign LUT_1[30182] = 32'b00000000000000001110111100110100;
assign LUT_1[30183] = 32'b00000000000000001000001110110000;
assign LUT_1[30184] = 32'b00000000000000001010100011000001;
assign LUT_1[30185] = 32'b00000000000000000011110100111101;
assign LUT_1[30186] = 32'b00000000000000000110010001010010;
assign LUT_1[30187] = 32'b11111111111111111111100011001110;
assign LUT_1[30188] = 32'b00000000000000010010011100011000;
assign LUT_1[30189] = 32'b00000000000000001011101110010100;
assign LUT_1[30190] = 32'b00000000000000001110001010101001;
assign LUT_1[30191] = 32'b00000000000000000111011100100101;
assign LUT_1[30192] = 32'b00000000000000001101010000101110;
assign LUT_1[30193] = 32'b00000000000000000110100010101010;
assign LUT_1[30194] = 32'b00000000000000001000111110111111;
assign LUT_1[30195] = 32'b00000000000000000010010000111011;
assign LUT_1[30196] = 32'b00000000000000010101001010000101;
assign LUT_1[30197] = 32'b00000000000000001110011100000001;
assign LUT_1[30198] = 32'b00000000000000010000111000010110;
assign LUT_1[30199] = 32'b00000000000000001010001010010010;
assign LUT_1[30200] = 32'b00000000000000001100011110100011;
assign LUT_1[30201] = 32'b00000000000000000101110000011111;
assign LUT_1[30202] = 32'b00000000000000001000001100110100;
assign LUT_1[30203] = 32'b00000000000000000001011110110000;
assign LUT_1[30204] = 32'b00000000000000010100010111111010;
assign LUT_1[30205] = 32'b00000000000000001101101001110110;
assign LUT_1[30206] = 32'b00000000000000010000000110001011;
assign LUT_1[30207] = 32'b00000000000000001001011000000111;
assign LUT_1[30208] = 32'b00000000000000000001010110110011;
assign LUT_1[30209] = 32'b11111111111111111010101000101111;
assign LUT_1[30210] = 32'b11111111111111111101000101000100;
assign LUT_1[30211] = 32'b11111111111111110110010111000000;
assign LUT_1[30212] = 32'b00000000000000001001010000001010;
assign LUT_1[30213] = 32'b00000000000000000010100010000110;
assign LUT_1[30214] = 32'b00000000000000000100111110011011;
assign LUT_1[30215] = 32'b11111111111111111110010000010111;
assign LUT_1[30216] = 32'b00000000000000000000100100101000;
assign LUT_1[30217] = 32'b11111111111111111001110110100100;
assign LUT_1[30218] = 32'b11111111111111111100010010111001;
assign LUT_1[30219] = 32'b11111111111111110101100100110101;
assign LUT_1[30220] = 32'b00000000000000001000011101111111;
assign LUT_1[30221] = 32'b00000000000000000001101111111011;
assign LUT_1[30222] = 32'b00000000000000000100001100010000;
assign LUT_1[30223] = 32'b11111111111111111101011110001100;
assign LUT_1[30224] = 32'b00000000000000000011010010010101;
assign LUT_1[30225] = 32'b11111111111111111100100100010001;
assign LUT_1[30226] = 32'b11111111111111111111000000100110;
assign LUT_1[30227] = 32'b11111111111111111000010010100010;
assign LUT_1[30228] = 32'b00000000000000001011001011101100;
assign LUT_1[30229] = 32'b00000000000000000100011101101000;
assign LUT_1[30230] = 32'b00000000000000000110111001111101;
assign LUT_1[30231] = 32'b00000000000000000000001011111001;
assign LUT_1[30232] = 32'b00000000000000000010100000001010;
assign LUT_1[30233] = 32'b11111111111111111011110010000110;
assign LUT_1[30234] = 32'b11111111111111111110001110011011;
assign LUT_1[30235] = 32'b11111111111111110111100000010111;
assign LUT_1[30236] = 32'b00000000000000001010011001100001;
assign LUT_1[30237] = 32'b00000000000000000011101011011101;
assign LUT_1[30238] = 32'b00000000000000000110000111110010;
assign LUT_1[30239] = 32'b11111111111111111111011001101110;
assign LUT_1[30240] = 32'b00000000000000000010010001110010;
assign LUT_1[30241] = 32'b11111111111111111011100011101110;
assign LUT_1[30242] = 32'b11111111111111111110000000000011;
assign LUT_1[30243] = 32'b11111111111111110111010001111111;
assign LUT_1[30244] = 32'b00000000000000001010001011001001;
assign LUT_1[30245] = 32'b00000000000000000011011101000101;
assign LUT_1[30246] = 32'b00000000000000000101111001011010;
assign LUT_1[30247] = 32'b11111111111111111111001011010110;
assign LUT_1[30248] = 32'b00000000000000000001011111100111;
assign LUT_1[30249] = 32'b11111111111111111010110001100011;
assign LUT_1[30250] = 32'b11111111111111111101001101111000;
assign LUT_1[30251] = 32'b11111111111111110110011111110100;
assign LUT_1[30252] = 32'b00000000000000001001011000111110;
assign LUT_1[30253] = 32'b00000000000000000010101010111010;
assign LUT_1[30254] = 32'b00000000000000000101000111001111;
assign LUT_1[30255] = 32'b11111111111111111110011001001011;
assign LUT_1[30256] = 32'b00000000000000000100001101010100;
assign LUT_1[30257] = 32'b11111111111111111101011111010000;
assign LUT_1[30258] = 32'b11111111111111111111111011100101;
assign LUT_1[30259] = 32'b11111111111111111001001101100001;
assign LUT_1[30260] = 32'b00000000000000001100000110101011;
assign LUT_1[30261] = 32'b00000000000000000101011000100111;
assign LUT_1[30262] = 32'b00000000000000000111110100111100;
assign LUT_1[30263] = 32'b00000000000000000001000110111000;
assign LUT_1[30264] = 32'b00000000000000000011011011001001;
assign LUT_1[30265] = 32'b11111111111111111100101101000101;
assign LUT_1[30266] = 32'b11111111111111111111001001011010;
assign LUT_1[30267] = 32'b11111111111111111000011011010110;
assign LUT_1[30268] = 32'b00000000000000001011010100100000;
assign LUT_1[30269] = 32'b00000000000000000100100110011100;
assign LUT_1[30270] = 32'b00000000000000000111000010110001;
assign LUT_1[30271] = 32'b00000000000000000000010100101101;
assign LUT_1[30272] = 32'b00000000000000000011010100011011;
assign LUT_1[30273] = 32'b11111111111111111100100110010111;
assign LUT_1[30274] = 32'b11111111111111111111000010101100;
assign LUT_1[30275] = 32'b11111111111111111000010100101000;
assign LUT_1[30276] = 32'b00000000000000001011001101110010;
assign LUT_1[30277] = 32'b00000000000000000100011111101110;
assign LUT_1[30278] = 32'b00000000000000000110111100000011;
assign LUT_1[30279] = 32'b00000000000000000000001101111111;
assign LUT_1[30280] = 32'b00000000000000000010100010010000;
assign LUT_1[30281] = 32'b11111111111111111011110100001100;
assign LUT_1[30282] = 32'b11111111111111111110010000100001;
assign LUT_1[30283] = 32'b11111111111111110111100010011101;
assign LUT_1[30284] = 32'b00000000000000001010011011100111;
assign LUT_1[30285] = 32'b00000000000000000011101101100011;
assign LUT_1[30286] = 32'b00000000000000000110001001111000;
assign LUT_1[30287] = 32'b11111111111111111111011011110100;
assign LUT_1[30288] = 32'b00000000000000000101001111111101;
assign LUT_1[30289] = 32'b11111111111111111110100001111001;
assign LUT_1[30290] = 32'b00000000000000000000111110001110;
assign LUT_1[30291] = 32'b11111111111111111010010000001010;
assign LUT_1[30292] = 32'b00000000000000001101001001010100;
assign LUT_1[30293] = 32'b00000000000000000110011011010000;
assign LUT_1[30294] = 32'b00000000000000001000110111100101;
assign LUT_1[30295] = 32'b00000000000000000010001001100001;
assign LUT_1[30296] = 32'b00000000000000000100011101110010;
assign LUT_1[30297] = 32'b11111111111111111101101111101110;
assign LUT_1[30298] = 32'b00000000000000000000001100000011;
assign LUT_1[30299] = 32'b11111111111111111001011101111111;
assign LUT_1[30300] = 32'b00000000000000001100010111001001;
assign LUT_1[30301] = 32'b00000000000000000101101001000101;
assign LUT_1[30302] = 32'b00000000000000001000000101011010;
assign LUT_1[30303] = 32'b00000000000000000001010111010110;
assign LUT_1[30304] = 32'b00000000000000000100001111011010;
assign LUT_1[30305] = 32'b11111111111111111101100001010110;
assign LUT_1[30306] = 32'b11111111111111111111111101101011;
assign LUT_1[30307] = 32'b11111111111111111001001111100111;
assign LUT_1[30308] = 32'b00000000000000001100001000110001;
assign LUT_1[30309] = 32'b00000000000000000101011010101101;
assign LUT_1[30310] = 32'b00000000000000000111110111000010;
assign LUT_1[30311] = 32'b00000000000000000001001000111110;
assign LUT_1[30312] = 32'b00000000000000000011011101001111;
assign LUT_1[30313] = 32'b11111111111111111100101111001011;
assign LUT_1[30314] = 32'b11111111111111111111001011100000;
assign LUT_1[30315] = 32'b11111111111111111000011101011100;
assign LUT_1[30316] = 32'b00000000000000001011010110100110;
assign LUT_1[30317] = 32'b00000000000000000100101000100010;
assign LUT_1[30318] = 32'b00000000000000000111000100110111;
assign LUT_1[30319] = 32'b00000000000000000000010110110011;
assign LUT_1[30320] = 32'b00000000000000000110001010111100;
assign LUT_1[30321] = 32'b11111111111111111111011100111000;
assign LUT_1[30322] = 32'b00000000000000000001111001001101;
assign LUT_1[30323] = 32'b11111111111111111011001011001001;
assign LUT_1[30324] = 32'b00000000000000001110000100010011;
assign LUT_1[30325] = 32'b00000000000000000111010110001111;
assign LUT_1[30326] = 32'b00000000000000001001110010100100;
assign LUT_1[30327] = 32'b00000000000000000011000100100000;
assign LUT_1[30328] = 32'b00000000000000000101011000110001;
assign LUT_1[30329] = 32'b11111111111111111110101010101101;
assign LUT_1[30330] = 32'b00000000000000000001000111000010;
assign LUT_1[30331] = 32'b11111111111111111010011000111110;
assign LUT_1[30332] = 32'b00000000000000001101010010001000;
assign LUT_1[30333] = 32'b00000000000000000110100100000100;
assign LUT_1[30334] = 32'b00000000000000001001000000011001;
assign LUT_1[30335] = 32'b00000000000000000010010010010101;
assign LUT_1[30336] = 32'b00000000000000000100010110110110;
assign LUT_1[30337] = 32'b11111111111111111101101000110010;
assign LUT_1[30338] = 32'b00000000000000000000000101000111;
assign LUT_1[30339] = 32'b11111111111111111001010111000011;
assign LUT_1[30340] = 32'b00000000000000001100010000001101;
assign LUT_1[30341] = 32'b00000000000000000101100010001001;
assign LUT_1[30342] = 32'b00000000000000000111111110011110;
assign LUT_1[30343] = 32'b00000000000000000001010000011010;
assign LUT_1[30344] = 32'b00000000000000000011100100101011;
assign LUT_1[30345] = 32'b11111111111111111100110110100111;
assign LUT_1[30346] = 32'b11111111111111111111010010111100;
assign LUT_1[30347] = 32'b11111111111111111000100100111000;
assign LUT_1[30348] = 32'b00000000000000001011011110000010;
assign LUT_1[30349] = 32'b00000000000000000100101111111110;
assign LUT_1[30350] = 32'b00000000000000000111001100010011;
assign LUT_1[30351] = 32'b00000000000000000000011110001111;
assign LUT_1[30352] = 32'b00000000000000000110010010011000;
assign LUT_1[30353] = 32'b11111111111111111111100100010100;
assign LUT_1[30354] = 32'b00000000000000000010000000101001;
assign LUT_1[30355] = 32'b11111111111111111011010010100101;
assign LUT_1[30356] = 32'b00000000000000001110001011101111;
assign LUT_1[30357] = 32'b00000000000000000111011101101011;
assign LUT_1[30358] = 32'b00000000000000001001111010000000;
assign LUT_1[30359] = 32'b00000000000000000011001011111100;
assign LUT_1[30360] = 32'b00000000000000000101100000001101;
assign LUT_1[30361] = 32'b11111111111111111110110010001001;
assign LUT_1[30362] = 32'b00000000000000000001001110011110;
assign LUT_1[30363] = 32'b11111111111111111010100000011010;
assign LUT_1[30364] = 32'b00000000000000001101011001100100;
assign LUT_1[30365] = 32'b00000000000000000110101011100000;
assign LUT_1[30366] = 32'b00000000000000001001000111110101;
assign LUT_1[30367] = 32'b00000000000000000010011001110001;
assign LUT_1[30368] = 32'b00000000000000000101010001110101;
assign LUT_1[30369] = 32'b11111111111111111110100011110001;
assign LUT_1[30370] = 32'b00000000000000000001000000000110;
assign LUT_1[30371] = 32'b11111111111111111010010010000010;
assign LUT_1[30372] = 32'b00000000000000001101001011001100;
assign LUT_1[30373] = 32'b00000000000000000110011101001000;
assign LUT_1[30374] = 32'b00000000000000001000111001011101;
assign LUT_1[30375] = 32'b00000000000000000010001011011001;
assign LUT_1[30376] = 32'b00000000000000000100011111101010;
assign LUT_1[30377] = 32'b11111111111111111101110001100110;
assign LUT_1[30378] = 32'b00000000000000000000001101111011;
assign LUT_1[30379] = 32'b11111111111111111001011111110111;
assign LUT_1[30380] = 32'b00000000000000001100011001000001;
assign LUT_1[30381] = 32'b00000000000000000101101010111101;
assign LUT_1[30382] = 32'b00000000000000001000000111010010;
assign LUT_1[30383] = 32'b00000000000000000001011001001110;
assign LUT_1[30384] = 32'b00000000000000000111001101010111;
assign LUT_1[30385] = 32'b00000000000000000000011111010011;
assign LUT_1[30386] = 32'b00000000000000000010111011101000;
assign LUT_1[30387] = 32'b11111111111111111100001101100100;
assign LUT_1[30388] = 32'b00000000000000001111000110101110;
assign LUT_1[30389] = 32'b00000000000000001000011000101010;
assign LUT_1[30390] = 32'b00000000000000001010110100111111;
assign LUT_1[30391] = 32'b00000000000000000100000110111011;
assign LUT_1[30392] = 32'b00000000000000000110011011001100;
assign LUT_1[30393] = 32'b11111111111111111111101101001000;
assign LUT_1[30394] = 32'b00000000000000000010001001011101;
assign LUT_1[30395] = 32'b11111111111111111011011011011001;
assign LUT_1[30396] = 32'b00000000000000001110010100100011;
assign LUT_1[30397] = 32'b00000000000000000111100110011111;
assign LUT_1[30398] = 32'b00000000000000001010000010110100;
assign LUT_1[30399] = 32'b00000000000000000011010100110000;
assign LUT_1[30400] = 32'b00000000000000000110010100011110;
assign LUT_1[30401] = 32'b11111111111111111111100110011010;
assign LUT_1[30402] = 32'b00000000000000000010000010101111;
assign LUT_1[30403] = 32'b11111111111111111011010100101011;
assign LUT_1[30404] = 32'b00000000000000001110001101110101;
assign LUT_1[30405] = 32'b00000000000000000111011111110001;
assign LUT_1[30406] = 32'b00000000000000001001111100000110;
assign LUT_1[30407] = 32'b00000000000000000011001110000010;
assign LUT_1[30408] = 32'b00000000000000000101100010010011;
assign LUT_1[30409] = 32'b11111111111111111110110100001111;
assign LUT_1[30410] = 32'b00000000000000000001010000100100;
assign LUT_1[30411] = 32'b11111111111111111010100010100000;
assign LUT_1[30412] = 32'b00000000000000001101011011101010;
assign LUT_1[30413] = 32'b00000000000000000110101101100110;
assign LUT_1[30414] = 32'b00000000000000001001001001111011;
assign LUT_1[30415] = 32'b00000000000000000010011011110111;
assign LUT_1[30416] = 32'b00000000000000001000010000000000;
assign LUT_1[30417] = 32'b00000000000000000001100001111100;
assign LUT_1[30418] = 32'b00000000000000000011111110010001;
assign LUT_1[30419] = 32'b11111111111111111101010000001101;
assign LUT_1[30420] = 32'b00000000000000010000001001010111;
assign LUT_1[30421] = 32'b00000000000000001001011011010011;
assign LUT_1[30422] = 32'b00000000000000001011110111101000;
assign LUT_1[30423] = 32'b00000000000000000101001001100100;
assign LUT_1[30424] = 32'b00000000000000000111011101110101;
assign LUT_1[30425] = 32'b00000000000000000000101111110001;
assign LUT_1[30426] = 32'b00000000000000000011001100000110;
assign LUT_1[30427] = 32'b11111111111111111100011110000010;
assign LUT_1[30428] = 32'b00000000000000001111010111001100;
assign LUT_1[30429] = 32'b00000000000000001000101001001000;
assign LUT_1[30430] = 32'b00000000000000001011000101011101;
assign LUT_1[30431] = 32'b00000000000000000100010111011001;
assign LUT_1[30432] = 32'b00000000000000000111001111011101;
assign LUT_1[30433] = 32'b00000000000000000000100001011001;
assign LUT_1[30434] = 32'b00000000000000000010111101101110;
assign LUT_1[30435] = 32'b11111111111111111100001111101010;
assign LUT_1[30436] = 32'b00000000000000001111001000110100;
assign LUT_1[30437] = 32'b00000000000000001000011010110000;
assign LUT_1[30438] = 32'b00000000000000001010110111000101;
assign LUT_1[30439] = 32'b00000000000000000100001001000001;
assign LUT_1[30440] = 32'b00000000000000000110011101010010;
assign LUT_1[30441] = 32'b11111111111111111111101111001110;
assign LUT_1[30442] = 32'b00000000000000000010001011100011;
assign LUT_1[30443] = 32'b11111111111111111011011101011111;
assign LUT_1[30444] = 32'b00000000000000001110010110101001;
assign LUT_1[30445] = 32'b00000000000000000111101000100101;
assign LUT_1[30446] = 32'b00000000000000001010000100111010;
assign LUT_1[30447] = 32'b00000000000000000011010110110110;
assign LUT_1[30448] = 32'b00000000000000001001001010111111;
assign LUT_1[30449] = 32'b00000000000000000010011100111011;
assign LUT_1[30450] = 32'b00000000000000000100111001010000;
assign LUT_1[30451] = 32'b11111111111111111110001011001100;
assign LUT_1[30452] = 32'b00000000000000010001000100010110;
assign LUT_1[30453] = 32'b00000000000000001010010110010010;
assign LUT_1[30454] = 32'b00000000000000001100110010100111;
assign LUT_1[30455] = 32'b00000000000000000110000100100011;
assign LUT_1[30456] = 32'b00000000000000001000011000110100;
assign LUT_1[30457] = 32'b00000000000000000001101010110000;
assign LUT_1[30458] = 32'b00000000000000000100000111000101;
assign LUT_1[30459] = 32'b11111111111111111101011001000001;
assign LUT_1[30460] = 32'b00000000000000010000010010001011;
assign LUT_1[30461] = 32'b00000000000000001001100100000111;
assign LUT_1[30462] = 32'b00000000000000001100000000011100;
assign LUT_1[30463] = 32'b00000000000000000101010010011000;
assign LUT_1[30464] = 32'b11111111111111111111001010111111;
assign LUT_1[30465] = 32'b11111111111111111000011100111011;
assign LUT_1[30466] = 32'b11111111111111111010111001010000;
assign LUT_1[30467] = 32'b11111111111111110100001011001100;
assign LUT_1[30468] = 32'b00000000000000000111000100010110;
assign LUT_1[30469] = 32'b00000000000000000000010110010010;
assign LUT_1[30470] = 32'b00000000000000000010110010100111;
assign LUT_1[30471] = 32'b11111111111111111100000100100011;
assign LUT_1[30472] = 32'b11111111111111111110011000110100;
assign LUT_1[30473] = 32'b11111111111111110111101010110000;
assign LUT_1[30474] = 32'b11111111111111111010000111000101;
assign LUT_1[30475] = 32'b11111111111111110011011001000001;
assign LUT_1[30476] = 32'b00000000000000000110010010001011;
assign LUT_1[30477] = 32'b11111111111111111111100100000111;
assign LUT_1[30478] = 32'b00000000000000000010000000011100;
assign LUT_1[30479] = 32'b11111111111111111011010010011000;
assign LUT_1[30480] = 32'b00000000000000000001000110100001;
assign LUT_1[30481] = 32'b11111111111111111010011000011101;
assign LUT_1[30482] = 32'b11111111111111111100110100110010;
assign LUT_1[30483] = 32'b11111111111111110110000110101110;
assign LUT_1[30484] = 32'b00000000000000001000111111111000;
assign LUT_1[30485] = 32'b00000000000000000010010001110100;
assign LUT_1[30486] = 32'b00000000000000000100101110001001;
assign LUT_1[30487] = 32'b11111111111111111110000000000101;
assign LUT_1[30488] = 32'b00000000000000000000010100010110;
assign LUT_1[30489] = 32'b11111111111111111001100110010010;
assign LUT_1[30490] = 32'b11111111111111111100000010100111;
assign LUT_1[30491] = 32'b11111111111111110101010100100011;
assign LUT_1[30492] = 32'b00000000000000001000001101101101;
assign LUT_1[30493] = 32'b00000000000000000001011111101001;
assign LUT_1[30494] = 32'b00000000000000000011111011111110;
assign LUT_1[30495] = 32'b11111111111111111101001101111010;
assign LUT_1[30496] = 32'b00000000000000000000000101111110;
assign LUT_1[30497] = 32'b11111111111111111001010111111010;
assign LUT_1[30498] = 32'b11111111111111111011110100001111;
assign LUT_1[30499] = 32'b11111111111111110101000110001011;
assign LUT_1[30500] = 32'b00000000000000000111111111010101;
assign LUT_1[30501] = 32'b00000000000000000001010001010001;
assign LUT_1[30502] = 32'b00000000000000000011101101100110;
assign LUT_1[30503] = 32'b11111111111111111100111111100010;
assign LUT_1[30504] = 32'b11111111111111111111010011110011;
assign LUT_1[30505] = 32'b11111111111111111000100101101111;
assign LUT_1[30506] = 32'b11111111111111111011000010000100;
assign LUT_1[30507] = 32'b11111111111111110100010100000000;
assign LUT_1[30508] = 32'b00000000000000000111001101001010;
assign LUT_1[30509] = 32'b00000000000000000000011111000110;
assign LUT_1[30510] = 32'b00000000000000000010111011011011;
assign LUT_1[30511] = 32'b11111111111111111100001101010111;
assign LUT_1[30512] = 32'b00000000000000000010000001100000;
assign LUT_1[30513] = 32'b11111111111111111011010011011100;
assign LUT_1[30514] = 32'b11111111111111111101101111110001;
assign LUT_1[30515] = 32'b11111111111111110111000001101101;
assign LUT_1[30516] = 32'b00000000000000001001111010110111;
assign LUT_1[30517] = 32'b00000000000000000011001100110011;
assign LUT_1[30518] = 32'b00000000000000000101101001001000;
assign LUT_1[30519] = 32'b11111111111111111110111011000100;
assign LUT_1[30520] = 32'b00000000000000000001001111010101;
assign LUT_1[30521] = 32'b11111111111111111010100001010001;
assign LUT_1[30522] = 32'b11111111111111111100111101100110;
assign LUT_1[30523] = 32'b11111111111111110110001111100010;
assign LUT_1[30524] = 32'b00000000000000001001001000101100;
assign LUT_1[30525] = 32'b00000000000000000010011010101000;
assign LUT_1[30526] = 32'b00000000000000000100110110111101;
assign LUT_1[30527] = 32'b11111111111111111110001000111001;
assign LUT_1[30528] = 32'b00000000000000000001001000100111;
assign LUT_1[30529] = 32'b11111111111111111010011010100011;
assign LUT_1[30530] = 32'b11111111111111111100110110111000;
assign LUT_1[30531] = 32'b11111111111111110110001000110100;
assign LUT_1[30532] = 32'b00000000000000001001000001111110;
assign LUT_1[30533] = 32'b00000000000000000010010011111010;
assign LUT_1[30534] = 32'b00000000000000000100110000001111;
assign LUT_1[30535] = 32'b11111111111111111110000010001011;
assign LUT_1[30536] = 32'b00000000000000000000010110011100;
assign LUT_1[30537] = 32'b11111111111111111001101000011000;
assign LUT_1[30538] = 32'b11111111111111111100000100101101;
assign LUT_1[30539] = 32'b11111111111111110101010110101001;
assign LUT_1[30540] = 32'b00000000000000001000001111110011;
assign LUT_1[30541] = 32'b00000000000000000001100001101111;
assign LUT_1[30542] = 32'b00000000000000000011111110000100;
assign LUT_1[30543] = 32'b11111111111111111101010000000000;
assign LUT_1[30544] = 32'b00000000000000000011000100001001;
assign LUT_1[30545] = 32'b11111111111111111100010110000101;
assign LUT_1[30546] = 32'b11111111111111111110110010011010;
assign LUT_1[30547] = 32'b11111111111111111000000100010110;
assign LUT_1[30548] = 32'b00000000000000001010111101100000;
assign LUT_1[30549] = 32'b00000000000000000100001111011100;
assign LUT_1[30550] = 32'b00000000000000000110101011110001;
assign LUT_1[30551] = 32'b11111111111111111111111101101101;
assign LUT_1[30552] = 32'b00000000000000000010010001111110;
assign LUT_1[30553] = 32'b11111111111111111011100011111010;
assign LUT_1[30554] = 32'b11111111111111111110000000001111;
assign LUT_1[30555] = 32'b11111111111111110111010010001011;
assign LUT_1[30556] = 32'b00000000000000001010001011010101;
assign LUT_1[30557] = 32'b00000000000000000011011101010001;
assign LUT_1[30558] = 32'b00000000000000000101111001100110;
assign LUT_1[30559] = 32'b11111111111111111111001011100010;
assign LUT_1[30560] = 32'b00000000000000000010000011100110;
assign LUT_1[30561] = 32'b11111111111111111011010101100010;
assign LUT_1[30562] = 32'b11111111111111111101110001110111;
assign LUT_1[30563] = 32'b11111111111111110111000011110011;
assign LUT_1[30564] = 32'b00000000000000001001111100111101;
assign LUT_1[30565] = 32'b00000000000000000011001110111001;
assign LUT_1[30566] = 32'b00000000000000000101101011001110;
assign LUT_1[30567] = 32'b11111111111111111110111101001010;
assign LUT_1[30568] = 32'b00000000000000000001010001011011;
assign LUT_1[30569] = 32'b11111111111111111010100011010111;
assign LUT_1[30570] = 32'b11111111111111111100111111101100;
assign LUT_1[30571] = 32'b11111111111111110110010001101000;
assign LUT_1[30572] = 32'b00000000000000001001001010110010;
assign LUT_1[30573] = 32'b00000000000000000010011100101110;
assign LUT_1[30574] = 32'b00000000000000000100111001000011;
assign LUT_1[30575] = 32'b11111111111111111110001010111111;
assign LUT_1[30576] = 32'b00000000000000000011111111001000;
assign LUT_1[30577] = 32'b11111111111111111101010001000100;
assign LUT_1[30578] = 32'b11111111111111111111101101011001;
assign LUT_1[30579] = 32'b11111111111111111000111111010101;
assign LUT_1[30580] = 32'b00000000000000001011111000011111;
assign LUT_1[30581] = 32'b00000000000000000101001010011011;
assign LUT_1[30582] = 32'b00000000000000000111100110110000;
assign LUT_1[30583] = 32'b00000000000000000000111000101100;
assign LUT_1[30584] = 32'b00000000000000000011001100111101;
assign LUT_1[30585] = 32'b11111111111111111100011110111001;
assign LUT_1[30586] = 32'b11111111111111111110111011001110;
assign LUT_1[30587] = 32'b11111111111111111000001101001010;
assign LUT_1[30588] = 32'b00000000000000001011000110010100;
assign LUT_1[30589] = 32'b00000000000000000100011000010000;
assign LUT_1[30590] = 32'b00000000000000000110110100100101;
assign LUT_1[30591] = 32'b00000000000000000000000110100001;
assign LUT_1[30592] = 32'b00000000000000000010001011000010;
assign LUT_1[30593] = 32'b11111111111111111011011100111110;
assign LUT_1[30594] = 32'b11111111111111111101111001010011;
assign LUT_1[30595] = 32'b11111111111111110111001011001111;
assign LUT_1[30596] = 32'b00000000000000001010000100011001;
assign LUT_1[30597] = 32'b00000000000000000011010110010101;
assign LUT_1[30598] = 32'b00000000000000000101110010101010;
assign LUT_1[30599] = 32'b11111111111111111111000100100110;
assign LUT_1[30600] = 32'b00000000000000000001011000110111;
assign LUT_1[30601] = 32'b11111111111111111010101010110011;
assign LUT_1[30602] = 32'b11111111111111111101000111001000;
assign LUT_1[30603] = 32'b11111111111111110110011001000100;
assign LUT_1[30604] = 32'b00000000000000001001010010001110;
assign LUT_1[30605] = 32'b00000000000000000010100100001010;
assign LUT_1[30606] = 32'b00000000000000000101000000011111;
assign LUT_1[30607] = 32'b11111111111111111110010010011011;
assign LUT_1[30608] = 32'b00000000000000000100000110100100;
assign LUT_1[30609] = 32'b11111111111111111101011000100000;
assign LUT_1[30610] = 32'b11111111111111111111110100110101;
assign LUT_1[30611] = 32'b11111111111111111001000110110001;
assign LUT_1[30612] = 32'b00000000000000001011111111111011;
assign LUT_1[30613] = 32'b00000000000000000101010001110111;
assign LUT_1[30614] = 32'b00000000000000000111101110001100;
assign LUT_1[30615] = 32'b00000000000000000001000000001000;
assign LUT_1[30616] = 32'b00000000000000000011010100011001;
assign LUT_1[30617] = 32'b11111111111111111100100110010101;
assign LUT_1[30618] = 32'b11111111111111111111000010101010;
assign LUT_1[30619] = 32'b11111111111111111000010100100110;
assign LUT_1[30620] = 32'b00000000000000001011001101110000;
assign LUT_1[30621] = 32'b00000000000000000100011111101100;
assign LUT_1[30622] = 32'b00000000000000000110111100000001;
assign LUT_1[30623] = 32'b00000000000000000000001101111101;
assign LUT_1[30624] = 32'b00000000000000000011000110000001;
assign LUT_1[30625] = 32'b11111111111111111100010111111101;
assign LUT_1[30626] = 32'b11111111111111111110110100010010;
assign LUT_1[30627] = 32'b11111111111111111000000110001110;
assign LUT_1[30628] = 32'b00000000000000001010111111011000;
assign LUT_1[30629] = 32'b00000000000000000100010001010100;
assign LUT_1[30630] = 32'b00000000000000000110101101101001;
assign LUT_1[30631] = 32'b11111111111111111111111111100101;
assign LUT_1[30632] = 32'b00000000000000000010010011110110;
assign LUT_1[30633] = 32'b11111111111111111011100101110010;
assign LUT_1[30634] = 32'b11111111111111111110000010000111;
assign LUT_1[30635] = 32'b11111111111111110111010100000011;
assign LUT_1[30636] = 32'b00000000000000001010001101001101;
assign LUT_1[30637] = 32'b00000000000000000011011111001001;
assign LUT_1[30638] = 32'b00000000000000000101111011011110;
assign LUT_1[30639] = 32'b11111111111111111111001101011010;
assign LUT_1[30640] = 32'b00000000000000000101000001100011;
assign LUT_1[30641] = 32'b11111111111111111110010011011111;
assign LUT_1[30642] = 32'b00000000000000000000101111110100;
assign LUT_1[30643] = 32'b11111111111111111010000001110000;
assign LUT_1[30644] = 32'b00000000000000001100111010111010;
assign LUT_1[30645] = 32'b00000000000000000110001100110110;
assign LUT_1[30646] = 32'b00000000000000001000101001001011;
assign LUT_1[30647] = 32'b00000000000000000001111011000111;
assign LUT_1[30648] = 32'b00000000000000000100001111011000;
assign LUT_1[30649] = 32'b11111111111111111101100001010100;
assign LUT_1[30650] = 32'b11111111111111111111111101101001;
assign LUT_1[30651] = 32'b11111111111111111001001111100101;
assign LUT_1[30652] = 32'b00000000000000001100001000101111;
assign LUT_1[30653] = 32'b00000000000000000101011010101011;
assign LUT_1[30654] = 32'b00000000000000000111110111000000;
assign LUT_1[30655] = 32'b00000000000000000001001000111100;
assign LUT_1[30656] = 32'b00000000000000000100001000101010;
assign LUT_1[30657] = 32'b11111111111111111101011010100110;
assign LUT_1[30658] = 32'b11111111111111111111110110111011;
assign LUT_1[30659] = 32'b11111111111111111001001000110111;
assign LUT_1[30660] = 32'b00000000000000001100000010000001;
assign LUT_1[30661] = 32'b00000000000000000101010011111101;
assign LUT_1[30662] = 32'b00000000000000000111110000010010;
assign LUT_1[30663] = 32'b00000000000000000001000010001110;
assign LUT_1[30664] = 32'b00000000000000000011010110011111;
assign LUT_1[30665] = 32'b11111111111111111100101000011011;
assign LUT_1[30666] = 32'b11111111111111111111000100110000;
assign LUT_1[30667] = 32'b11111111111111111000010110101100;
assign LUT_1[30668] = 32'b00000000000000001011001111110110;
assign LUT_1[30669] = 32'b00000000000000000100100001110010;
assign LUT_1[30670] = 32'b00000000000000000110111110000111;
assign LUT_1[30671] = 32'b00000000000000000000010000000011;
assign LUT_1[30672] = 32'b00000000000000000110000100001100;
assign LUT_1[30673] = 32'b11111111111111111111010110001000;
assign LUT_1[30674] = 32'b00000000000000000001110010011101;
assign LUT_1[30675] = 32'b11111111111111111011000100011001;
assign LUT_1[30676] = 32'b00000000000000001101111101100011;
assign LUT_1[30677] = 32'b00000000000000000111001111011111;
assign LUT_1[30678] = 32'b00000000000000001001101011110100;
assign LUT_1[30679] = 32'b00000000000000000010111101110000;
assign LUT_1[30680] = 32'b00000000000000000101010010000001;
assign LUT_1[30681] = 32'b11111111111111111110100011111101;
assign LUT_1[30682] = 32'b00000000000000000001000000010010;
assign LUT_1[30683] = 32'b11111111111111111010010010001110;
assign LUT_1[30684] = 32'b00000000000000001101001011011000;
assign LUT_1[30685] = 32'b00000000000000000110011101010100;
assign LUT_1[30686] = 32'b00000000000000001000111001101001;
assign LUT_1[30687] = 32'b00000000000000000010001011100101;
assign LUT_1[30688] = 32'b00000000000000000101000011101001;
assign LUT_1[30689] = 32'b11111111111111111110010101100101;
assign LUT_1[30690] = 32'b00000000000000000000110001111010;
assign LUT_1[30691] = 32'b11111111111111111010000011110110;
assign LUT_1[30692] = 32'b00000000000000001100111101000000;
assign LUT_1[30693] = 32'b00000000000000000110001110111100;
assign LUT_1[30694] = 32'b00000000000000001000101011010001;
assign LUT_1[30695] = 32'b00000000000000000001111101001101;
assign LUT_1[30696] = 32'b00000000000000000100010001011110;
assign LUT_1[30697] = 32'b11111111111111111101100011011010;
assign LUT_1[30698] = 32'b11111111111111111111111111101111;
assign LUT_1[30699] = 32'b11111111111111111001010001101011;
assign LUT_1[30700] = 32'b00000000000000001100001010110101;
assign LUT_1[30701] = 32'b00000000000000000101011100110001;
assign LUT_1[30702] = 32'b00000000000000000111111001000110;
assign LUT_1[30703] = 32'b00000000000000000001001011000010;
assign LUT_1[30704] = 32'b00000000000000000110111111001011;
assign LUT_1[30705] = 32'b00000000000000000000010001000111;
assign LUT_1[30706] = 32'b00000000000000000010101101011100;
assign LUT_1[30707] = 32'b11111111111111111011111111011000;
assign LUT_1[30708] = 32'b00000000000000001110111000100010;
assign LUT_1[30709] = 32'b00000000000000001000001010011110;
assign LUT_1[30710] = 32'b00000000000000001010100110110011;
assign LUT_1[30711] = 32'b00000000000000000011111000101111;
assign LUT_1[30712] = 32'b00000000000000000110001101000000;
assign LUT_1[30713] = 32'b11111111111111111111011110111100;
assign LUT_1[30714] = 32'b00000000000000000001111011010001;
assign LUT_1[30715] = 32'b11111111111111111011001101001101;
assign LUT_1[30716] = 32'b00000000000000001110000110010111;
assign LUT_1[30717] = 32'b00000000000000000111011000010011;
assign LUT_1[30718] = 32'b00000000000000001001110100101000;
assign LUT_1[30719] = 32'b00000000000000000011000110100100;
assign LUT_1[30720] = 32'b00000000000000000010010011100001;
assign LUT_1[30721] = 32'b11111111111111111011100101011101;
assign LUT_1[30722] = 32'b11111111111111111110000001110010;
assign LUT_1[30723] = 32'b11111111111111110111010011101110;
assign LUT_1[30724] = 32'b00000000000000001010001100111000;
assign LUT_1[30725] = 32'b00000000000000000011011110110100;
assign LUT_1[30726] = 32'b00000000000000000101111011001001;
assign LUT_1[30727] = 32'b11111111111111111111001101000101;
assign LUT_1[30728] = 32'b00000000000000000001100001010110;
assign LUT_1[30729] = 32'b11111111111111111010110011010010;
assign LUT_1[30730] = 32'b11111111111111111101001111100111;
assign LUT_1[30731] = 32'b11111111111111110110100001100011;
assign LUT_1[30732] = 32'b00000000000000001001011010101101;
assign LUT_1[30733] = 32'b00000000000000000010101100101001;
assign LUT_1[30734] = 32'b00000000000000000101001000111110;
assign LUT_1[30735] = 32'b11111111111111111110011010111010;
assign LUT_1[30736] = 32'b00000000000000000100001111000011;
assign LUT_1[30737] = 32'b11111111111111111101100000111111;
assign LUT_1[30738] = 32'b11111111111111111111111101010100;
assign LUT_1[30739] = 32'b11111111111111111001001111010000;
assign LUT_1[30740] = 32'b00000000000000001100001000011010;
assign LUT_1[30741] = 32'b00000000000000000101011010010110;
assign LUT_1[30742] = 32'b00000000000000000111110110101011;
assign LUT_1[30743] = 32'b00000000000000000001001000100111;
assign LUT_1[30744] = 32'b00000000000000000011011100111000;
assign LUT_1[30745] = 32'b11111111111111111100101110110100;
assign LUT_1[30746] = 32'b11111111111111111111001011001001;
assign LUT_1[30747] = 32'b11111111111111111000011101000101;
assign LUT_1[30748] = 32'b00000000000000001011010110001111;
assign LUT_1[30749] = 32'b00000000000000000100101000001011;
assign LUT_1[30750] = 32'b00000000000000000111000100100000;
assign LUT_1[30751] = 32'b00000000000000000000010110011100;
assign LUT_1[30752] = 32'b00000000000000000011001110100000;
assign LUT_1[30753] = 32'b11111111111111111100100000011100;
assign LUT_1[30754] = 32'b11111111111111111110111100110001;
assign LUT_1[30755] = 32'b11111111111111111000001110101101;
assign LUT_1[30756] = 32'b00000000000000001011000111110111;
assign LUT_1[30757] = 32'b00000000000000000100011001110011;
assign LUT_1[30758] = 32'b00000000000000000110110110001000;
assign LUT_1[30759] = 32'b00000000000000000000001000000100;
assign LUT_1[30760] = 32'b00000000000000000010011100010101;
assign LUT_1[30761] = 32'b11111111111111111011101110010001;
assign LUT_1[30762] = 32'b11111111111111111110001010100110;
assign LUT_1[30763] = 32'b11111111111111110111011100100010;
assign LUT_1[30764] = 32'b00000000000000001010010101101100;
assign LUT_1[30765] = 32'b00000000000000000011100111101000;
assign LUT_1[30766] = 32'b00000000000000000110000011111101;
assign LUT_1[30767] = 32'b11111111111111111111010101111001;
assign LUT_1[30768] = 32'b00000000000000000101001010000010;
assign LUT_1[30769] = 32'b11111111111111111110011011111110;
assign LUT_1[30770] = 32'b00000000000000000000111000010011;
assign LUT_1[30771] = 32'b11111111111111111010001010001111;
assign LUT_1[30772] = 32'b00000000000000001101000011011001;
assign LUT_1[30773] = 32'b00000000000000000110010101010101;
assign LUT_1[30774] = 32'b00000000000000001000110001101010;
assign LUT_1[30775] = 32'b00000000000000000010000011100110;
assign LUT_1[30776] = 32'b00000000000000000100010111110111;
assign LUT_1[30777] = 32'b11111111111111111101101001110011;
assign LUT_1[30778] = 32'b00000000000000000000000110001000;
assign LUT_1[30779] = 32'b11111111111111111001011000000100;
assign LUT_1[30780] = 32'b00000000000000001100010001001110;
assign LUT_1[30781] = 32'b00000000000000000101100011001010;
assign LUT_1[30782] = 32'b00000000000000000111111111011111;
assign LUT_1[30783] = 32'b00000000000000000001010001011011;
assign LUT_1[30784] = 32'b00000000000000000100010001001001;
assign LUT_1[30785] = 32'b11111111111111111101100011000101;
assign LUT_1[30786] = 32'b11111111111111111111111111011010;
assign LUT_1[30787] = 32'b11111111111111111001010001010110;
assign LUT_1[30788] = 32'b00000000000000001100001010100000;
assign LUT_1[30789] = 32'b00000000000000000101011100011100;
assign LUT_1[30790] = 32'b00000000000000000111111000110001;
assign LUT_1[30791] = 32'b00000000000000000001001010101101;
assign LUT_1[30792] = 32'b00000000000000000011011110111110;
assign LUT_1[30793] = 32'b11111111111111111100110000111010;
assign LUT_1[30794] = 32'b11111111111111111111001101001111;
assign LUT_1[30795] = 32'b11111111111111111000011111001011;
assign LUT_1[30796] = 32'b00000000000000001011011000010101;
assign LUT_1[30797] = 32'b00000000000000000100101010010001;
assign LUT_1[30798] = 32'b00000000000000000111000110100110;
assign LUT_1[30799] = 32'b00000000000000000000011000100010;
assign LUT_1[30800] = 32'b00000000000000000110001100101011;
assign LUT_1[30801] = 32'b11111111111111111111011110100111;
assign LUT_1[30802] = 32'b00000000000000000001111010111100;
assign LUT_1[30803] = 32'b11111111111111111011001100111000;
assign LUT_1[30804] = 32'b00000000000000001110000110000010;
assign LUT_1[30805] = 32'b00000000000000000111010111111110;
assign LUT_1[30806] = 32'b00000000000000001001110100010011;
assign LUT_1[30807] = 32'b00000000000000000011000110001111;
assign LUT_1[30808] = 32'b00000000000000000101011010100000;
assign LUT_1[30809] = 32'b11111111111111111110101100011100;
assign LUT_1[30810] = 32'b00000000000000000001001000110001;
assign LUT_1[30811] = 32'b11111111111111111010011010101101;
assign LUT_1[30812] = 32'b00000000000000001101010011110111;
assign LUT_1[30813] = 32'b00000000000000000110100101110011;
assign LUT_1[30814] = 32'b00000000000000001001000010001000;
assign LUT_1[30815] = 32'b00000000000000000010010100000100;
assign LUT_1[30816] = 32'b00000000000000000101001100001000;
assign LUT_1[30817] = 32'b11111111111111111110011110000100;
assign LUT_1[30818] = 32'b00000000000000000000111010011001;
assign LUT_1[30819] = 32'b11111111111111111010001100010101;
assign LUT_1[30820] = 32'b00000000000000001101000101011111;
assign LUT_1[30821] = 32'b00000000000000000110010111011011;
assign LUT_1[30822] = 32'b00000000000000001000110011110000;
assign LUT_1[30823] = 32'b00000000000000000010000101101100;
assign LUT_1[30824] = 32'b00000000000000000100011001111101;
assign LUT_1[30825] = 32'b11111111111111111101101011111001;
assign LUT_1[30826] = 32'b00000000000000000000001000001110;
assign LUT_1[30827] = 32'b11111111111111111001011010001010;
assign LUT_1[30828] = 32'b00000000000000001100010011010100;
assign LUT_1[30829] = 32'b00000000000000000101100101010000;
assign LUT_1[30830] = 32'b00000000000000001000000001100101;
assign LUT_1[30831] = 32'b00000000000000000001010011100001;
assign LUT_1[30832] = 32'b00000000000000000111000111101010;
assign LUT_1[30833] = 32'b00000000000000000000011001100110;
assign LUT_1[30834] = 32'b00000000000000000010110101111011;
assign LUT_1[30835] = 32'b11111111111111111100000111110111;
assign LUT_1[30836] = 32'b00000000000000001111000001000001;
assign LUT_1[30837] = 32'b00000000000000001000010010111101;
assign LUT_1[30838] = 32'b00000000000000001010101111010010;
assign LUT_1[30839] = 32'b00000000000000000100000001001110;
assign LUT_1[30840] = 32'b00000000000000000110010101011111;
assign LUT_1[30841] = 32'b11111111111111111111100111011011;
assign LUT_1[30842] = 32'b00000000000000000010000011110000;
assign LUT_1[30843] = 32'b11111111111111111011010101101100;
assign LUT_1[30844] = 32'b00000000000000001110001110110110;
assign LUT_1[30845] = 32'b00000000000000000111100000110010;
assign LUT_1[30846] = 32'b00000000000000001001111101000111;
assign LUT_1[30847] = 32'b00000000000000000011001111000011;
assign LUT_1[30848] = 32'b00000000000000000101010011100100;
assign LUT_1[30849] = 32'b11111111111111111110100101100000;
assign LUT_1[30850] = 32'b00000000000000000001000001110101;
assign LUT_1[30851] = 32'b11111111111111111010010011110001;
assign LUT_1[30852] = 32'b00000000000000001101001100111011;
assign LUT_1[30853] = 32'b00000000000000000110011110110111;
assign LUT_1[30854] = 32'b00000000000000001000111011001100;
assign LUT_1[30855] = 32'b00000000000000000010001101001000;
assign LUT_1[30856] = 32'b00000000000000000100100001011001;
assign LUT_1[30857] = 32'b11111111111111111101110011010101;
assign LUT_1[30858] = 32'b00000000000000000000001111101010;
assign LUT_1[30859] = 32'b11111111111111111001100001100110;
assign LUT_1[30860] = 32'b00000000000000001100011010110000;
assign LUT_1[30861] = 32'b00000000000000000101101100101100;
assign LUT_1[30862] = 32'b00000000000000001000001001000001;
assign LUT_1[30863] = 32'b00000000000000000001011010111101;
assign LUT_1[30864] = 32'b00000000000000000111001111000110;
assign LUT_1[30865] = 32'b00000000000000000000100001000010;
assign LUT_1[30866] = 32'b00000000000000000010111101010111;
assign LUT_1[30867] = 32'b11111111111111111100001111010011;
assign LUT_1[30868] = 32'b00000000000000001111001000011101;
assign LUT_1[30869] = 32'b00000000000000001000011010011001;
assign LUT_1[30870] = 32'b00000000000000001010110110101110;
assign LUT_1[30871] = 32'b00000000000000000100001000101010;
assign LUT_1[30872] = 32'b00000000000000000110011100111011;
assign LUT_1[30873] = 32'b11111111111111111111101110110111;
assign LUT_1[30874] = 32'b00000000000000000010001011001100;
assign LUT_1[30875] = 32'b11111111111111111011011101001000;
assign LUT_1[30876] = 32'b00000000000000001110010110010010;
assign LUT_1[30877] = 32'b00000000000000000111101000001110;
assign LUT_1[30878] = 32'b00000000000000001010000100100011;
assign LUT_1[30879] = 32'b00000000000000000011010110011111;
assign LUT_1[30880] = 32'b00000000000000000110001110100011;
assign LUT_1[30881] = 32'b11111111111111111111100000011111;
assign LUT_1[30882] = 32'b00000000000000000001111100110100;
assign LUT_1[30883] = 32'b11111111111111111011001110110000;
assign LUT_1[30884] = 32'b00000000000000001110000111111010;
assign LUT_1[30885] = 32'b00000000000000000111011001110110;
assign LUT_1[30886] = 32'b00000000000000001001110110001011;
assign LUT_1[30887] = 32'b00000000000000000011001000000111;
assign LUT_1[30888] = 32'b00000000000000000101011100011000;
assign LUT_1[30889] = 32'b11111111111111111110101110010100;
assign LUT_1[30890] = 32'b00000000000000000001001010101001;
assign LUT_1[30891] = 32'b11111111111111111010011100100101;
assign LUT_1[30892] = 32'b00000000000000001101010101101111;
assign LUT_1[30893] = 32'b00000000000000000110100111101011;
assign LUT_1[30894] = 32'b00000000000000001001000100000000;
assign LUT_1[30895] = 32'b00000000000000000010010101111100;
assign LUT_1[30896] = 32'b00000000000000001000001010000101;
assign LUT_1[30897] = 32'b00000000000000000001011100000001;
assign LUT_1[30898] = 32'b00000000000000000011111000010110;
assign LUT_1[30899] = 32'b11111111111111111101001010010010;
assign LUT_1[30900] = 32'b00000000000000010000000011011100;
assign LUT_1[30901] = 32'b00000000000000001001010101011000;
assign LUT_1[30902] = 32'b00000000000000001011110001101101;
assign LUT_1[30903] = 32'b00000000000000000101000011101001;
assign LUT_1[30904] = 32'b00000000000000000111010111111010;
assign LUT_1[30905] = 32'b00000000000000000000101001110110;
assign LUT_1[30906] = 32'b00000000000000000011000110001011;
assign LUT_1[30907] = 32'b11111111111111111100011000000111;
assign LUT_1[30908] = 32'b00000000000000001111010001010001;
assign LUT_1[30909] = 32'b00000000000000001000100011001101;
assign LUT_1[30910] = 32'b00000000000000001010111111100010;
assign LUT_1[30911] = 32'b00000000000000000100010001011110;
assign LUT_1[30912] = 32'b00000000000000000111010001001100;
assign LUT_1[30913] = 32'b00000000000000000000100011001000;
assign LUT_1[30914] = 32'b00000000000000000010111111011101;
assign LUT_1[30915] = 32'b11111111111111111100010001011001;
assign LUT_1[30916] = 32'b00000000000000001111001010100011;
assign LUT_1[30917] = 32'b00000000000000001000011100011111;
assign LUT_1[30918] = 32'b00000000000000001010111000110100;
assign LUT_1[30919] = 32'b00000000000000000100001010110000;
assign LUT_1[30920] = 32'b00000000000000000110011111000001;
assign LUT_1[30921] = 32'b11111111111111111111110000111101;
assign LUT_1[30922] = 32'b00000000000000000010001101010010;
assign LUT_1[30923] = 32'b11111111111111111011011111001110;
assign LUT_1[30924] = 32'b00000000000000001110011000011000;
assign LUT_1[30925] = 32'b00000000000000000111101010010100;
assign LUT_1[30926] = 32'b00000000000000001010000110101001;
assign LUT_1[30927] = 32'b00000000000000000011011000100101;
assign LUT_1[30928] = 32'b00000000000000001001001100101110;
assign LUT_1[30929] = 32'b00000000000000000010011110101010;
assign LUT_1[30930] = 32'b00000000000000000100111010111111;
assign LUT_1[30931] = 32'b11111111111111111110001100111011;
assign LUT_1[30932] = 32'b00000000000000010001000110000101;
assign LUT_1[30933] = 32'b00000000000000001010011000000001;
assign LUT_1[30934] = 32'b00000000000000001100110100010110;
assign LUT_1[30935] = 32'b00000000000000000110000110010010;
assign LUT_1[30936] = 32'b00000000000000001000011010100011;
assign LUT_1[30937] = 32'b00000000000000000001101100011111;
assign LUT_1[30938] = 32'b00000000000000000100001000110100;
assign LUT_1[30939] = 32'b11111111111111111101011010110000;
assign LUT_1[30940] = 32'b00000000000000010000010011111010;
assign LUT_1[30941] = 32'b00000000000000001001100101110110;
assign LUT_1[30942] = 32'b00000000000000001100000010001011;
assign LUT_1[30943] = 32'b00000000000000000101010100000111;
assign LUT_1[30944] = 32'b00000000000000001000001100001011;
assign LUT_1[30945] = 32'b00000000000000000001011110000111;
assign LUT_1[30946] = 32'b00000000000000000011111010011100;
assign LUT_1[30947] = 32'b11111111111111111101001100011000;
assign LUT_1[30948] = 32'b00000000000000010000000101100010;
assign LUT_1[30949] = 32'b00000000000000001001010111011110;
assign LUT_1[30950] = 32'b00000000000000001011110011110011;
assign LUT_1[30951] = 32'b00000000000000000101000101101111;
assign LUT_1[30952] = 32'b00000000000000000111011010000000;
assign LUT_1[30953] = 32'b00000000000000000000101011111100;
assign LUT_1[30954] = 32'b00000000000000000011001000010001;
assign LUT_1[30955] = 32'b11111111111111111100011010001101;
assign LUT_1[30956] = 32'b00000000000000001111010011010111;
assign LUT_1[30957] = 32'b00000000000000001000100101010011;
assign LUT_1[30958] = 32'b00000000000000001011000001101000;
assign LUT_1[30959] = 32'b00000000000000000100010011100100;
assign LUT_1[30960] = 32'b00000000000000001010000111101101;
assign LUT_1[30961] = 32'b00000000000000000011011001101001;
assign LUT_1[30962] = 32'b00000000000000000101110101111110;
assign LUT_1[30963] = 32'b11111111111111111111000111111010;
assign LUT_1[30964] = 32'b00000000000000010010000001000100;
assign LUT_1[30965] = 32'b00000000000000001011010011000000;
assign LUT_1[30966] = 32'b00000000000000001101101111010101;
assign LUT_1[30967] = 32'b00000000000000000111000001010001;
assign LUT_1[30968] = 32'b00000000000000001001010101100010;
assign LUT_1[30969] = 32'b00000000000000000010100111011110;
assign LUT_1[30970] = 32'b00000000000000000101000011110011;
assign LUT_1[30971] = 32'b11111111111111111110010101101111;
assign LUT_1[30972] = 32'b00000000000000010001001110111001;
assign LUT_1[30973] = 32'b00000000000000001010100000110101;
assign LUT_1[30974] = 32'b00000000000000001100111101001010;
assign LUT_1[30975] = 32'b00000000000000000110001111000110;
assign LUT_1[30976] = 32'b00000000000000000000000111101101;
assign LUT_1[30977] = 32'b11111111111111111001011001101001;
assign LUT_1[30978] = 32'b11111111111111111011110101111110;
assign LUT_1[30979] = 32'b11111111111111110101000111111010;
assign LUT_1[30980] = 32'b00000000000000001000000001000100;
assign LUT_1[30981] = 32'b00000000000000000001010011000000;
assign LUT_1[30982] = 32'b00000000000000000011101111010101;
assign LUT_1[30983] = 32'b11111111111111111101000001010001;
assign LUT_1[30984] = 32'b11111111111111111111010101100010;
assign LUT_1[30985] = 32'b11111111111111111000100111011110;
assign LUT_1[30986] = 32'b11111111111111111011000011110011;
assign LUT_1[30987] = 32'b11111111111111110100010101101111;
assign LUT_1[30988] = 32'b00000000000000000111001110111001;
assign LUT_1[30989] = 32'b00000000000000000000100000110101;
assign LUT_1[30990] = 32'b00000000000000000010111101001010;
assign LUT_1[30991] = 32'b11111111111111111100001111000110;
assign LUT_1[30992] = 32'b00000000000000000010000011001111;
assign LUT_1[30993] = 32'b11111111111111111011010101001011;
assign LUT_1[30994] = 32'b11111111111111111101110001100000;
assign LUT_1[30995] = 32'b11111111111111110111000011011100;
assign LUT_1[30996] = 32'b00000000000000001001111100100110;
assign LUT_1[30997] = 32'b00000000000000000011001110100010;
assign LUT_1[30998] = 32'b00000000000000000101101010110111;
assign LUT_1[30999] = 32'b11111111111111111110111100110011;
assign LUT_1[31000] = 32'b00000000000000000001010001000100;
assign LUT_1[31001] = 32'b11111111111111111010100011000000;
assign LUT_1[31002] = 32'b11111111111111111100111111010101;
assign LUT_1[31003] = 32'b11111111111111110110010001010001;
assign LUT_1[31004] = 32'b00000000000000001001001010011011;
assign LUT_1[31005] = 32'b00000000000000000010011100010111;
assign LUT_1[31006] = 32'b00000000000000000100111000101100;
assign LUT_1[31007] = 32'b11111111111111111110001010101000;
assign LUT_1[31008] = 32'b00000000000000000001000010101100;
assign LUT_1[31009] = 32'b11111111111111111010010100101000;
assign LUT_1[31010] = 32'b11111111111111111100110000111101;
assign LUT_1[31011] = 32'b11111111111111110110000010111001;
assign LUT_1[31012] = 32'b00000000000000001000111100000011;
assign LUT_1[31013] = 32'b00000000000000000010001101111111;
assign LUT_1[31014] = 32'b00000000000000000100101010010100;
assign LUT_1[31015] = 32'b11111111111111111101111100010000;
assign LUT_1[31016] = 32'b00000000000000000000010000100001;
assign LUT_1[31017] = 32'b11111111111111111001100010011101;
assign LUT_1[31018] = 32'b11111111111111111011111110110010;
assign LUT_1[31019] = 32'b11111111111111110101010000101110;
assign LUT_1[31020] = 32'b00000000000000001000001001111000;
assign LUT_1[31021] = 32'b00000000000000000001011011110100;
assign LUT_1[31022] = 32'b00000000000000000011111000001001;
assign LUT_1[31023] = 32'b11111111111111111101001010000101;
assign LUT_1[31024] = 32'b00000000000000000010111110001110;
assign LUT_1[31025] = 32'b11111111111111111100010000001010;
assign LUT_1[31026] = 32'b11111111111111111110101100011111;
assign LUT_1[31027] = 32'b11111111111111110111111110011011;
assign LUT_1[31028] = 32'b00000000000000001010110111100101;
assign LUT_1[31029] = 32'b00000000000000000100001001100001;
assign LUT_1[31030] = 32'b00000000000000000110100101110110;
assign LUT_1[31031] = 32'b11111111111111111111110111110010;
assign LUT_1[31032] = 32'b00000000000000000010001100000011;
assign LUT_1[31033] = 32'b11111111111111111011011101111111;
assign LUT_1[31034] = 32'b11111111111111111101111010010100;
assign LUT_1[31035] = 32'b11111111111111110111001100010000;
assign LUT_1[31036] = 32'b00000000000000001010000101011010;
assign LUT_1[31037] = 32'b00000000000000000011010111010110;
assign LUT_1[31038] = 32'b00000000000000000101110011101011;
assign LUT_1[31039] = 32'b11111111111111111111000101100111;
assign LUT_1[31040] = 32'b00000000000000000010000101010101;
assign LUT_1[31041] = 32'b11111111111111111011010111010001;
assign LUT_1[31042] = 32'b11111111111111111101110011100110;
assign LUT_1[31043] = 32'b11111111111111110111000101100010;
assign LUT_1[31044] = 32'b00000000000000001001111110101100;
assign LUT_1[31045] = 32'b00000000000000000011010000101000;
assign LUT_1[31046] = 32'b00000000000000000101101100111101;
assign LUT_1[31047] = 32'b11111111111111111110111110111001;
assign LUT_1[31048] = 32'b00000000000000000001010011001010;
assign LUT_1[31049] = 32'b11111111111111111010100101000110;
assign LUT_1[31050] = 32'b11111111111111111101000001011011;
assign LUT_1[31051] = 32'b11111111111111110110010011010111;
assign LUT_1[31052] = 32'b00000000000000001001001100100001;
assign LUT_1[31053] = 32'b00000000000000000010011110011101;
assign LUT_1[31054] = 32'b00000000000000000100111010110010;
assign LUT_1[31055] = 32'b11111111111111111110001100101110;
assign LUT_1[31056] = 32'b00000000000000000100000000110111;
assign LUT_1[31057] = 32'b11111111111111111101010010110011;
assign LUT_1[31058] = 32'b11111111111111111111101111001000;
assign LUT_1[31059] = 32'b11111111111111111001000001000100;
assign LUT_1[31060] = 32'b00000000000000001011111010001110;
assign LUT_1[31061] = 32'b00000000000000000101001100001010;
assign LUT_1[31062] = 32'b00000000000000000111101000011111;
assign LUT_1[31063] = 32'b00000000000000000000111010011011;
assign LUT_1[31064] = 32'b00000000000000000011001110101100;
assign LUT_1[31065] = 32'b11111111111111111100100000101000;
assign LUT_1[31066] = 32'b11111111111111111110111100111101;
assign LUT_1[31067] = 32'b11111111111111111000001110111001;
assign LUT_1[31068] = 32'b00000000000000001011001000000011;
assign LUT_1[31069] = 32'b00000000000000000100011001111111;
assign LUT_1[31070] = 32'b00000000000000000110110110010100;
assign LUT_1[31071] = 32'b00000000000000000000001000010000;
assign LUT_1[31072] = 32'b00000000000000000011000000010100;
assign LUT_1[31073] = 32'b11111111111111111100010010010000;
assign LUT_1[31074] = 32'b11111111111111111110101110100101;
assign LUT_1[31075] = 32'b11111111111111111000000000100001;
assign LUT_1[31076] = 32'b00000000000000001010111001101011;
assign LUT_1[31077] = 32'b00000000000000000100001011100111;
assign LUT_1[31078] = 32'b00000000000000000110100111111100;
assign LUT_1[31079] = 32'b11111111111111111111111001111000;
assign LUT_1[31080] = 32'b00000000000000000010001110001001;
assign LUT_1[31081] = 32'b11111111111111111011100000000101;
assign LUT_1[31082] = 32'b11111111111111111101111100011010;
assign LUT_1[31083] = 32'b11111111111111110111001110010110;
assign LUT_1[31084] = 32'b00000000000000001010000111100000;
assign LUT_1[31085] = 32'b00000000000000000011011001011100;
assign LUT_1[31086] = 32'b00000000000000000101110101110001;
assign LUT_1[31087] = 32'b11111111111111111111000111101101;
assign LUT_1[31088] = 32'b00000000000000000100111011110110;
assign LUT_1[31089] = 32'b11111111111111111110001101110010;
assign LUT_1[31090] = 32'b00000000000000000000101010000111;
assign LUT_1[31091] = 32'b11111111111111111001111100000011;
assign LUT_1[31092] = 32'b00000000000000001100110101001101;
assign LUT_1[31093] = 32'b00000000000000000110000111001001;
assign LUT_1[31094] = 32'b00000000000000001000100011011110;
assign LUT_1[31095] = 32'b00000000000000000001110101011010;
assign LUT_1[31096] = 32'b00000000000000000100001001101011;
assign LUT_1[31097] = 32'b11111111111111111101011011100111;
assign LUT_1[31098] = 32'b11111111111111111111110111111100;
assign LUT_1[31099] = 32'b11111111111111111001001001111000;
assign LUT_1[31100] = 32'b00000000000000001100000011000010;
assign LUT_1[31101] = 32'b00000000000000000101010100111110;
assign LUT_1[31102] = 32'b00000000000000000111110001010011;
assign LUT_1[31103] = 32'b00000000000000000001000011001111;
assign LUT_1[31104] = 32'b00000000000000000011000111110000;
assign LUT_1[31105] = 32'b11111111111111111100011001101100;
assign LUT_1[31106] = 32'b11111111111111111110110110000001;
assign LUT_1[31107] = 32'b11111111111111111000000111111101;
assign LUT_1[31108] = 32'b00000000000000001011000001000111;
assign LUT_1[31109] = 32'b00000000000000000100010011000011;
assign LUT_1[31110] = 32'b00000000000000000110101111011000;
assign LUT_1[31111] = 32'b00000000000000000000000001010100;
assign LUT_1[31112] = 32'b00000000000000000010010101100101;
assign LUT_1[31113] = 32'b11111111111111111011100111100001;
assign LUT_1[31114] = 32'b11111111111111111110000011110110;
assign LUT_1[31115] = 32'b11111111111111110111010101110010;
assign LUT_1[31116] = 32'b00000000000000001010001110111100;
assign LUT_1[31117] = 32'b00000000000000000011100000111000;
assign LUT_1[31118] = 32'b00000000000000000101111101001101;
assign LUT_1[31119] = 32'b11111111111111111111001111001001;
assign LUT_1[31120] = 32'b00000000000000000101000011010010;
assign LUT_1[31121] = 32'b11111111111111111110010101001110;
assign LUT_1[31122] = 32'b00000000000000000000110001100011;
assign LUT_1[31123] = 32'b11111111111111111010000011011111;
assign LUT_1[31124] = 32'b00000000000000001100111100101001;
assign LUT_1[31125] = 32'b00000000000000000110001110100101;
assign LUT_1[31126] = 32'b00000000000000001000101010111010;
assign LUT_1[31127] = 32'b00000000000000000001111100110110;
assign LUT_1[31128] = 32'b00000000000000000100010001000111;
assign LUT_1[31129] = 32'b11111111111111111101100011000011;
assign LUT_1[31130] = 32'b11111111111111111111111111011000;
assign LUT_1[31131] = 32'b11111111111111111001010001010100;
assign LUT_1[31132] = 32'b00000000000000001100001010011110;
assign LUT_1[31133] = 32'b00000000000000000101011100011010;
assign LUT_1[31134] = 32'b00000000000000000111111000101111;
assign LUT_1[31135] = 32'b00000000000000000001001010101011;
assign LUT_1[31136] = 32'b00000000000000000100000010101111;
assign LUT_1[31137] = 32'b11111111111111111101010100101011;
assign LUT_1[31138] = 32'b11111111111111111111110001000000;
assign LUT_1[31139] = 32'b11111111111111111001000010111100;
assign LUT_1[31140] = 32'b00000000000000001011111100000110;
assign LUT_1[31141] = 32'b00000000000000000101001110000010;
assign LUT_1[31142] = 32'b00000000000000000111101010010111;
assign LUT_1[31143] = 32'b00000000000000000000111100010011;
assign LUT_1[31144] = 32'b00000000000000000011010000100100;
assign LUT_1[31145] = 32'b11111111111111111100100010100000;
assign LUT_1[31146] = 32'b11111111111111111110111110110101;
assign LUT_1[31147] = 32'b11111111111111111000010000110001;
assign LUT_1[31148] = 32'b00000000000000001011001001111011;
assign LUT_1[31149] = 32'b00000000000000000100011011110111;
assign LUT_1[31150] = 32'b00000000000000000110111000001100;
assign LUT_1[31151] = 32'b00000000000000000000001010001000;
assign LUT_1[31152] = 32'b00000000000000000101111110010001;
assign LUT_1[31153] = 32'b11111111111111111111010000001101;
assign LUT_1[31154] = 32'b00000000000000000001101100100010;
assign LUT_1[31155] = 32'b11111111111111111010111110011110;
assign LUT_1[31156] = 32'b00000000000000001101110111101000;
assign LUT_1[31157] = 32'b00000000000000000111001001100100;
assign LUT_1[31158] = 32'b00000000000000001001100101111001;
assign LUT_1[31159] = 32'b00000000000000000010110111110101;
assign LUT_1[31160] = 32'b00000000000000000101001100000110;
assign LUT_1[31161] = 32'b11111111111111111110011110000010;
assign LUT_1[31162] = 32'b00000000000000000000111010010111;
assign LUT_1[31163] = 32'b11111111111111111010001100010011;
assign LUT_1[31164] = 32'b00000000000000001101000101011101;
assign LUT_1[31165] = 32'b00000000000000000110010111011001;
assign LUT_1[31166] = 32'b00000000000000001000110011101110;
assign LUT_1[31167] = 32'b00000000000000000010000101101010;
assign LUT_1[31168] = 32'b00000000000000000101000101011000;
assign LUT_1[31169] = 32'b11111111111111111110010111010100;
assign LUT_1[31170] = 32'b00000000000000000000110011101001;
assign LUT_1[31171] = 32'b11111111111111111010000101100101;
assign LUT_1[31172] = 32'b00000000000000001100111110101111;
assign LUT_1[31173] = 32'b00000000000000000110010000101011;
assign LUT_1[31174] = 32'b00000000000000001000101101000000;
assign LUT_1[31175] = 32'b00000000000000000001111110111100;
assign LUT_1[31176] = 32'b00000000000000000100010011001101;
assign LUT_1[31177] = 32'b11111111111111111101100101001001;
assign LUT_1[31178] = 32'b00000000000000000000000001011110;
assign LUT_1[31179] = 32'b11111111111111111001010011011010;
assign LUT_1[31180] = 32'b00000000000000001100001100100100;
assign LUT_1[31181] = 32'b00000000000000000101011110100000;
assign LUT_1[31182] = 32'b00000000000000000111111010110101;
assign LUT_1[31183] = 32'b00000000000000000001001100110001;
assign LUT_1[31184] = 32'b00000000000000000111000000111010;
assign LUT_1[31185] = 32'b00000000000000000000010010110110;
assign LUT_1[31186] = 32'b00000000000000000010101111001011;
assign LUT_1[31187] = 32'b11111111111111111100000001000111;
assign LUT_1[31188] = 32'b00000000000000001110111010010001;
assign LUT_1[31189] = 32'b00000000000000001000001100001101;
assign LUT_1[31190] = 32'b00000000000000001010101000100010;
assign LUT_1[31191] = 32'b00000000000000000011111010011110;
assign LUT_1[31192] = 32'b00000000000000000110001110101111;
assign LUT_1[31193] = 32'b11111111111111111111100000101011;
assign LUT_1[31194] = 32'b00000000000000000001111101000000;
assign LUT_1[31195] = 32'b11111111111111111011001110111100;
assign LUT_1[31196] = 32'b00000000000000001110001000000110;
assign LUT_1[31197] = 32'b00000000000000000111011010000010;
assign LUT_1[31198] = 32'b00000000000000001001110110010111;
assign LUT_1[31199] = 32'b00000000000000000011001000010011;
assign LUT_1[31200] = 32'b00000000000000000110000000010111;
assign LUT_1[31201] = 32'b11111111111111111111010010010011;
assign LUT_1[31202] = 32'b00000000000000000001101110101000;
assign LUT_1[31203] = 32'b11111111111111111011000000100100;
assign LUT_1[31204] = 32'b00000000000000001101111001101110;
assign LUT_1[31205] = 32'b00000000000000000111001011101010;
assign LUT_1[31206] = 32'b00000000000000001001100111111111;
assign LUT_1[31207] = 32'b00000000000000000010111001111011;
assign LUT_1[31208] = 32'b00000000000000000101001110001100;
assign LUT_1[31209] = 32'b11111111111111111110100000001000;
assign LUT_1[31210] = 32'b00000000000000000000111100011101;
assign LUT_1[31211] = 32'b11111111111111111010001110011001;
assign LUT_1[31212] = 32'b00000000000000001101000111100011;
assign LUT_1[31213] = 32'b00000000000000000110011001011111;
assign LUT_1[31214] = 32'b00000000000000001000110101110100;
assign LUT_1[31215] = 32'b00000000000000000010000111110000;
assign LUT_1[31216] = 32'b00000000000000000111111011111001;
assign LUT_1[31217] = 32'b00000000000000000001001101110101;
assign LUT_1[31218] = 32'b00000000000000000011101010001010;
assign LUT_1[31219] = 32'b11111111111111111100111100000110;
assign LUT_1[31220] = 32'b00000000000000001111110101010000;
assign LUT_1[31221] = 32'b00000000000000001001000111001100;
assign LUT_1[31222] = 32'b00000000000000001011100011100001;
assign LUT_1[31223] = 32'b00000000000000000100110101011101;
assign LUT_1[31224] = 32'b00000000000000000111001001101110;
assign LUT_1[31225] = 32'b00000000000000000000011011101010;
assign LUT_1[31226] = 32'b00000000000000000010110111111111;
assign LUT_1[31227] = 32'b11111111111111111100001001111011;
assign LUT_1[31228] = 32'b00000000000000001111000011000101;
assign LUT_1[31229] = 32'b00000000000000001000010101000001;
assign LUT_1[31230] = 32'b00000000000000001010110001010110;
assign LUT_1[31231] = 32'b00000000000000000100000011010010;
assign LUT_1[31232] = 32'b11111111111111111100000001111110;
assign LUT_1[31233] = 32'b11111111111111110101010011111010;
assign LUT_1[31234] = 32'b11111111111111110111110000001111;
assign LUT_1[31235] = 32'b11111111111111110001000010001011;
assign LUT_1[31236] = 32'b00000000000000000011111011010101;
assign LUT_1[31237] = 32'b11111111111111111101001101010001;
assign LUT_1[31238] = 32'b11111111111111111111101001100110;
assign LUT_1[31239] = 32'b11111111111111111000111011100010;
assign LUT_1[31240] = 32'b11111111111111111011001111110011;
assign LUT_1[31241] = 32'b11111111111111110100100001101111;
assign LUT_1[31242] = 32'b11111111111111110110111110000100;
assign LUT_1[31243] = 32'b11111111111111110000010000000000;
assign LUT_1[31244] = 32'b00000000000000000011001001001010;
assign LUT_1[31245] = 32'b11111111111111111100011011000110;
assign LUT_1[31246] = 32'b11111111111111111110110111011011;
assign LUT_1[31247] = 32'b11111111111111111000001001010111;
assign LUT_1[31248] = 32'b11111111111111111101111101100000;
assign LUT_1[31249] = 32'b11111111111111110111001111011100;
assign LUT_1[31250] = 32'b11111111111111111001101011110001;
assign LUT_1[31251] = 32'b11111111111111110010111101101101;
assign LUT_1[31252] = 32'b00000000000000000101110110110111;
assign LUT_1[31253] = 32'b11111111111111111111001000110011;
assign LUT_1[31254] = 32'b00000000000000000001100101001000;
assign LUT_1[31255] = 32'b11111111111111111010110111000100;
assign LUT_1[31256] = 32'b11111111111111111101001011010101;
assign LUT_1[31257] = 32'b11111111111111110110011101010001;
assign LUT_1[31258] = 32'b11111111111111111000111001100110;
assign LUT_1[31259] = 32'b11111111111111110010001011100010;
assign LUT_1[31260] = 32'b00000000000000000101000100101100;
assign LUT_1[31261] = 32'b11111111111111111110010110101000;
assign LUT_1[31262] = 32'b00000000000000000000110010111101;
assign LUT_1[31263] = 32'b11111111111111111010000100111001;
assign LUT_1[31264] = 32'b11111111111111111100111100111101;
assign LUT_1[31265] = 32'b11111111111111110110001110111001;
assign LUT_1[31266] = 32'b11111111111111111000101011001110;
assign LUT_1[31267] = 32'b11111111111111110001111101001010;
assign LUT_1[31268] = 32'b00000000000000000100110110010100;
assign LUT_1[31269] = 32'b11111111111111111110001000010000;
assign LUT_1[31270] = 32'b00000000000000000000100100100101;
assign LUT_1[31271] = 32'b11111111111111111001110110100001;
assign LUT_1[31272] = 32'b11111111111111111100001010110010;
assign LUT_1[31273] = 32'b11111111111111110101011100101110;
assign LUT_1[31274] = 32'b11111111111111110111111001000011;
assign LUT_1[31275] = 32'b11111111111111110001001010111111;
assign LUT_1[31276] = 32'b00000000000000000100000100001001;
assign LUT_1[31277] = 32'b11111111111111111101010110000101;
assign LUT_1[31278] = 32'b11111111111111111111110010011010;
assign LUT_1[31279] = 32'b11111111111111111001000100010110;
assign LUT_1[31280] = 32'b11111111111111111110111000011111;
assign LUT_1[31281] = 32'b11111111111111111000001010011011;
assign LUT_1[31282] = 32'b11111111111111111010100110110000;
assign LUT_1[31283] = 32'b11111111111111110011111000101100;
assign LUT_1[31284] = 32'b00000000000000000110110001110110;
assign LUT_1[31285] = 32'b00000000000000000000000011110010;
assign LUT_1[31286] = 32'b00000000000000000010100000000111;
assign LUT_1[31287] = 32'b11111111111111111011110010000011;
assign LUT_1[31288] = 32'b11111111111111111110000110010100;
assign LUT_1[31289] = 32'b11111111111111110111011000010000;
assign LUT_1[31290] = 32'b11111111111111111001110100100101;
assign LUT_1[31291] = 32'b11111111111111110011000110100001;
assign LUT_1[31292] = 32'b00000000000000000101111111101011;
assign LUT_1[31293] = 32'b11111111111111111111010001100111;
assign LUT_1[31294] = 32'b00000000000000000001101101111100;
assign LUT_1[31295] = 32'b11111111111111111010111111111000;
assign LUT_1[31296] = 32'b11111111111111111101111111100110;
assign LUT_1[31297] = 32'b11111111111111110111010001100010;
assign LUT_1[31298] = 32'b11111111111111111001101101110111;
assign LUT_1[31299] = 32'b11111111111111110010111111110011;
assign LUT_1[31300] = 32'b00000000000000000101111000111101;
assign LUT_1[31301] = 32'b11111111111111111111001010111001;
assign LUT_1[31302] = 32'b00000000000000000001100111001110;
assign LUT_1[31303] = 32'b11111111111111111010111001001010;
assign LUT_1[31304] = 32'b11111111111111111101001101011011;
assign LUT_1[31305] = 32'b11111111111111110110011111010111;
assign LUT_1[31306] = 32'b11111111111111111000111011101100;
assign LUT_1[31307] = 32'b11111111111111110010001101101000;
assign LUT_1[31308] = 32'b00000000000000000101000110110010;
assign LUT_1[31309] = 32'b11111111111111111110011000101110;
assign LUT_1[31310] = 32'b00000000000000000000110101000011;
assign LUT_1[31311] = 32'b11111111111111111010000110111111;
assign LUT_1[31312] = 32'b11111111111111111111111011001000;
assign LUT_1[31313] = 32'b11111111111111111001001101000100;
assign LUT_1[31314] = 32'b11111111111111111011101001011001;
assign LUT_1[31315] = 32'b11111111111111110100111011010101;
assign LUT_1[31316] = 32'b00000000000000000111110100011111;
assign LUT_1[31317] = 32'b00000000000000000001000110011011;
assign LUT_1[31318] = 32'b00000000000000000011100010110000;
assign LUT_1[31319] = 32'b11111111111111111100110100101100;
assign LUT_1[31320] = 32'b11111111111111111111001000111101;
assign LUT_1[31321] = 32'b11111111111111111000011010111001;
assign LUT_1[31322] = 32'b11111111111111111010110111001110;
assign LUT_1[31323] = 32'b11111111111111110100001001001010;
assign LUT_1[31324] = 32'b00000000000000000111000010010100;
assign LUT_1[31325] = 32'b00000000000000000000010100010000;
assign LUT_1[31326] = 32'b00000000000000000010110000100101;
assign LUT_1[31327] = 32'b11111111111111111100000010100001;
assign LUT_1[31328] = 32'b11111111111111111110111010100101;
assign LUT_1[31329] = 32'b11111111111111111000001100100001;
assign LUT_1[31330] = 32'b11111111111111111010101000110110;
assign LUT_1[31331] = 32'b11111111111111110011111010110010;
assign LUT_1[31332] = 32'b00000000000000000110110011111100;
assign LUT_1[31333] = 32'b00000000000000000000000101111000;
assign LUT_1[31334] = 32'b00000000000000000010100010001101;
assign LUT_1[31335] = 32'b11111111111111111011110100001001;
assign LUT_1[31336] = 32'b11111111111111111110001000011010;
assign LUT_1[31337] = 32'b11111111111111110111011010010110;
assign LUT_1[31338] = 32'b11111111111111111001110110101011;
assign LUT_1[31339] = 32'b11111111111111110011001000100111;
assign LUT_1[31340] = 32'b00000000000000000110000001110001;
assign LUT_1[31341] = 32'b11111111111111111111010011101101;
assign LUT_1[31342] = 32'b00000000000000000001110000000010;
assign LUT_1[31343] = 32'b11111111111111111011000001111110;
assign LUT_1[31344] = 32'b00000000000000000000110110000111;
assign LUT_1[31345] = 32'b11111111111111111010001000000011;
assign LUT_1[31346] = 32'b11111111111111111100100100011000;
assign LUT_1[31347] = 32'b11111111111111110101110110010100;
assign LUT_1[31348] = 32'b00000000000000001000101111011110;
assign LUT_1[31349] = 32'b00000000000000000010000001011010;
assign LUT_1[31350] = 32'b00000000000000000100011101101111;
assign LUT_1[31351] = 32'b11111111111111111101101111101011;
assign LUT_1[31352] = 32'b00000000000000000000000011111100;
assign LUT_1[31353] = 32'b11111111111111111001010101111000;
assign LUT_1[31354] = 32'b11111111111111111011110010001101;
assign LUT_1[31355] = 32'b11111111111111110101000100001001;
assign LUT_1[31356] = 32'b00000000000000000111111101010011;
assign LUT_1[31357] = 32'b00000000000000000001001111001111;
assign LUT_1[31358] = 32'b00000000000000000011101011100100;
assign LUT_1[31359] = 32'b11111111111111111100111101100000;
assign LUT_1[31360] = 32'b11111111111111111111000010000001;
assign LUT_1[31361] = 32'b11111111111111111000010011111101;
assign LUT_1[31362] = 32'b11111111111111111010110000010010;
assign LUT_1[31363] = 32'b11111111111111110100000010001110;
assign LUT_1[31364] = 32'b00000000000000000110111011011000;
assign LUT_1[31365] = 32'b00000000000000000000001101010100;
assign LUT_1[31366] = 32'b00000000000000000010101001101001;
assign LUT_1[31367] = 32'b11111111111111111011111011100101;
assign LUT_1[31368] = 32'b11111111111111111110001111110110;
assign LUT_1[31369] = 32'b11111111111111110111100001110010;
assign LUT_1[31370] = 32'b11111111111111111001111110000111;
assign LUT_1[31371] = 32'b11111111111111110011010000000011;
assign LUT_1[31372] = 32'b00000000000000000110001001001101;
assign LUT_1[31373] = 32'b11111111111111111111011011001001;
assign LUT_1[31374] = 32'b00000000000000000001110111011110;
assign LUT_1[31375] = 32'b11111111111111111011001001011010;
assign LUT_1[31376] = 32'b00000000000000000000111101100011;
assign LUT_1[31377] = 32'b11111111111111111010001111011111;
assign LUT_1[31378] = 32'b11111111111111111100101011110100;
assign LUT_1[31379] = 32'b11111111111111110101111101110000;
assign LUT_1[31380] = 32'b00000000000000001000110110111010;
assign LUT_1[31381] = 32'b00000000000000000010001000110110;
assign LUT_1[31382] = 32'b00000000000000000100100101001011;
assign LUT_1[31383] = 32'b11111111111111111101110111000111;
assign LUT_1[31384] = 32'b00000000000000000000001011011000;
assign LUT_1[31385] = 32'b11111111111111111001011101010100;
assign LUT_1[31386] = 32'b11111111111111111011111001101001;
assign LUT_1[31387] = 32'b11111111111111110101001011100101;
assign LUT_1[31388] = 32'b00000000000000001000000100101111;
assign LUT_1[31389] = 32'b00000000000000000001010110101011;
assign LUT_1[31390] = 32'b00000000000000000011110011000000;
assign LUT_1[31391] = 32'b11111111111111111101000100111100;
assign LUT_1[31392] = 32'b11111111111111111111111101000000;
assign LUT_1[31393] = 32'b11111111111111111001001110111100;
assign LUT_1[31394] = 32'b11111111111111111011101011010001;
assign LUT_1[31395] = 32'b11111111111111110100111101001101;
assign LUT_1[31396] = 32'b00000000000000000111110110010111;
assign LUT_1[31397] = 32'b00000000000000000001001000010011;
assign LUT_1[31398] = 32'b00000000000000000011100100101000;
assign LUT_1[31399] = 32'b11111111111111111100110110100100;
assign LUT_1[31400] = 32'b11111111111111111111001010110101;
assign LUT_1[31401] = 32'b11111111111111111000011100110001;
assign LUT_1[31402] = 32'b11111111111111111010111001000110;
assign LUT_1[31403] = 32'b11111111111111110100001011000010;
assign LUT_1[31404] = 32'b00000000000000000111000100001100;
assign LUT_1[31405] = 32'b00000000000000000000010110001000;
assign LUT_1[31406] = 32'b00000000000000000010110010011101;
assign LUT_1[31407] = 32'b11111111111111111100000100011001;
assign LUT_1[31408] = 32'b00000000000000000001111000100010;
assign LUT_1[31409] = 32'b11111111111111111011001010011110;
assign LUT_1[31410] = 32'b11111111111111111101100110110011;
assign LUT_1[31411] = 32'b11111111111111110110111000101111;
assign LUT_1[31412] = 32'b00000000000000001001110001111001;
assign LUT_1[31413] = 32'b00000000000000000011000011110101;
assign LUT_1[31414] = 32'b00000000000000000101100000001010;
assign LUT_1[31415] = 32'b11111111111111111110110010000110;
assign LUT_1[31416] = 32'b00000000000000000001000110010111;
assign LUT_1[31417] = 32'b11111111111111111010011000010011;
assign LUT_1[31418] = 32'b11111111111111111100110100101000;
assign LUT_1[31419] = 32'b11111111111111110110000110100100;
assign LUT_1[31420] = 32'b00000000000000001000111111101110;
assign LUT_1[31421] = 32'b00000000000000000010010001101010;
assign LUT_1[31422] = 32'b00000000000000000100101101111111;
assign LUT_1[31423] = 32'b11111111111111111101111111111011;
assign LUT_1[31424] = 32'b00000000000000000000111111101001;
assign LUT_1[31425] = 32'b11111111111111111010010001100101;
assign LUT_1[31426] = 32'b11111111111111111100101101111010;
assign LUT_1[31427] = 32'b11111111111111110101111111110110;
assign LUT_1[31428] = 32'b00000000000000001000111001000000;
assign LUT_1[31429] = 32'b00000000000000000010001010111100;
assign LUT_1[31430] = 32'b00000000000000000100100111010001;
assign LUT_1[31431] = 32'b11111111111111111101111001001101;
assign LUT_1[31432] = 32'b00000000000000000000001101011110;
assign LUT_1[31433] = 32'b11111111111111111001011111011010;
assign LUT_1[31434] = 32'b11111111111111111011111011101111;
assign LUT_1[31435] = 32'b11111111111111110101001101101011;
assign LUT_1[31436] = 32'b00000000000000001000000110110101;
assign LUT_1[31437] = 32'b00000000000000000001011000110001;
assign LUT_1[31438] = 32'b00000000000000000011110101000110;
assign LUT_1[31439] = 32'b11111111111111111101000111000010;
assign LUT_1[31440] = 32'b00000000000000000010111011001011;
assign LUT_1[31441] = 32'b11111111111111111100001101000111;
assign LUT_1[31442] = 32'b11111111111111111110101001011100;
assign LUT_1[31443] = 32'b11111111111111110111111011011000;
assign LUT_1[31444] = 32'b00000000000000001010110100100010;
assign LUT_1[31445] = 32'b00000000000000000100000110011110;
assign LUT_1[31446] = 32'b00000000000000000110100010110011;
assign LUT_1[31447] = 32'b11111111111111111111110100101111;
assign LUT_1[31448] = 32'b00000000000000000010001001000000;
assign LUT_1[31449] = 32'b11111111111111111011011010111100;
assign LUT_1[31450] = 32'b11111111111111111101110111010001;
assign LUT_1[31451] = 32'b11111111111111110111001001001101;
assign LUT_1[31452] = 32'b00000000000000001010000010010111;
assign LUT_1[31453] = 32'b00000000000000000011010100010011;
assign LUT_1[31454] = 32'b00000000000000000101110000101000;
assign LUT_1[31455] = 32'b11111111111111111111000010100100;
assign LUT_1[31456] = 32'b00000000000000000001111010101000;
assign LUT_1[31457] = 32'b11111111111111111011001100100100;
assign LUT_1[31458] = 32'b11111111111111111101101000111001;
assign LUT_1[31459] = 32'b11111111111111110110111010110101;
assign LUT_1[31460] = 32'b00000000000000001001110011111111;
assign LUT_1[31461] = 32'b00000000000000000011000101111011;
assign LUT_1[31462] = 32'b00000000000000000101100010010000;
assign LUT_1[31463] = 32'b11111111111111111110110100001100;
assign LUT_1[31464] = 32'b00000000000000000001001000011101;
assign LUT_1[31465] = 32'b11111111111111111010011010011001;
assign LUT_1[31466] = 32'b11111111111111111100110110101110;
assign LUT_1[31467] = 32'b11111111111111110110001000101010;
assign LUT_1[31468] = 32'b00000000000000001001000001110100;
assign LUT_1[31469] = 32'b00000000000000000010010011110000;
assign LUT_1[31470] = 32'b00000000000000000100110000000101;
assign LUT_1[31471] = 32'b11111111111111111110000010000001;
assign LUT_1[31472] = 32'b00000000000000000011110110001010;
assign LUT_1[31473] = 32'b11111111111111111101001000000110;
assign LUT_1[31474] = 32'b11111111111111111111100100011011;
assign LUT_1[31475] = 32'b11111111111111111000110110010111;
assign LUT_1[31476] = 32'b00000000000000001011101111100001;
assign LUT_1[31477] = 32'b00000000000000000101000001011101;
assign LUT_1[31478] = 32'b00000000000000000111011101110010;
assign LUT_1[31479] = 32'b00000000000000000000101111101110;
assign LUT_1[31480] = 32'b00000000000000000011000011111111;
assign LUT_1[31481] = 32'b11111111111111111100010101111011;
assign LUT_1[31482] = 32'b11111111111111111110110010010000;
assign LUT_1[31483] = 32'b11111111111111111000000100001100;
assign LUT_1[31484] = 32'b00000000000000001010111101010110;
assign LUT_1[31485] = 32'b00000000000000000100001111010010;
assign LUT_1[31486] = 32'b00000000000000000110101011100111;
assign LUT_1[31487] = 32'b11111111111111111111111101100011;
assign LUT_1[31488] = 32'b11111111111111111001110110001010;
assign LUT_1[31489] = 32'b11111111111111110011001000000110;
assign LUT_1[31490] = 32'b11111111111111110101100100011011;
assign LUT_1[31491] = 32'b11111111111111101110110110010111;
assign LUT_1[31492] = 32'b00000000000000000001101111100001;
assign LUT_1[31493] = 32'b11111111111111111011000001011101;
assign LUT_1[31494] = 32'b11111111111111111101011101110010;
assign LUT_1[31495] = 32'b11111111111111110110101111101110;
assign LUT_1[31496] = 32'b11111111111111111001000011111111;
assign LUT_1[31497] = 32'b11111111111111110010010101111011;
assign LUT_1[31498] = 32'b11111111111111110100110010010000;
assign LUT_1[31499] = 32'b11111111111111101110000100001100;
assign LUT_1[31500] = 32'b00000000000000000000111101010110;
assign LUT_1[31501] = 32'b11111111111111111010001111010010;
assign LUT_1[31502] = 32'b11111111111111111100101011100111;
assign LUT_1[31503] = 32'b11111111111111110101111101100011;
assign LUT_1[31504] = 32'b11111111111111111011110001101100;
assign LUT_1[31505] = 32'b11111111111111110101000011101000;
assign LUT_1[31506] = 32'b11111111111111110111011111111101;
assign LUT_1[31507] = 32'b11111111111111110000110001111001;
assign LUT_1[31508] = 32'b00000000000000000011101011000011;
assign LUT_1[31509] = 32'b11111111111111111100111100111111;
assign LUT_1[31510] = 32'b11111111111111111111011001010100;
assign LUT_1[31511] = 32'b11111111111111111000101011010000;
assign LUT_1[31512] = 32'b11111111111111111010111111100001;
assign LUT_1[31513] = 32'b11111111111111110100010001011101;
assign LUT_1[31514] = 32'b11111111111111110110101101110010;
assign LUT_1[31515] = 32'b11111111111111101111111111101110;
assign LUT_1[31516] = 32'b00000000000000000010111000111000;
assign LUT_1[31517] = 32'b11111111111111111100001010110100;
assign LUT_1[31518] = 32'b11111111111111111110100111001001;
assign LUT_1[31519] = 32'b11111111111111110111111001000101;
assign LUT_1[31520] = 32'b11111111111111111010110001001001;
assign LUT_1[31521] = 32'b11111111111111110100000011000101;
assign LUT_1[31522] = 32'b11111111111111110110011111011010;
assign LUT_1[31523] = 32'b11111111111111101111110001010110;
assign LUT_1[31524] = 32'b00000000000000000010101010100000;
assign LUT_1[31525] = 32'b11111111111111111011111100011100;
assign LUT_1[31526] = 32'b11111111111111111110011000110001;
assign LUT_1[31527] = 32'b11111111111111110111101010101101;
assign LUT_1[31528] = 32'b11111111111111111001111110111110;
assign LUT_1[31529] = 32'b11111111111111110011010000111010;
assign LUT_1[31530] = 32'b11111111111111110101101101001111;
assign LUT_1[31531] = 32'b11111111111111101110111111001011;
assign LUT_1[31532] = 32'b00000000000000000001111000010101;
assign LUT_1[31533] = 32'b11111111111111111011001010010001;
assign LUT_1[31534] = 32'b11111111111111111101100110100110;
assign LUT_1[31535] = 32'b11111111111111110110111000100010;
assign LUT_1[31536] = 32'b11111111111111111100101100101011;
assign LUT_1[31537] = 32'b11111111111111110101111110100111;
assign LUT_1[31538] = 32'b11111111111111111000011010111100;
assign LUT_1[31539] = 32'b11111111111111110001101100111000;
assign LUT_1[31540] = 32'b00000000000000000100100110000010;
assign LUT_1[31541] = 32'b11111111111111111101110111111110;
assign LUT_1[31542] = 32'b00000000000000000000010100010011;
assign LUT_1[31543] = 32'b11111111111111111001100110001111;
assign LUT_1[31544] = 32'b11111111111111111011111010100000;
assign LUT_1[31545] = 32'b11111111111111110101001100011100;
assign LUT_1[31546] = 32'b11111111111111110111101000110001;
assign LUT_1[31547] = 32'b11111111111111110000111010101101;
assign LUT_1[31548] = 32'b00000000000000000011110011110111;
assign LUT_1[31549] = 32'b11111111111111111101000101110011;
assign LUT_1[31550] = 32'b11111111111111111111100010001000;
assign LUT_1[31551] = 32'b11111111111111111000110100000100;
assign LUT_1[31552] = 32'b11111111111111111011110011110010;
assign LUT_1[31553] = 32'b11111111111111110101000101101110;
assign LUT_1[31554] = 32'b11111111111111110111100010000011;
assign LUT_1[31555] = 32'b11111111111111110000110011111111;
assign LUT_1[31556] = 32'b00000000000000000011101101001001;
assign LUT_1[31557] = 32'b11111111111111111100111111000101;
assign LUT_1[31558] = 32'b11111111111111111111011011011010;
assign LUT_1[31559] = 32'b11111111111111111000101101010110;
assign LUT_1[31560] = 32'b11111111111111111011000001100111;
assign LUT_1[31561] = 32'b11111111111111110100010011100011;
assign LUT_1[31562] = 32'b11111111111111110110101111111000;
assign LUT_1[31563] = 32'b11111111111111110000000001110100;
assign LUT_1[31564] = 32'b00000000000000000010111010111110;
assign LUT_1[31565] = 32'b11111111111111111100001100111010;
assign LUT_1[31566] = 32'b11111111111111111110101001001111;
assign LUT_1[31567] = 32'b11111111111111110111111011001011;
assign LUT_1[31568] = 32'b11111111111111111101101111010100;
assign LUT_1[31569] = 32'b11111111111111110111000001010000;
assign LUT_1[31570] = 32'b11111111111111111001011101100101;
assign LUT_1[31571] = 32'b11111111111111110010101111100001;
assign LUT_1[31572] = 32'b00000000000000000101101000101011;
assign LUT_1[31573] = 32'b11111111111111111110111010100111;
assign LUT_1[31574] = 32'b00000000000000000001010110111100;
assign LUT_1[31575] = 32'b11111111111111111010101000111000;
assign LUT_1[31576] = 32'b11111111111111111100111101001001;
assign LUT_1[31577] = 32'b11111111111111110110001111000101;
assign LUT_1[31578] = 32'b11111111111111111000101011011010;
assign LUT_1[31579] = 32'b11111111111111110001111101010110;
assign LUT_1[31580] = 32'b00000000000000000100110110100000;
assign LUT_1[31581] = 32'b11111111111111111110001000011100;
assign LUT_1[31582] = 32'b00000000000000000000100100110001;
assign LUT_1[31583] = 32'b11111111111111111001110110101101;
assign LUT_1[31584] = 32'b11111111111111111100101110110001;
assign LUT_1[31585] = 32'b11111111111111110110000000101101;
assign LUT_1[31586] = 32'b11111111111111111000011101000010;
assign LUT_1[31587] = 32'b11111111111111110001101110111110;
assign LUT_1[31588] = 32'b00000000000000000100101000001000;
assign LUT_1[31589] = 32'b11111111111111111101111010000100;
assign LUT_1[31590] = 32'b00000000000000000000010110011001;
assign LUT_1[31591] = 32'b11111111111111111001101000010101;
assign LUT_1[31592] = 32'b11111111111111111011111100100110;
assign LUT_1[31593] = 32'b11111111111111110101001110100010;
assign LUT_1[31594] = 32'b11111111111111110111101010110111;
assign LUT_1[31595] = 32'b11111111111111110000111100110011;
assign LUT_1[31596] = 32'b00000000000000000011110101111101;
assign LUT_1[31597] = 32'b11111111111111111101000111111001;
assign LUT_1[31598] = 32'b11111111111111111111100100001110;
assign LUT_1[31599] = 32'b11111111111111111000110110001010;
assign LUT_1[31600] = 32'b11111111111111111110101010010011;
assign LUT_1[31601] = 32'b11111111111111110111111100001111;
assign LUT_1[31602] = 32'b11111111111111111010011000100100;
assign LUT_1[31603] = 32'b11111111111111110011101010100000;
assign LUT_1[31604] = 32'b00000000000000000110100011101010;
assign LUT_1[31605] = 32'b11111111111111111111110101100110;
assign LUT_1[31606] = 32'b00000000000000000010010001111011;
assign LUT_1[31607] = 32'b11111111111111111011100011110111;
assign LUT_1[31608] = 32'b11111111111111111101111000001000;
assign LUT_1[31609] = 32'b11111111111111110111001010000100;
assign LUT_1[31610] = 32'b11111111111111111001100110011001;
assign LUT_1[31611] = 32'b11111111111111110010111000010101;
assign LUT_1[31612] = 32'b00000000000000000101110001011111;
assign LUT_1[31613] = 32'b11111111111111111111000011011011;
assign LUT_1[31614] = 32'b00000000000000000001011111110000;
assign LUT_1[31615] = 32'b11111111111111111010110001101100;
assign LUT_1[31616] = 32'b11111111111111111100110110001101;
assign LUT_1[31617] = 32'b11111111111111110110001000001001;
assign LUT_1[31618] = 32'b11111111111111111000100100011110;
assign LUT_1[31619] = 32'b11111111111111110001110110011010;
assign LUT_1[31620] = 32'b00000000000000000100101111100100;
assign LUT_1[31621] = 32'b11111111111111111110000001100000;
assign LUT_1[31622] = 32'b00000000000000000000011101110101;
assign LUT_1[31623] = 32'b11111111111111111001101111110001;
assign LUT_1[31624] = 32'b11111111111111111100000100000010;
assign LUT_1[31625] = 32'b11111111111111110101010101111110;
assign LUT_1[31626] = 32'b11111111111111110111110010010011;
assign LUT_1[31627] = 32'b11111111111111110001000100001111;
assign LUT_1[31628] = 32'b00000000000000000011111101011001;
assign LUT_1[31629] = 32'b11111111111111111101001111010101;
assign LUT_1[31630] = 32'b11111111111111111111101011101010;
assign LUT_1[31631] = 32'b11111111111111111000111101100110;
assign LUT_1[31632] = 32'b11111111111111111110110001101111;
assign LUT_1[31633] = 32'b11111111111111111000000011101011;
assign LUT_1[31634] = 32'b11111111111111111010100000000000;
assign LUT_1[31635] = 32'b11111111111111110011110001111100;
assign LUT_1[31636] = 32'b00000000000000000110101011000110;
assign LUT_1[31637] = 32'b11111111111111111111111101000010;
assign LUT_1[31638] = 32'b00000000000000000010011001010111;
assign LUT_1[31639] = 32'b11111111111111111011101011010011;
assign LUT_1[31640] = 32'b11111111111111111101111111100100;
assign LUT_1[31641] = 32'b11111111111111110111010001100000;
assign LUT_1[31642] = 32'b11111111111111111001101101110101;
assign LUT_1[31643] = 32'b11111111111111110010111111110001;
assign LUT_1[31644] = 32'b00000000000000000101111000111011;
assign LUT_1[31645] = 32'b11111111111111111111001010110111;
assign LUT_1[31646] = 32'b00000000000000000001100111001100;
assign LUT_1[31647] = 32'b11111111111111111010111001001000;
assign LUT_1[31648] = 32'b11111111111111111101110001001100;
assign LUT_1[31649] = 32'b11111111111111110111000011001000;
assign LUT_1[31650] = 32'b11111111111111111001011111011101;
assign LUT_1[31651] = 32'b11111111111111110010110001011001;
assign LUT_1[31652] = 32'b00000000000000000101101010100011;
assign LUT_1[31653] = 32'b11111111111111111110111100011111;
assign LUT_1[31654] = 32'b00000000000000000001011000110100;
assign LUT_1[31655] = 32'b11111111111111111010101010110000;
assign LUT_1[31656] = 32'b11111111111111111100111111000001;
assign LUT_1[31657] = 32'b11111111111111110110010000111101;
assign LUT_1[31658] = 32'b11111111111111111000101101010010;
assign LUT_1[31659] = 32'b11111111111111110001111111001110;
assign LUT_1[31660] = 32'b00000000000000000100111000011000;
assign LUT_1[31661] = 32'b11111111111111111110001010010100;
assign LUT_1[31662] = 32'b00000000000000000000100110101001;
assign LUT_1[31663] = 32'b11111111111111111001111000100101;
assign LUT_1[31664] = 32'b11111111111111111111101100101110;
assign LUT_1[31665] = 32'b11111111111111111000111110101010;
assign LUT_1[31666] = 32'b11111111111111111011011010111111;
assign LUT_1[31667] = 32'b11111111111111110100101100111011;
assign LUT_1[31668] = 32'b00000000000000000111100110000101;
assign LUT_1[31669] = 32'b00000000000000000000111000000001;
assign LUT_1[31670] = 32'b00000000000000000011010100010110;
assign LUT_1[31671] = 32'b11111111111111111100100110010010;
assign LUT_1[31672] = 32'b11111111111111111110111010100011;
assign LUT_1[31673] = 32'b11111111111111111000001100011111;
assign LUT_1[31674] = 32'b11111111111111111010101000110100;
assign LUT_1[31675] = 32'b11111111111111110011111010110000;
assign LUT_1[31676] = 32'b00000000000000000110110011111010;
assign LUT_1[31677] = 32'b00000000000000000000000101110110;
assign LUT_1[31678] = 32'b00000000000000000010100010001011;
assign LUT_1[31679] = 32'b11111111111111111011110100000111;
assign LUT_1[31680] = 32'b11111111111111111110110011110101;
assign LUT_1[31681] = 32'b11111111111111111000000101110001;
assign LUT_1[31682] = 32'b11111111111111111010100010000110;
assign LUT_1[31683] = 32'b11111111111111110011110100000010;
assign LUT_1[31684] = 32'b00000000000000000110101101001100;
assign LUT_1[31685] = 32'b11111111111111111111111111001000;
assign LUT_1[31686] = 32'b00000000000000000010011011011101;
assign LUT_1[31687] = 32'b11111111111111111011101101011001;
assign LUT_1[31688] = 32'b11111111111111111110000001101010;
assign LUT_1[31689] = 32'b11111111111111110111010011100110;
assign LUT_1[31690] = 32'b11111111111111111001101111111011;
assign LUT_1[31691] = 32'b11111111111111110011000001110111;
assign LUT_1[31692] = 32'b00000000000000000101111011000001;
assign LUT_1[31693] = 32'b11111111111111111111001100111101;
assign LUT_1[31694] = 32'b00000000000000000001101001010010;
assign LUT_1[31695] = 32'b11111111111111111010111011001110;
assign LUT_1[31696] = 32'b00000000000000000000101111010111;
assign LUT_1[31697] = 32'b11111111111111111010000001010011;
assign LUT_1[31698] = 32'b11111111111111111100011101101000;
assign LUT_1[31699] = 32'b11111111111111110101101111100100;
assign LUT_1[31700] = 32'b00000000000000001000101000101110;
assign LUT_1[31701] = 32'b00000000000000000001111010101010;
assign LUT_1[31702] = 32'b00000000000000000100010110111111;
assign LUT_1[31703] = 32'b11111111111111111101101000111011;
assign LUT_1[31704] = 32'b11111111111111111111111101001100;
assign LUT_1[31705] = 32'b11111111111111111001001111001000;
assign LUT_1[31706] = 32'b11111111111111111011101011011101;
assign LUT_1[31707] = 32'b11111111111111110100111101011001;
assign LUT_1[31708] = 32'b00000000000000000111110110100011;
assign LUT_1[31709] = 32'b00000000000000000001001000011111;
assign LUT_1[31710] = 32'b00000000000000000011100100110100;
assign LUT_1[31711] = 32'b11111111111111111100110110110000;
assign LUT_1[31712] = 32'b11111111111111111111101110110100;
assign LUT_1[31713] = 32'b11111111111111111001000000110000;
assign LUT_1[31714] = 32'b11111111111111111011011101000101;
assign LUT_1[31715] = 32'b11111111111111110100101111000001;
assign LUT_1[31716] = 32'b00000000000000000111101000001011;
assign LUT_1[31717] = 32'b00000000000000000000111010000111;
assign LUT_1[31718] = 32'b00000000000000000011010110011100;
assign LUT_1[31719] = 32'b11111111111111111100101000011000;
assign LUT_1[31720] = 32'b11111111111111111110111100101001;
assign LUT_1[31721] = 32'b11111111111111111000001110100101;
assign LUT_1[31722] = 32'b11111111111111111010101010111010;
assign LUT_1[31723] = 32'b11111111111111110011111100110110;
assign LUT_1[31724] = 32'b00000000000000000110110110000000;
assign LUT_1[31725] = 32'b00000000000000000000000111111100;
assign LUT_1[31726] = 32'b00000000000000000010100100010001;
assign LUT_1[31727] = 32'b11111111111111111011110110001101;
assign LUT_1[31728] = 32'b00000000000000000001101010010110;
assign LUT_1[31729] = 32'b11111111111111111010111100010010;
assign LUT_1[31730] = 32'b11111111111111111101011000100111;
assign LUT_1[31731] = 32'b11111111111111110110101010100011;
assign LUT_1[31732] = 32'b00000000000000001001100011101101;
assign LUT_1[31733] = 32'b00000000000000000010110101101001;
assign LUT_1[31734] = 32'b00000000000000000101010001111110;
assign LUT_1[31735] = 32'b11111111111111111110100011111010;
assign LUT_1[31736] = 32'b00000000000000000000111000001011;
assign LUT_1[31737] = 32'b11111111111111111010001010000111;
assign LUT_1[31738] = 32'b11111111111111111100100110011100;
assign LUT_1[31739] = 32'b11111111111111110101111000011000;
assign LUT_1[31740] = 32'b00000000000000001000110001100010;
assign LUT_1[31741] = 32'b00000000000000000010000011011110;
assign LUT_1[31742] = 32'b00000000000000000100011111110011;
assign LUT_1[31743] = 32'b11111111111111111101110001101111;
assign LUT_1[31744] = 32'b00000000000000001000101010010001;
assign LUT_1[31745] = 32'b00000000000000000001111100001101;
assign LUT_1[31746] = 32'b00000000000000000100011000100010;
assign LUT_1[31747] = 32'b11111111111111111101101010011110;
assign LUT_1[31748] = 32'b00000000000000010000100011101000;
assign LUT_1[31749] = 32'b00000000000000001001110101100100;
assign LUT_1[31750] = 32'b00000000000000001100010001111001;
assign LUT_1[31751] = 32'b00000000000000000101100011110101;
assign LUT_1[31752] = 32'b00000000000000000111111000000110;
assign LUT_1[31753] = 32'b00000000000000000001001010000010;
assign LUT_1[31754] = 32'b00000000000000000011100110010111;
assign LUT_1[31755] = 32'b11111111111111111100111000010011;
assign LUT_1[31756] = 32'b00000000000000001111110001011101;
assign LUT_1[31757] = 32'b00000000000000001001000011011001;
assign LUT_1[31758] = 32'b00000000000000001011011111101110;
assign LUT_1[31759] = 32'b00000000000000000100110001101010;
assign LUT_1[31760] = 32'b00000000000000001010100101110011;
assign LUT_1[31761] = 32'b00000000000000000011110111101111;
assign LUT_1[31762] = 32'b00000000000000000110010100000100;
assign LUT_1[31763] = 32'b11111111111111111111100110000000;
assign LUT_1[31764] = 32'b00000000000000010010011111001010;
assign LUT_1[31765] = 32'b00000000000000001011110001000110;
assign LUT_1[31766] = 32'b00000000000000001110001101011011;
assign LUT_1[31767] = 32'b00000000000000000111011111010111;
assign LUT_1[31768] = 32'b00000000000000001001110011101000;
assign LUT_1[31769] = 32'b00000000000000000011000101100100;
assign LUT_1[31770] = 32'b00000000000000000101100001111001;
assign LUT_1[31771] = 32'b11111111111111111110110011110101;
assign LUT_1[31772] = 32'b00000000000000010001101100111111;
assign LUT_1[31773] = 32'b00000000000000001010111110111011;
assign LUT_1[31774] = 32'b00000000000000001101011011010000;
assign LUT_1[31775] = 32'b00000000000000000110101101001100;
assign LUT_1[31776] = 32'b00000000000000001001100101010000;
assign LUT_1[31777] = 32'b00000000000000000010110111001100;
assign LUT_1[31778] = 32'b00000000000000000101010011100001;
assign LUT_1[31779] = 32'b11111111111111111110100101011101;
assign LUT_1[31780] = 32'b00000000000000010001011110100111;
assign LUT_1[31781] = 32'b00000000000000001010110000100011;
assign LUT_1[31782] = 32'b00000000000000001101001100111000;
assign LUT_1[31783] = 32'b00000000000000000110011110110100;
assign LUT_1[31784] = 32'b00000000000000001000110011000101;
assign LUT_1[31785] = 32'b00000000000000000010000101000001;
assign LUT_1[31786] = 32'b00000000000000000100100001010110;
assign LUT_1[31787] = 32'b11111111111111111101110011010010;
assign LUT_1[31788] = 32'b00000000000000010000101100011100;
assign LUT_1[31789] = 32'b00000000000000001001111110011000;
assign LUT_1[31790] = 32'b00000000000000001100011010101101;
assign LUT_1[31791] = 32'b00000000000000000101101100101001;
assign LUT_1[31792] = 32'b00000000000000001011100000110010;
assign LUT_1[31793] = 32'b00000000000000000100110010101110;
assign LUT_1[31794] = 32'b00000000000000000111001111000011;
assign LUT_1[31795] = 32'b00000000000000000000100000111111;
assign LUT_1[31796] = 32'b00000000000000010011011010001001;
assign LUT_1[31797] = 32'b00000000000000001100101100000101;
assign LUT_1[31798] = 32'b00000000000000001111001000011010;
assign LUT_1[31799] = 32'b00000000000000001000011010010110;
assign LUT_1[31800] = 32'b00000000000000001010101110100111;
assign LUT_1[31801] = 32'b00000000000000000100000000100011;
assign LUT_1[31802] = 32'b00000000000000000110011100111000;
assign LUT_1[31803] = 32'b11111111111111111111101110110100;
assign LUT_1[31804] = 32'b00000000000000010010100111111110;
assign LUT_1[31805] = 32'b00000000000000001011111001111010;
assign LUT_1[31806] = 32'b00000000000000001110010110001111;
assign LUT_1[31807] = 32'b00000000000000000111101000001011;
assign LUT_1[31808] = 32'b00000000000000001010100111111001;
assign LUT_1[31809] = 32'b00000000000000000011111001110101;
assign LUT_1[31810] = 32'b00000000000000000110010110001010;
assign LUT_1[31811] = 32'b11111111111111111111101000000110;
assign LUT_1[31812] = 32'b00000000000000010010100001010000;
assign LUT_1[31813] = 32'b00000000000000001011110011001100;
assign LUT_1[31814] = 32'b00000000000000001110001111100001;
assign LUT_1[31815] = 32'b00000000000000000111100001011101;
assign LUT_1[31816] = 32'b00000000000000001001110101101110;
assign LUT_1[31817] = 32'b00000000000000000011000111101010;
assign LUT_1[31818] = 32'b00000000000000000101100011111111;
assign LUT_1[31819] = 32'b11111111111111111110110101111011;
assign LUT_1[31820] = 32'b00000000000000010001101111000101;
assign LUT_1[31821] = 32'b00000000000000001011000001000001;
assign LUT_1[31822] = 32'b00000000000000001101011101010110;
assign LUT_1[31823] = 32'b00000000000000000110101111010010;
assign LUT_1[31824] = 32'b00000000000000001100100011011011;
assign LUT_1[31825] = 32'b00000000000000000101110101010111;
assign LUT_1[31826] = 32'b00000000000000001000010001101100;
assign LUT_1[31827] = 32'b00000000000000000001100011101000;
assign LUT_1[31828] = 32'b00000000000000010100011100110010;
assign LUT_1[31829] = 32'b00000000000000001101101110101110;
assign LUT_1[31830] = 32'b00000000000000010000001011000011;
assign LUT_1[31831] = 32'b00000000000000001001011100111111;
assign LUT_1[31832] = 32'b00000000000000001011110001010000;
assign LUT_1[31833] = 32'b00000000000000000101000011001100;
assign LUT_1[31834] = 32'b00000000000000000111011111100001;
assign LUT_1[31835] = 32'b00000000000000000000110001011101;
assign LUT_1[31836] = 32'b00000000000000010011101010100111;
assign LUT_1[31837] = 32'b00000000000000001100111100100011;
assign LUT_1[31838] = 32'b00000000000000001111011000111000;
assign LUT_1[31839] = 32'b00000000000000001000101010110100;
assign LUT_1[31840] = 32'b00000000000000001011100010111000;
assign LUT_1[31841] = 32'b00000000000000000100110100110100;
assign LUT_1[31842] = 32'b00000000000000000111010001001001;
assign LUT_1[31843] = 32'b00000000000000000000100011000101;
assign LUT_1[31844] = 32'b00000000000000010011011100001111;
assign LUT_1[31845] = 32'b00000000000000001100101110001011;
assign LUT_1[31846] = 32'b00000000000000001111001010100000;
assign LUT_1[31847] = 32'b00000000000000001000011100011100;
assign LUT_1[31848] = 32'b00000000000000001010110000101101;
assign LUT_1[31849] = 32'b00000000000000000100000010101001;
assign LUT_1[31850] = 32'b00000000000000000110011110111110;
assign LUT_1[31851] = 32'b11111111111111111111110000111010;
assign LUT_1[31852] = 32'b00000000000000010010101010000100;
assign LUT_1[31853] = 32'b00000000000000001011111100000000;
assign LUT_1[31854] = 32'b00000000000000001110011000010101;
assign LUT_1[31855] = 32'b00000000000000000111101010010001;
assign LUT_1[31856] = 32'b00000000000000001101011110011010;
assign LUT_1[31857] = 32'b00000000000000000110110000010110;
assign LUT_1[31858] = 32'b00000000000000001001001100101011;
assign LUT_1[31859] = 32'b00000000000000000010011110100111;
assign LUT_1[31860] = 32'b00000000000000010101010111110001;
assign LUT_1[31861] = 32'b00000000000000001110101001101101;
assign LUT_1[31862] = 32'b00000000000000010001000110000010;
assign LUT_1[31863] = 32'b00000000000000001010010111111110;
assign LUT_1[31864] = 32'b00000000000000001100101100001111;
assign LUT_1[31865] = 32'b00000000000000000101111110001011;
assign LUT_1[31866] = 32'b00000000000000001000011010100000;
assign LUT_1[31867] = 32'b00000000000000000001101100011100;
assign LUT_1[31868] = 32'b00000000000000010100100101100110;
assign LUT_1[31869] = 32'b00000000000000001101110111100010;
assign LUT_1[31870] = 32'b00000000000000010000010011110111;
assign LUT_1[31871] = 32'b00000000000000001001100101110011;
assign LUT_1[31872] = 32'b00000000000000001011101010010100;
assign LUT_1[31873] = 32'b00000000000000000100111100010000;
assign LUT_1[31874] = 32'b00000000000000000111011000100101;
assign LUT_1[31875] = 32'b00000000000000000000101010100001;
assign LUT_1[31876] = 32'b00000000000000010011100011101011;
assign LUT_1[31877] = 32'b00000000000000001100110101100111;
assign LUT_1[31878] = 32'b00000000000000001111010001111100;
assign LUT_1[31879] = 32'b00000000000000001000100011111000;
assign LUT_1[31880] = 32'b00000000000000001010111000001001;
assign LUT_1[31881] = 32'b00000000000000000100001010000101;
assign LUT_1[31882] = 32'b00000000000000000110100110011010;
assign LUT_1[31883] = 32'b11111111111111111111111000010110;
assign LUT_1[31884] = 32'b00000000000000010010110001100000;
assign LUT_1[31885] = 32'b00000000000000001100000011011100;
assign LUT_1[31886] = 32'b00000000000000001110011111110001;
assign LUT_1[31887] = 32'b00000000000000000111110001101101;
assign LUT_1[31888] = 32'b00000000000000001101100101110110;
assign LUT_1[31889] = 32'b00000000000000000110110111110010;
assign LUT_1[31890] = 32'b00000000000000001001010100000111;
assign LUT_1[31891] = 32'b00000000000000000010100110000011;
assign LUT_1[31892] = 32'b00000000000000010101011111001101;
assign LUT_1[31893] = 32'b00000000000000001110110001001001;
assign LUT_1[31894] = 32'b00000000000000010001001101011110;
assign LUT_1[31895] = 32'b00000000000000001010011111011010;
assign LUT_1[31896] = 32'b00000000000000001100110011101011;
assign LUT_1[31897] = 32'b00000000000000000110000101100111;
assign LUT_1[31898] = 32'b00000000000000001000100001111100;
assign LUT_1[31899] = 32'b00000000000000000001110011111000;
assign LUT_1[31900] = 32'b00000000000000010100101101000010;
assign LUT_1[31901] = 32'b00000000000000001101111110111110;
assign LUT_1[31902] = 32'b00000000000000010000011011010011;
assign LUT_1[31903] = 32'b00000000000000001001101101001111;
assign LUT_1[31904] = 32'b00000000000000001100100101010011;
assign LUT_1[31905] = 32'b00000000000000000101110111001111;
assign LUT_1[31906] = 32'b00000000000000001000010011100100;
assign LUT_1[31907] = 32'b00000000000000000001100101100000;
assign LUT_1[31908] = 32'b00000000000000010100011110101010;
assign LUT_1[31909] = 32'b00000000000000001101110000100110;
assign LUT_1[31910] = 32'b00000000000000010000001100111011;
assign LUT_1[31911] = 32'b00000000000000001001011110110111;
assign LUT_1[31912] = 32'b00000000000000001011110011001000;
assign LUT_1[31913] = 32'b00000000000000000101000101000100;
assign LUT_1[31914] = 32'b00000000000000000111100001011001;
assign LUT_1[31915] = 32'b00000000000000000000110011010101;
assign LUT_1[31916] = 32'b00000000000000010011101100011111;
assign LUT_1[31917] = 32'b00000000000000001100111110011011;
assign LUT_1[31918] = 32'b00000000000000001111011010110000;
assign LUT_1[31919] = 32'b00000000000000001000101100101100;
assign LUT_1[31920] = 32'b00000000000000001110100000110101;
assign LUT_1[31921] = 32'b00000000000000000111110010110001;
assign LUT_1[31922] = 32'b00000000000000001010001111000110;
assign LUT_1[31923] = 32'b00000000000000000011100001000010;
assign LUT_1[31924] = 32'b00000000000000010110011010001100;
assign LUT_1[31925] = 32'b00000000000000001111101100001000;
assign LUT_1[31926] = 32'b00000000000000010010001000011101;
assign LUT_1[31927] = 32'b00000000000000001011011010011001;
assign LUT_1[31928] = 32'b00000000000000001101101110101010;
assign LUT_1[31929] = 32'b00000000000000000111000000100110;
assign LUT_1[31930] = 32'b00000000000000001001011100111011;
assign LUT_1[31931] = 32'b00000000000000000010101110110111;
assign LUT_1[31932] = 32'b00000000000000010101101000000001;
assign LUT_1[31933] = 32'b00000000000000001110111001111101;
assign LUT_1[31934] = 32'b00000000000000010001010110010010;
assign LUT_1[31935] = 32'b00000000000000001010101000001110;
assign LUT_1[31936] = 32'b00000000000000001101100111111100;
assign LUT_1[31937] = 32'b00000000000000000110111001111000;
assign LUT_1[31938] = 32'b00000000000000001001010110001101;
assign LUT_1[31939] = 32'b00000000000000000010101000001001;
assign LUT_1[31940] = 32'b00000000000000010101100001010011;
assign LUT_1[31941] = 32'b00000000000000001110110011001111;
assign LUT_1[31942] = 32'b00000000000000010001001111100100;
assign LUT_1[31943] = 32'b00000000000000001010100001100000;
assign LUT_1[31944] = 32'b00000000000000001100110101110001;
assign LUT_1[31945] = 32'b00000000000000000110000111101101;
assign LUT_1[31946] = 32'b00000000000000001000100100000010;
assign LUT_1[31947] = 32'b00000000000000000001110101111110;
assign LUT_1[31948] = 32'b00000000000000010100101111001000;
assign LUT_1[31949] = 32'b00000000000000001110000001000100;
assign LUT_1[31950] = 32'b00000000000000010000011101011001;
assign LUT_1[31951] = 32'b00000000000000001001101111010101;
assign LUT_1[31952] = 32'b00000000000000001111100011011110;
assign LUT_1[31953] = 32'b00000000000000001000110101011010;
assign LUT_1[31954] = 32'b00000000000000001011010001101111;
assign LUT_1[31955] = 32'b00000000000000000100100011101011;
assign LUT_1[31956] = 32'b00000000000000010111011100110101;
assign LUT_1[31957] = 32'b00000000000000010000101110110001;
assign LUT_1[31958] = 32'b00000000000000010011001011000110;
assign LUT_1[31959] = 32'b00000000000000001100011101000010;
assign LUT_1[31960] = 32'b00000000000000001110110001010011;
assign LUT_1[31961] = 32'b00000000000000001000000011001111;
assign LUT_1[31962] = 32'b00000000000000001010011111100100;
assign LUT_1[31963] = 32'b00000000000000000011110001100000;
assign LUT_1[31964] = 32'b00000000000000010110101010101010;
assign LUT_1[31965] = 32'b00000000000000001111111100100110;
assign LUT_1[31966] = 32'b00000000000000010010011000111011;
assign LUT_1[31967] = 32'b00000000000000001011101010110111;
assign LUT_1[31968] = 32'b00000000000000001110100010111011;
assign LUT_1[31969] = 32'b00000000000000000111110100110111;
assign LUT_1[31970] = 32'b00000000000000001010010001001100;
assign LUT_1[31971] = 32'b00000000000000000011100011001000;
assign LUT_1[31972] = 32'b00000000000000010110011100010010;
assign LUT_1[31973] = 32'b00000000000000001111101110001110;
assign LUT_1[31974] = 32'b00000000000000010010001010100011;
assign LUT_1[31975] = 32'b00000000000000001011011100011111;
assign LUT_1[31976] = 32'b00000000000000001101110000110000;
assign LUT_1[31977] = 32'b00000000000000000111000010101100;
assign LUT_1[31978] = 32'b00000000000000001001011111000001;
assign LUT_1[31979] = 32'b00000000000000000010110000111101;
assign LUT_1[31980] = 32'b00000000000000010101101010000111;
assign LUT_1[31981] = 32'b00000000000000001110111100000011;
assign LUT_1[31982] = 32'b00000000000000010001011000011000;
assign LUT_1[31983] = 32'b00000000000000001010101010010100;
assign LUT_1[31984] = 32'b00000000000000010000011110011101;
assign LUT_1[31985] = 32'b00000000000000001001110000011001;
assign LUT_1[31986] = 32'b00000000000000001100001100101110;
assign LUT_1[31987] = 32'b00000000000000000101011110101010;
assign LUT_1[31988] = 32'b00000000000000011000010111110100;
assign LUT_1[31989] = 32'b00000000000000010001101001110000;
assign LUT_1[31990] = 32'b00000000000000010100000110000101;
assign LUT_1[31991] = 32'b00000000000000001101011000000001;
assign LUT_1[31992] = 32'b00000000000000001111101100010010;
assign LUT_1[31993] = 32'b00000000000000001000111110001110;
assign LUT_1[31994] = 32'b00000000000000001011011010100011;
assign LUT_1[31995] = 32'b00000000000000000100101100011111;
assign LUT_1[31996] = 32'b00000000000000010111100101101001;
assign LUT_1[31997] = 32'b00000000000000010000110111100101;
assign LUT_1[31998] = 32'b00000000000000010011010011111010;
assign LUT_1[31999] = 32'b00000000000000001100100101110110;
assign LUT_1[32000] = 32'b00000000000000000110011110011101;
assign LUT_1[32001] = 32'b11111111111111111111110000011001;
assign LUT_1[32002] = 32'b00000000000000000010001100101110;
assign LUT_1[32003] = 32'b11111111111111111011011110101010;
assign LUT_1[32004] = 32'b00000000000000001110010111110100;
assign LUT_1[32005] = 32'b00000000000000000111101001110000;
assign LUT_1[32006] = 32'b00000000000000001010000110000101;
assign LUT_1[32007] = 32'b00000000000000000011011000000001;
assign LUT_1[32008] = 32'b00000000000000000101101100010010;
assign LUT_1[32009] = 32'b11111111111111111110111110001110;
assign LUT_1[32010] = 32'b00000000000000000001011010100011;
assign LUT_1[32011] = 32'b11111111111111111010101100011111;
assign LUT_1[32012] = 32'b00000000000000001101100101101001;
assign LUT_1[32013] = 32'b00000000000000000110110111100101;
assign LUT_1[32014] = 32'b00000000000000001001010011111010;
assign LUT_1[32015] = 32'b00000000000000000010100101110110;
assign LUT_1[32016] = 32'b00000000000000001000011001111111;
assign LUT_1[32017] = 32'b00000000000000000001101011111011;
assign LUT_1[32018] = 32'b00000000000000000100001000010000;
assign LUT_1[32019] = 32'b11111111111111111101011010001100;
assign LUT_1[32020] = 32'b00000000000000010000010011010110;
assign LUT_1[32021] = 32'b00000000000000001001100101010010;
assign LUT_1[32022] = 32'b00000000000000001100000001100111;
assign LUT_1[32023] = 32'b00000000000000000101010011100011;
assign LUT_1[32024] = 32'b00000000000000000111100111110100;
assign LUT_1[32025] = 32'b00000000000000000000111001110000;
assign LUT_1[32026] = 32'b00000000000000000011010110000101;
assign LUT_1[32027] = 32'b11111111111111111100101000000001;
assign LUT_1[32028] = 32'b00000000000000001111100001001011;
assign LUT_1[32029] = 32'b00000000000000001000110011000111;
assign LUT_1[32030] = 32'b00000000000000001011001111011100;
assign LUT_1[32031] = 32'b00000000000000000100100001011000;
assign LUT_1[32032] = 32'b00000000000000000111011001011100;
assign LUT_1[32033] = 32'b00000000000000000000101011011000;
assign LUT_1[32034] = 32'b00000000000000000011000111101101;
assign LUT_1[32035] = 32'b11111111111111111100011001101001;
assign LUT_1[32036] = 32'b00000000000000001111010010110011;
assign LUT_1[32037] = 32'b00000000000000001000100100101111;
assign LUT_1[32038] = 32'b00000000000000001011000001000100;
assign LUT_1[32039] = 32'b00000000000000000100010011000000;
assign LUT_1[32040] = 32'b00000000000000000110100111010001;
assign LUT_1[32041] = 32'b11111111111111111111111001001101;
assign LUT_1[32042] = 32'b00000000000000000010010101100010;
assign LUT_1[32043] = 32'b11111111111111111011100111011110;
assign LUT_1[32044] = 32'b00000000000000001110100000101000;
assign LUT_1[32045] = 32'b00000000000000000111110010100100;
assign LUT_1[32046] = 32'b00000000000000001010001110111001;
assign LUT_1[32047] = 32'b00000000000000000011100000110101;
assign LUT_1[32048] = 32'b00000000000000001001010100111110;
assign LUT_1[32049] = 32'b00000000000000000010100110111010;
assign LUT_1[32050] = 32'b00000000000000000101000011001111;
assign LUT_1[32051] = 32'b11111111111111111110010101001011;
assign LUT_1[32052] = 32'b00000000000000010001001110010101;
assign LUT_1[32053] = 32'b00000000000000001010100000010001;
assign LUT_1[32054] = 32'b00000000000000001100111100100110;
assign LUT_1[32055] = 32'b00000000000000000110001110100010;
assign LUT_1[32056] = 32'b00000000000000001000100010110011;
assign LUT_1[32057] = 32'b00000000000000000001110100101111;
assign LUT_1[32058] = 32'b00000000000000000100010001000100;
assign LUT_1[32059] = 32'b11111111111111111101100011000000;
assign LUT_1[32060] = 32'b00000000000000010000011100001010;
assign LUT_1[32061] = 32'b00000000000000001001101110000110;
assign LUT_1[32062] = 32'b00000000000000001100001010011011;
assign LUT_1[32063] = 32'b00000000000000000101011100010111;
assign LUT_1[32064] = 32'b00000000000000001000011100000101;
assign LUT_1[32065] = 32'b00000000000000000001101110000001;
assign LUT_1[32066] = 32'b00000000000000000100001010010110;
assign LUT_1[32067] = 32'b11111111111111111101011100010010;
assign LUT_1[32068] = 32'b00000000000000010000010101011100;
assign LUT_1[32069] = 32'b00000000000000001001100111011000;
assign LUT_1[32070] = 32'b00000000000000001100000011101101;
assign LUT_1[32071] = 32'b00000000000000000101010101101001;
assign LUT_1[32072] = 32'b00000000000000000111101001111010;
assign LUT_1[32073] = 32'b00000000000000000000111011110110;
assign LUT_1[32074] = 32'b00000000000000000011011000001011;
assign LUT_1[32075] = 32'b11111111111111111100101010000111;
assign LUT_1[32076] = 32'b00000000000000001111100011010001;
assign LUT_1[32077] = 32'b00000000000000001000110101001101;
assign LUT_1[32078] = 32'b00000000000000001011010001100010;
assign LUT_1[32079] = 32'b00000000000000000100100011011110;
assign LUT_1[32080] = 32'b00000000000000001010010111100111;
assign LUT_1[32081] = 32'b00000000000000000011101001100011;
assign LUT_1[32082] = 32'b00000000000000000110000101111000;
assign LUT_1[32083] = 32'b11111111111111111111010111110100;
assign LUT_1[32084] = 32'b00000000000000010010010000111110;
assign LUT_1[32085] = 32'b00000000000000001011100010111010;
assign LUT_1[32086] = 32'b00000000000000001101111111001111;
assign LUT_1[32087] = 32'b00000000000000000111010001001011;
assign LUT_1[32088] = 32'b00000000000000001001100101011100;
assign LUT_1[32089] = 32'b00000000000000000010110111011000;
assign LUT_1[32090] = 32'b00000000000000000101010011101101;
assign LUT_1[32091] = 32'b11111111111111111110100101101001;
assign LUT_1[32092] = 32'b00000000000000010001011110110011;
assign LUT_1[32093] = 32'b00000000000000001010110000101111;
assign LUT_1[32094] = 32'b00000000000000001101001101000100;
assign LUT_1[32095] = 32'b00000000000000000110011111000000;
assign LUT_1[32096] = 32'b00000000000000001001010111000100;
assign LUT_1[32097] = 32'b00000000000000000010101001000000;
assign LUT_1[32098] = 32'b00000000000000000101000101010101;
assign LUT_1[32099] = 32'b11111111111111111110010111010001;
assign LUT_1[32100] = 32'b00000000000000010001010000011011;
assign LUT_1[32101] = 32'b00000000000000001010100010010111;
assign LUT_1[32102] = 32'b00000000000000001100111110101100;
assign LUT_1[32103] = 32'b00000000000000000110010000101000;
assign LUT_1[32104] = 32'b00000000000000001000100100111001;
assign LUT_1[32105] = 32'b00000000000000000001110110110101;
assign LUT_1[32106] = 32'b00000000000000000100010011001010;
assign LUT_1[32107] = 32'b11111111111111111101100101000110;
assign LUT_1[32108] = 32'b00000000000000010000011110010000;
assign LUT_1[32109] = 32'b00000000000000001001110000001100;
assign LUT_1[32110] = 32'b00000000000000001100001100100001;
assign LUT_1[32111] = 32'b00000000000000000101011110011101;
assign LUT_1[32112] = 32'b00000000000000001011010010100110;
assign LUT_1[32113] = 32'b00000000000000000100100100100010;
assign LUT_1[32114] = 32'b00000000000000000111000000110111;
assign LUT_1[32115] = 32'b00000000000000000000010010110011;
assign LUT_1[32116] = 32'b00000000000000010011001011111101;
assign LUT_1[32117] = 32'b00000000000000001100011101111001;
assign LUT_1[32118] = 32'b00000000000000001110111010001110;
assign LUT_1[32119] = 32'b00000000000000001000001100001010;
assign LUT_1[32120] = 32'b00000000000000001010100000011011;
assign LUT_1[32121] = 32'b00000000000000000011110010010111;
assign LUT_1[32122] = 32'b00000000000000000110001110101100;
assign LUT_1[32123] = 32'b11111111111111111111100000101000;
assign LUT_1[32124] = 32'b00000000000000010010011001110010;
assign LUT_1[32125] = 32'b00000000000000001011101011101110;
assign LUT_1[32126] = 32'b00000000000000001110001000000011;
assign LUT_1[32127] = 32'b00000000000000000111011001111111;
assign LUT_1[32128] = 32'b00000000000000001001011110100000;
assign LUT_1[32129] = 32'b00000000000000000010110000011100;
assign LUT_1[32130] = 32'b00000000000000000101001100110001;
assign LUT_1[32131] = 32'b11111111111111111110011110101101;
assign LUT_1[32132] = 32'b00000000000000010001010111110111;
assign LUT_1[32133] = 32'b00000000000000001010101001110011;
assign LUT_1[32134] = 32'b00000000000000001101000110001000;
assign LUT_1[32135] = 32'b00000000000000000110011000000100;
assign LUT_1[32136] = 32'b00000000000000001000101100010101;
assign LUT_1[32137] = 32'b00000000000000000001111110010001;
assign LUT_1[32138] = 32'b00000000000000000100011010100110;
assign LUT_1[32139] = 32'b11111111111111111101101100100010;
assign LUT_1[32140] = 32'b00000000000000010000100101101100;
assign LUT_1[32141] = 32'b00000000000000001001110111101000;
assign LUT_1[32142] = 32'b00000000000000001100010011111101;
assign LUT_1[32143] = 32'b00000000000000000101100101111001;
assign LUT_1[32144] = 32'b00000000000000001011011010000010;
assign LUT_1[32145] = 32'b00000000000000000100101011111110;
assign LUT_1[32146] = 32'b00000000000000000111001000010011;
assign LUT_1[32147] = 32'b00000000000000000000011010001111;
assign LUT_1[32148] = 32'b00000000000000010011010011011001;
assign LUT_1[32149] = 32'b00000000000000001100100101010101;
assign LUT_1[32150] = 32'b00000000000000001111000001101010;
assign LUT_1[32151] = 32'b00000000000000001000010011100110;
assign LUT_1[32152] = 32'b00000000000000001010100111110111;
assign LUT_1[32153] = 32'b00000000000000000011111001110011;
assign LUT_1[32154] = 32'b00000000000000000110010110001000;
assign LUT_1[32155] = 32'b11111111111111111111101000000100;
assign LUT_1[32156] = 32'b00000000000000010010100001001110;
assign LUT_1[32157] = 32'b00000000000000001011110011001010;
assign LUT_1[32158] = 32'b00000000000000001110001111011111;
assign LUT_1[32159] = 32'b00000000000000000111100001011011;
assign LUT_1[32160] = 32'b00000000000000001010011001011111;
assign LUT_1[32161] = 32'b00000000000000000011101011011011;
assign LUT_1[32162] = 32'b00000000000000000110000111110000;
assign LUT_1[32163] = 32'b11111111111111111111011001101100;
assign LUT_1[32164] = 32'b00000000000000010010010010110110;
assign LUT_1[32165] = 32'b00000000000000001011100100110010;
assign LUT_1[32166] = 32'b00000000000000001110000001000111;
assign LUT_1[32167] = 32'b00000000000000000111010011000011;
assign LUT_1[32168] = 32'b00000000000000001001100111010100;
assign LUT_1[32169] = 32'b00000000000000000010111001010000;
assign LUT_1[32170] = 32'b00000000000000000101010101100101;
assign LUT_1[32171] = 32'b11111111111111111110100111100001;
assign LUT_1[32172] = 32'b00000000000000010001100000101011;
assign LUT_1[32173] = 32'b00000000000000001010110010100111;
assign LUT_1[32174] = 32'b00000000000000001101001110111100;
assign LUT_1[32175] = 32'b00000000000000000110100000111000;
assign LUT_1[32176] = 32'b00000000000000001100010101000001;
assign LUT_1[32177] = 32'b00000000000000000101100110111101;
assign LUT_1[32178] = 32'b00000000000000001000000011010010;
assign LUT_1[32179] = 32'b00000000000000000001010101001110;
assign LUT_1[32180] = 32'b00000000000000010100001110011000;
assign LUT_1[32181] = 32'b00000000000000001101100000010100;
assign LUT_1[32182] = 32'b00000000000000001111111100101001;
assign LUT_1[32183] = 32'b00000000000000001001001110100101;
assign LUT_1[32184] = 32'b00000000000000001011100010110110;
assign LUT_1[32185] = 32'b00000000000000000100110100110010;
assign LUT_1[32186] = 32'b00000000000000000111010001000111;
assign LUT_1[32187] = 32'b00000000000000000000100011000011;
assign LUT_1[32188] = 32'b00000000000000010011011100001101;
assign LUT_1[32189] = 32'b00000000000000001100101110001001;
assign LUT_1[32190] = 32'b00000000000000001111001010011110;
assign LUT_1[32191] = 32'b00000000000000001000011100011010;
assign LUT_1[32192] = 32'b00000000000000001011011100001000;
assign LUT_1[32193] = 32'b00000000000000000100101110000100;
assign LUT_1[32194] = 32'b00000000000000000111001010011001;
assign LUT_1[32195] = 32'b00000000000000000000011100010101;
assign LUT_1[32196] = 32'b00000000000000010011010101011111;
assign LUT_1[32197] = 32'b00000000000000001100100111011011;
assign LUT_1[32198] = 32'b00000000000000001111000011110000;
assign LUT_1[32199] = 32'b00000000000000001000010101101100;
assign LUT_1[32200] = 32'b00000000000000001010101001111101;
assign LUT_1[32201] = 32'b00000000000000000011111011111001;
assign LUT_1[32202] = 32'b00000000000000000110011000001110;
assign LUT_1[32203] = 32'b11111111111111111111101010001010;
assign LUT_1[32204] = 32'b00000000000000010010100011010100;
assign LUT_1[32205] = 32'b00000000000000001011110101010000;
assign LUT_1[32206] = 32'b00000000000000001110010001100101;
assign LUT_1[32207] = 32'b00000000000000000111100011100001;
assign LUT_1[32208] = 32'b00000000000000001101010111101010;
assign LUT_1[32209] = 32'b00000000000000000110101001100110;
assign LUT_1[32210] = 32'b00000000000000001001000101111011;
assign LUT_1[32211] = 32'b00000000000000000010010111110111;
assign LUT_1[32212] = 32'b00000000000000010101010001000001;
assign LUT_1[32213] = 32'b00000000000000001110100010111101;
assign LUT_1[32214] = 32'b00000000000000010000111111010010;
assign LUT_1[32215] = 32'b00000000000000001010010001001110;
assign LUT_1[32216] = 32'b00000000000000001100100101011111;
assign LUT_1[32217] = 32'b00000000000000000101110111011011;
assign LUT_1[32218] = 32'b00000000000000001000010011110000;
assign LUT_1[32219] = 32'b00000000000000000001100101101100;
assign LUT_1[32220] = 32'b00000000000000010100011110110110;
assign LUT_1[32221] = 32'b00000000000000001101110000110010;
assign LUT_1[32222] = 32'b00000000000000010000001101000111;
assign LUT_1[32223] = 32'b00000000000000001001011111000011;
assign LUT_1[32224] = 32'b00000000000000001100010111000111;
assign LUT_1[32225] = 32'b00000000000000000101101001000011;
assign LUT_1[32226] = 32'b00000000000000001000000101011000;
assign LUT_1[32227] = 32'b00000000000000000001010111010100;
assign LUT_1[32228] = 32'b00000000000000010100010000011110;
assign LUT_1[32229] = 32'b00000000000000001101100010011010;
assign LUT_1[32230] = 32'b00000000000000001111111110101111;
assign LUT_1[32231] = 32'b00000000000000001001010000101011;
assign LUT_1[32232] = 32'b00000000000000001011100100111100;
assign LUT_1[32233] = 32'b00000000000000000100110110111000;
assign LUT_1[32234] = 32'b00000000000000000111010011001101;
assign LUT_1[32235] = 32'b00000000000000000000100101001001;
assign LUT_1[32236] = 32'b00000000000000010011011110010011;
assign LUT_1[32237] = 32'b00000000000000001100110000001111;
assign LUT_1[32238] = 32'b00000000000000001111001100100100;
assign LUT_1[32239] = 32'b00000000000000001000011110100000;
assign LUT_1[32240] = 32'b00000000000000001110010010101001;
assign LUT_1[32241] = 32'b00000000000000000111100100100101;
assign LUT_1[32242] = 32'b00000000000000001010000000111010;
assign LUT_1[32243] = 32'b00000000000000000011010010110110;
assign LUT_1[32244] = 32'b00000000000000010110001100000000;
assign LUT_1[32245] = 32'b00000000000000001111011101111100;
assign LUT_1[32246] = 32'b00000000000000010001111010010001;
assign LUT_1[32247] = 32'b00000000000000001011001100001101;
assign LUT_1[32248] = 32'b00000000000000001101100000011110;
assign LUT_1[32249] = 32'b00000000000000000110110010011010;
assign LUT_1[32250] = 32'b00000000000000001001001110101111;
assign LUT_1[32251] = 32'b00000000000000000010100000101011;
assign LUT_1[32252] = 32'b00000000000000010101011001110101;
assign LUT_1[32253] = 32'b00000000000000001110101011110001;
assign LUT_1[32254] = 32'b00000000000000010001001000000110;
assign LUT_1[32255] = 32'b00000000000000001010011010000010;
assign LUT_1[32256] = 32'b00000000000000000010011000101110;
assign LUT_1[32257] = 32'b11111111111111111011101010101010;
assign LUT_1[32258] = 32'b11111111111111111110000110111111;
assign LUT_1[32259] = 32'b11111111111111110111011000111011;
assign LUT_1[32260] = 32'b00000000000000001010010010000101;
assign LUT_1[32261] = 32'b00000000000000000011100100000001;
assign LUT_1[32262] = 32'b00000000000000000110000000010110;
assign LUT_1[32263] = 32'b11111111111111111111010010010010;
assign LUT_1[32264] = 32'b00000000000000000001100110100011;
assign LUT_1[32265] = 32'b11111111111111111010111000011111;
assign LUT_1[32266] = 32'b11111111111111111101010100110100;
assign LUT_1[32267] = 32'b11111111111111110110100110110000;
assign LUT_1[32268] = 32'b00000000000000001001011111111010;
assign LUT_1[32269] = 32'b00000000000000000010110001110110;
assign LUT_1[32270] = 32'b00000000000000000101001110001011;
assign LUT_1[32271] = 32'b11111111111111111110100000000111;
assign LUT_1[32272] = 32'b00000000000000000100010100010000;
assign LUT_1[32273] = 32'b11111111111111111101100110001100;
assign LUT_1[32274] = 32'b00000000000000000000000010100001;
assign LUT_1[32275] = 32'b11111111111111111001010100011101;
assign LUT_1[32276] = 32'b00000000000000001100001101100111;
assign LUT_1[32277] = 32'b00000000000000000101011111100011;
assign LUT_1[32278] = 32'b00000000000000000111111011111000;
assign LUT_1[32279] = 32'b00000000000000000001001101110100;
assign LUT_1[32280] = 32'b00000000000000000011100010000101;
assign LUT_1[32281] = 32'b11111111111111111100110100000001;
assign LUT_1[32282] = 32'b11111111111111111111010000010110;
assign LUT_1[32283] = 32'b11111111111111111000100010010010;
assign LUT_1[32284] = 32'b00000000000000001011011011011100;
assign LUT_1[32285] = 32'b00000000000000000100101101011000;
assign LUT_1[32286] = 32'b00000000000000000111001001101101;
assign LUT_1[32287] = 32'b00000000000000000000011011101001;
assign LUT_1[32288] = 32'b00000000000000000011010011101101;
assign LUT_1[32289] = 32'b11111111111111111100100101101001;
assign LUT_1[32290] = 32'b11111111111111111111000001111110;
assign LUT_1[32291] = 32'b11111111111111111000010011111010;
assign LUT_1[32292] = 32'b00000000000000001011001101000100;
assign LUT_1[32293] = 32'b00000000000000000100011111000000;
assign LUT_1[32294] = 32'b00000000000000000110111011010101;
assign LUT_1[32295] = 32'b00000000000000000000001101010001;
assign LUT_1[32296] = 32'b00000000000000000010100001100010;
assign LUT_1[32297] = 32'b11111111111111111011110011011110;
assign LUT_1[32298] = 32'b11111111111111111110001111110011;
assign LUT_1[32299] = 32'b11111111111111110111100001101111;
assign LUT_1[32300] = 32'b00000000000000001010011010111001;
assign LUT_1[32301] = 32'b00000000000000000011101100110101;
assign LUT_1[32302] = 32'b00000000000000000110001001001010;
assign LUT_1[32303] = 32'b11111111111111111111011011000110;
assign LUT_1[32304] = 32'b00000000000000000101001111001111;
assign LUT_1[32305] = 32'b11111111111111111110100001001011;
assign LUT_1[32306] = 32'b00000000000000000000111101100000;
assign LUT_1[32307] = 32'b11111111111111111010001111011100;
assign LUT_1[32308] = 32'b00000000000000001101001000100110;
assign LUT_1[32309] = 32'b00000000000000000110011010100010;
assign LUT_1[32310] = 32'b00000000000000001000110110110111;
assign LUT_1[32311] = 32'b00000000000000000010001000110011;
assign LUT_1[32312] = 32'b00000000000000000100011101000100;
assign LUT_1[32313] = 32'b11111111111111111101101111000000;
assign LUT_1[32314] = 32'b00000000000000000000001011010101;
assign LUT_1[32315] = 32'b11111111111111111001011101010001;
assign LUT_1[32316] = 32'b00000000000000001100010110011011;
assign LUT_1[32317] = 32'b00000000000000000101101000010111;
assign LUT_1[32318] = 32'b00000000000000001000000100101100;
assign LUT_1[32319] = 32'b00000000000000000001010110101000;
assign LUT_1[32320] = 32'b00000000000000000100010110010110;
assign LUT_1[32321] = 32'b11111111111111111101101000010010;
assign LUT_1[32322] = 32'b00000000000000000000000100100111;
assign LUT_1[32323] = 32'b11111111111111111001010110100011;
assign LUT_1[32324] = 32'b00000000000000001100001111101101;
assign LUT_1[32325] = 32'b00000000000000000101100001101001;
assign LUT_1[32326] = 32'b00000000000000000111111101111110;
assign LUT_1[32327] = 32'b00000000000000000001001111111010;
assign LUT_1[32328] = 32'b00000000000000000011100100001011;
assign LUT_1[32329] = 32'b11111111111111111100110110000111;
assign LUT_1[32330] = 32'b11111111111111111111010010011100;
assign LUT_1[32331] = 32'b11111111111111111000100100011000;
assign LUT_1[32332] = 32'b00000000000000001011011101100010;
assign LUT_1[32333] = 32'b00000000000000000100101111011110;
assign LUT_1[32334] = 32'b00000000000000000111001011110011;
assign LUT_1[32335] = 32'b00000000000000000000011101101111;
assign LUT_1[32336] = 32'b00000000000000000110010001111000;
assign LUT_1[32337] = 32'b11111111111111111111100011110100;
assign LUT_1[32338] = 32'b00000000000000000010000000001001;
assign LUT_1[32339] = 32'b11111111111111111011010010000101;
assign LUT_1[32340] = 32'b00000000000000001110001011001111;
assign LUT_1[32341] = 32'b00000000000000000111011101001011;
assign LUT_1[32342] = 32'b00000000000000001001111001100000;
assign LUT_1[32343] = 32'b00000000000000000011001011011100;
assign LUT_1[32344] = 32'b00000000000000000101011111101101;
assign LUT_1[32345] = 32'b11111111111111111110110001101001;
assign LUT_1[32346] = 32'b00000000000000000001001101111110;
assign LUT_1[32347] = 32'b11111111111111111010011111111010;
assign LUT_1[32348] = 32'b00000000000000001101011001000100;
assign LUT_1[32349] = 32'b00000000000000000110101011000000;
assign LUT_1[32350] = 32'b00000000000000001001000111010101;
assign LUT_1[32351] = 32'b00000000000000000010011001010001;
assign LUT_1[32352] = 32'b00000000000000000101010001010101;
assign LUT_1[32353] = 32'b11111111111111111110100011010001;
assign LUT_1[32354] = 32'b00000000000000000000111111100110;
assign LUT_1[32355] = 32'b11111111111111111010010001100010;
assign LUT_1[32356] = 32'b00000000000000001101001010101100;
assign LUT_1[32357] = 32'b00000000000000000110011100101000;
assign LUT_1[32358] = 32'b00000000000000001000111000111101;
assign LUT_1[32359] = 32'b00000000000000000010001010111001;
assign LUT_1[32360] = 32'b00000000000000000100011111001010;
assign LUT_1[32361] = 32'b11111111111111111101110001000110;
assign LUT_1[32362] = 32'b00000000000000000000001101011011;
assign LUT_1[32363] = 32'b11111111111111111001011111010111;
assign LUT_1[32364] = 32'b00000000000000001100011000100001;
assign LUT_1[32365] = 32'b00000000000000000101101010011101;
assign LUT_1[32366] = 32'b00000000000000001000000110110010;
assign LUT_1[32367] = 32'b00000000000000000001011000101110;
assign LUT_1[32368] = 32'b00000000000000000111001100110111;
assign LUT_1[32369] = 32'b00000000000000000000011110110011;
assign LUT_1[32370] = 32'b00000000000000000010111011001000;
assign LUT_1[32371] = 32'b11111111111111111100001101000100;
assign LUT_1[32372] = 32'b00000000000000001111000110001110;
assign LUT_1[32373] = 32'b00000000000000001000011000001010;
assign LUT_1[32374] = 32'b00000000000000001010110100011111;
assign LUT_1[32375] = 32'b00000000000000000100000110011011;
assign LUT_1[32376] = 32'b00000000000000000110011010101100;
assign LUT_1[32377] = 32'b11111111111111111111101100101000;
assign LUT_1[32378] = 32'b00000000000000000010001000111101;
assign LUT_1[32379] = 32'b11111111111111111011011010111001;
assign LUT_1[32380] = 32'b00000000000000001110010100000011;
assign LUT_1[32381] = 32'b00000000000000000111100101111111;
assign LUT_1[32382] = 32'b00000000000000001010000010010100;
assign LUT_1[32383] = 32'b00000000000000000011010100010000;
assign LUT_1[32384] = 32'b00000000000000000101011000110001;
assign LUT_1[32385] = 32'b11111111111111111110101010101101;
assign LUT_1[32386] = 32'b00000000000000000001000111000010;
assign LUT_1[32387] = 32'b11111111111111111010011000111110;
assign LUT_1[32388] = 32'b00000000000000001101010010001000;
assign LUT_1[32389] = 32'b00000000000000000110100100000100;
assign LUT_1[32390] = 32'b00000000000000001001000000011001;
assign LUT_1[32391] = 32'b00000000000000000010010010010101;
assign LUT_1[32392] = 32'b00000000000000000100100110100110;
assign LUT_1[32393] = 32'b11111111111111111101111000100010;
assign LUT_1[32394] = 32'b00000000000000000000010100110111;
assign LUT_1[32395] = 32'b11111111111111111001100110110011;
assign LUT_1[32396] = 32'b00000000000000001100011111111101;
assign LUT_1[32397] = 32'b00000000000000000101110001111001;
assign LUT_1[32398] = 32'b00000000000000001000001110001110;
assign LUT_1[32399] = 32'b00000000000000000001100000001010;
assign LUT_1[32400] = 32'b00000000000000000111010100010011;
assign LUT_1[32401] = 32'b00000000000000000000100110001111;
assign LUT_1[32402] = 32'b00000000000000000011000010100100;
assign LUT_1[32403] = 32'b11111111111111111100010100100000;
assign LUT_1[32404] = 32'b00000000000000001111001101101010;
assign LUT_1[32405] = 32'b00000000000000001000011111100110;
assign LUT_1[32406] = 32'b00000000000000001010111011111011;
assign LUT_1[32407] = 32'b00000000000000000100001101110111;
assign LUT_1[32408] = 32'b00000000000000000110100010001000;
assign LUT_1[32409] = 32'b11111111111111111111110100000100;
assign LUT_1[32410] = 32'b00000000000000000010010000011001;
assign LUT_1[32411] = 32'b11111111111111111011100010010101;
assign LUT_1[32412] = 32'b00000000000000001110011011011111;
assign LUT_1[32413] = 32'b00000000000000000111101101011011;
assign LUT_1[32414] = 32'b00000000000000001010001001110000;
assign LUT_1[32415] = 32'b00000000000000000011011011101100;
assign LUT_1[32416] = 32'b00000000000000000110010011110000;
assign LUT_1[32417] = 32'b11111111111111111111100101101100;
assign LUT_1[32418] = 32'b00000000000000000010000010000001;
assign LUT_1[32419] = 32'b11111111111111111011010011111101;
assign LUT_1[32420] = 32'b00000000000000001110001101000111;
assign LUT_1[32421] = 32'b00000000000000000111011111000011;
assign LUT_1[32422] = 32'b00000000000000001001111011011000;
assign LUT_1[32423] = 32'b00000000000000000011001101010100;
assign LUT_1[32424] = 32'b00000000000000000101100001100101;
assign LUT_1[32425] = 32'b11111111111111111110110011100001;
assign LUT_1[32426] = 32'b00000000000000000001001111110110;
assign LUT_1[32427] = 32'b11111111111111111010100001110010;
assign LUT_1[32428] = 32'b00000000000000001101011010111100;
assign LUT_1[32429] = 32'b00000000000000000110101100111000;
assign LUT_1[32430] = 32'b00000000000000001001001001001101;
assign LUT_1[32431] = 32'b00000000000000000010011011001001;
assign LUT_1[32432] = 32'b00000000000000001000001111010010;
assign LUT_1[32433] = 32'b00000000000000000001100001001110;
assign LUT_1[32434] = 32'b00000000000000000011111101100011;
assign LUT_1[32435] = 32'b11111111111111111101001111011111;
assign LUT_1[32436] = 32'b00000000000000010000001000101001;
assign LUT_1[32437] = 32'b00000000000000001001011010100101;
assign LUT_1[32438] = 32'b00000000000000001011110110111010;
assign LUT_1[32439] = 32'b00000000000000000101001000110110;
assign LUT_1[32440] = 32'b00000000000000000111011101000111;
assign LUT_1[32441] = 32'b00000000000000000000101111000011;
assign LUT_1[32442] = 32'b00000000000000000011001011011000;
assign LUT_1[32443] = 32'b11111111111111111100011101010100;
assign LUT_1[32444] = 32'b00000000000000001111010110011110;
assign LUT_1[32445] = 32'b00000000000000001000101000011010;
assign LUT_1[32446] = 32'b00000000000000001011000100101111;
assign LUT_1[32447] = 32'b00000000000000000100010110101011;
assign LUT_1[32448] = 32'b00000000000000000111010110011001;
assign LUT_1[32449] = 32'b00000000000000000000101000010101;
assign LUT_1[32450] = 32'b00000000000000000011000100101010;
assign LUT_1[32451] = 32'b11111111111111111100010110100110;
assign LUT_1[32452] = 32'b00000000000000001111001111110000;
assign LUT_1[32453] = 32'b00000000000000001000100001101100;
assign LUT_1[32454] = 32'b00000000000000001010111110000001;
assign LUT_1[32455] = 32'b00000000000000000100001111111101;
assign LUT_1[32456] = 32'b00000000000000000110100100001110;
assign LUT_1[32457] = 32'b11111111111111111111110110001010;
assign LUT_1[32458] = 32'b00000000000000000010010010011111;
assign LUT_1[32459] = 32'b11111111111111111011100100011011;
assign LUT_1[32460] = 32'b00000000000000001110011101100101;
assign LUT_1[32461] = 32'b00000000000000000111101111100001;
assign LUT_1[32462] = 32'b00000000000000001010001011110110;
assign LUT_1[32463] = 32'b00000000000000000011011101110010;
assign LUT_1[32464] = 32'b00000000000000001001010001111011;
assign LUT_1[32465] = 32'b00000000000000000010100011110111;
assign LUT_1[32466] = 32'b00000000000000000101000000001100;
assign LUT_1[32467] = 32'b11111111111111111110010010001000;
assign LUT_1[32468] = 32'b00000000000000010001001011010010;
assign LUT_1[32469] = 32'b00000000000000001010011101001110;
assign LUT_1[32470] = 32'b00000000000000001100111001100011;
assign LUT_1[32471] = 32'b00000000000000000110001011011111;
assign LUT_1[32472] = 32'b00000000000000001000011111110000;
assign LUT_1[32473] = 32'b00000000000000000001110001101100;
assign LUT_1[32474] = 32'b00000000000000000100001110000001;
assign LUT_1[32475] = 32'b11111111111111111101011111111101;
assign LUT_1[32476] = 32'b00000000000000010000011001000111;
assign LUT_1[32477] = 32'b00000000000000001001101011000011;
assign LUT_1[32478] = 32'b00000000000000001100000111011000;
assign LUT_1[32479] = 32'b00000000000000000101011001010100;
assign LUT_1[32480] = 32'b00000000000000001000010001011000;
assign LUT_1[32481] = 32'b00000000000000000001100011010100;
assign LUT_1[32482] = 32'b00000000000000000011111111101001;
assign LUT_1[32483] = 32'b11111111111111111101010001100101;
assign LUT_1[32484] = 32'b00000000000000010000001010101111;
assign LUT_1[32485] = 32'b00000000000000001001011100101011;
assign LUT_1[32486] = 32'b00000000000000001011111001000000;
assign LUT_1[32487] = 32'b00000000000000000101001010111100;
assign LUT_1[32488] = 32'b00000000000000000111011111001101;
assign LUT_1[32489] = 32'b00000000000000000000110001001001;
assign LUT_1[32490] = 32'b00000000000000000011001101011110;
assign LUT_1[32491] = 32'b11111111111111111100011111011010;
assign LUT_1[32492] = 32'b00000000000000001111011000100100;
assign LUT_1[32493] = 32'b00000000000000001000101010100000;
assign LUT_1[32494] = 32'b00000000000000001011000110110101;
assign LUT_1[32495] = 32'b00000000000000000100011000110001;
assign LUT_1[32496] = 32'b00000000000000001010001100111010;
assign LUT_1[32497] = 32'b00000000000000000011011110110110;
assign LUT_1[32498] = 32'b00000000000000000101111011001011;
assign LUT_1[32499] = 32'b11111111111111111111001101000111;
assign LUT_1[32500] = 32'b00000000000000010010000110010001;
assign LUT_1[32501] = 32'b00000000000000001011011000001101;
assign LUT_1[32502] = 32'b00000000000000001101110100100010;
assign LUT_1[32503] = 32'b00000000000000000111000110011110;
assign LUT_1[32504] = 32'b00000000000000001001011010101111;
assign LUT_1[32505] = 32'b00000000000000000010101100101011;
assign LUT_1[32506] = 32'b00000000000000000101001001000000;
assign LUT_1[32507] = 32'b11111111111111111110011010111100;
assign LUT_1[32508] = 32'b00000000000000010001010100000110;
assign LUT_1[32509] = 32'b00000000000000001010100110000010;
assign LUT_1[32510] = 32'b00000000000000001101000010010111;
assign LUT_1[32511] = 32'b00000000000000000110010100010011;
assign LUT_1[32512] = 32'b00000000000000000000001100111010;
assign LUT_1[32513] = 32'b11111111111111111001011110110110;
assign LUT_1[32514] = 32'b11111111111111111011111011001011;
assign LUT_1[32515] = 32'b11111111111111110101001101000111;
assign LUT_1[32516] = 32'b00000000000000001000000110010001;
assign LUT_1[32517] = 32'b00000000000000000001011000001101;
assign LUT_1[32518] = 32'b00000000000000000011110100100010;
assign LUT_1[32519] = 32'b11111111111111111101000110011110;
assign LUT_1[32520] = 32'b11111111111111111111011010101111;
assign LUT_1[32521] = 32'b11111111111111111000101100101011;
assign LUT_1[32522] = 32'b11111111111111111011001001000000;
assign LUT_1[32523] = 32'b11111111111111110100011010111100;
assign LUT_1[32524] = 32'b00000000000000000111010100000110;
assign LUT_1[32525] = 32'b00000000000000000000100110000010;
assign LUT_1[32526] = 32'b00000000000000000011000010010111;
assign LUT_1[32527] = 32'b11111111111111111100010100010011;
assign LUT_1[32528] = 32'b00000000000000000010001000011100;
assign LUT_1[32529] = 32'b11111111111111111011011010011000;
assign LUT_1[32530] = 32'b11111111111111111101110110101101;
assign LUT_1[32531] = 32'b11111111111111110111001000101001;
assign LUT_1[32532] = 32'b00000000000000001010000001110011;
assign LUT_1[32533] = 32'b00000000000000000011010011101111;
assign LUT_1[32534] = 32'b00000000000000000101110000000100;
assign LUT_1[32535] = 32'b11111111111111111111000010000000;
assign LUT_1[32536] = 32'b00000000000000000001010110010001;
assign LUT_1[32537] = 32'b11111111111111111010101000001101;
assign LUT_1[32538] = 32'b11111111111111111101000100100010;
assign LUT_1[32539] = 32'b11111111111111110110010110011110;
assign LUT_1[32540] = 32'b00000000000000001001001111101000;
assign LUT_1[32541] = 32'b00000000000000000010100001100100;
assign LUT_1[32542] = 32'b00000000000000000100111101111001;
assign LUT_1[32543] = 32'b11111111111111111110001111110101;
assign LUT_1[32544] = 32'b00000000000000000001000111111001;
assign LUT_1[32545] = 32'b11111111111111111010011001110101;
assign LUT_1[32546] = 32'b11111111111111111100110110001010;
assign LUT_1[32547] = 32'b11111111111111110110001000000110;
assign LUT_1[32548] = 32'b00000000000000001001000001010000;
assign LUT_1[32549] = 32'b00000000000000000010010011001100;
assign LUT_1[32550] = 32'b00000000000000000100101111100001;
assign LUT_1[32551] = 32'b11111111111111111110000001011101;
assign LUT_1[32552] = 32'b00000000000000000000010101101110;
assign LUT_1[32553] = 32'b11111111111111111001100111101010;
assign LUT_1[32554] = 32'b11111111111111111100000011111111;
assign LUT_1[32555] = 32'b11111111111111110101010101111011;
assign LUT_1[32556] = 32'b00000000000000001000001111000101;
assign LUT_1[32557] = 32'b00000000000000000001100001000001;
assign LUT_1[32558] = 32'b00000000000000000011111101010110;
assign LUT_1[32559] = 32'b11111111111111111101001111010010;
assign LUT_1[32560] = 32'b00000000000000000011000011011011;
assign LUT_1[32561] = 32'b11111111111111111100010101010111;
assign LUT_1[32562] = 32'b11111111111111111110110001101100;
assign LUT_1[32563] = 32'b11111111111111111000000011101000;
assign LUT_1[32564] = 32'b00000000000000001010111100110010;
assign LUT_1[32565] = 32'b00000000000000000100001110101110;
assign LUT_1[32566] = 32'b00000000000000000110101011000011;
assign LUT_1[32567] = 32'b11111111111111111111111100111111;
assign LUT_1[32568] = 32'b00000000000000000010010001010000;
assign LUT_1[32569] = 32'b11111111111111111011100011001100;
assign LUT_1[32570] = 32'b11111111111111111101111111100001;
assign LUT_1[32571] = 32'b11111111111111110111010001011101;
assign LUT_1[32572] = 32'b00000000000000001010001010100111;
assign LUT_1[32573] = 32'b00000000000000000011011100100011;
assign LUT_1[32574] = 32'b00000000000000000101111000111000;
assign LUT_1[32575] = 32'b11111111111111111111001010110100;
assign LUT_1[32576] = 32'b00000000000000000010001010100010;
assign LUT_1[32577] = 32'b11111111111111111011011100011110;
assign LUT_1[32578] = 32'b11111111111111111101111000110011;
assign LUT_1[32579] = 32'b11111111111111110111001010101111;
assign LUT_1[32580] = 32'b00000000000000001010000011111001;
assign LUT_1[32581] = 32'b00000000000000000011010101110101;
assign LUT_1[32582] = 32'b00000000000000000101110010001010;
assign LUT_1[32583] = 32'b11111111111111111111000100000110;
assign LUT_1[32584] = 32'b00000000000000000001011000010111;
assign LUT_1[32585] = 32'b11111111111111111010101010010011;
assign LUT_1[32586] = 32'b11111111111111111101000110101000;
assign LUT_1[32587] = 32'b11111111111111110110011000100100;
assign LUT_1[32588] = 32'b00000000000000001001010001101110;
assign LUT_1[32589] = 32'b00000000000000000010100011101010;
assign LUT_1[32590] = 32'b00000000000000000100111111111111;
assign LUT_1[32591] = 32'b11111111111111111110010001111011;
assign LUT_1[32592] = 32'b00000000000000000100000110000100;
assign LUT_1[32593] = 32'b11111111111111111101011000000000;
assign LUT_1[32594] = 32'b11111111111111111111110100010101;
assign LUT_1[32595] = 32'b11111111111111111001000110010001;
assign LUT_1[32596] = 32'b00000000000000001011111111011011;
assign LUT_1[32597] = 32'b00000000000000000101010001010111;
assign LUT_1[32598] = 32'b00000000000000000111101101101100;
assign LUT_1[32599] = 32'b00000000000000000000111111101000;
assign LUT_1[32600] = 32'b00000000000000000011010011111001;
assign LUT_1[32601] = 32'b11111111111111111100100101110101;
assign LUT_1[32602] = 32'b11111111111111111111000010001010;
assign LUT_1[32603] = 32'b11111111111111111000010100000110;
assign LUT_1[32604] = 32'b00000000000000001011001101010000;
assign LUT_1[32605] = 32'b00000000000000000100011111001100;
assign LUT_1[32606] = 32'b00000000000000000110111011100001;
assign LUT_1[32607] = 32'b00000000000000000000001101011101;
assign LUT_1[32608] = 32'b00000000000000000011000101100001;
assign LUT_1[32609] = 32'b11111111111111111100010111011101;
assign LUT_1[32610] = 32'b11111111111111111110110011110010;
assign LUT_1[32611] = 32'b11111111111111111000000101101110;
assign LUT_1[32612] = 32'b00000000000000001010111110111000;
assign LUT_1[32613] = 32'b00000000000000000100010000110100;
assign LUT_1[32614] = 32'b00000000000000000110101101001001;
assign LUT_1[32615] = 32'b11111111111111111111111111000101;
assign LUT_1[32616] = 32'b00000000000000000010010011010110;
assign LUT_1[32617] = 32'b11111111111111111011100101010010;
assign LUT_1[32618] = 32'b11111111111111111110000001100111;
assign LUT_1[32619] = 32'b11111111111111110111010011100011;
assign LUT_1[32620] = 32'b00000000000000001010001100101101;
assign LUT_1[32621] = 32'b00000000000000000011011110101001;
assign LUT_1[32622] = 32'b00000000000000000101111010111110;
assign LUT_1[32623] = 32'b11111111111111111111001100111010;
assign LUT_1[32624] = 32'b00000000000000000101000001000011;
assign LUT_1[32625] = 32'b11111111111111111110010010111111;
assign LUT_1[32626] = 32'b00000000000000000000101111010100;
assign LUT_1[32627] = 32'b11111111111111111010000001010000;
assign LUT_1[32628] = 32'b00000000000000001100111010011010;
assign LUT_1[32629] = 32'b00000000000000000110001100010110;
assign LUT_1[32630] = 32'b00000000000000001000101000101011;
assign LUT_1[32631] = 32'b00000000000000000001111010100111;
assign LUT_1[32632] = 32'b00000000000000000100001110111000;
assign LUT_1[32633] = 32'b11111111111111111101100000110100;
assign LUT_1[32634] = 32'b11111111111111111111111101001001;
assign LUT_1[32635] = 32'b11111111111111111001001111000101;
assign LUT_1[32636] = 32'b00000000000000001100001000001111;
assign LUT_1[32637] = 32'b00000000000000000101011010001011;
assign LUT_1[32638] = 32'b00000000000000000111110110100000;
assign LUT_1[32639] = 32'b00000000000000000001001000011100;
assign LUT_1[32640] = 32'b00000000000000000011001100111101;
assign LUT_1[32641] = 32'b11111111111111111100011110111001;
assign LUT_1[32642] = 32'b11111111111111111110111011001110;
assign LUT_1[32643] = 32'b11111111111111111000001101001010;
assign LUT_1[32644] = 32'b00000000000000001011000110010100;
assign LUT_1[32645] = 32'b00000000000000000100011000010000;
assign LUT_1[32646] = 32'b00000000000000000110110100100101;
assign LUT_1[32647] = 32'b00000000000000000000000110100001;
assign LUT_1[32648] = 32'b00000000000000000010011010110010;
assign LUT_1[32649] = 32'b11111111111111111011101100101110;
assign LUT_1[32650] = 32'b11111111111111111110001001000011;
assign LUT_1[32651] = 32'b11111111111111110111011010111111;
assign LUT_1[32652] = 32'b00000000000000001010010100001001;
assign LUT_1[32653] = 32'b00000000000000000011100110000101;
assign LUT_1[32654] = 32'b00000000000000000110000010011010;
assign LUT_1[32655] = 32'b11111111111111111111010100010110;
assign LUT_1[32656] = 32'b00000000000000000101001000011111;
assign LUT_1[32657] = 32'b11111111111111111110011010011011;
assign LUT_1[32658] = 32'b00000000000000000000110110110000;
assign LUT_1[32659] = 32'b11111111111111111010001000101100;
assign LUT_1[32660] = 32'b00000000000000001101000001110110;
assign LUT_1[32661] = 32'b00000000000000000110010011110010;
assign LUT_1[32662] = 32'b00000000000000001000110000000111;
assign LUT_1[32663] = 32'b00000000000000000010000010000011;
assign LUT_1[32664] = 32'b00000000000000000100010110010100;
assign LUT_1[32665] = 32'b11111111111111111101101000010000;
assign LUT_1[32666] = 32'b00000000000000000000000100100101;
assign LUT_1[32667] = 32'b11111111111111111001010110100001;
assign LUT_1[32668] = 32'b00000000000000001100001111101011;
assign LUT_1[32669] = 32'b00000000000000000101100001100111;
assign LUT_1[32670] = 32'b00000000000000000111111101111100;
assign LUT_1[32671] = 32'b00000000000000000001001111111000;
assign LUT_1[32672] = 32'b00000000000000000100000111111100;
assign LUT_1[32673] = 32'b11111111111111111101011001111000;
assign LUT_1[32674] = 32'b11111111111111111111110110001101;
assign LUT_1[32675] = 32'b11111111111111111001001000001001;
assign LUT_1[32676] = 32'b00000000000000001100000001010011;
assign LUT_1[32677] = 32'b00000000000000000101010011001111;
assign LUT_1[32678] = 32'b00000000000000000111101111100100;
assign LUT_1[32679] = 32'b00000000000000000001000001100000;
assign LUT_1[32680] = 32'b00000000000000000011010101110001;
assign LUT_1[32681] = 32'b11111111111111111100100111101101;
assign LUT_1[32682] = 32'b11111111111111111111000100000010;
assign LUT_1[32683] = 32'b11111111111111111000010101111110;
assign LUT_1[32684] = 32'b00000000000000001011001111001000;
assign LUT_1[32685] = 32'b00000000000000000100100001000100;
assign LUT_1[32686] = 32'b00000000000000000110111101011001;
assign LUT_1[32687] = 32'b00000000000000000000001111010101;
assign LUT_1[32688] = 32'b00000000000000000110000011011110;
assign LUT_1[32689] = 32'b11111111111111111111010101011010;
assign LUT_1[32690] = 32'b00000000000000000001110001101111;
assign LUT_1[32691] = 32'b11111111111111111011000011101011;
assign LUT_1[32692] = 32'b00000000000000001101111100110101;
assign LUT_1[32693] = 32'b00000000000000000111001110110001;
assign LUT_1[32694] = 32'b00000000000000001001101011000110;
assign LUT_1[32695] = 32'b00000000000000000010111101000010;
assign LUT_1[32696] = 32'b00000000000000000101010001010011;
assign LUT_1[32697] = 32'b11111111111111111110100011001111;
assign LUT_1[32698] = 32'b00000000000000000000111111100100;
assign LUT_1[32699] = 32'b11111111111111111010010001100000;
assign LUT_1[32700] = 32'b00000000000000001101001010101010;
assign LUT_1[32701] = 32'b00000000000000000110011100100110;
assign LUT_1[32702] = 32'b00000000000000001000111000111011;
assign LUT_1[32703] = 32'b00000000000000000010001010110111;
assign LUT_1[32704] = 32'b00000000000000000101001010100101;
assign LUT_1[32705] = 32'b11111111111111111110011100100001;
assign LUT_1[32706] = 32'b00000000000000000000111000110110;
assign LUT_1[32707] = 32'b11111111111111111010001010110010;
assign LUT_1[32708] = 32'b00000000000000001101000011111100;
assign LUT_1[32709] = 32'b00000000000000000110010101111000;
assign LUT_1[32710] = 32'b00000000000000001000110010001101;
assign LUT_1[32711] = 32'b00000000000000000010000100001001;
assign LUT_1[32712] = 32'b00000000000000000100011000011010;
assign LUT_1[32713] = 32'b11111111111111111101101010010110;
assign LUT_1[32714] = 32'b00000000000000000000000110101011;
assign LUT_1[32715] = 32'b11111111111111111001011000100111;
assign LUT_1[32716] = 32'b00000000000000001100010001110001;
assign LUT_1[32717] = 32'b00000000000000000101100011101101;
assign LUT_1[32718] = 32'b00000000000000001000000000000010;
assign LUT_1[32719] = 32'b00000000000000000001010001111110;
assign LUT_1[32720] = 32'b00000000000000000111000110000111;
assign LUT_1[32721] = 32'b00000000000000000000011000000011;
assign LUT_1[32722] = 32'b00000000000000000010110100011000;
assign LUT_1[32723] = 32'b11111111111111111100000110010100;
assign LUT_1[32724] = 32'b00000000000000001110111111011110;
assign LUT_1[32725] = 32'b00000000000000001000010001011010;
assign LUT_1[32726] = 32'b00000000000000001010101101101111;
assign LUT_1[32727] = 32'b00000000000000000011111111101011;
assign LUT_1[32728] = 32'b00000000000000000110010011111100;
assign LUT_1[32729] = 32'b11111111111111111111100101111000;
assign LUT_1[32730] = 32'b00000000000000000010000010001101;
assign LUT_1[32731] = 32'b11111111111111111011010100001001;
assign LUT_1[32732] = 32'b00000000000000001110001101010011;
assign LUT_1[32733] = 32'b00000000000000000111011111001111;
assign LUT_1[32734] = 32'b00000000000000001001111011100100;
assign LUT_1[32735] = 32'b00000000000000000011001101100000;
assign LUT_1[32736] = 32'b00000000000000000110000101100100;
assign LUT_1[32737] = 32'b11111111111111111111010111100000;
assign LUT_1[32738] = 32'b00000000000000000001110011110101;
assign LUT_1[32739] = 32'b11111111111111111011000101110001;
assign LUT_1[32740] = 32'b00000000000000001101111110111011;
assign LUT_1[32741] = 32'b00000000000000000111010000110111;
assign LUT_1[32742] = 32'b00000000000000001001101101001100;
assign LUT_1[32743] = 32'b00000000000000000010111111001000;
assign LUT_1[32744] = 32'b00000000000000000101010011011001;
assign LUT_1[32745] = 32'b11111111111111111110100101010101;
assign LUT_1[32746] = 32'b00000000000000000001000001101010;
assign LUT_1[32747] = 32'b11111111111111111010010011100110;
assign LUT_1[32748] = 32'b00000000000000001101001100110000;
assign LUT_1[32749] = 32'b00000000000000000110011110101100;
assign LUT_1[32750] = 32'b00000000000000001000111011000001;
assign LUT_1[32751] = 32'b00000000000000000010001100111101;
assign LUT_1[32752] = 32'b00000000000000001000000001000110;
assign LUT_1[32753] = 32'b00000000000000000001010011000010;
assign LUT_1[32754] = 32'b00000000000000000011101111010111;
assign LUT_1[32755] = 32'b11111111111111111101000001010011;
assign LUT_1[32756] = 32'b00000000000000001111111010011101;
assign LUT_1[32757] = 32'b00000000000000001001001100011001;
assign LUT_1[32758] = 32'b00000000000000001011101000101110;
assign LUT_1[32759] = 32'b00000000000000000100111010101010;
assign LUT_1[32760] = 32'b00000000000000000111001110111011;
assign LUT_1[32761] = 32'b00000000000000000000100000110111;
assign LUT_1[32762] = 32'b00000000000000000010111101001100;
assign LUT_1[32763] = 32'b11111111111111111100001111001000;
assign LUT_1[32764] = 32'b00000000000000001111001000010010;
assign LUT_1[32765] = 32'b00000000000000001000011010001110;
assign LUT_1[32766] = 32'b00000000000000001010110110100011;
assign LUT_1[32767] = 32'b00000000000000000100001000011111;
assign LUT_1[32768] = 32'b00000000000000000000110110010100;
assign LUT_1[32769] = 32'b11111111111111111010001000010000;
assign LUT_1[32770] = 32'b11111111111111111100100100100101;
assign LUT_1[32771] = 32'b11111111111111110101110110100001;
assign LUT_1[32772] = 32'b00000000000000001000101111101011;
assign LUT_1[32773] = 32'b00000000000000000010000001100111;
assign LUT_1[32774] = 32'b00000000000000000100011101111100;
assign LUT_1[32775] = 32'b11111111111111111101101111111000;
assign LUT_1[32776] = 32'b00000000000000000000000100001001;
assign LUT_1[32777] = 32'b11111111111111111001010110000101;
assign LUT_1[32778] = 32'b11111111111111111011110010011010;
assign LUT_1[32779] = 32'b11111111111111110101000100010110;
assign LUT_1[32780] = 32'b00000000000000000111111101100000;
assign LUT_1[32781] = 32'b00000000000000000001001111011100;
assign LUT_1[32782] = 32'b00000000000000000011101011110001;
assign LUT_1[32783] = 32'b11111111111111111100111101101101;
assign LUT_1[32784] = 32'b00000000000000000010110001110110;
assign LUT_1[32785] = 32'b11111111111111111100000011110010;
assign LUT_1[32786] = 32'b11111111111111111110100000000111;
assign LUT_1[32787] = 32'b11111111111111110111110010000011;
assign LUT_1[32788] = 32'b00000000000000001010101011001101;
assign LUT_1[32789] = 32'b00000000000000000011111101001001;
assign LUT_1[32790] = 32'b00000000000000000110011001011110;
assign LUT_1[32791] = 32'b11111111111111111111101011011010;
assign LUT_1[32792] = 32'b00000000000000000001111111101011;
assign LUT_1[32793] = 32'b11111111111111111011010001100111;
assign LUT_1[32794] = 32'b11111111111111111101101101111100;
assign LUT_1[32795] = 32'b11111111111111110110111111111000;
assign LUT_1[32796] = 32'b00000000000000001001111001000010;
assign LUT_1[32797] = 32'b00000000000000000011001010111110;
assign LUT_1[32798] = 32'b00000000000000000101100111010011;
assign LUT_1[32799] = 32'b11111111111111111110111001001111;
assign LUT_1[32800] = 32'b00000000000000000001110001010011;
assign LUT_1[32801] = 32'b11111111111111111011000011001111;
assign LUT_1[32802] = 32'b11111111111111111101011111100100;
assign LUT_1[32803] = 32'b11111111111111110110110001100000;
assign LUT_1[32804] = 32'b00000000000000001001101010101010;
assign LUT_1[32805] = 32'b00000000000000000010111100100110;
assign LUT_1[32806] = 32'b00000000000000000101011000111011;
assign LUT_1[32807] = 32'b11111111111111111110101010110111;
assign LUT_1[32808] = 32'b00000000000000000000111111001000;
assign LUT_1[32809] = 32'b11111111111111111010010001000100;
assign LUT_1[32810] = 32'b11111111111111111100101101011001;
assign LUT_1[32811] = 32'b11111111111111110101111111010101;
assign LUT_1[32812] = 32'b00000000000000001000111000011111;
assign LUT_1[32813] = 32'b00000000000000000010001010011011;
assign LUT_1[32814] = 32'b00000000000000000100100110110000;
assign LUT_1[32815] = 32'b11111111111111111101111000101100;
assign LUT_1[32816] = 32'b00000000000000000011101100110101;
assign LUT_1[32817] = 32'b11111111111111111100111110110001;
assign LUT_1[32818] = 32'b11111111111111111111011011000110;
assign LUT_1[32819] = 32'b11111111111111111000101101000010;
assign LUT_1[32820] = 32'b00000000000000001011100110001100;
assign LUT_1[32821] = 32'b00000000000000000100111000001000;
assign LUT_1[32822] = 32'b00000000000000000111010100011101;
assign LUT_1[32823] = 32'b00000000000000000000100110011001;
assign LUT_1[32824] = 32'b00000000000000000010111010101010;
assign LUT_1[32825] = 32'b11111111111111111100001100100110;
assign LUT_1[32826] = 32'b11111111111111111110101000111011;
assign LUT_1[32827] = 32'b11111111111111110111111010110111;
assign LUT_1[32828] = 32'b00000000000000001010110100000001;
assign LUT_1[32829] = 32'b00000000000000000100000101111101;
assign LUT_1[32830] = 32'b00000000000000000110100010010010;
assign LUT_1[32831] = 32'b11111111111111111111110100001110;
assign LUT_1[32832] = 32'b00000000000000000010110011111100;
assign LUT_1[32833] = 32'b11111111111111111100000101111000;
assign LUT_1[32834] = 32'b11111111111111111110100010001101;
assign LUT_1[32835] = 32'b11111111111111110111110100001001;
assign LUT_1[32836] = 32'b00000000000000001010101101010011;
assign LUT_1[32837] = 32'b00000000000000000011111111001111;
assign LUT_1[32838] = 32'b00000000000000000110011011100100;
assign LUT_1[32839] = 32'b11111111111111111111101101100000;
assign LUT_1[32840] = 32'b00000000000000000010000001110001;
assign LUT_1[32841] = 32'b11111111111111111011010011101101;
assign LUT_1[32842] = 32'b11111111111111111101110000000010;
assign LUT_1[32843] = 32'b11111111111111110111000001111110;
assign LUT_1[32844] = 32'b00000000000000001001111011001000;
assign LUT_1[32845] = 32'b00000000000000000011001101000100;
assign LUT_1[32846] = 32'b00000000000000000101101001011001;
assign LUT_1[32847] = 32'b11111111111111111110111011010101;
assign LUT_1[32848] = 32'b00000000000000000100101111011110;
assign LUT_1[32849] = 32'b11111111111111111110000001011010;
assign LUT_1[32850] = 32'b00000000000000000000011101101111;
assign LUT_1[32851] = 32'b11111111111111111001101111101011;
assign LUT_1[32852] = 32'b00000000000000001100101000110101;
assign LUT_1[32853] = 32'b00000000000000000101111010110001;
assign LUT_1[32854] = 32'b00000000000000001000010111000110;
assign LUT_1[32855] = 32'b00000000000000000001101001000010;
assign LUT_1[32856] = 32'b00000000000000000011111101010011;
assign LUT_1[32857] = 32'b11111111111111111101001111001111;
assign LUT_1[32858] = 32'b11111111111111111111101011100100;
assign LUT_1[32859] = 32'b11111111111111111000111101100000;
assign LUT_1[32860] = 32'b00000000000000001011110110101010;
assign LUT_1[32861] = 32'b00000000000000000101001000100110;
assign LUT_1[32862] = 32'b00000000000000000111100100111011;
assign LUT_1[32863] = 32'b00000000000000000000110110110111;
assign LUT_1[32864] = 32'b00000000000000000011101110111011;
assign LUT_1[32865] = 32'b11111111111111111101000000110111;
assign LUT_1[32866] = 32'b11111111111111111111011101001100;
assign LUT_1[32867] = 32'b11111111111111111000101111001000;
assign LUT_1[32868] = 32'b00000000000000001011101000010010;
assign LUT_1[32869] = 32'b00000000000000000100111010001110;
assign LUT_1[32870] = 32'b00000000000000000111010110100011;
assign LUT_1[32871] = 32'b00000000000000000000101000011111;
assign LUT_1[32872] = 32'b00000000000000000010111100110000;
assign LUT_1[32873] = 32'b11111111111111111100001110101100;
assign LUT_1[32874] = 32'b11111111111111111110101011000001;
assign LUT_1[32875] = 32'b11111111111111110111111100111101;
assign LUT_1[32876] = 32'b00000000000000001010110110000111;
assign LUT_1[32877] = 32'b00000000000000000100001000000011;
assign LUT_1[32878] = 32'b00000000000000000110100100011000;
assign LUT_1[32879] = 32'b11111111111111111111110110010100;
assign LUT_1[32880] = 32'b00000000000000000101101010011101;
assign LUT_1[32881] = 32'b11111111111111111110111100011001;
assign LUT_1[32882] = 32'b00000000000000000001011000101110;
assign LUT_1[32883] = 32'b11111111111111111010101010101010;
assign LUT_1[32884] = 32'b00000000000000001101100011110100;
assign LUT_1[32885] = 32'b00000000000000000110110101110000;
assign LUT_1[32886] = 32'b00000000000000001001010010000101;
assign LUT_1[32887] = 32'b00000000000000000010100100000001;
assign LUT_1[32888] = 32'b00000000000000000100111000010010;
assign LUT_1[32889] = 32'b11111111111111111110001010001110;
assign LUT_1[32890] = 32'b00000000000000000000100110100011;
assign LUT_1[32891] = 32'b11111111111111111001111000011111;
assign LUT_1[32892] = 32'b00000000000000001100110001101001;
assign LUT_1[32893] = 32'b00000000000000000110000011100101;
assign LUT_1[32894] = 32'b00000000000000001000011111111010;
assign LUT_1[32895] = 32'b00000000000000000001110001110110;
assign LUT_1[32896] = 32'b00000000000000000011110110010111;
assign LUT_1[32897] = 32'b11111111111111111101001000010011;
assign LUT_1[32898] = 32'b11111111111111111111100100101000;
assign LUT_1[32899] = 32'b11111111111111111000110110100100;
assign LUT_1[32900] = 32'b00000000000000001011101111101110;
assign LUT_1[32901] = 32'b00000000000000000101000001101010;
assign LUT_1[32902] = 32'b00000000000000000111011101111111;
assign LUT_1[32903] = 32'b00000000000000000000101111111011;
assign LUT_1[32904] = 32'b00000000000000000011000100001100;
assign LUT_1[32905] = 32'b11111111111111111100010110001000;
assign LUT_1[32906] = 32'b11111111111111111110110010011101;
assign LUT_1[32907] = 32'b11111111111111111000000100011001;
assign LUT_1[32908] = 32'b00000000000000001010111101100011;
assign LUT_1[32909] = 32'b00000000000000000100001111011111;
assign LUT_1[32910] = 32'b00000000000000000110101011110100;
assign LUT_1[32911] = 32'b11111111111111111111111101110000;
assign LUT_1[32912] = 32'b00000000000000000101110001111001;
assign LUT_1[32913] = 32'b11111111111111111111000011110101;
assign LUT_1[32914] = 32'b00000000000000000001100000001010;
assign LUT_1[32915] = 32'b11111111111111111010110010000110;
assign LUT_1[32916] = 32'b00000000000000001101101011010000;
assign LUT_1[32917] = 32'b00000000000000000110111101001100;
assign LUT_1[32918] = 32'b00000000000000001001011001100001;
assign LUT_1[32919] = 32'b00000000000000000010101011011101;
assign LUT_1[32920] = 32'b00000000000000000100111111101110;
assign LUT_1[32921] = 32'b11111111111111111110010001101010;
assign LUT_1[32922] = 32'b00000000000000000000101101111111;
assign LUT_1[32923] = 32'b11111111111111111001111111111011;
assign LUT_1[32924] = 32'b00000000000000001100111001000101;
assign LUT_1[32925] = 32'b00000000000000000110001011000001;
assign LUT_1[32926] = 32'b00000000000000001000100111010110;
assign LUT_1[32927] = 32'b00000000000000000001111001010010;
assign LUT_1[32928] = 32'b00000000000000000100110001010110;
assign LUT_1[32929] = 32'b11111111111111111110000011010010;
assign LUT_1[32930] = 32'b00000000000000000000011111100111;
assign LUT_1[32931] = 32'b11111111111111111001110001100011;
assign LUT_1[32932] = 32'b00000000000000001100101010101101;
assign LUT_1[32933] = 32'b00000000000000000101111100101001;
assign LUT_1[32934] = 32'b00000000000000001000011000111110;
assign LUT_1[32935] = 32'b00000000000000000001101010111010;
assign LUT_1[32936] = 32'b00000000000000000011111111001011;
assign LUT_1[32937] = 32'b11111111111111111101010001000111;
assign LUT_1[32938] = 32'b11111111111111111111101101011100;
assign LUT_1[32939] = 32'b11111111111111111000111111011000;
assign LUT_1[32940] = 32'b00000000000000001011111000100010;
assign LUT_1[32941] = 32'b00000000000000000101001010011110;
assign LUT_1[32942] = 32'b00000000000000000111100110110011;
assign LUT_1[32943] = 32'b00000000000000000000111000101111;
assign LUT_1[32944] = 32'b00000000000000000110101100111000;
assign LUT_1[32945] = 32'b11111111111111111111111110110100;
assign LUT_1[32946] = 32'b00000000000000000010011011001001;
assign LUT_1[32947] = 32'b11111111111111111011101101000101;
assign LUT_1[32948] = 32'b00000000000000001110100110001111;
assign LUT_1[32949] = 32'b00000000000000000111111000001011;
assign LUT_1[32950] = 32'b00000000000000001010010100100000;
assign LUT_1[32951] = 32'b00000000000000000011100110011100;
assign LUT_1[32952] = 32'b00000000000000000101111010101101;
assign LUT_1[32953] = 32'b11111111111111111111001100101001;
assign LUT_1[32954] = 32'b00000000000000000001101000111110;
assign LUT_1[32955] = 32'b11111111111111111010111010111010;
assign LUT_1[32956] = 32'b00000000000000001101110100000100;
assign LUT_1[32957] = 32'b00000000000000000111000110000000;
assign LUT_1[32958] = 32'b00000000000000001001100010010101;
assign LUT_1[32959] = 32'b00000000000000000010110100010001;
assign LUT_1[32960] = 32'b00000000000000000101110011111111;
assign LUT_1[32961] = 32'b11111111111111111111000101111011;
assign LUT_1[32962] = 32'b00000000000000000001100010010000;
assign LUT_1[32963] = 32'b11111111111111111010110100001100;
assign LUT_1[32964] = 32'b00000000000000001101101101010110;
assign LUT_1[32965] = 32'b00000000000000000110111111010010;
assign LUT_1[32966] = 32'b00000000000000001001011011100111;
assign LUT_1[32967] = 32'b00000000000000000010101101100011;
assign LUT_1[32968] = 32'b00000000000000000101000001110100;
assign LUT_1[32969] = 32'b11111111111111111110010011110000;
assign LUT_1[32970] = 32'b00000000000000000000110000000101;
assign LUT_1[32971] = 32'b11111111111111111010000010000001;
assign LUT_1[32972] = 32'b00000000000000001100111011001011;
assign LUT_1[32973] = 32'b00000000000000000110001101000111;
assign LUT_1[32974] = 32'b00000000000000001000101001011100;
assign LUT_1[32975] = 32'b00000000000000000001111011011000;
assign LUT_1[32976] = 32'b00000000000000000111101111100001;
assign LUT_1[32977] = 32'b00000000000000000001000001011101;
assign LUT_1[32978] = 32'b00000000000000000011011101110010;
assign LUT_1[32979] = 32'b11111111111111111100101111101110;
assign LUT_1[32980] = 32'b00000000000000001111101000111000;
assign LUT_1[32981] = 32'b00000000000000001000111010110100;
assign LUT_1[32982] = 32'b00000000000000001011010111001001;
assign LUT_1[32983] = 32'b00000000000000000100101001000101;
assign LUT_1[32984] = 32'b00000000000000000110111101010110;
assign LUT_1[32985] = 32'b00000000000000000000001111010010;
assign LUT_1[32986] = 32'b00000000000000000010101011100111;
assign LUT_1[32987] = 32'b11111111111111111011111101100011;
assign LUT_1[32988] = 32'b00000000000000001110110110101101;
assign LUT_1[32989] = 32'b00000000000000001000001000101001;
assign LUT_1[32990] = 32'b00000000000000001010100100111110;
assign LUT_1[32991] = 32'b00000000000000000011110110111010;
assign LUT_1[32992] = 32'b00000000000000000110101110111110;
assign LUT_1[32993] = 32'b00000000000000000000000000111010;
assign LUT_1[32994] = 32'b00000000000000000010011101001111;
assign LUT_1[32995] = 32'b11111111111111111011101111001011;
assign LUT_1[32996] = 32'b00000000000000001110101000010101;
assign LUT_1[32997] = 32'b00000000000000000111111010010001;
assign LUT_1[32998] = 32'b00000000000000001010010110100110;
assign LUT_1[32999] = 32'b00000000000000000011101000100010;
assign LUT_1[33000] = 32'b00000000000000000101111100110011;
assign LUT_1[33001] = 32'b11111111111111111111001110101111;
assign LUT_1[33002] = 32'b00000000000000000001101011000100;
assign LUT_1[33003] = 32'b11111111111111111010111101000000;
assign LUT_1[33004] = 32'b00000000000000001101110110001010;
assign LUT_1[33005] = 32'b00000000000000000111001000000110;
assign LUT_1[33006] = 32'b00000000000000001001100100011011;
assign LUT_1[33007] = 32'b00000000000000000010110110010111;
assign LUT_1[33008] = 32'b00000000000000001000101010100000;
assign LUT_1[33009] = 32'b00000000000000000001111100011100;
assign LUT_1[33010] = 32'b00000000000000000100011000110001;
assign LUT_1[33011] = 32'b11111111111111111101101010101101;
assign LUT_1[33012] = 32'b00000000000000010000100011110111;
assign LUT_1[33013] = 32'b00000000000000001001110101110011;
assign LUT_1[33014] = 32'b00000000000000001100010010001000;
assign LUT_1[33015] = 32'b00000000000000000101100100000100;
assign LUT_1[33016] = 32'b00000000000000000111111000010101;
assign LUT_1[33017] = 32'b00000000000000000001001010010001;
assign LUT_1[33018] = 32'b00000000000000000011100110100110;
assign LUT_1[33019] = 32'b11111111111111111100111000100010;
assign LUT_1[33020] = 32'b00000000000000001111110001101100;
assign LUT_1[33021] = 32'b00000000000000001001000011101000;
assign LUT_1[33022] = 32'b00000000000000001011011111111101;
assign LUT_1[33023] = 32'b00000000000000000100110001111001;
assign LUT_1[33024] = 32'b11111111111111111110101010100000;
assign LUT_1[33025] = 32'b11111111111111110111111100011100;
assign LUT_1[33026] = 32'b11111111111111111010011000110001;
assign LUT_1[33027] = 32'b11111111111111110011101010101101;
assign LUT_1[33028] = 32'b00000000000000000110100011110111;
assign LUT_1[33029] = 32'b11111111111111111111110101110011;
assign LUT_1[33030] = 32'b00000000000000000010010010001000;
assign LUT_1[33031] = 32'b11111111111111111011100100000100;
assign LUT_1[33032] = 32'b11111111111111111101111000010101;
assign LUT_1[33033] = 32'b11111111111111110111001010010001;
assign LUT_1[33034] = 32'b11111111111111111001100110100110;
assign LUT_1[33035] = 32'b11111111111111110010111000100010;
assign LUT_1[33036] = 32'b00000000000000000101110001101100;
assign LUT_1[33037] = 32'b11111111111111111111000011101000;
assign LUT_1[33038] = 32'b00000000000000000001011111111101;
assign LUT_1[33039] = 32'b11111111111111111010110001111001;
assign LUT_1[33040] = 32'b00000000000000000000100110000010;
assign LUT_1[33041] = 32'b11111111111111111001110111111110;
assign LUT_1[33042] = 32'b11111111111111111100010100010011;
assign LUT_1[33043] = 32'b11111111111111110101100110001111;
assign LUT_1[33044] = 32'b00000000000000001000011111011001;
assign LUT_1[33045] = 32'b00000000000000000001110001010101;
assign LUT_1[33046] = 32'b00000000000000000100001101101010;
assign LUT_1[33047] = 32'b11111111111111111101011111100110;
assign LUT_1[33048] = 32'b11111111111111111111110011110111;
assign LUT_1[33049] = 32'b11111111111111111001000101110011;
assign LUT_1[33050] = 32'b11111111111111111011100010001000;
assign LUT_1[33051] = 32'b11111111111111110100110100000100;
assign LUT_1[33052] = 32'b00000000000000000111101101001110;
assign LUT_1[33053] = 32'b00000000000000000000111111001010;
assign LUT_1[33054] = 32'b00000000000000000011011011011111;
assign LUT_1[33055] = 32'b11111111111111111100101101011011;
assign LUT_1[33056] = 32'b11111111111111111111100101011111;
assign LUT_1[33057] = 32'b11111111111111111000110111011011;
assign LUT_1[33058] = 32'b11111111111111111011010011110000;
assign LUT_1[33059] = 32'b11111111111111110100100101101100;
assign LUT_1[33060] = 32'b00000000000000000111011110110110;
assign LUT_1[33061] = 32'b00000000000000000000110000110010;
assign LUT_1[33062] = 32'b00000000000000000011001101000111;
assign LUT_1[33063] = 32'b11111111111111111100011111000011;
assign LUT_1[33064] = 32'b11111111111111111110110011010100;
assign LUT_1[33065] = 32'b11111111111111111000000101010000;
assign LUT_1[33066] = 32'b11111111111111111010100001100101;
assign LUT_1[33067] = 32'b11111111111111110011110011100001;
assign LUT_1[33068] = 32'b00000000000000000110101100101011;
assign LUT_1[33069] = 32'b11111111111111111111111110100111;
assign LUT_1[33070] = 32'b00000000000000000010011010111100;
assign LUT_1[33071] = 32'b11111111111111111011101100111000;
assign LUT_1[33072] = 32'b00000000000000000001100001000001;
assign LUT_1[33073] = 32'b11111111111111111010110010111101;
assign LUT_1[33074] = 32'b11111111111111111101001111010010;
assign LUT_1[33075] = 32'b11111111111111110110100001001110;
assign LUT_1[33076] = 32'b00000000000000001001011010011000;
assign LUT_1[33077] = 32'b00000000000000000010101100010100;
assign LUT_1[33078] = 32'b00000000000000000101001000101001;
assign LUT_1[33079] = 32'b11111111111111111110011010100101;
assign LUT_1[33080] = 32'b00000000000000000000101110110110;
assign LUT_1[33081] = 32'b11111111111111111010000000110010;
assign LUT_1[33082] = 32'b11111111111111111100011101000111;
assign LUT_1[33083] = 32'b11111111111111110101101111000011;
assign LUT_1[33084] = 32'b00000000000000001000101000001101;
assign LUT_1[33085] = 32'b00000000000000000001111010001001;
assign LUT_1[33086] = 32'b00000000000000000100010110011110;
assign LUT_1[33087] = 32'b11111111111111111101101000011010;
assign LUT_1[33088] = 32'b00000000000000000000101000001000;
assign LUT_1[33089] = 32'b11111111111111111001111010000100;
assign LUT_1[33090] = 32'b11111111111111111100010110011001;
assign LUT_1[33091] = 32'b11111111111111110101101000010101;
assign LUT_1[33092] = 32'b00000000000000001000100001011111;
assign LUT_1[33093] = 32'b00000000000000000001110011011011;
assign LUT_1[33094] = 32'b00000000000000000100001111110000;
assign LUT_1[33095] = 32'b11111111111111111101100001101100;
assign LUT_1[33096] = 32'b11111111111111111111110101111101;
assign LUT_1[33097] = 32'b11111111111111111001000111111001;
assign LUT_1[33098] = 32'b11111111111111111011100100001110;
assign LUT_1[33099] = 32'b11111111111111110100110110001010;
assign LUT_1[33100] = 32'b00000000000000000111101111010100;
assign LUT_1[33101] = 32'b00000000000000000001000001010000;
assign LUT_1[33102] = 32'b00000000000000000011011101100101;
assign LUT_1[33103] = 32'b11111111111111111100101111100001;
assign LUT_1[33104] = 32'b00000000000000000010100011101010;
assign LUT_1[33105] = 32'b11111111111111111011110101100110;
assign LUT_1[33106] = 32'b11111111111111111110010001111011;
assign LUT_1[33107] = 32'b11111111111111110111100011110111;
assign LUT_1[33108] = 32'b00000000000000001010011101000001;
assign LUT_1[33109] = 32'b00000000000000000011101110111101;
assign LUT_1[33110] = 32'b00000000000000000110001011010010;
assign LUT_1[33111] = 32'b11111111111111111111011101001110;
assign LUT_1[33112] = 32'b00000000000000000001110001011111;
assign LUT_1[33113] = 32'b11111111111111111011000011011011;
assign LUT_1[33114] = 32'b11111111111111111101011111110000;
assign LUT_1[33115] = 32'b11111111111111110110110001101100;
assign LUT_1[33116] = 32'b00000000000000001001101010110110;
assign LUT_1[33117] = 32'b00000000000000000010111100110010;
assign LUT_1[33118] = 32'b00000000000000000101011001000111;
assign LUT_1[33119] = 32'b11111111111111111110101011000011;
assign LUT_1[33120] = 32'b00000000000000000001100011000111;
assign LUT_1[33121] = 32'b11111111111111111010110101000011;
assign LUT_1[33122] = 32'b11111111111111111101010001011000;
assign LUT_1[33123] = 32'b11111111111111110110100011010100;
assign LUT_1[33124] = 32'b00000000000000001001011100011110;
assign LUT_1[33125] = 32'b00000000000000000010101110011010;
assign LUT_1[33126] = 32'b00000000000000000101001010101111;
assign LUT_1[33127] = 32'b11111111111111111110011100101011;
assign LUT_1[33128] = 32'b00000000000000000000110000111100;
assign LUT_1[33129] = 32'b11111111111111111010000010111000;
assign LUT_1[33130] = 32'b11111111111111111100011111001101;
assign LUT_1[33131] = 32'b11111111111111110101110001001001;
assign LUT_1[33132] = 32'b00000000000000001000101010010011;
assign LUT_1[33133] = 32'b00000000000000000001111100001111;
assign LUT_1[33134] = 32'b00000000000000000100011000100100;
assign LUT_1[33135] = 32'b11111111111111111101101010100000;
assign LUT_1[33136] = 32'b00000000000000000011011110101001;
assign LUT_1[33137] = 32'b11111111111111111100110000100101;
assign LUT_1[33138] = 32'b11111111111111111111001100111010;
assign LUT_1[33139] = 32'b11111111111111111000011110110110;
assign LUT_1[33140] = 32'b00000000000000001011011000000000;
assign LUT_1[33141] = 32'b00000000000000000100101001111100;
assign LUT_1[33142] = 32'b00000000000000000111000110010001;
assign LUT_1[33143] = 32'b00000000000000000000011000001101;
assign LUT_1[33144] = 32'b00000000000000000010101100011110;
assign LUT_1[33145] = 32'b11111111111111111011111110011010;
assign LUT_1[33146] = 32'b11111111111111111110011010101111;
assign LUT_1[33147] = 32'b11111111111111110111101100101011;
assign LUT_1[33148] = 32'b00000000000000001010100101110101;
assign LUT_1[33149] = 32'b00000000000000000011110111110001;
assign LUT_1[33150] = 32'b00000000000000000110010100000110;
assign LUT_1[33151] = 32'b11111111111111111111100110000010;
assign LUT_1[33152] = 32'b00000000000000000001101010100011;
assign LUT_1[33153] = 32'b11111111111111111010111100011111;
assign LUT_1[33154] = 32'b11111111111111111101011000110100;
assign LUT_1[33155] = 32'b11111111111111110110101010110000;
assign LUT_1[33156] = 32'b00000000000000001001100011111010;
assign LUT_1[33157] = 32'b00000000000000000010110101110110;
assign LUT_1[33158] = 32'b00000000000000000101010010001011;
assign LUT_1[33159] = 32'b11111111111111111110100100000111;
assign LUT_1[33160] = 32'b00000000000000000000111000011000;
assign LUT_1[33161] = 32'b11111111111111111010001010010100;
assign LUT_1[33162] = 32'b11111111111111111100100110101001;
assign LUT_1[33163] = 32'b11111111111111110101111000100101;
assign LUT_1[33164] = 32'b00000000000000001000110001101111;
assign LUT_1[33165] = 32'b00000000000000000010000011101011;
assign LUT_1[33166] = 32'b00000000000000000100100000000000;
assign LUT_1[33167] = 32'b11111111111111111101110001111100;
assign LUT_1[33168] = 32'b00000000000000000011100110000101;
assign LUT_1[33169] = 32'b11111111111111111100111000000001;
assign LUT_1[33170] = 32'b11111111111111111111010100010110;
assign LUT_1[33171] = 32'b11111111111111111000100110010010;
assign LUT_1[33172] = 32'b00000000000000001011011111011100;
assign LUT_1[33173] = 32'b00000000000000000100110001011000;
assign LUT_1[33174] = 32'b00000000000000000111001101101101;
assign LUT_1[33175] = 32'b00000000000000000000011111101001;
assign LUT_1[33176] = 32'b00000000000000000010110011111010;
assign LUT_1[33177] = 32'b11111111111111111100000101110110;
assign LUT_1[33178] = 32'b11111111111111111110100010001011;
assign LUT_1[33179] = 32'b11111111111111110111110100000111;
assign LUT_1[33180] = 32'b00000000000000001010101101010001;
assign LUT_1[33181] = 32'b00000000000000000011111111001101;
assign LUT_1[33182] = 32'b00000000000000000110011011100010;
assign LUT_1[33183] = 32'b11111111111111111111101101011110;
assign LUT_1[33184] = 32'b00000000000000000010100101100010;
assign LUT_1[33185] = 32'b11111111111111111011110111011110;
assign LUT_1[33186] = 32'b11111111111111111110010011110011;
assign LUT_1[33187] = 32'b11111111111111110111100101101111;
assign LUT_1[33188] = 32'b00000000000000001010011110111001;
assign LUT_1[33189] = 32'b00000000000000000011110000110101;
assign LUT_1[33190] = 32'b00000000000000000110001101001010;
assign LUT_1[33191] = 32'b11111111111111111111011111000110;
assign LUT_1[33192] = 32'b00000000000000000001110011010111;
assign LUT_1[33193] = 32'b11111111111111111011000101010011;
assign LUT_1[33194] = 32'b11111111111111111101100001101000;
assign LUT_1[33195] = 32'b11111111111111110110110011100100;
assign LUT_1[33196] = 32'b00000000000000001001101100101110;
assign LUT_1[33197] = 32'b00000000000000000010111110101010;
assign LUT_1[33198] = 32'b00000000000000000101011010111111;
assign LUT_1[33199] = 32'b11111111111111111110101100111011;
assign LUT_1[33200] = 32'b00000000000000000100100001000100;
assign LUT_1[33201] = 32'b11111111111111111101110011000000;
assign LUT_1[33202] = 32'b00000000000000000000001111010101;
assign LUT_1[33203] = 32'b11111111111111111001100001010001;
assign LUT_1[33204] = 32'b00000000000000001100011010011011;
assign LUT_1[33205] = 32'b00000000000000000101101100010111;
assign LUT_1[33206] = 32'b00000000000000001000001000101100;
assign LUT_1[33207] = 32'b00000000000000000001011010101000;
assign LUT_1[33208] = 32'b00000000000000000011101110111001;
assign LUT_1[33209] = 32'b11111111111111111101000000110101;
assign LUT_1[33210] = 32'b11111111111111111111011101001010;
assign LUT_1[33211] = 32'b11111111111111111000101111000110;
assign LUT_1[33212] = 32'b00000000000000001011101000010000;
assign LUT_1[33213] = 32'b00000000000000000100111010001100;
assign LUT_1[33214] = 32'b00000000000000000111010110100001;
assign LUT_1[33215] = 32'b00000000000000000000101000011101;
assign LUT_1[33216] = 32'b00000000000000000011101000001011;
assign LUT_1[33217] = 32'b11111111111111111100111010000111;
assign LUT_1[33218] = 32'b11111111111111111111010110011100;
assign LUT_1[33219] = 32'b11111111111111111000101000011000;
assign LUT_1[33220] = 32'b00000000000000001011100001100010;
assign LUT_1[33221] = 32'b00000000000000000100110011011110;
assign LUT_1[33222] = 32'b00000000000000000111001111110011;
assign LUT_1[33223] = 32'b00000000000000000000100001101111;
assign LUT_1[33224] = 32'b00000000000000000010110110000000;
assign LUT_1[33225] = 32'b11111111111111111100000111111100;
assign LUT_1[33226] = 32'b11111111111111111110100100010001;
assign LUT_1[33227] = 32'b11111111111111110111110110001101;
assign LUT_1[33228] = 32'b00000000000000001010101111010111;
assign LUT_1[33229] = 32'b00000000000000000100000001010011;
assign LUT_1[33230] = 32'b00000000000000000110011101101000;
assign LUT_1[33231] = 32'b11111111111111111111101111100100;
assign LUT_1[33232] = 32'b00000000000000000101100011101101;
assign LUT_1[33233] = 32'b11111111111111111110110101101001;
assign LUT_1[33234] = 32'b00000000000000000001010001111110;
assign LUT_1[33235] = 32'b11111111111111111010100011111010;
assign LUT_1[33236] = 32'b00000000000000001101011101000100;
assign LUT_1[33237] = 32'b00000000000000000110101111000000;
assign LUT_1[33238] = 32'b00000000000000001001001011010101;
assign LUT_1[33239] = 32'b00000000000000000010011101010001;
assign LUT_1[33240] = 32'b00000000000000000100110001100010;
assign LUT_1[33241] = 32'b11111111111111111110000011011110;
assign LUT_1[33242] = 32'b00000000000000000000011111110011;
assign LUT_1[33243] = 32'b11111111111111111001110001101111;
assign LUT_1[33244] = 32'b00000000000000001100101010111001;
assign LUT_1[33245] = 32'b00000000000000000101111100110101;
assign LUT_1[33246] = 32'b00000000000000001000011001001010;
assign LUT_1[33247] = 32'b00000000000000000001101011000110;
assign LUT_1[33248] = 32'b00000000000000000100100011001010;
assign LUT_1[33249] = 32'b11111111111111111101110101000110;
assign LUT_1[33250] = 32'b00000000000000000000010001011011;
assign LUT_1[33251] = 32'b11111111111111111001100011010111;
assign LUT_1[33252] = 32'b00000000000000001100011100100001;
assign LUT_1[33253] = 32'b00000000000000000101101110011101;
assign LUT_1[33254] = 32'b00000000000000001000001010110010;
assign LUT_1[33255] = 32'b00000000000000000001011100101110;
assign LUT_1[33256] = 32'b00000000000000000011110000111111;
assign LUT_1[33257] = 32'b11111111111111111101000010111011;
assign LUT_1[33258] = 32'b11111111111111111111011111010000;
assign LUT_1[33259] = 32'b11111111111111111000110001001100;
assign LUT_1[33260] = 32'b00000000000000001011101010010110;
assign LUT_1[33261] = 32'b00000000000000000100111100010010;
assign LUT_1[33262] = 32'b00000000000000000111011000100111;
assign LUT_1[33263] = 32'b00000000000000000000101010100011;
assign LUT_1[33264] = 32'b00000000000000000110011110101100;
assign LUT_1[33265] = 32'b11111111111111111111110000101000;
assign LUT_1[33266] = 32'b00000000000000000010001100111101;
assign LUT_1[33267] = 32'b11111111111111111011011110111001;
assign LUT_1[33268] = 32'b00000000000000001110011000000011;
assign LUT_1[33269] = 32'b00000000000000000111101001111111;
assign LUT_1[33270] = 32'b00000000000000001010000110010100;
assign LUT_1[33271] = 32'b00000000000000000011011000010000;
assign LUT_1[33272] = 32'b00000000000000000101101100100001;
assign LUT_1[33273] = 32'b11111111111111111110111110011101;
assign LUT_1[33274] = 32'b00000000000000000001011010110010;
assign LUT_1[33275] = 32'b11111111111111111010101100101110;
assign LUT_1[33276] = 32'b00000000000000001101100101111000;
assign LUT_1[33277] = 32'b00000000000000000110110111110100;
assign LUT_1[33278] = 32'b00000000000000001001010100001001;
assign LUT_1[33279] = 32'b00000000000000000010100110000101;
assign LUT_1[33280] = 32'b11111111111111111010100100110001;
assign LUT_1[33281] = 32'b11111111111111110011110110101101;
assign LUT_1[33282] = 32'b11111111111111110110010011000010;
assign LUT_1[33283] = 32'b11111111111111101111100100111110;
assign LUT_1[33284] = 32'b00000000000000000010011110001000;
assign LUT_1[33285] = 32'b11111111111111111011110000000100;
assign LUT_1[33286] = 32'b11111111111111111110001100011001;
assign LUT_1[33287] = 32'b11111111111111110111011110010101;
assign LUT_1[33288] = 32'b11111111111111111001110010100110;
assign LUT_1[33289] = 32'b11111111111111110011000100100010;
assign LUT_1[33290] = 32'b11111111111111110101100000110111;
assign LUT_1[33291] = 32'b11111111111111101110110010110011;
assign LUT_1[33292] = 32'b00000000000000000001101011111101;
assign LUT_1[33293] = 32'b11111111111111111010111101111001;
assign LUT_1[33294] = 32'b11111111111111111101011010001110;
assign LUT_1[33295] = 32'b11111111111111110110101100001010;
assign LUT_1[33296] = 32'b11111111111111111100100000010011;
assign LUT_1[33297] = 32'b11111111111111110101110010001111;
assign LUT_1[33298] = 32'b11111111111111111000001110100100;
assign LUT_1[33299] = 32'b11111111111111110001100000100000;
assign LUT_1[33300] = 32'b00000000000000000100011001101010;
assign LUT_1[33301] = 32'b11111111111111111101101011100110;
assign LUT_1[33302] = 32'b00000000000000000000000111111011;
assign LUT_1[33303] = 32'b11111111111111111001011001110111;
assign LUT_1[33304] = 32'b11111111111111111011101110001000;
assign LUT_1[33305] = 32'b11111111111111110101000000000100;
assign LUT_1[33306] = 32'b11111111111111110111011100011001;
assign LUT_1[33307] = 32'b11111111111111110000101110010101;
assign LUT_1[33308] = 32'b00000000000000000011100111011111;
assign LUT_1[33309] = 32'b11111111111111111100111001011011;
assign LUT_1[33310] = 32'b11111111111111111111010101110000;
assign LUT_1[33311] = 32'b11111111111111111000100111101100;
assign LUT_1[33312] = 32'b11111111111111111011011111110000;
assign LUT_1[33313] = 32'b11111111111111110100110001101100;
assign LUT_1[33314] = 32'b11111111111111110111001110000001;
assign LUT_1[33315] = 32'b11111111111111110000011111111101;
assign LUT_1[33316] = 32'b00000000000000000011011001000111;
assign LUT_1[33317] = 32'b11111111111111111100101011000011;
assign LUT_1[33318] = 32'b11111111111111111111000111011000;
assign LUT_1[33319] = 32'b11111111111111111000011001010100;
assign LUT_1[33320] = 32'b11111111111111111010101101100101;
assign LUT_1[33321] = 32'b11111111111111110011111111100001;
assign LUT_1[33322] = 32'b11111111111111110110011011110110;
assign LUT_1[33323] = 32'b11111111111111101111101101110010;
assign LUT_1[33324] = 32'b00000000000000000010100110111100;
assign LUT_1[33325] = 32'b11111111111111111011111000111000;
assign LUT_1[33326] = 32'b11111111111111111110010101001101;
assign LUT_1[33327] = 32'b11111111111111110111100111001001;
assign LUT_1[33328] = 32'b11111111111111111101011011010010;
assign LUT_1[33329] = 32'b11111111111111110110101101001110;
assign LUT_1[33330] = 32'b11111111111111111001001001100011;
assign LUT_1[33331] = 32'b11111111111111110010011011011111;
assign LUT_1[33332] = 32'b00000000000000000101010100101001;
assign LUT_1[33333] = 32'b11111111111111111110100110100101;
assign LUT_1[33334] = 32'b00000000000000000001000010111010;
assign LUT_1[33335] = 32'b11111111111111111010010100110110;
assign LUT_1[33336] = 32'b11111111111111111100101001000111;
assign LUT_1[33337] = 32'b11111111111111110101111011000011;
assign LUT_1[33338] = 32'b11111111111111111000010111011000;
assign LUT_1[33339] = 32'b11111111111111110001101001010100;
assign LUT_1[33340] = 32'b00000000000000000100100010011110;
assign LUT_1[33341] = 32'b11111111111111111101110100011010;
assign LUT_1[33342] = 32'b00000000000000000000010000101111;
assign LUT_1[33343] = 32'b11111111111111111001100010101011;
assign LUT_1[33344] = 32'b11111111111111111100100010011001;
assign LUT_1[33345] = 32'b11111111111111110101110100010101;
assign LUT_1[33346] = 32'b11111111111111111000010000101010;
assign LUT_1[33347] = 32'b11111111111111110001100010100110;
assign LUT_1[33348] = 32'b00000000000000000100011011110000;
assign LUT_1[33349] = 32'b11111111111111111101101101101100;
assign LUT_1[33350] = 32'b00000000000000000000001010000001;
assign LUT_1[33351] = 32'b11111111111111111001011011111101;
assign LUT_1[33352] = 32'b11111111111111111011110000001110;
assign LUT_1[33353] = 32'b11111111111111110101000010001010;
assign LUT_1[33354] = 32'b11111111111111110111011110011111;
assign LUT_1[33355] = 32'b11111111111111110000110000011011;
assign LUT_1[33356] = 32'b00000000000000000011101001100101;
assign LUT_1[33357] = 32'b11111111111111111100111011100001;
assign LUT_1[33358] = 32'b11111111111111111111010111110110;
assign LUT_1[33359] = 32'b11111111111111111000101001110010;
assign LUT_1[33360] = 32'b11111111111111111110011101111011;
assign LUT_1[33361] = 32'b11111111111111110111101111110111;
assign LUT_1[33362] = 32'b11111111111111111010001100001100;
assign LUT_1[33363] = 32'b11111111111111110011011110001000;
assign LUT_1[33364] = 32'b00000000000000000110010111010010;
assign LUT_1[33365] = 32'b11111111111111111111101001001110;
assign LUT_1[33366] = 32'b00000000000000000010000101100011;
assign LUT_1[33367] = 32'b11111111111111111011010111011111;
assign LUT_1[33368] = 32'b11111111111111111101101011110000;
assign LUT_1[33369] = 32'b11111111111111110110111101101100;
assign LUT_1[33370] = 32'b11111111111111111001011010000001;
assign LUT_1[33371] = 32'b11111111111111110010101011111101;
assign LUT_1[33372] = 32'b00000000000000000101100101000111;
assign LUT_1[33373] = 32'b11111111111111111110110111000011;
assign LUT_1[33374] = 32'b00000000000000000001010011011000;
assign LUT_1[33375] = 32'b11111111111111111010100101010100;
assign LUT_1[33376] = 32'b11111111111111111101011101011000;
assign LUT_1[33377] = 32'b11111111111111110110101111010100;
assign LUT_1[33378] = 32'b11111111111111111001001011101001;
assign LUT_1[33379] = 32'b11111111111111110010011101100101;
assign LUT_1[33380] = 32'b00000000000000000101010110101111;
assign LUT_1[33381] = 32'b11111111111111111110101000101011;
assign LUT_1[33382] = 32'b00000000000000000001000101000000;
assign LUT_1[33383] = 32'b11111111111111111010010110111100;
assign LUT_1[33384] = 32'b11111111111111111100101011001101;
assign LUT_1[33385] = 32'b11111111111111110101111101001001;
assign LUT_1[33386] = 32'b11111111111111111000011001011110;
assign LUT_1[33387] = 32'b11111111111111110001101011011010;
assign LUT_1[33388] = 32'b00000000000000000100100100100100;
assign LUT_1[33389] = 32'b11111111111111111101110110100000;
assign LUT_1[33390] = 32'b00000000000000000000010010110101;
assign LUT_1[33391] = 32'b11111111111111111001100100110001;
assign LUT_1[33392] = 32'b11111111111111111111011000111010;
assign LUT_1[33393] = 32'b11111111111111111000101010110110;
assign LUT_1[33394] = 32'b11111111111111111011000111001011;
assign LUT_1[33395] = 32'b11111111111111110100011001000111;
assign LUT_1[33396] = 32'b00000000000000000111010010010001;
assign LUT_1[33397] = 32'b00000000000000000000100100001101;
assign LUT_1[33398] = 32'b00000000000000000011000000100010;
assign LUT_1[33399] = 32'b11111111111111111100010010011110;
assign LUT_1[33400] = 32'b11111111111111111110100110101111;
assign LUT_1[33401] = 32'b11111111111111110111111000101011;
assign LUT_1[33402] = 32'b11111111111111111010010101000000;
assign LUT_1[33403] = 32'b11111111111111110011100110111100;
assign LUT_1[33404] = 32'b00000000000000000110100000000110;
assign LUT_1[33405] = 32'b11111111111111111111110010000010;
assign LUT_1[33406] = 32'b00000000000000000010001110010111;
assign LUT_1[33407] = 32'b11111111111111111011100000010011;
assign LUT_1[33408] = 32'b11111111111111111101100100110100;
assign LUT_1[33409] = 32'b11111111111111110110110110110000;
assign LUT_1[33410] = 32'b11111111111111111001010011000101;
assign LUT_1[33411] = 32'b11111111111111110010100101000001;
assign LUT_1[33412] = 32'b00000000000000000101011110001011;
assign LUT_1[33413] = 32'b11111111111111111110110000000111;
assign LUT_1[33414] = 32'b00000000000000000001001100011100;
assign LUT_1[33415] = 32'b11111111111111111010011110011000;
assign LUT_1[33416] = 32'b11111111111111111100110010101001;
assign LUT_1[33417] = 32'b11111111111111110110000100100101;
assign LUT_1[33418] = 32'b11111111111111111000100000111010;
assign LUT_1[33419] = 32'b11111111111111110001110010110110;
assign LUT_1[33420] = 32'b00000000000000000100101100000000;
assign LUT_1[33421] = 32'b11111111111111111101111101111100;
assign LUT_1[33422] = 32'b00000000000000000000011010010001;
assign LUT_1[33423] = 32'b11111111111111111001101100001101;
assign LUT_1[33424] = 32'b11111111111111111111100000010110;
assign LUT_1[33425] = 32'b11111111111111111000110010010010;
assign LUT_1[33426] = 32'b11111111111111111011001110100111;
assign LUT_1[33427] = 32'b11111111111111110100100000100011;
assign LUT_1[33428] = 32'b00000000000000000111011001101101;
assign LUT_1[33429] = 32'b00000000000000000000101011101001;
assign LUT_1[33430] = 32'b00000000000000000011000111111110;
assign LUT_1[33431] = 32'b11111111111111111100011001111010;
assign LUT_1[33432] = 32'b11111111111111111110101110001011;
assign LUT_1[33433] = 32'b11111111111111111000000000000111;
assign LUT_1[33434] = 32'b11111111111111111010011100011100;
assign LUT_1[33435] = 32'b11111111111111110011101110011000;
assign LUT_1[33436] = 32'b00000000000000000110100111100010;
assign LUT_1[33437] = 32'b11111111111111111111111001011110;
assign LUT_1[33438] = 32'b00000000000000000010010101110011;
assign LUT_1[33439] = 32'b11111111111111111011100111101111;
assign LUT_1[33440] = 32'b11111111111111111110011111110011;
assign LUT_1[33441] = 32'b11111111111111110111110001101111;
assign LUT_1[33442] = 32'b11111111111111111010001110000100;
assign LUT_1[33443] = 32'b11111111111111110011100000000000;
assign LUT_1[33444] = 32'b00000000000000000110011001001010;
assign LUT_1[33445] = 32'b11111111111111111111101011000110;
assign LUT_1[33446] = 32'b00000000000000000010000111011011;
assign LUT_1[33447] = 32'b11111111111111111011011001010111;
assign LUT_1[33448] = 32'b11111111111111111101101101101000;
assign LUT_1[33449] = 32'b11111111111111110110111111100100;
assign LUT_1[33450] = 32'b11111111111111111001011011111001;
assign LUT_1[33451] = 32'b11111111111111110010101101110101;
assign LUT_1[33452] = 32'b00000000000000000101100110111111;
assign LUT_1[33453] = 32'b11111111111111111110111000111011;
assign LUT_1[33454] = 32'b00000000000000000001010101010000;
assign LUT_1[33455] = 32'b11111111111111111010100111001100;
assign LUT_1[33456] = 32'b00000000000000000000011011010101;
assign LUT_1[33457] = 32'b11111111111111111001101101010001;
assign LUT_1[33458] = 32'b11111111111111111100001001100110;
assign LUT_1[33459] = 32'b11111111111111110101011011100010;
assign LUT_1[33460] = 32'b00000000000000001000010100101100;
assign LUT_1[33461] = 32'b00000000000000000001100110101000;
assign LUT_1[33462] = 32'b00000000000000000100000010111101;
assign LUT_1[33463] = 32'b11111111111111111101010100111001;
assign LUT_1[33464] = 32'b11111111111111111111101001001010;
assign LUT_1[33465] = 32'b11111111111111111000111011000110;
assign LUT_1[33466] = 32'b11111111111111111011010111011011;
assign LUT_1[33467] = 32'b11111111111111110100101001010111;
assign LUT_1[33468] = 32'b00000000000000000111100010100001;
assign LUT_1[33469] = 32'b00000000000000000000110100011101;
assign LUT_1[33470] = 32'b00000000000000000011010000110010;
assign LUT_1[33471] = 32'b11111111111111111100100010101110;
assign LUT_1[33472] = 32'b11111111111111111111100010011100;
assign LUT_1[33473] = 32'b11111111111111111000110100011000;
assign LUT_1[33474] = 32'b11111111111111111011010000101101;
assign LUT_1[33475] = 32'b11111111111111110100100010101001;
assign LUT_1[33476] = 32'b00000000000000000111011011110011;
assign LUT_1[33477] = 32'b00000000000000000000101101101111;
assign LUT_1[33478] = 32'b00000000000000000011001010000100;
assign LUT_1[33479] = 32'b11111111111111111100011100000000;
assign LUT_1[33480] = 32'b11111111111111111110110000010001;
assign LUT_1[33481] = 32'b11111111111111111000000010001101;
assign LUT_1[33482] = 32'b11111111111111111010011110100010;
assign LUT_1[33483] = 32'b11111111111111110011110000011110;
assign LUT_1[33484] = 32'b00000000000000000110101001101000;
assign LUT_1[33485] = 32'b11111111111111111111111011100100;
assign LUT_1[33486] = 32'b00000000000000000010010111111001;
assign LUT_1[33487] = 32'b11111111111111111011101001110101;
assign LUT_1[33488] = 32'b00000000000000000001011101111110;
assign LUT_1[33489] = 32'b11111111111111111010101111111010;
assign LUT_1[33490] = 32'b11111111111111111101001100001111;
assign LUT_1[33491] = 32'b11111111111111110110011110001011;
assign LUT_1[33492] = 32'b00000000000000001001010111010101;
assign LUT_1[33493] = 32'b00000000000000000010101001010001;
assign LUT_1[33494] = 32'b00000000000000000101000101100110;
assign LUT_1[33495] = 32'b11111111111111111110010111100010;
assign LUT_1[33496] = 32'b00000000000000000000101011110011;
assign LUT_1[33497] = 32'b11111111111111111001111101101111;
assign LUT_1[33498] = 32'b11111111111111111100011010000100;
assign LUT_1[33499] = 32'b11111111111111110101101100000000;
assign LUT_1[33500] = 32'b00000000000000001000100101001010;
assign LUT_1[33501] = 32'b00000000000000000001110111000110;
assign LUT_1[33502] = 32'b00000000000000000100010011011011;
assign LUT_1[33503] = 32'b11111111111111111101100101010111;
assign LUT_1[33504] = 32'b00000000000000000000011101011011;
assign LUT_1[33505] = 32'b11111111111111111001101111010111;
assign LUT_1[33506] = 32'b11111111111111111100001011101100;
assign LUT_1[33507] = 32'b11111111111111110101011101101000;
assign LUT_1[33508] = 32'b00000000000000001000010110110010;
assign LUT_1[33509] = 32'b00000000000000000001101000101110;
assign LUT_1[33510] = 32'b00000000000000000100000101000011;
assign LUT_1[33511] = 32'b11111111111111111101010110111111;
assign LUT_1[33512] = 32'b11111111111111111111101011010000;
assign LUT_1[33513] = 32'b11111111111111111000111101001100;
assign LUT_1[33514] = 32'b11111111111111111011011001100001;
assign LUT_1[33515] = 32'b11111111111111110100101011011101;
assign LUT_1[33516] = 32'b00000000000000000111100100100111;
assign LUT_1[33517] = 32'b00000000000000000000110110100011;
assign LUT_1[33518] = 32'b00000000000000000011010010111000;
assign LUT_1[33519] = 32'b11111111111111111100100100110100;
assign LUT_1[33520] = 32'b00000000000000000010011000111101;
assign LUT_1[33521] = 32'b11111111111111111011101010111001;
assign LUT_1[33522] = 32'b11111111111111111110000111001110;
assign LUT_1[33523] = 32'b11111111111111110111011001001010;
assign LUT_1[33524] = 32'b00000000000000001010010010010100;
assign LUT_1[33525] = 32'b00000000000000000011100100010000;
assign LUT_1[33526] = 32'b00000000000000000110000000100101;
assign LUT_1[33527] = 32'b11111111111111111111010010100001;
assign LUT_1[33528] = 32'b00000000000000000001100110110010;
assign LUT_1[33529] = 32'b11111111111111111010111000101110;
assign LUT_1[33530] = 32'b11111111111111111101010101000011;
assign LUT_1[33531] = 32'b11111111111111110110100110111111;
assign LUT_1[33532] = 32'b00000000000000001001100000001001;
assign LUT_1[33533] = 32'b00000000000000000010110010000101;
assign LUT_1[33534] = 32'b00000000000000000101001110011010;
assign LUT_1[33535] = 32'b11111111111111111110100000010110;
assign LUT_1[33536] = 32'b11111111111111111000011000111101;
assign LUT_1[33537] = 32'b11111111111111110001101010111001;
assign LUT_1[33538] = 32'b11111111111111110100000111001110;
assign LUT_1[33539] = 32'b11111111111111101101011001001010;
assign LUT_1[33540] = 32'b00000000000000000000010010010100;
assign LUT_1[33541] = 32'b11111111111111111001100100010000;
assign LUT_1[33542] = 32'b11111111111111111100000000100101;
assign LUT_1[33543] = 32'b11111111111111110101010010100001;
assign LUT_1[33544] = 32'b11111111111111110111100110110010;
assign LUT_1[33545] = 32'b11111111111111110000111000101110;
assign LUT_1[33546] = 32'b11111111111111110011010101000011;
assign LUT_1[33547] = 32'b11111111111111101100100110111111;
assign LUT_1[33548] = 32'b11111111111111111111100000001001;
assign LUT_1[33549] = 32'b11111111111111111000110010000101;
assign LUT_1[33550] = 32'b11111111111111111011001110011010;
assign LUT_1[33551] = 32'b11111111111111110100100000010110;
assign LUT_1[33552] = 32'b11111111111111111010010100011111;
assign LUT_1[33553] = 32'b11111111111111110011100110011011;
assign LUT_1[33554] = 32'b11111111111111110110000010110000;
assign LUT_1[33555] = 32'b11111111111111101111010100101100;
assign LUT_1[33556] = 32'b00000000000000000010001101110110;
assign LUT_1[33557] = 32'b11111111111111111011011111110010;
assign LUT_1[33558] = 32'b11111111111111111101111100000111;
assign LUT_1[33559] = 32'b11111111111111110111001110000011;
assign LUT_1[33560] = 32'b11111111111111111001100010010100;
assign LUT_1[33561] = 32'b11111111111111110010110100010000;
assign LUT_1[33562] = 32'b11111111111111110101010000100101;
assign LUT_1[33563] = 32'b11111111111111101110100010100001;
assign LUT_1[33564] = 32'b00000000000000000001011011101011;
assign LUT_1[33565] = 32'b11111111111111111010101101100111;
assign LUT_1[33566] = 32'b11111111111111111101001001111100;
assign LUT_1[33567] = 32'b11111111111111110110011011111000;
assign LUT_1[33568] = 32'b11111111111111111001010011111100;
assign LUT_1[33569] = 32'b11111111111111110010100101111000;
assign LUT_1[33570] = 32'b11111111111111110101000010001101;
assign LUT_1[33571] = 32'b11111111111111101110010100001001;
assign LUT_1[33572] = 32'b00000000000000000001001101010011;
assign LUT_1[33573] = 32'b11111111111111111010011111001111;
assign LUT_1[33574] = 32'b11111111111111111100111011100100;
assign LUT_1[33575] = 32'b11111111111111110110001101100000;
assign LUT_1[33576] = 32'b11111111111111111000100001110001;
assign LUT_1[33577] = 32'b11111111111111110001110011101101;
assign LUT_1[33578] = 32'b11111111111111110100010000000010;
assign LUT_1[33579] = 32'b11111111111111101101100001111110;
assign LUT_1[33580] = 32'b00000000000000000000011011001000;
assign LUT_1[33581] = 32'b11111111111111111001101101000100;
assign LUT_1[33582] = 32'b11111111111111111100001001011001;
assign LUT_1[33583] = 32'b11111111111111110101011011010101;
assign LUT_1[33584] = 32'b11111111111111111011001111011110;
assign LUT_1[33585] = 32'b11111111111111110100100001011010;
assign LUT_1[33586] = 32'b11111111111111110110111101101111;
assign LUT_1[33587] = 32'b11111111111111110000001111101011;
assign LUT_1[33588] = 32'b00000000000000000011001000110101;
assign LUT_1[33589] = 32'b11111111111111111100011010110001;
assign LUT_1[33590] = 32'b11111111111111111110110111000110;
assign LUT_1[33591] = 32'b11111111111111111000001001000010;
assign LUT_1[33592] = 32'b11111111111111111010011101010011;
assign LUT_1[33593] = 32'b11111111111111110011101111001111;
assign LUT_1[33594] = 32'b11111111111111110110001011100100;
assign LUT_1[33595] = 32'b11111111111111101111011101100000;
assign LUT_1[33596] = 32'b00000000000000000010010110101010;
assign LUT_1[33597] = 32'b11111111111111111011101000100110;
assign LUT_1[33598] = 32'b11111111111111111110000100111011;
assign LUT_1[33599] = 32'b11111111111111110111010110110111;
assign LUT_1[33600] = 32'b11111111111111111010010110100101;
assign LUT_1[33601] = 32'b11111111111111110011101000100001;
assign LUT_1[33602] = 32'b11111111111111110110000100110110;
assign LUT_1[33603] = 32'b11111111111111101111010110110010;
assign LUT_1[33604] = 32'b00000000000000000010001111111100;
assign LUT_1[33605] = 32'b11111111111111111011100001111000;
assign LUT_1[33606] = 32'b11111111111111111101111110001101;
assign LUT_1[33607] = 32'b11111111111111110111010000001001;
assign LUT_1[33608] = 32'b11111111111111111001100100011010;
assign LUT_1[33609] = 32'b11111111111111110010110110010110;
assign LUT_1[33610] = 32'b11111111111111110101010010101011;
assign LUT_1[33611] = 32'b11111111111111101110100100100111;
assign LUT_1[33612] = 32'b00000000000000000001011101110001;
assign LUT_1[33613] = 32'b11111111111111111010101111101101;
assign LUT_1[33614] = 32'b11111111111111111101001100000010;
assign LUT_1[33615] = 32'b11111111111111110110011101111110;
assign LUT_1[33616] = 32'b11111111111111111100010010000111;
assign LUT_1[33617] = 32'b11111111111111110101100100000011;
assign LUT_1[33618] = 32'b11111111111111111000000000011000;
assign LUT_1[33619] = 32'b11111111111111110001010010010100;
assign LUT_1[33620] = 32'b00000000000000000100001011011110;
assign LUT_1[33621] = 32'b11111111111111111101011101011010;
assign LUT_1[33622] = 32'b11111111111111111111111001101111;
assign LUT_1[33623] = 32'b11111111111111111001001011101011;
assign LUT_1[33624] = 32'b11111111111111111011011111111100;
assign LUT_1[33625] = 32'b11111111111111110100110001111000;
assign LUT_1[33626] = 32'b11111111111111110111001110001101;
assign LUT_1[33627] = 32'b11111111111111110000100000001001;
assign LUT_1[33628] = 32'b00000000000000000011011001010011;
assign LUT_1[33629] = 32'b11111111111111111100101011001111;
assign LUT_1[33630] = 32'b11111111111111111111000111100100;
assign LUT_1[33631] = 32'b11111111111111111000011001100000;
assign LUT_1[33632] = 32'b11111111111111111011010001100100;
assign LUT_1[33633] = 32'b11111111111111110100100011100000;
assign LUT_1[33634] = 32'b11111111111111110110111111110101;
assign LUT_1[33635] = 32'b11111111111111110000010001110001;
assign LUT_1[33636] = 32'b00000000000000000011001010111011;
assign LUT_1[33637] = 32'b11111111111111111100011100110111;
assign LUT_1[33638] = 32'b11111111111111111110111001001100;
assign LUT_1[33639] = 32'b11111111111111111000001011001000;
assign LUT_1[33640] = 32'b11111111111111111010011111011001;
assign LUT_1[33641] = 32'b11111111111111110011110001010101;
assign LUT_1[33642] = 32'b11111111111111110110001101101010;
assign LUT_1[33643] = 32'b11111111111111101111011111100110;
assign LUT_1[33644] = 32'b00000000000000000010011000110000;
assign LUT_1[33645] = 32'b11111111111111111011101010101100;
assign LUT_1[33646] = 32'b11111111111111111110000111000001;
assign LUT_1[33647] = 32'b11111111111111110111011000111101;
assign LUT_1[33648] = 32'b11111111111111111101001101000110;
assign LUT_1[33649] = 32'b11111111111111110110011111000010;
assign LUT_1[33650] = 32'b11111111111111111000111011010111;
assign LUT_1[33651] = 32'b11111111111111110010001101010011;
assign LUT_1[33652] = 32'b00000000000000000101000110011101;
assign LUT_1[33653] = 32'b11111111111111111110011000011001;
assign LUT_1[33654] = 32'b00000000000000000000110100101110;
assign LUT_1[33655] = 32'b11111111111111111010000110101010;
assign LUT_1[33656] = 32'b11111111111111111100011010111011;
assign LUT_1[33657] = 32'b11111111111111110101101100110111;
assign LUT_1[33658] = 32'b11111111111111111000001001001100;
assign LUT_1[33659] = 32'b11111111111111110001011011001000;
assign LUT_1[33660] = 32'b00000000000000000100010100010010;
assign LUT_1[33661] = 32'b11111111111111111101100110001110;
assign LUT_1[33662] = 32'b00000000000000000000000010100011;
assign LUT_1[33663] = 32'b11111111111111111001010100011111;
assign LUT_1[33664] = 32'b11111111111111111011011001000000;
assign LUT_1[33665] = 32'b11111111111111110100101010111100;
assign LUT_1[33666] = 32'b11111111111111110111000111010001;
assign LUT_1[33667] = 32'b11111111111111110000011001001101;
assign LUT_1[33668] = 32'b00000000000000000011010010010111;
assign LUT_1[33669] = 32'b11111111111111111100100100010011;
assign LUT_1[33670] = 32'b11111111111111111111000000101000;
assign LUT_1[33671] = 32'b11111111111111111000010010100100;
assign LUT_1[33672] = 32'b11111111111111111010100110110101;
assign LUT_1[33673] = 32'b11111111111111110011111000110001;
assign LUT_1[33674] = 32'b11111111111111110110010101000110;
assign LUT_1[33675] = 32'b11111111111111101111100111000010;
assign LUT_1[33676] = 32'b00000000000000000010100000001100;
assign LUT_1[33677] = 32'b11111111111111111011110010001000;
assign LUT_1[33678] = 32'b11111111111111111110001110011101;
assign LUT_1[33679] = 32'b11111111111111110111100000011001;
assign LUT_1[33680] = 32'b11111111111111111101010100100010;
assign LUT_1[33681] = 32'b11111111111111110110100110011110;
assign LUT_1[33682] = 32'b11111111111111111001000010110011;
assign LUT_1[33683] = 32'b11111111111111110010010100101111;
assign LUT_1[33684] = 32'b00000000000000000101001101111001;
assign LUT_1[33685] = 32'b11111111111111111110011111110101;
assign LUT_1[33686] = 32'b00000000000000000000111100001010;
assign LUT_1[33687] = 32'b11111111111111111010001110000110;
assign LUT_1[33688] = 32'b11111111111111111100100010010111;
assign LUT_1[33689] = 32'b11111111111111110101110100010011;
assign LUT_1[33690] = 32'b11111111111111111000010000101000;
assign LUT_1[33691] = 32'b11111111111111110001100010100100;
assign LUT_1[33692] = 32'b00000000000000000100011011101110;
assign LUT_1[33693] = 32'b11111111111111111101101101101010;
assign LUT_1[33694] = 32'b00000000000000000000001001111111;
assign LUT_1[33695] = 32'b11111111111111111001011011111011;
assign LUT_1[33696] = 32'b11111111111111111100010011111111;
assign LUT_1[33697] = 32'b11111111111111110101100101111011;
assign LUT_1[33698] = 32'b11111111111111111000000010010000;
assign LUT_1[33699] = 32'b11111111111111110001010100001100;
assign LUT_1[33700] = 32'b00000000000000000100001101010110;
assign LUT_1[33701] = 32'b11111111111111111101011111010010;
assign LUT_1[33702] = 32'b11111111111111111111111011100111;
assign LUT_1[33703] = 32'b11111111111111111001001101100011;
assign LUT_1[33704] = 32'b11111111111111111011100001110100;
assign LUT_1[33705] = 32'b11111111111111110100110011110000;
assign LUT_1[33706] = 32'b11111111111111110111010000000101;
assign LUT_1[33707] = 32'b11111111111111110000100010000001;
assign LUT_1[33708] = 32'b00000000000000000011011011001011;
assign LUT_1[33709] = 32'b11111111111111111100101101000111;
assign LUT_1[33710] = 32'b11111111111111111111001001011100;
assign LUT_1[33711] = 32'b11111111111111111000011011011000;
assign LUT_1[33712] = 32'b11111111111111111110001111100001;
assign LUT_1[33713] = 32'b11111111111111110111100001011101;
assign LUT_1[33714] = 32'b11111111111111111001111101110010;
assign LUT_1[33715] = 32'b11111111111111110011001111101110;
assign LUT_1[33716] = 32'b00000000000000000110001000111000;
assign LUT_1[33717] = 32'b11111111111111111111011010110100;
assign LUT_1[33718] = 32'b00000000000000000001110111001001;
assign LUT_1[33719] = 32'b11111111111111111011001001000101;
assign LUT_1[33720] = 32'b11111111111111111101011101010110;
assign LUT_1[33721] = 32'b11111111111111110110101111010010;
assign LUT_1[33722] = 32'b11111111111111111001001011100111;
assign LUT_1[33723] = 32'b11111111111111110010011101100011;
assign LUT_1[33724] = 32'b00000000000000000101010110101101;
assign LUT_1[33725] = 32'b11111111111111111110101000101001;
assign LUT_1[33726] = 32'b00000000000000000001000100111110;
assign LUT_1[33727] = 32'b11111111111111111010010110111010;
assign LUT_1[33728] = 32'b11111111111111111101010110101000;
assign LUT_1[33729] = 32'b11111111111111110110101000100100;
assign LUT_1[33730] = 32'b11111111111111111001000100111001;
assign LUT_1[33731] = 32'b11111111111111110010010110110101;
assign LUT_1[33732] = 32'b00000000000000000101001111111111;
assign LUT_1[33733] = 32'b11111111111111111110100001111011;
assign LUT_1[33734] = 32'b00000000000000000000111110010000;
assign LUT_1[33735] = 32'b11111111111111111010010000001100;
assign LUT_1[33736] = 32'b11111111111111111100100100011101;
assign LUT_1[33737] = 32'b11111111111111110101110110011001;
assign LUT_1[33738] = 32'b11111111111111111000010010101110;
assign LUT_1[33739] = 32'b11111111111111110001100100101010;
assign LUT_1[33740] = 32'b00000000000000000100011101110100;
assign LUT_1[33741] = 32'b11111111111111111101101111110000;
assign LUT_1[33742] = 32'b00000000000000000000001100000101;
assign LUT_1[33743] = 32'b11111111111111111001011110000001;
assign LUT_1[33744] = 32'b11111111111111111111010010001010;
assign LUT_1[33745] = 32'b11111111111111111000100100000110;
assign LUT_1[33746] = 32'b11111111111111111011000000011011;
assign LUT_1[33747] = 32'b11111111111111110100010010010111;
assign LUT_1[33748] = 32'b00000000000000000111001011100001;
assign LUT_1[33749] = 32'b00000000000000000000011101011101;
assign LUT_1[33750] = 32'b00000000000000000010111001110010;
assign LUT_1[33751] = 32'b11111111111111111100001011101110;
assign LUT_1[33752] = 32'b11111111111111111110011111111111;
assign LUT_1[33753] = 32'b11111111111111110111110001111011;
assign LUT_1[33754] = 32'b11111111111111111010001110010000;
assign LUT_1[33755] = 32'b11111111111111110011100000001100;
assign LUT_1[33756] = 32'b00000000000000000110011001010110;
assign LUT_1[33757] = 32'b11111111111111111111101011010010;
assign LUT_1[33758] = 32'b00000000000000000010000111100111;
assign LUT_1[33759] = 32'b11111111111111111011011001100011;
assign LUT_1[33760] = 32'b11111111111111111110010001100111;
assign LUT_1[33761] = 32'b11111111111111110111100011100011;
assign LUT_1[33762] = 32'b11111111111111111001111111111000;
assign LUT_1[33763] = 32'b11111111111111110011010001110100;
assign LUT_1[33764] = 32'b00000000000000000110001010111110;
assign LUT_1[33765] = 32'b11111111111111111111011100111010;
assign LUT_1[33766] = 32'b00000000000000000001111001001111;
assign LUT_1[33767] = 32'b11111111111111111011001011001011;
assign LUT_1[33768] = 32'b11111111111111111101011111011100;
assign LUT_1[33769] = 32'b11111111111111110110110001011000;
assign LUT_1[33770] = 32'b11111111111111111001001101101101;
assign LUT_1[33771] = 32'b11111111111111110010011111101001;
assign LUT_1[33772] = 32'b00000000000000000101011000110011;
assign LUT_1[33773] = 32'b11111111111111111110101010101111;
assign LUT_1[33774] = 32'b00000000000000000001000111000100;
assign LUT_1[33775] = 32'b11111111111111111010011001000000;
assign LUT_1[33776] = 32'b00000000000000000000001101001001;
assign LUT_1[33777] = 32'b11111111111111111001011111000101;
assign LUT_1[33778] = 32'b11111111111111111011111011011010;
assign LUT_1[33779] = 32'b11111111111111110101001101010110;
assign LUT_1[33780] = 32'b00000000000000001000000110100000;
assign LUT_1[33781] = 32'b00000000000000000001011000011100;
assign LUT_1[33782] = 32'b00000000000000000011110100110001;
assign LUT_1[33783] = 32'b11111111111111111101000110101101;
assign LUT_1[33784] = 32'b11111111111111111111011010111110;
assign LUT_1[33785] = 32'b11111111111111111000101100111010;
assign LUT_1[33786] = 32'b11111111111111111011001001001111;
assign LUT_1[33787] = 32'b11111111111111110100011011001011;
assign LUT_1[33788] = 32'b00000000000000000111010100010101;
assign LUT_1[33789] = 32'b00000000000000000000100110010001;
assign LUT_1[33790] = 32'b00000000000000000011000010100110;
assign LUT_1[33791] = 32'b11111111111111111100010100100010;
assign LUT_1[33792] = 32'b00000000000000000111001101000100;
assign LUT_1[33793] = 32'b00000000000000000000011111000000;
assign LUT_1[33794] = 32'b00000000000000000010111011010101;
assign LUT_1[33795] = 32'b11111111111111111100001101010001;
assign LUT_1[33796] = 32'b00000000000000001111000110011011;
assign LUT_1[33797] = 32'b00000000000000001000011000010111;
assign LUT_1[33798] = 32'b00000000000000001010110100101100;
assign LUT_1[33799] = 32'b00000000000000000100000110101000;
assign LUT_1[33800] = 32'b00000000000000000110011010111001;
assign LUT_1[33801] = 32'b11111111111111111111101100110101;
assign LUT_1[33802] = 32'b00000000000000000010001001001010;
assign LUT_1[33803] = 32'b11111111111111111011011011000110;
assign LUT_1[33804] = 32'b00000000000000001110010100010000;
assign LUT_1[33805] = 32'b00000000000000000111100110001100;
assign LUT_1[33806] = 32'b00000000000000001010000010100001;
assign LUT_1[33807] = 32'b00000000000000000011010100011101;
assign LUT_1[33808] = 32'b00000000000000001001001000100110;
assign LUT_1[33809] = 32'b00000000000000000010011010100010;
assign LUT_1[33810] = 32'b00000000000000000100110110110111;
assign LUT_1[33811] = 32'b11111111111111111110001000110011;
assign LUT_1[33812] = 32'b00000000000000010001000001111101;
assign LUT_1[33813] = 32'b00000000000000001010010011111001;
assign LUT_1[33814] = 32'b00000000000000001100110000001110;
assign LUT_1[33815] = 32'b00000000000000000110000010001010;
assign LUT_1[33816] = 32'b00000000000000001000010110011011;
assign LUT_1[33817] = 32'b00000000000000000001101000010111;
assign LUT_1[33818] = 32'b00000000000000000100000100101100;
assign LUT_1[33819] = 32'b11111111111111111101010110101000;
assign LUT_1[33820] = 32'b00000000000000010000001111110010;
assign LUT_1[33821] = 32'b00000000000000001001100001101110;
assign LUT_1[33822] = 32'b00000000000000001011111110000011;
assign LUT_1[33823] = 32'b00000000000000000101001111111111;
assign LUT_1[33824] = 32'b00000000000000001000001000000011;
assign LUT_1[33825] = 32'b00000000000000000001011001111111;
assign LUT_1[33826] = 32'b00000000000000000011110110010100;
assign LUT_1[33827] = 32'b11111111111111111101001000010000;
assign LUT_1[33828] = 32'b00000000000000010000000001011010;
assign LUT_1[33829] = 32'b00000000000000001001010011010110;
assign LUT_1[33830] = 32'b00000000000000001011101111101011;
assign LUT_1[33831] = 32'b00000000000000000101000001100111;
assign LUT_1[33832] = 32'b00000000000000000111010101111000;
assign LUT_1[33833] = 32'b00000000000000000000100111110100;
assign LUT_1[33834] = 32'b00000000000000000011000100001001;
assign LUT_1[33835] = 32'b11111111111111111100010110000101;
assign LUT_1[33836] = 32'b00000000000000001111001111001111;
assign LUT_1[33837] = 32'b00000000000000001000100001001011;
assign LUT_1[33838] = 32'b00000000000000001010111101100000;
assign LUT_1[33839] = 32'b00000000000000000100001111011100;
assign LUT_1[33840] = 32'b00000000000000001010000011100101;
assign LUT_1[33841] = 32'b00000000000000000011010101100001;
assign LUT_1[33842] = 32'b00000000000000000101110001110110;
assign LUT_1[33843] = 32'b11111111111111111111000011110010;
assign LUT_1[33844] = 32'b00000000000000010001111100111100;
assign LUT_1[33845] = 32'b00000000000000001011001110111000;
assign LUT_1[33846] = 32'b00000000000000001101101011001101;
assign LUT_1[33847] = 32'b00000000000000000110111101001001;
assign LUT_1[33848] = 32'b00000000000000001001010001011010;
assign LUT_1[33849] = 32'b00000000000000000010100011010110;
assign LUT_1[33850] = 32'b00000000000000000100111111101011;
assign LUT_1[33851] = 32'b11111111111111111110010001100111;
assign LUT_1[33852] = 32'b00000000000000010001001010110001;
assign LUT_1[33853] = 32'b00000000000000001010011100101101;
assign LUT_1[33854] = 32'b00000000000000001100111001000010;
assign LUT_1[33855] = 32'b00000000000000000110001010111110;
assign LUT_1[33856] = 32'b00000000000000001001001010101100;
assign LUT_1[33857] = 32'b00000000000000000010011100101000;
assign LUT_1[33858] = 32'b00000000000000000100111000111101;
assign LUT_1[33859] = 32'b11111111111111111110001010111001;
assign LUT_1[33860] = 32'b00000000000000010001000100000011;
assign LUT_1[33861] = 32'b00000000000000001010010101111111;
assign LUT_1[33862] = 32'b00000000000000001100110010010100;
assign LUT_1[33863] = 32'b00000000000000000110000100010000;
assign LUT_1[33864] = 32'b00000000000000001000011000100001;
assign LUT_1[33865] = 32'b00000000000000000001101010011101;
assign LUT_1[33866] = 32'b00000000000000000100000110110010;
assign LUT_1[33867] = 32'b11111111111111111101011000101110;
assign LUT_1[33868] = 32'b00000000000000010000010001111000;
assign LUT_1[33869] = 32'b00000000000000001001100011110100;
assign LUT_1[33870] = 32'b00000000000000001100000000001001;
assign LUT_1[33871] = 32'b00000000000000000101010010000101;
assign LUT_1[33872] = 32'b00000000000000001011000110001110;
assign LUT_1[33873] = 32'b00000000000000000100011000001010;
assign LUT_1[33874] = 32'b00000000000000000110110100011111;
assign LUT_1[33875] = 32'b00000000000000000000000110011011;
assign LUT_1[33876] = 32'b00000000000000010010111111100101;
assign LUT_1[33877] = 32'b00000000000000001100010001100001;
assign LUT_1[33878] = 32'b00000000000000001110101101110110;
assign LUT_1[33879] = 32'b00000000000000000111111111110010;
assign LUT_1[33880] = 32'b00000000000000001010010100000011;
assign LUT_1[33881] = 32'b00000000000000000011100101111111;
assign LUT_1[33882] = 32'b00000000000000000110000010010100;
assign LUT_1[33883] = 32'b11111111111111111111010100010000;
assign LUT_1[33884] = 32'b00000000000000010010001101011010;
assign LUT_1[33885] = 32'b00000000000000001011011111010110;
assign LUT_1[33886] = 32'b00000000000000001101111011101011;
assign LUT_1[33887] = 32'b00000000000000000111001101100111;
assign LUT_1[33888] = 32'b00000000000000001010000101101011;
assign LUT_1[33889] = 32'b00000000000000000011010111100111;
assign LUT_1[33890] = 32'b00000000000000000101110011111100;
assign LUT_1[33891] = 32'b11111111111111111111000101111000;
assign LUT_1[33892] = 32'b00000000000000010001111111000010;
assign LUT_1[33893] = 32'b00000000000000001011010000111110;
assign LUT_1[33894] = 32'b00000000000000001101101101010011;
assign LUT_1[33895] = 32'b00000000000000000110111111001111;
assign LUT_1[33896] = 32'b00000000000000001001010011100000;
assign LUT_1[33897] = 32'b00000000000000000010100101011100;
assign LUT_1[33898] = 32'b00000000000000000101000001110001;
assign LUT_1[33899] = 32'b11111111111111111110010011101101;
assign LUT_1[33900] = 32'b00000000000000010001001100110111;
assign LUT_1[33901] = 32'b00000000000000001010011110110011;
assign LUT_1[33902] = 32'b00000000000000001100111011001000;
assign LUT_1[33903] = 32'b00000000000000000110001101000100;
assign LUT_1[33904] = 32'b00000000000000001100000001001101;
assign LUT_1[33905] = 32'b00000000000000000101010011001001;
assign LUT_1[33906] = 32'b00000000000000000111101111011110;
assign LUT_1[33907] = 32'b00000000000000000001000001011010;
assign LUT_1[33908] = 32'b00000000000000010011111010100100;
assign LUT_1[33909] = 32'b00000000000000001101001100100000;
assign LUT_1[33910] = 32'b00000000000000001111101000110101;
assign LUT_1[33911] = 32'b00000000000000001000111010110001;
assign LUT_1[33912] = 32'b00000000000000001011001111000010;
assign LUT_1[33913] = 32'b00000000000000000100100000111110;
assign LUT_1[33914] = 32'b00000000000000000110111101010011;
assign LUT_1[33915] = 32'b00000000000000000000001111001111;
assign LUT_1[33916] = 32'b00000000000000010011001000011001;
assign LUT_1[33917] = 32'b00000000000000001100011010010101;
assign LUT_1[33918] = 32'b00000000000000001110110110101010;
assign LUT_1[33919] = 32'b00000000000000001000001000100110;
assign LUT_1[33920] = 32'b00000000000000001010001101000111;
assign LUT_1[33921] = 32'b00000000000000000011011111000011;
assign LUT_1[33922] = 32'b00000000000000000101111011011000;
assign LUT_1[33923] = 32'b11111111111111111111001101010100;
assign LUT_1[33924] = 32'b00000000000000010010000110011110;
assign LUT_1[33925] = 32'b00000000000000001011011000011010;
assign LUT_1[33926] = 32'b00000000000000001101110100101111;
assign LUT_1[33927] = 32'b00000000000000000111000110101011;
assign LUT_1[33928] = 32'b00000000000000001001011010111100;
assign LUT_1[33929] = 32'b00000000000000000010101100111000;
assign LUT_1[33930] = 32'b00000000000000000101001001001101;
assign LUT_1[33931] = 32'b11111111111111111110011011001001;
assign LUT_1[33932] = 32'b00000000000000010001010100010011;
assign LUT_1[33933] = 32'b00000000000000001010100110001111;
assign LUT_1[33934] = 32'b00000000000000001101000010100100;
assign LUT_1[33935] = 32'b00000000000000000110010100100000;
assign LUT_1[33936] = 32'b00000000000000001100001000101001;
assign LUT_1[33937] = 32'b00000000000000000101011010100101;
assign LUT_1[33938] = 32'b00000000000000000111110110111010;
assign LUT_1[33939] = 32'b00000000000000000001001000110110;
assign LUT_1[33940] = 32'b00000000000000010100000010000000;
assign LUT_1[33941] = 32'b00000000000000001101010011111100;
assign LUT_1[33942] = 32'b00000000000000001111110000010001;
assign LUT_1[33943] = 32'b00000000000000001001000010001101;
assign LUT_1[33944] = 32'b00000000000000001011010110011110;
assign LUT_1[33945] = 32'b00000000000000000100101000011010;
assign LUT_1[33946] = 32'b00000000000000000111000100101111;
assign LUT_1[33947] = 32'b00000000000000000000010110101011;
assign LUT_1[33948] = 32'b00000000000000010011001111110101;
assign LUT_1[33949] = 32'b00000000000000001100100001110001;
assign LUT_1[33950] = 32'b00000000000000001110111110000110;
assign LUT_1[33951] = 32'b00000000000000001000010000000010;
assign LUT_1[33952] = 32'b00000000000000001011001000000110;
assign LUT_1[33953] = 32'b00000000000000000100011010000010;
assign LUT_1[33954] = 32'b00000000000000000110110110010111;
assign LUT_1[33955] = 32'b00000000000000000000001000010011;
assign LUT_1[33956] = 32'b00000000000000010011000001011101;
assign LUT_1[33957] = 32'b00000000000000001100010011011001;
assign LUT_1[33958] = 32'b00000000000000001110101111101110;
assign LUT_1[33959] = 32'b00000000000000001000000001101010;
assign LUT_1[33960] = 32'b00000000000000001010010101111011;
assign LUT_1[33961] = 32'b00000000000000000011100111110111;
assign LUT_1[33962] = 32'b00000000000000000110000100001100;
assign LUT_1[33963] = 32'b11111111111111111111010110001000;
assign LUT_1[33964] = 32'b00000000000000010010001111010010;
assign LUT_1[33965] = 32'b00000000000000001011100001001110;
assign LUT_1[33966] = 32'b00000000000000001101111101100011;
assign LUT_1[33967] = 32'b00000000000000000111001111011111;
assign LUT_1[33968] = 32'b00000000000000001101000011101000;
assign LUT_1[33969] = 32'b00000000000000000110010101100100;
assign LUT_1[33970] = 32'b00000000000000001000110001111001;
assign LUT_1[33971] = 32'b00000000000000000010000011110101;
assign LUT_1[33972] = 32'b00000000000000010100111100111111;
assign LUT_1[33973] = 32'b00000000000000001110001110111011;
assign LUT_1[33974] = 32'b00000000000000010000101011010000;
assign LUT_1[33975] = 32'b00000000000000001001111101001100;
assign LUT_1[33976] = 32'b00000000000000001100010001011101;
assign LUT_1[33977] = 32'b00000000000000000101100011011001;
assign LUT_1[33978] = 32'b00000000000000000111111111101110;
assign LUT_1[33979] = 32'b00000000000000000001010001101010;
assign LUT_1[33980] = 32'b00000000000000010100001010110100;
assign LUT_1[33981] = 32'b00000000000000001101011100110000;
assign LUT_1[33982] = 32'b00000000000000001111111001000101;
assign LUT_1[33983] = 32'b00000000000000001001001011000001;
assign LUT_1[33984] = 32'b00000000000000001100001010101111;
assign LUT_1[33985] = 32'b00000000000000000101011100101011;
assign LUT_1[33986] = 32'b00000000000000000111111001000000;
assign LUT_1[33987] = 32'b00000000000000000001001010111100;
assign LUT_1[33988] = 32'b00000000000000010100000100000110;
assign LUT_1[33989] = 32'b00000000000000001101010110000010;
assign LUT_1[33990] = 32'b00000000000000001111110010010111;
assign LUT_1[33991] = 32'b00000000000000001001000100010011;
assign LUT_1[33992] = 32'b00000000000000001011011000100100;
assign LUT_1[33993] = 32'b00000000000000000100101010100000;
assign LUT_1[33994] = 32'b00000000000000000111000110110101;
assign LUT_1[33995] = 32'b00000000000000000000011000110001;
assign LUT_1[33996] = 32'b00000000000000010011010001111011;
assign LUT_1[33997] = 32'b00000000000000001100100011110111;
assign LUT_1[33998] = 32'b00000000000000001111000000001100;
assign LUT_1[33999] = 32'b00000000000000001000010010001000;
assign LUT_1[34000] = 32'b00000000000000001110000110010001;
assign LUT_1[34001] = 32'b00000000000000000111011000001101;
assign LUT_1[34002] = 32'b00000000000000001001110100100010;
assign LUT_1[34003] = 32'b00000000000000000011000110011110;
assign LUT_1[34004] = 32'b00000000000000010101111111101000;
assign LUT_1[34005] = 32'b00000000000000001111010001100100;
assign LUT_1[34006] = 32'b00000000000000010001101101111001;
assign LUT_1[34007] = 32'b00000000000000001010111111110101;
assign LUT_1[34008] = 32'b00000000000000001101010100000110;
assign LUT_1[34009] = 32'b00000000000000000110100110000010;
assign LUT_1[34010] = 32'b00000000000000001001000010010111;
assign LUT_1[34011] = 32'b00000000000000000010010100010011;
assign LUT_1[34012] = 32'b00000000000000010101001101011101;
assign LUT_1[34013] = 32'b00000000000000001110011111011001;
assign LUT_1[34014] = 32'b00000000000000010000111011101110;
assign LUT_1[34015] = 32'b00000000000000001010001101101010;
assign LUT_1[34016] = 32'b00000000000000001101000101101110;
assign LUT_1[34017] = 32'b00000000000000000110010111101010;
assign LUT_1[34018] = 32'b00000000000000001000110011111111;
assign LUT_1[34019] = 32'b00000000000000000010000101111011;
assign LUT_1[34020] = 32'b00000000000000010100111111000101;
assign LUT_1[34021] = 32'b00000000000000001110010001000001;
assign LUT_1[34022] = 32'b00000000000000010000101101010110;
assign LUT_1[34023] = 32'b00000000000000001001111111010010;
assign LUT_1[34024] = 32'b00000000000000001100010011100011;
assign LUT_1[34025] = 32'b00000000000000000101100101011111;
assign LUT_1[34026] = 32'b00000000000000001000000001110100;
assign LUT_1[34027] = 32'b00000000000000000001010011110000;
assign LUT_1[34028] = 32'b00000000000000010100001100111010;
assign LUT_1[34029] = 32'b00000000000000001101011110110110;
assign LUT_1[34030] = 32'b00000000000000001111111011001011;
assign LUT_1[34031] = 32'b00000000000000001001001101000111;
assign LUT_1[34032] = 32'b00000000000000001111000001010000;
assign LUT_1[34033] = 32'b00000000000000001000010011001100;
assign LUT_1[34034] = 32'b00000000000000001010101111100001;
assign LUT_1[34035] = 32'b00000000000000000100000001011101;
assign LUT_1[34036] = 32'b00000000000000010110111010100111;
assign LUT_1[34037] = 32'b00000000000000010000001100100011;
assign LUT_1[34038] = 32'b00000000000000010010101000111000;
assign LUT_1[34039] = 32'b00000000000000001011111010110100;
assign LUT_1[34040] = 32'b00000000000000001110001111000101;
assign LUT_1[34041] = 32'b00000000000000000111100001000001;
assign LUT_1[34042] = 32'b00000000000000001001111101010110;
assign LUT_1[34043] = 32'b00000000000000000011001111010010;
assign LUT_1[34044] = 32'b00000000000000010110001000011100;
assign LUT_1[34045] = 32'b00000000000000001111011010011000;
assign LUT_1[34046] = 32'b00000000000000010001110110101101;
assign LUT_1[34047] = 32'b00000000000000001011001000101001;
assign LUT_1[34048] = 32'b00000000000000000101000001010000;
assign LUT_1[34049] = 32'b11111111111111111110010011001100;
assign LUT_1[34050] = 32'b00000000000000000000101111100001;
assign LUT_1[34051] = 32'b11111111111111111010000001011101;
assign LUT_1[34052] = 32'b00000000000000001100111010100111;
assign LUT_1[34053] = 32'b00000000000000000110001100100011;
assign LUT_1[34054] = 32'b00000000000000001000101000111000;
assign LUT_1[34055] = 32'b00000000000000000001111010110100;
assign LUT_1[34056] = 32'b00000000000000000100001111000101;
assign LUT_1[34057] = 32'b11111111111111111101100001000001;
assign LUT_1[34058] = 32'b11111111111111111111111101010110;
assign LUT_1[34059] = 32'b11111111111111111001001111010010;
assign LUT_1[34060] = 32'b00000000000000001100001000011100;
assign LUT_1[34061] = 32'b00000000000000000101011010011000;
assign LUT_1[34062] = 32'b00000000000000000111110110101101;
assign LUT_1[34063] = 32'b00000000000000000001001000101001;
assign LUT_1[34064] = 32'b00000000000000000110111100110010;
assign LUT_1[34065] = 32'b00000000000000000000001110101110;
assign LUT_1[34066] = 32'b00000000000000000010101011000011;
assign LUT_1[34067] = 32'b11111111111111111011111100111111;
assign LUT_1[34068] = 32'b00000000000000001110110110001001;
assign LUT_1[34069] = 32'b00000000000000001000001000000101;
assign LUT_1[34070] = 32'b00000000000000001010100100011010;
assign LUT_1[34071] = 32'b00000000000000000011110110010110;
assign LUT_1[34072] = 32'b00000000000000000110001010100111;
assign LUT_1[34073] = 32'b11111111111111111111011100100011;
assign LUT_1[34074] = 32'b00000000000000000001111000111000;
assign LUT_1[34075] = 32'b11111111111111111011001010110100;
assign LUT_1[34076] = 32'b00000000000000001110000011111110;
assign LUT_1[34077] = 32'b00000000000000000111010101111010;
assign LUT_1[34078] = 32'b00000000000000001001110010001111;
assign LUT_1[34079] = 32'b00000000000000000011000100001011;
assign LUT_1[34080] = 32'b00000000000000000101111100001111;
assign LUT_1[34081] = 32'b11111111111111111111001110001011;
assign LUT_1[34082] = 32'b00000000000000000001101010100000;
assign LUT_1[34083] = 32'b11111111111111111010111100011100;
assign LUT_1[34084] = 32'b00000000000000001101110101100110;
assign LUT_1[34085] = 32'b00000000000000000111000111100010;
assign LUT_1[34086] = 32'b00000000000000001001100011110111;
assign LUT_1[34087] = 32'b00000000000000000010110101110011;
assign LUT_1[34088] = 32'b00000000000000000101001010000100;
assign LUT_1[34089] = 32'b11111111111111111110011100000000;
assign LUT_1[34090] = 32'b00000000000000000000111000010101;
assign LUT_1[34091] = 32'b11111111111111111010001010010001;
assign LUT_1[34092] = 32'b00000000000000001101000011011011;
assign LUT_1[34093] = 32'b00000000000000000110010101010111;
assign LUT_1[34094] = 32'b00000000000000001000110001101100;
assign LUT_1[34095] = 32'b00000000000000000010000011101000;
assign LUT_1[34096] = 32'b00000000000000000111110111110001;
assign LUT_1[34097] = 32'b00000000000000000001001001101101;
assign LUT_1[34098] = 32'b00000000000000000011100110000010;
assign LUT_1[34099] = 32'b11111111111111111100110111111110;
assign LUT_1[34100] = 32'b00000000000000001111110001001000;
assign LUT_1[34101] = 32'b00000000000000001001000011000100;
assign LUT_1[34102] = 32'b00000000000000001011011111011001;
assign LUT_1[34103] = 32'b00000000000000000100110001010101;
assign LUT_1[34104] = 32'b00000000000000000111000101100110;
assign LUT_1[34105] = 32'b00000000000000000000010111100010;
assign LUT_1[34106] = 32'b00000000000000000010110011110111;
assign LUT_1[34107] = 32'b11111111111111111100000101110011;
assign LUT_1[34108] = 32'b00000000000000001110111110111101;
assign LUT_1[34109] = 32'b00000000000000001000010000111001;
assign LUT_1[34110] = 32'b00000000000000001010101101001110;
assign LUT_1[34111] = 32'b00000000000000000011111111001010;
assign LUT_1[34112] = 32'b00000000000000000110111110111000;
assign LUT_1[34113] = 32'b00000000000000000000010000110100;
assign LUT_1[34114] = 32'b00000000000000000010101101001001;
assign LUT_1[34115] = 32'b11111111111111111011111111000101;
assign LUT_1[34116] = 32'b00000000000000001110111000001111;
assign LUT_1[34117] = 32'b00000000000000001000001010001011;
assign LUT_1[34118] = 32'b00000000000000001010100110100000;
assign LUT_1[34119] = 32'b00000000000000000011111000011100;
assign LUT_1[34120] = 32'b00000000000000000110001100101101;
assign LUT_1[34121] = 32'b11111111111111111111011110101001;
assign LUT_1[34122] = 32'b00000000000000000001111010111110;
assign LUT_1[34123] = 32'b11111111111111111011001100111010;
assign LUT_1[34124] = 32'b00000000000000001110000110000100;
assign LUT_1[34125] = 32'b00000000000000000111011000000000;
assign LUT_1[34126] = 32'b00000000000000001001110100010101;
assign LUT_1[34127] = 32'b00000000000000000011000110010001;
assign LUT_1[34128] = 32'b00000000000000001000111010011010;
assign LUT_1[34129] = 32'b00000000000000000010001100010110;
assign LUT_1[34130] = 32'b00000000000000000100101000101011;
assign LUT_1[34131] = 32'b11111111111111111101111010100111;
assign LUT_1[34132] = 32'b00000000000000010000110011110001;
assign LUT_1[34133] = 32'b00000000000000001010000101101101;
assign LUT_1[34134] = 32'b00000000000000001100100010000010;
assign LUT_1[34135] = 32'b00000000000000000101110011111110;
assign LUT_1[34136] = 32'b00000000000000001000001000001111;
assign LUT_1[34137] = 32'b00000000000000000001011010001011;
assign LUT_1[34138] = 32'b00000000000000000011110110100000;
assign LUT_1[34139] = 32'b11111111111111111101001000011100;
assign LUT_1[34140] = 32'b00000000000000010000000001100110;
assign LUT_1[34141] = 32'b00000000000000001001010011100010;
assign LUT_1[34142] = 32'b00000000000000001011101111110111;
assign LUT_1[34143] = 32'b00000000000000000101000001110011;
assign LUT_1[34144] = 32'b00000000000000000111111001110111;
assign LUT_1[34145] = 32'b00000000000000000001001011110011;
assign LUT_1[34146] = 32'b00000000000000000011101000001000;
assign LUT_1[34147] = 32'b11111111111111111100111010000100;
assign LUT_1[34148] = 32'b00000000000000001111110011001110;
assign LUT_1[34149] = 32'b00000000000000001001000101001010;
assign LUT_1[34150] = 32'b00000000000000001011100001011111;
assign LUT_1[34151] = 32'b00000000000000000100110011011011;
assign LUT_1[34152] = 32'b00000000000000000111000111101100;
assign LUT_1[34153] = 32'b00000000000000000000011001101000;
assign LUT_1[34154] = 32'b00000000000000000010110101111101;
assign LUT_1[34155] = 32'b11111111111111111100000111111001;
assign LUT_1[34156] = 32'b00000000000000001111000001000011;
assign LUT_1[34157] = 32'b00000000000000001000010010111111;
assign LUT_1[34158] = 32'b00000000000000001010101111010100;
assign LUT_1[34159] = 32'b00000000000000000100000001010000;
assign LUT_1[34160] = 32'b00000000000000001001110101011001;
assign LUT_1[34161] = 32'b00000000000000000011000111010101;
assign LUT_1[34162] = 32'b00000000000000000101100011101010;
assign LUT_1[34163] = 32'b11111111111111111110110101100110;
assign LUT_1[34164] = 32'b00000000000000010001101110110000;
assign LUT_1[34165] = 32'b00000000000000001011000000101100;
assign LUT_1[34166] = 32'b00000000000000001101011101000001;
assign LUT_1[34167] = 32'b00000000000000000110101110111101;
assign LUT_1[34168] = 32'b00000000000000001001000011001110;
assign LUT_1[34169] = 32'b00000000000000000010010101001010;
assign LUT_1[34170] = 32'b00000000000000000100110001011111;
assign LUT_1[34171] = 32'b11111111111111111110000011011011;
assign LUT_1[34172] = 32'b00000000000000010000111100100101;
assign LUT_1[34173] = 32'b00000000000000001010001110100001;
assign LUT_1[34174] = 32'b00000000000000001100101010110110;
assign LUT_1[34175] = 32'b00000000000000000101111100110010;
assign LUT_1[34176] = 32'b00000000000000001000000001010011;
assign LUT_1[34177] = 32'b00000000000000000001010011001111;
assign LUT_1[34178] = 32'b00000000000000000011101111100100;
assign LUT_1[34179] = 32'b11111111111111111101000001100000;
assign LUT_1[34180] = 32'b00000000000000001111111010101010;
assign LUT_1[34181] = 32'b00000000000000001001001100100110;
assign LUT_1[34182] = 32'b00000000000000001011101000111011;
assign LUT_1[34183] = 32'b00000000000000000100111010110111;
assign LUT_1[34184] = 32'b00000000000000000111001111001000;
assign LUT_1[34185] = 32'b00000000000000000000100001000100;
assign LUT_1[34186] = 32'b00000000000000000010111101011001;
assign LUT_1[34187] = 32'b11111111111111111100001111010101;
assign LUT_1[34188] = 32'b00000000000000001111001000011111;
assign LUT_1[34189] = 32'b00000000000000001000011010011011;
assign LUT_1[34190] = 32'b00000000000000001010110110110000;
assign LUT_1[34191] = 32'b00000000000000000100001000101100;
assign LUT_1[34192] = 32'b00000000000000001001111100110101;
assign LUT_1[34193] = 32'b00000000000000000011001110110001;
assign LUT_1[34194] = 32'b00000000000000000101101011000110;
assign LUT_1[34195] = 32'b11111111111111111110111101000010;
assign LUT_1[34196] = 32'b00000000000000010001110110001100;
assign LUT_1[34197] = 32'b00000000000000001011001000001000;
assign LUT_1[34198] = 32'b00000000000000001101100100011101;
assign LUT_1[34199] = 32'b00000000000000000110110110011001;
assign LUT_1[34200] = 32'b00000000000000001001001010101010;
assign LUT_1[34201] = 32'b00000000000000000010011100100110;
assign LUT_1[34202] = 32'b00000000000000000100111000111011;
assign LUT_1[34203] = 32'b11111111111111111110001010110111;
assign LUT_1[34204] = 32'b00000000000000010001000100000001;
assign LUT_1[34205] = 32'b00000000000000001010010101111101;
assign LUT_1[34206] = 32'b00000000000000001100110010010010;
assign LUT_1[34207] = 32'b00000000000000000110000100001110;
assign LUT_1[34208] = 32'b00000000000000001000111100010010;
assign LUT_1[34209] = 32'b00000000000000000010001110001110;
assign LUT_1[34210] = 32'b00000000000000000100101010100011;
assign LUT_1[34211] = 32'b11111111111111111101111100011111;
assign LUT_1[34212] = 32'b00000000000000010000110101101001;
assign LUT_1[34213] = 32'b00000000000000001010000111100101;
assign LUT_1[34214] = 32'b00000000000000001100100011111010;
assign LUT_1[34215] = 32'b00000000000000000101110101110110;
assign LUT_1[34216] = 32'b00000000000000001000001010000111;
assign LUT_1[34217] = 32'b00000000000000000001011100000011;
assign LUT_1[34218] = 32'b00000000000000000011111000011000;
assign LUT_1[34219] = 32'b11111111111111111101001010010100;
assign LUT_1[34220] = 32'b00000000000000010000000011011110;
assign LUT_1[34221] = 32'b00000000000000001001010101011010;
assign LUT_1[34222] = 32'b00000000000000001011110001101111;
assign LUT_1[34223] = 32'b00000000000000000101000011101011;
assign LUT_1[34224] = 32'b00000000000000001010110111110100;
assign LUT_1[34225] = 32'b00000000000000000100001001110000;
assign LUT_1[34226] = 32'b00000000000000000110100110000101;
assign LUT_1[34227] = 32'b11111111111111111111111000000001;
assign LUT_1[34228] = 32'b00000000000000010010110001001011;
assign LUT_1[34229] = 32'b00000000000000001100000011000111;
assign LUT_1[34230] = 32'b00000000000000001110011111011100;
assign LUT_1[34231] = 32'b00000000000000000111110001011000;
assign LUT_1[34232] = 32'b00000000000000001010000101101001;
assign LUT_1[34233] = 32'b00000000000000000011010111100101;
assign LUT_1[34234] = 32'b00000000000000000101110011111010;
assign LUT_1[34235] = 32'b11111111111111111111000101110110;
assign LUT_1[34236] = 32'b00000000000000010001111111000000;
assign LUT_1[34237] = 32'b00000000000000001011010000111100;
assign LUT_1[34238] = 32'b00000000000000001101101101010001;
assign LUT_1[34239] = 32'b00000000000000000110111111001101;
assign LUT_1[34240] = 32'b00000000000000001001111110111011;
assign LUT_1[34241] = 32'b00000000000000000011010000110111;
assign LUT_1[34242] = 32'b00000000000000000101101101001100;
assign LUT_1[34243] = 32'b11111111111111111110111111001000;
assign LUT_1[34244] = 32'b00000000000000010001111000010010;
assign LUT_1[34245] = 32'b00000000000000001011001010001110;
assign LUT_1[34246] = 32'b00000000000000001101100110100011;
assign LUT_1[34247] = 32'b00000000000000000110111000011111;
assign LUT_1[34248] = 32'b00000000000000001001001100110000;
assign LUT_1[34249] = 32'b00000000000000000010011110101100;
assign LUT_1[34250] = 32'b00000000000000000100111011000001;
assign LUT_1[34251] = 32'b11111111111111111110001100111101;
assign LUT_1[34252] = 32'b00000000000000010001000110000111;
assign LUT_1[34253] = 32'b00000000000000001010011000000011;
assign LUT_1[34254] = 32'b00000000000000001100110100011000;
assign LUT_1[34255] = 32'b00000000000000000110000110010100;
assign LUT_1[34256] = 32'b00000000000000001011111010011101;
assign LUT_1[34257] = 32'b00000000000000000101001100011001;
assign LUT_1[34258] = 32'b00000000000000000111101000101110;
assign LUT_1[34259] = 32'b00000000000000000000111010101010;
assign LUT_1[34260] = 32'b00000000000000010011110011110100;
assign LUT_1[34261] = 32'b00000000000000001101000101110000;
assign LUT_1[34262] = 32'b00000000000000001111100010000101;
assign LUT_1[34263] = 32'b00000000000000001000110100000001;
assign LUT_1[34264] = 32'b00000000000000001011001000010010;
assign LUT_1[34265] = 32'b00000000000000000100011010001110;
assign LUT_1[34266] = 32'b00000000000000000110110110100011;
assign LUT_1[34267] = 32'b00000000000000000000001000011111;
assign LUT_1[34268] = 32'b00000000000000010011000001101001;
assign LUT_1[34269] = 32'b00000000000000001100010011100101;
assign LUT_1[34270] = 32'b00000000000000001110101111111010;
assign LUT_1[34271] = 32'b00000000000000001000000001110110;
assign LUT_1[34272] = 32'b00000000000000001010111001111010;
assign LUT_1[34273] = 32'b00000000000000000100001011110110;
assign LUT_1[34274] = 32'b00000000000000000110101000001011;
assign LUT_1[34275] = 32'b11111111111111111111111010000111;
assign LUT_1[34276] = 32'b00000000000000010010110011010001;
assign LUT_1[34277] = 32'b00000000000000001100000101001101;
assign LUT_1[34278] = 32'b00000000000000001110100001100010;
assign LUT_1[34279] = 32'b00000000000000000111110011011110;
assign LUT_1[34280] = 32'b00000000000000001010000111101111;
assign LUT_1[34281] = 32'b00000000000000000011011001101011;
assign LUT_1[34282] = 32'b00000000000000000101110110000000;
assign LUT_1[34283] = 32'b11111111111111111111000111111100;
assign LUT_1[34284] = 32'b00000000000000010010000001000110;
assign LUT_1[34285] = 32'b00000000000000001011010011000010;
assign LUT_1[34286] = 32'b00000000000000001101101111010111;
assign LUT_1[34287] = 32'b00000000000000000111000001010011;
assign LUT_1[34288] = 32'b00000000000000001100110101011100;
assign LUT_1[34289] = 32'b00000000000000000110000111011000;
assign LUT_1[34290] = 32'b00000000000000001000100011101101;
assign LUT_1[34291] = 32'b00000000000000000001110101101001;
assign LUT_1[34292] = 32'b00000000000000010100101110110011;
assign LUT_1[34293] = 32'b00000000000000001110000000101111;
assign LUT_1[34294] = 32'b00000000000000010000011101000100;
assign LUT_1[34295] = 32'b00000000000000001001101111000000;
assign LUT_1[34296] = 32'b00000000000000001100000011010001;
assign LUT_1[34297] = 32'b00000000000000000101010101001101;
assign LUT_1[34298] = 32'b00000000000000000111110001100010;
assign LUT_1[34299] = 32'b00000000000000000001000011011110;
assign LUT_1[34300] = 32'b00000000000000010011111100101000;
assign LUT_1[34301] = 32'b00000000000000001101001110100100;
assign LUT_1[34302] = 32'b00000000000000001111101010111001;
assign LUT_1[34303] = 32'b00000000000000001000111100110101;
assign LUT_1[34304] = 32'b00000000000000000000111011100001;
assign LUT_1[34305] = 32'b11111111111111111010001101011101;
assign LUT_1[34306] = 32'b11111111111111111100101001110010;
assign LUT_1[34307] = 32'b11111111111111110101111011101110;
assign LUT_1[34308] = 32'b00000000000000001000110100111000;
assign LUT_1[34309] = 32'b00000000000000000010000110110100;
assign LUT_1[34310] = 32'b00000000000000000100100011001001;
assign LUT_1[34311] = 32'b11111111111111111101110101000101;
assign LUT_1[34312] = 32'b00000000000000000000001001010110;
assign LUT_1[34313] = 32'b11111111111111111001011011010010;
assign LUT_1[34314] = 32'b11111111111111111011110111100111;
assign LUT_1[34315] = 32'b11111111111111110101001001100011;
assign LUT_1[34316] = 32'b00000000000000001000000010101101;
assign LUT_1[34317] = 32'b00000000000000000001010100101001;
assign LUT_1[34318] = 32'b00000000000000000011110000111110;
assign LUT_1[34319] = 32'b11111111111111111101000010111010;
assign LUT_1[34320] = 32'b00000000000000000010110111000011;
assign LUT_1[34321] = 32'b11111111111111111100001000111111;
assign LUT_1[34322] = 32'b11111111111111111110100101010100;
assign LUT_1[34323] = 32'b11111111111111110111110111010000;
assign LUT_1[34324] = 32'b00000000000000001010110000011010;
assign LUT_1[34325] = 32'b00000000000000000100000010010110;
assign LUT_1[34326] = 32'b00000000000000000110011110101011;
assign LUT_1[34327] = 32'b11111111111111111111110000100111;
assign LUT_1[34328] = 32'b00000000000000000010000100111000;
assign LUT_1[34329] = 32'b11111111111111111011010110110100;
assign LUT_1[34330] = 32'b11111111111111111101110011001001;
assign LUT_1[34331] = 32'b11111111111111110111000101000101;
assign LUT_1[34332] = 32'b00000000000000001001111110001111;
assign LUT_1[34333] = 32'b00000000000000000011010000001011;
assign LUT_1[34334] = 32'b00000000000000000101101100100000;
assign LUT_1[34335] = 32'b11111111111111111110111110011100;
assign LUT_1[34336] = 32'b00000000000000000001110110100000;
assign LUT_1[34337] = 32'b11111111111111111011001000011100;
assign LUT_1[34338] = 32'b11111111111111111101100100110001;
assign LUT_1[34339] = 32'b11111111111111110110110110101101;
assign LUT_1[34340] = 32'b00000000000000001001101111110111;
assign LUT_1[34341] = 32'b00000000000000000011000001110011;
assign LUT_1[34342] = 32'b00000000000000000101011110001000;
assign LUT_1[34343] = 32'b11111111111111111110110000000100;
assign LUT_1[34344] = 32'b00000000000000000001000100010101;
assign LUT_1[34345] = 32'b11111111111111111010010110010001;
assign LUT_1[34346] = 32'b11111111111111111100110010100110;
assign LUT_1[34347] = 32'b11111111111111110110000100100010;
assign LUT_1[34348] = 32'b00000000000000001000111101101100;
assign LUT_1[34349] = 32'b00000000000000000010001111101000;
assign LUT_1[34350] = 32'b00000000000000000100101011111101;
assign LUT_1[34351] = 32'b11111111111111111101111101111001;
assign LUT_1[34352] = 32'b00000000000000000011110010000010;
assign LUT_1[34353] = 32'b11111111111111111101000011111110;
assign LUT_1[34354] = 32'b11111111111111111111100000010011;
assign LUT_1[34355] = 32'b11111111111111111000110010001111;
assign LUT_1[34356] = 32'b00000000000000001011101011011001;
assign LUT_1[34357] = 32'b00000000000000000100111101010101;
assign LUT_1[34358] = 32'b00000000000000000111011001101010;
assign LUT_1[34359] = 32'b00000000000000000000101011100110;
assign LUT_1[34360] = 32'b00000000000000000010111111110111;
assign LUT_1[34361] = 32'b11111111111111111100010001110011;
assign LUT_1[34362] = 32'b11111111111111111110101110001000;
assign LUT_1[34363] = 32'b11111111111111111000000000000100;
assign LUT_1[34364] = 32'b00000000000000001010111001001110;
assign LUT_1[34365] = 32'b00000000000000000100001011001010;
assign LUT_1[34366] = 32'b00000000000000000110100111011111;
assign LUT_1[34367] = 32'b11111111111111111111111001011011;
assign LUT_1[34368] = 32'b00000000000000000010111001001001;
assign LUT_1[34369] = 32'b11111111111111111100001011000101;
assign LUT_1[34370] = 32'b11111111111111111110100111011010;
assign LUT_1[34371] = 32'b11111111111111110111111001010110;
assign LUT_1[34372] = 32'b00000000000000001010110010100000;
assign LUT_1[34373] = 32'b00000000000000000100000100011100;
assign LUT_1[34374] = 32'b00000000000000000110100000110001;
assign LUT_1[34375] = 32'b11111111111111111111110010101101;
assign LUT_1[34376] = 32'b00000000000000000010000110111110;
assign LUT_1[34377] = 32'b11111111111111111011011000111010;
assign LUT_1[34378] = 32'b11111111111111111101110101001111;
assign LUT_1[34379] = 32'b11111111111111110111000111001011;
assign LUT_1[34380] = 32'b00000000000000001010000000010101;
assign LUT_1[34381] = 32'b00000000000000000011010010010001;
assign LUT_1[34382] = 32'b00000000000000000101101110100110;
assign LUT_1[34383] = 32'b11111111111111111111000000100010;
assign LUT_1[34384] = 32'b00000000000000000100110100101011;
assign LUT_1[34385] = 32'b11111111111111111110000110100111;
assign LUT_1[34386] = 32'b00000000000000000000100010111100;
assign LUT_1[34387] = 32'b11111111111111111001110100111000;
assign LUT_1[34388] = 32'b00000000000000001100101110000010;
assign LUT_1[34389] = 32'b00000000000000000101111111111110;
assign LUT_1[34390] = 32'b00000000000000001000011100010011;
assign LUT_1[34391] = 32'b00000000000000000001101110001111;
assign LUT_1[34392] = 32'b00000000000000000100000010100000;
assign LUT_1[34393] = 32'b11111111111111111101010100011100;
assign LUT_1[34394] = 32'b11111111111111111111110000110001;
assign LUT_1[34395] = 32'b11111111111111111001000010101101;
assign LUT_1[34396] = 32'b00000000000000001011111011110111;
assign LUT_1[34397] = 32'b00000000000000000101001101110011;
assign LUT_1[34398] = 32'b00000000000000000111101010001000;
assign LUT_1[34399] = 32'b00000000000000000000111100000100;
assign LUT_1[34400] = 32'b00000000000000000011110100001000;
assign LUT_1[34401] = 32'b11111111111111111101000110000100;
assign LUT_1[34402] = 32'b11111111111111111111100010011001;
assign LUT_1[34403] = 32'b11111111111111111000110100010101;
assign LUT_1[34404] = 32'b00000000000000001011101101011111;
assign LUT_1[34405] = 32'b00000000000000000100111111011011;
assign LUT_1[34406] = 32'b00000000000000000111011011110000;
assign LUT_1[34407] = 32'b00000000000000000000101101101100;
assign LUT_1[34408] = 32'b00000000000000000011000001111101;
assign LUT_1[34409] = 32'b11111111111111111100010011111001;
assign LUT_1[34410] = 32'b11111111111111111110110000001110;
assign LUT_1[34411] = 32'b11111111111111111000000010001010;
assign LUT_1[34412] = 32'b00000000000000001010111011010100;
assign LUT_1[34413] = 32'b00000000000000000100001101010000;
assign LUT_1[34414] = 32'b00000000000000000110101001100101;
assign LUT_1[34415] = 32'b11111111111111111111111011100001;
assign LUT_1[34416] = 32'b00000000000000000101101111101010;
assign LUT_1[34417] = 32'b11111111111111111111000001100110;
assign LUT_1[34418] = 32'b00000000000000000001011101111011;
assign LUT_1[34419] = 32'b11111111111111111010101111110111;
assign LUT_1[34420] = 32'b00000000000000001101101001000001;
assign LUT_1[34421] = 32'b00000000000000000110111010111101;
assign LUT_1[34422] = 32'b00000000000000001001010111010010;
assign LUT_1[34423] = 32'b00000000000000000010101001001110;
assign LUT_1[34424] = 32'b00000000000000000100111101011111;
assign LUT_1[34425] = 32'b11111111111111111110001111011011;
assign LUT_1[34426] = 32'b00000000000000000000101011110000;
assign LUT_1[34427] = 32'b11111111111111111001111101101100;
assign LUT_1[34428] = 32'b00000000000000001100110110110110;
assign LUT_1[34429] = 32'b00000000000000000110001000110010;
assign LUT_1[34430] = 32'b00000000000000001000100101000111;
assign LUT_1[34431] = 32'b00000000000000000001110111000011;
assign LUT_1[34432] = 32'b00000000000000000011111011100100;
assign LUT_1[34433] = 32'b11111111111111111101001101100000;
assign LUT_1[34434] = 32'b11111111111111111111101001110101;
assign LUT_1[34435] = 32'b11111111111111111000111011110001;
assign LUT_1[34436] = 32'b00000000000000001011110100111011;
assign LUT_1[34437] = 32'b00000000000000000101000110110111;
assign LUT_1[34438] = 32'b00000000000000000111100011001100;
assign LUT_1[34439] = 32'b00000000000000000000110101001000;
assign LUT_1[34440] = 32'b00000000000000000011001001011001;
assign LUT_1[34441] = 32'b11111111111111111100011011010101;
assign LUT_1[34442] = 32'b11111111111111111110110111101010;
assign LUT_1[34443] = 32'b11111111111111111000001001100110;
assign LUT_1[34444] = 32'b00000000000000001011000010110000;
assign LUT_1[34445] = 32'b00000000000000000100010100101100;
assign LUT_1[34446] = 32'b00000000000000000110110001000001;
assign LUT_1[34447] = 32'b00000000000000000000000010111101;
assign LUT_1[34448] = 32'b00000000000000000101110111000110;
assign LUT_1[34449] = 32'b11111111111111111111001001000010;
assign LUT_1[34450] = 32'b00000000000000000001100101010111;
assign LUT_1[34451] = 32'b11111111111111111010110111010011;
assign LUT_1[34452] = 32'b00000000000000001101110000011101;
assign LUT_1[34453] = 32'b00000000000000000111000010011001;
assign LUT_1[34454] = 32'b00000000000000001001011110101110;
assign LUT_1[34455] = 32'b00000000000000000010110000101010;
assign LUT_1[34456] = 32'b00000000000000000101000100111011;
assign LUT_1[34457] = 32'b11111111111111111110010110110111;
assign LUT_1[34458] = 32'b00000000000000000000110011001100;
assign LUT_1[34459] = 32'b11111111111111111010000101001000;
assign LUT_1[34460] = 32'b00000000000000001100111110010010;
assign LUT_1[34461] = 32'b00000000000000000110010000001110;
assign LUT_1[34462] = 32'b00000000000000001000101100100011;
assign LUT_1[34463] = 32'b00000000000000000001111110011111;
assign LUT_1[34464] = 32'b00000000000000000100110110100011;
assign LUT_1[34465] = 32'b11111111111111111110001000011111;
assign LUT_1[34466] = 32'b00000000000000000000100100110100;
assign LUT_1[34467] = 32'b11111111111111111001110110110000;
assign LUT_1[34468] = 32'b00000000000000001100101111111010;
assign LUT_1[34469] = 32'b00000000000000000110000001110110;
assign LUT_1[34470] = 32'b00000000000000001000011110001011;
assign LUT_1[34471] = 32'b00000000000000000001110000000111;
assign LUT_1[34472] = 32'b00000000000000000100000100011000;
assign LUT_1[34473] = 32'b11111111111111111101010110010100;
assign LUT_1[34474] = 32'b11111111111111111111110010101001;
assign LUT_1[34475] = 32'b11111111111111111001000100100101;
assign LUT_1[34476] = 32'b00000000000000001011111101101111;
assign LUT_1[34477] = 32'b00000000000000000101001111101011;
assign LUT_1[34478] = 32'b00000000000000000111101100000000;
assign LUT_1[34479] = 32'b00000000000000000000111101111100;
assign LUT_1[34480] = 32'b00000000000000000110110010000101;
assign LUT_1[34481] = 32'b00000000000000000000000100000001;
assign LUT_1[34482] = 32'b00000000000000000010100000010110;
assign LUT_1[34483] = 32'b11111111111111111011110010010010;
assign LUT_1[34484] = 32'b00000000000000001110101011011100;
assign LUT_1[34485] = 32'b00000000000000000111111101011000;
assign LUT_1[34486] = 32'b00000000000000001010011001101101;
assign LUT_1[34487] = 32'b00000000000000000011101011101001;
assign LUT_1[34488] = 32'b00000000000000000101111111111010;
assign LUT_1[34489] = 32'b11111111111111111111010001110110;
assign LUT_1[34490] = 32'b00000000000000000001101110001011;
assign LUT_1[34491] = 32'b11111111111111111011000000000111;
assign LUT_1[34492] = 32'b00000000000000001101111001010001;
assign LUT_1[34493] = 32'b00000000000000000111001011001101;
assign LUT_1[34494] = 32'b00000000000000001001100111100010;
assign LUT_1[34495] = 32'b00000000000000000010111001011110;
assign LUT_1[34496] = 32'b00000000000000000101111001001100;
assign LUT_1[34497] = 32'b11111111111111111111001011001000;
assign LUT_1[34498] = 32'b00000000000000000001100111011101;
assign LUT_1[34499] = 32'b11111111111111111010111001011001;
assign LUT_1[34500] = 32'b00000000000000001101110010100011;
assign LUT_1[34501] = 32'b00000000000000000111000100011111;
assign LUT_1[34502] = 32'b00000000000000001001100000110100;
assign LUT_1[34503] = 32'b00000000000000000010110010110000;
assign LUT_1[34504] = 32'b00000000000000000101000111000001;
assign LUT_1[34505] = 32'b11111111111111111110011000111101;
assign LUT_1[34506] = 32'b00000000000000000000110101010010;
assign LUT_1[34507] = 32'b11111111111111111010000111001110;
assign LUT_1[34508] = 32'b00000000000000001101000000011000;
assign LUT_1[34509] = 32'b00000000000000000110010010010100;
assign LUT_1[34510] = 32'b00000000000000001000101110101001;
assign LUT_1[34511] = 32'b00000000000000000010000000100101;
assign LUT_1[34512] = 32'b00000000000000000111110100101110;
assign LUT_1[34513] = 32'b00000000000000000001000110101010;
assign LUT_1[34514] = 32'b00000000000000000011100010111111;
assign LUT_1[34515] = 32'b11111111111111111100110100111011;
assign LUT_1[34516] = 32'b00000000000000001111101110000101;
assign LUT_1[34517] = 32'b00000000000000001001000000000001;
assign LUT_1[34518] = 32'b00000000000000001011011100010110;
assign LUT_1[34519] = 32'b00000000000000000100101110010010;
assign LUT_1[34520] = 32'b00000000000000000111000010100011;
assign LUT_1[34521] = 32'b00000000000000000000010100011111;
assign LUT_1[34522] = 32'b00000000000000000010110000110100;
assign LUT_1[34523] = 32'b11111111111111111100000010110000;
assign LUT_1[34524] = 32'b00000000000000001110111011111010;
assign LUT_1[34525] = 32'b00000000000000001000001101110110;
assign LUT_1[34526] = 32'b00000000000000001010101010001011;
assign LUT_1[34527] = 32'b00000000000000000011111100000111;
assign LUT_1[34528] = 32'b00000000000000000110110100001011;
assign LUT_1[34529] = 32'b00000000000000000000000110000111;
assign LUT_1[34530] = 32'b00000000000000000010100010011100;
assign LUT_1[34531] = 32'b11111111111111111011110100011000;
assign LUT_1[34532] = 32'b00000000000000001110101101100010;
assign LUT_1[34533] = 32'b00000000000000000111111111011110;
assign LUT_1[34534] = 32'b00000000000000001010011011110011;
assign LUT_1[34535] = 32'b00000000000000000011101101101111;
assign LUT_1[34536] = 32'b00000000000000000110000010000000;
assign LUT_1[34537] = 32'b11111111111111111111010011111100;
assign LUT_1[34538] = 32'b00000000000000000001110000010001;
assign LUT_1[34539] = 32'b11111111111111111011000010001101;
assign LUT_1[34540] = 32'b00000000000000001101111011010111;
assign LUT_1[34541] = 32'b00000000000000000111001101010011;
assign LUT_1[34542] = 32'b00000000000000001001101001101000;
assign LUT_1[34543] = 32'b00000000000000000010111011100100;
assign LUT_1[34544] = 32'b00000000000000001000101111101101;
assign LUT_1[34545] = 32'b00000000000000000010000001101001;
assign LUT_1[34546] = 32'b00000000000000000100011101111110;
assign LUT_1[34547] = 32'b11111111111111111101101111111010;
assign LUT_1[34548] = 32'b00000000000000010000101001000100;
assign LUT_1[34549] = 32'b00000000000000001001111011000000;
assign LUT_1[34550] = 32'b00000000000000001100010111010101;
assign LUT_1[34551] = 32'b00000000000000000101101001010001;
assign LUT_1[34552] = 32'b00000000000000000111111101100010;
assign LUT_1[34553] = 32'b00000000000000000001001111011110;
assign LUT_1[34554] = 32'b00000000000000000011101011110011;
assign LUT_1[34555] = 32'b11111111111111111100111101101111;
assign LUT_1[34556] = 32'b00000000000000001111110110111001;
assign LUT_1[34557] = 32'b00000000000000001001001000110101;
assign LUT_1[34558] = 32'b00000000000000001011100101001010;
assign LUT_1[34559] = 32'b00000000000000000100110111000110;
assign LUT_1[34560] = 32'b11111111111111111110101111101101;
assign LUT_1[34561] = 32'b11111111111111111000000001101001;
assign LUT_1[34562] = 32'b11111111111111111010011101111110;
assign LUT_1[34563] = 32'b11111111111111110011101111111010;
assign LUT_1[34564] = 32'b00000000000000000110101001000100;
assign LUT_1[34565] = 32'b11111111111111111111111011000000;
assign LUT_1[34566] = 32'b00000000000000000010010111010101;
assign LUT_1[34567] = 32'b11111111111111111011101001010001;
assign LUT_1[34568] = 32'b11111111111111111101111101100010;
assign LUT_1[34569] = 32'b11111111111111110111001111011110;
assign LUT_1[34570] = 32'b11111111111111111001101011110011;
assign LUT_1[34571] = 32'b11111111111111110010111101101111;
assign LUT_1[34572] = 32'b00000000000000000101110110111001;
assign LUT_1[34573] = 32'b11111111111111111111001000110101;
assign LUT_1[34574] = 32'b00000000000000000001100101001010;
assign LUT_1[34575] = 32'b11111111111111111010110111000110;
assign LUT_1[34576] = 32'b00000000000000000000101011001111;
assign LUT_1[34577] = 32'b11111111111111111001111101001011;
assign LUT_1[34578] = 32'b11111111111111111100011001100000;
assign LUT_1[34579] = 32'b11111111111111110101101011011100;
assign LUT_1[34580] = 32'b00000000000000001000100100100110;
assign LUT_1[34581] = 32'b00000000000000000001110110100010;
assign LUT_1[34582] = 32'b00000000000000000100010010110111;
assign LUT_1[34583] = 32'b11111111111111111101100100110011;
assign LUT_1[34584] = 32'b11111111111111111111111001000100;
assign LUT_1[34585] = 32'b11111111111111111001001011000000;
assign LUT_1[34586] = 32'b11111111111111111011100111010101;
assign LUT_1[34587] = 32'b11111111111111110100111001010001;
assign LUT_1[34588] = 32'b00000000000000000111110010011011;
assign LUT_1[34589] = 32'b00000000000000000001000100010111;
assign LUT_1[34590] = 32'b00000000000000000011100000101100;
assign LUT_1[34591] = 32'b11111111111111111100110010101000;
assign LUT_1[34592] = 32'b11111111111111111111101010101100;
assign LUT_1[34593] = 32'b11111111111111111000111100101000;
assign LUT_1[34594] = 32'b11111111111111111011011000111101;
assign LUT_1[34595] = 32'b11111111111111110100101010111001;
assign LUT_1[34596] = 32'b00000000000000000111100100000011;
assign LUT_1[34597] = 32'b00000000000000000000110101111111;
assign LUT_1[34598] = 32'b00000000000000000011010010010100;
assign LUT_1[34599] = 32'b11111111111111111100100100010000;
assign LUT_1[34600] = 32'b11111111111111111110111000100001;
assign LUT_1[34601] = 32'b11111111111111111000001010011101;
assign LUT_1[34602] = 32'b11111111111111111010100110110010;
assign LUT_1[34603] = 32'b11111111111111110011111000101110;
assign LUT_1[34604] = 32'b00000000000000000110110001111000;
assign LUT_1[34605] = 32'b00000000000000000000000011110100;
assign LUT_1[34606] = 32'b00000000000000000010100000001001;
assign LUT_1[34607] = 32'b11111111111111111011110010000101;
assign LUT_1[34608] = 32'b00000000000000000001100110001110;
assign LUT_1[34609] = 32'b11111111111111111010111000001010;
assign LUT_1[34610] = 32'b11111111111111111101010100011111;
assign LUT_1[34611] = 32'b11111111111111110110100110011011;
assign LUT_1[34612] = 32'b00000000000000001001011111100101;
assign LUT_1[34613] = 32'b00000000000000000010110001100001;
assign LUT_1[34614] = 32'b00000000000000000101001101110110;
assign LUT_1[34615] = 32'b11111111111111111110011111110010;
assign LUT_1[34616] = 32'b00000000000000000000110100000011;
assign LUT_1[34617] = 32'b11111111111111111010000101111111;
assign LUT_1[34618] = 32'b11111111111111111100100010010100;
assign LUT_1[34619] = 32'b11111111111111110101110100010000;
assign LUT_1[34620] = 32'b00000000000000001000101101011010;
assign LUT_1[34621] = 32'b00000000000000000001111111010110;
assign LUT_1[34622] = 32'b00000000000000000100011011101011;
assign LUT_1[34623] = 32'b11111111111111111101101101100111;
assign LUT_1[34624] = 32'b00000000000000000000101101010101;
assign LUT_1[34625] = 32'b11111111111111111001111111010001;
assign LUT_1[34626] = 32'b11111111111111111100011011100110;
assign LUT_1[34627] = 32'b11111111111111110101101101100010;
assign LUT_1[34628] = 32'b00000000000000001000100110101100;
assign LUT_1[34629] = 32'b00000000000000000001111000101000;
assign LUT_1[34630] = 32'b00000000000000000100010100111101;
assign LUT_1[34631] = 32'b11111111111111111101100110111001;
assign LUT_1[34632] = 32'b11111111111111111111111011001010;
assign LUT_1[34633] = 32'b11111111111111111001001101000110;
assign LUT_1[34634] = 32'b11111111111111111011101001011011;
assign LUT_1[34635] = 32'b11111111111111110100111011010111;
assign LUT_1[34636] = 32'b00000000000000000111110100100001;
assign LUT_1[34637] = 32'b00000000000000000001000110011101;
assign LUT_1[34638] = 32'b00000000000000000011100010110010;
assign LUT_1[34639] = 32'b11111111111111111100110100101110;
assign LUT_1[34640] = 32'b00000000000000000010101000110111;
assign LUT_1[34641] = 32'b11111111111111111011111010110011;
assign LUT_1[34642] = 32'b11111111111111111110010111001000;
assign LUT_1[34643] = 32'b11111111111111110111101001000100;
assign LUT_1[34644] = 32'b00000000000000001010100010001110;
assign LUT_1[34645] = 32'b00000000000000000011110100001010;
assign LUT_1[34646] = 32'b00000000000000000110010000011111;
assign LUT_1[34647] = 32'b11111111111111111111100010011011;
assign LUT_1[34648] = 32'b00000000000000000001110110101100;
assign LUT_1[34649] = 32'b11111111111111111011001000101000;
assign LUT_1[34650] = 32'b11111111111111111101100100111101;
assign LUT_1[34651] = 32'b11111111111111110110110110111001;
assign LUT_1[34652] = 32'b00000000000000001001110000000011;
assign LUT_1[34653] = 32'b00000000000000000011000001111111;
assign LUT_1[34654] = 32'b00000000000000000101011110010100;
assign LUT_1[34655] = 32'b11111111111111111110110000010000;
assign LUT_1[34656] = 32'b00000000000000000001101000010100;
assign LUT_1[34657] = 32'b11111111111111111010111010010000;
assign LUT_1[34658] = 32'b11111111111111111101010110100101;
assign LUT_1[34659] = 32'b11111111111111110110101000100001;
assign LUT_1[34660] = 32'b00000000000000001001100001101011;
assign LUT_1[34661] = 32'b00000000000000000010110011100111;
assign LUT_1[34662] = 32'b00000000000000000101001111111100;
assign LUT_1[34663] = 32'b11111111111111111110100001111000;
assign LUT_1[34664] = 32'b00000000000000000000110110001001;
assign LUT_1[34665] = 32'b11111111111111111010001000000101;
assign LUT_1[34666] = 32'b11111111111111111100100100011010;
assign LUT_1[34667] = 32'b11111111111111110101110110010110;
assign LUT_1[34668] = 32'b00000000000000001000101111100000;
assign LUT_1[34669] = 32'b00000000000000000010000001011100;
assign LUT_1[34670] = 32'b00000000000000000100011101110001;
assign LUT_1[34671] = 32'b11111111111111111101101111101101;
assign LUT_1[34672] = 32'b00000000000000000011100011110110;
assign LUT_1[34673] = 32'b11111111111111111100110101110010;
assign LUT_1[34674] = 32'b11111111111111111111010010000111;
assign LUT_1[34675] = 32'b11111111111111111000100100000011;
assign LUT_1[34676] = 32'b00000000000000001011011101001101;
assign LUT_1[34677] = 32'b00000000000000000100101111001001;
assign LUT_1[34678] = 32'b00000000000000000111001011011110;
assign LUT_1[34679] = 32'b00000000000000000000011101011010;
assign LUT_1[34680] = 32'b00000000000000000010110001101011;
assign LUT_1[34681] = 32'b11111111111111111100000011100111;
assign LUT_1[34682] = 32'b11111111111111111110011111111100;
assign LUT_1[34683] = 32'b11111111111111110111110001111000;
assign LUT_1[34684] = 32'b00000000000000001010101011000010;
assign LUT_1[34685] = 32'b00000000000000000011111100111110;
assign LUT_1[34686] = 32'b00000000000000000110011001010011;
assign LUT_1[34687] = 32'b11111111111111111111101011001111;
assign LUT_1[34688] = 32'b00000000000000000001101111110000;
assign LUT_1[34689] = 32'b11111111111111111011000001101100;
assign LUT_1[34690] = 32'b11111111111111111101011110000001;
assign LUT_1[34691] = 32'b11111111111111110110101111111101;
assign LUT_1[34692] = 32'b00000000000000001001101001000111;
assign LUT_1[34693] = 32'b00000000000000000010111011000011;
assign LUT_1[34694] = 32'b00000000000000000101010111011000;
assign LUT_1[34695] = 32'b11111111111111111110101001010100;
assign LUT_1[34696] = 32'b00000000000000000000111101100101;
assign LUT_1[34697] = 32'b11111111111111111010001111100001;
assign LUT_1[34698] = 32'b11111111111111111100101011110110;
assign LUT_1[34699] = 32'b11111111111111110101111101110010;
assign LUT_1[34700] = 32'b00000000000000001000110110111100;
assign LUT_1[34701] = 32'b00000000000000000010001000111000;
assign LUT_1[34702] = 32'b00000000000000000100100101001101;
assign LUT_1[34703] = 32'b11111111111111111101110111001001;
assign LUT_1[34704] = 32'b00000000000000000011101011010010;
assign LUT_1[34705] = 32'b11111111111111111100111101001110;
assign LUT_1[34706] = 32'b11111111111111111111011001100011;
assign LUT_1[34707] = 32'b11111111111111111000101011011111;
assign LUT_1[34708] = 32'b00000000000000001011100100101001;
assign LUT_1[34709] = 32'b00000000000000000100110110100101;
assign LUT_1[34710] = 32'b00000000000000000111010010111010;
assign LUT_1[34711] = 32'b00000000000000000000100100110110;
assign LUT_1[34712] = 32'b00000000000000000010111001000111;
assign LUT_1[34713] = 32'b11111111111111111100001011000011;
assign LUT_1[34714] = 32'b11111111111111111110100111011000;
assign LUT_1[34715] = 32'b11111111111111110111111001010100;
assign LUT_1[34716] = 32'b00000000000000001010110010011110;
assign LUT_1[34717] = 32'b00000000000000000100000100011010;
assign LUT_1[34718] = 32'b00000000000000000110100000101111;
assign LUT_1[34719] = 32'b11111111111111111111110010101011;
assign LUT_1[34720] = 32'b00000000000000000010101010101111;
assign LUT_1[34721] = 32'b11111111111111111011111100101011;
assign LUT_1[34722] = 32'b11111111111111111110011001000000;
assign LUT_1[34723] = 32'b11111111111111110111101010111100;
assign LUT_1[34724] = 32'b00000000000000001010100100000110;
assign LUT_1[34725] = 32'b00000000000000000011110110000010;
assign LUT_1[34726] = 32'b00000000000000000110010010010111;
assign LUT_1[34727] = 32'b11111111111111111111100100010011;
assign LUT_1[34728] = 32'b00000000000000000001111000100100;
assign LUT_1[34729] = 32'b11111111111111111011001010100000;
assign LUT_1[34730] = 32'b11111111111111111101100110110101;
assign LUT_1[34731] = 32'b11111111111111110110111000110001;
assign LUT_1[34732] = 32'b00000000000000001001110001111011;
assign LUT_1[34733] = 32'b00000000000000000011000011110111;
assign LUT_1[34734] = 32'b00000000000000000101100000001100;
assign LUT_1[34735] = 32'b11111111111111111110110010001000;
assign LUT_1[34736] = 32'b00000000000000000100100110010001;
assign LUT_1[34737] = 32'b11111111111111111101111000001101;
assign LUT_1[34738] = 32'b00000000000000000000010100100010;
assign LUT_1[34739] = 32'b11111111111111111001100110011110;
assign LUT_1[34740] = 32'b00000000000000001100011111101000;
assign LUT_1[34741] = 32'b00000000000000000101110001100100;
assign LUT_1[34742] = 32'b00000000000000001000001101111001;
assign LUT_1[34743] = 32'b00000000000000000001011111110101;
assign LUT_1[34744] = 32'b00000000000000000011110100000110;
assign LUT_1[34745] = 32'b11111111111111111101000110000010;
assign LUT_1[34746] = 32'b11111111111111111111100010010111;
assign LUT_1[34747] = 32'b11111111111111111000110100010011;
assign LUT_1[34748] = 32'b00000000000000001011101101011101;
assign LUT_1[34749] = 32'b00000000000000000100111111011001;
assign LUT_1[34750] = 32'b00000000000000000111011011101110;
assign LUT_1[34751] = 32'b00000000000000000000101101101010;
assign LUT_1[34752] = 32'b00000000000000000011101101011000;
assign LUT_1[34753] = 32'b11111111111111111100111111010100;
assign LUT_1[34754] = 32'b11111111111111111111011011101001;
assign LUT_1[34755] = 32'b11111111111111111000101101100101;
assign LUT_1[34756] = 32'b00000000000000001011100110101111;
assign LUT_1[34757] = 32'b00000000000000000100111000101011;
assign LUT_1[34758] = 32'b00000000000000000111010101000000;
assign LUT_1[34759] = 32'b00000000000000000000100110111100;
assign LUT_1[34760] = 32'b00000000000000000010111011001101;
assign LUT_1[34761] = 32'b11111111111111111100001101001001;
assign LUT_1[34762] = 32'b11111111111111111110101001011110;
assign LUT_1[34763] = 32'b11111111111111110111111011011010;
assign LUT_1[34764] = 32'b00000000000000001010110100100100;
assign LUT_1[34765] = 32'b00000000000000000100000110100000;
assign LUT_1[34766] = 32'b00000000000000000110100010110101;
assign LUT_1[34767] = 32'b11111111111111111111110100110001;
assign LUT_1[34768] = 32'b00000000000000000101101000111010;
assign LUT_1[34769] = 32'b11111111111111111110111010110110;
assign LUT_1[34770] = 32'b00000000000000000001010111001011;
assign LUT_1[34771] = 32'b11111111111111111010101001000111;
assign LUT_1[34772] = 32'b00000000000000001101100010010001;
assign LUT_1[34773] = 32'b00000000000000000110110100001101;
assign LUT_1[34774] = 32'b00000000000000001001010000100010;
assign LUT_1[34775] = 32'b00000000000000000010100010011110;
assign LUT_1[34776] = 32'b00000000000000000100110110101111;
assign LUT_1[34777] = 32'b11111111111111111110001000101011;
assign LUT_1[34778] = 32'b00000000000000000000100101000000;
assign LUT_1[34779] = 32'b11111111111111111001110110111100;
assign LUT_1[34780] = 32'b00000000000000001100110000000110;
assign LUT_1[34781] = 32'b00000000000000000110000010000010;
assign LUT_1[34782] = 32'b00000000000000001000011110010111;
assign LUT_1[34783] = 32'b00000000000000000001110000010011;
assign LUT_1[34784] = 32'b00000000000000000100101000010111;
assign LUT_1[34785] = 32'b11111111111111111101111010010011;
assign LUT_1[34786] = 32'b00000000000000000000010110101000;
assign LUT_1[34787] = 32'b11111111111111111001101000100100;
assign LUT_1[34788] = 32'b00000000000000001100100001101110;
assign LUT_1[34789] = 32'b00000000000000000101110011101010;
assign LUT_1[34790] = 32'b00000000000000001000001111111111;
assign LUT_1[34791] = 32'b00000000000000000001100001111011;
assign LUT_1[34792] = 32'b00000000000000000011110110001100;
assign LUT_1[34793] = 32'b11111111111111111101001000001000;
assign LUT_1[34794] = 32'b11111111111111111111100100011101;
assign LUT_1[34795] = 32'b11111111111111111000110110011001;
assign LUT_1[34796] = 32'b00000000000000001011101111100011;
assign LUT_1[34797] = 32'b00000000000000000101000001011111;
assign LUT_1[34798] = 32'b00000000000000000111011101110100;
assign LUT_1[34799] = 32'b00000000000000000000101111110000;
assign LUT_1[34800] = 32'b00000000000000000110100011111001;
assign LUT_1[34801] = 32'b11111111111111111111110101110101;
assign LUT_1[34802] = 32'b00000000000000000010010010001010;
assign LUT_1[34803] = 32'b11111111111111111011100100000110;
assign LUT_1[34804] = 32'b00000000000000001110011101010000;
assign LUT_1[34805] = 32'b00000000000000000111101111001100;
assign LUT_1[34806] = 32'b00000000000000001010001011100001;
assign LUT_1[34807] = 32'b00000000000000000011011101011101;
assign LUT_1[34808] = 32'b00000000000000000101110001101110;
assign LUT_1[34809] = 32'b11111111111111111111000011101010;
assign LUT_1[34810] = 32'b00000000000000000001011111111111;
assign LUT_1[34811] = 32'b11111111111111111010110001111011;
assign LUT_1[34812] = 32'b00000000000000001101101011000101;
assign LUT_1[34813] = 32'b00000000000000000110111101000001;
assign LUT_1[34814] = 32'b00000000000000001001011001010110;
assign LUT_1[34815] = 32'b00000000000000000010101011010010;
assign LUT_1[34816] = 32'b00000000000000000001111000001111;
assign LUT_1[34817] = 32'b11111111111111111011001010001011;
assign LUT_1[34818] = 32'b11111111111111111101100110100000;
assign LUT_1[34819] = 32'b11111111111111110110111000011100;
assign LUT_1[34820] = 32'b00000000000000001001110001100110;
assign LUT_1[34821] = 32'b00000000000000000011000011100010;
assign LUT_1[34822] = 32'b00000000000000000101011111110111;
assign LUT_1[34823] = 32'b11111111111111111110110001110011;
assign LUT_1[34824] = 32'b00000000000000000001000110000100;
assign LUT_1[34825] = 32'b11111111111111111010011000000000;
assign LUT_1[34826] = 32'b11111111111111111100110100010101;
assign LUT_1[34827] = 32'b11111111111111110110000110010001;
assign LUT_1[34828] = 32'b00000000000000001000111111011011;
assign LUT_1[34829] = 32'b00000000000000000010010001010111;
assign LUT_1[34830] = 32'b00000000000000000100101101101100;
assign LUT_1[34831] = 32'b11111111111111111101111111101000;
assign LUT_1[34832] = 32'b00000000000000000011110011110001;
assign LUT_1[34833] = 32'b11111111111111111101000101101101;
assign LUT_1[34834] = 32'b11111111111111111111100010000010;
assign LUT_1[34835] = 32'b11111111111111111000110011111110;
assign LUT_1[34836] = 32'b00000000000000001011101101001000;
assign LUT_1[34837] = 32'b00000000000000000100111111000100;
assign LUT_1[34838] = 32'b00000000000000000111011011011001;
assign LUT_1[34839] = 32'b00000000000000000000101101010101;
assign LUT_1[34840] = 32'b00000000000000000011000001100110;
assign LUT_1[34841] = 32'b11111111111111111100010011100010;
assign LUT_1[34842] = 32'b11111111111111111110101111110111;
assign LUT_1[34843] = 32'b11111111111111111000000001110011;
assign LUT_1[34844] = 32'b00000000000000001010111010111101;
assign LUT_1[34845] = 32'b00000000000000000100001100111001;
assign LUT_1[34846] = 32'b00000000000000000110101001001110;
assign LUT_1[34847] = 32'b11111111111111111111111011001010;
assign LUT_1[34848] = 32'b00000000000000000010110011001110;
assign LUT_1[34849] = 32'b11111111111111111100000101001010;
assign LUT_1[34850] = 32'b11111111111111111110100001011111;
assign LUT_1[34851] = 32'b11111111111111110111110011011011;
assign LUT_1[34852] = 32'b00000000000000001010101100100101;
assign LUT_1[34853] = 32'b00000000000000000011111110100001;
assign LUT_1[34854] = 32'b00000000000000000110011010110110;
assign LUT_1[34855] = 32'b11111111111111111111101100110010;
assign LUT_1[34856] = 32'b00000000000000000010000001000011;
assign LUT_1[34857] = 32'b11111111111111111011010010111111;
assign LUT_1[34858] = 32'b11111111111111111101101111010100;
assign LUT_1[34859] = 32'b11111111111111110111000001010000;
assign LUT_1[34860] = 32'b00000000000000001001111010011010;
assign LUT_1[34861] = 32'b00000000000000000011001100010110;
assign LUT_1[34862] = 32'b00000000000000000101101000101011;
assign LUT_1[34863] = 32'b11111111111111111110111010100111;
assign LUT_1[34864] = 32'b00000000000000000100101110110000;
assign LUT_1[34865] = 32'b11111111111111111110000000101100;
assign LUT_1[34866] = 32'b00000000000000000000011101000001;
assign LUT_1[34867] = 32'b11111111111111111001101110111101;
assign LUT_1[34868] = 32'b00000000000000001100101000000111;
assign LUT_1[34869] = 32'b00000000000000000101111010000011;
assign LUT_1[34870] = 32'b00000000000000001000010110011000;
assign LUT_1[34871] = 32'b00000000000000000001101000010100;
assign LUT_1[34872] = 32'b00000000000000000011111100100101;
assign LUT_1[34873] = 32'b11111111111111111101001110100001;
assign LUT_1[34874] = 32'b11111111111111111111101010110110;
assign LUT_1[34875] = 32'b11111111111111111000111100110010;
assign LUT_1[34876] = 32'b00000000000000001011110101111100;
assign LUT_1[34877] = 32'b00000000000000000101000111111000;
assign LUT_1[34878] = 32'b00000000000000000111100100001101;
assign LUT_1[34879] = 32'b00000000000000000000110110001001;
assign LUT_1[34880] = 32'b00000000000000000011110101110111;
assign LUT_1[34881] = 32'b11111111111111111101000111110011;
assign LUT_1[34882] = 32'b11111111111111111111100100001000;
assign LUT_1[34883] = 32'b11111111111111111000110110000100;
assign LUT_1[34884] = 32'b00000000000000001011101111001110;
assign LUT_1[34885] = 32'b00000000000000000101000001001010;
assign LUT_1[34886] = 32'b00000000000000000111011101011111;
assign LUT_1[34887] = 32'b00000000000000000000101111011011;
assign LUT_1[34888] = 32'b00000000000000000011000011101100;
assign LUT_1[34889] = 32'b11111111111111111100010101101000;
assign LUT_1[34890] = 32'b11111111111111111110110001111101;
assign LUT_1[34891] = 32'b11111111111111111000000011111001;
assign LUT_1[34892] = 32'b00000000000000001010111101000011;
assign LUT_1[34893] = 32'b00000000000000000100001110111111;
assign LUT_1[34894] = 32'b00000000000000000110101011010100;
assign LUT_1[34895] = 32'b11111111111111111111111101010000;
assign LUT_1[34896] = 32'b00000000000000000101110001011001;
assign LUT_1[34897] = 32'b11111111111111111111000011010101;
assign LUT_1[34898] = 32'b00000000000000000001011111101010;
assign LUT_1[34899] = 32'b11111111111111111010110001100110;
assign LUT_1[34900] = 32'b00000000000000001101101010110000;
assign LUT_1[34901] = 32'b00000000000000000110111100101100;
assign LUT_1[34902] = 32'b00000000000000001001011001000001;
assign LUT_1[34903] = 32'b00000000000000000010101010111101;
assign LUT_1[34904] = 32'b00000000000000000100111111001110;
assign LUT_1[34905] = 32'b11111111111111111110010001001010;
assign LUT_1[34906] = 32'b00000000000000000000101101011111;
assign LUT_1[34907] = 32'b11111111111111111001111111011011;
assign LUT_1[34908] = 32'b00000000000000001100111000100101;
assign LUT_1[34909] = 32'b00000000000000000110001010100001;
assign LUT_1[34910] = 32'b00000000000000001000100110110110;
assign LUT_1[34911] = 32'b00000000000000000001111000110010;
assign LUT_1[34912] = 32'b00000000000000000100110000110110;
assign LUT_1[34913] = 32'b11111111111111111110000010110010;
assign LUT_1[34914] = 32'b00000000000000000000011111000111;
assign LUT_1[34915] = 32'b11111111111111111001110001000011;
assign LUT_1[34916] = 32'b00000000000000001100101010001101;
assign LUT_1[34917] = 32'b00000000000000000101111100001001;
assign LUT_1[34918] = 32'b00000000000000001000011000011110;
assign LUT_1[34919] = 32'b00000000000000000001101010011010;
assign LUT_1[34920] = 32'b00000000000000000011111110101011;
assign LUT_1[34921] = 32'b11111111111111111101010000100111;
assign LUT_1[34922] = 32'b11111111111111111111101100111100;
assign LUT_1[34923] = 32'b11111111111111111000111110111000;
assign LUT_1[34924] = 32'b00000000000000001011111000000010;
assign LUT_1[34925] = 32'b00000000000000000101001001111110;
assign LUT_1[34926] = 32'b00000000000000000111100110010011;
assign LUT_1[34927] = 32'b00000000000000000000111000001111;
assign LUT_1[34928] = 32'b00000000000000000110101100011000;
assign LUT_1[34929] = 32'b11111111111111111111111110010100;
assign LUT_1[34930] = 32'b00000000000000000010011010101001;
assign LUT_1[34931] = 32'b11111111111111111011101100100101;
assign LUT_1[34932] = 32'b00000000000000001110100101101111;
assign LUT_1[34933] = 32'b00000000000000000111110111101011;
assign LUT_1[34934] = 32'b00000000000000001010010100000000;
assign LUT_1[34935] = 32'b00000000000000000011100101111100;
assign LUT_1[34936] = 32'b00000000000000000101111010001101;
assign LUT_1[34937] = 32'b11111111111111111111001100001001;
assign LUT_1[34938] = 32'b00000000000000000001101000011110;
assign LUT_1[34939] = 32'b11111111111111111010111010011010;
assign LUT_1[34940] = 32'b00000000000000001101110011100100;
assign LUT_1[34941] = 32'b00000000000000000111000101100000;
assign LUT_1[34942] = 32'b00000000000000001001100001110101;
assign LUT_1[34943] = 32'b00000000000000000010110011110001;
assign LUT_1[34944] = 32'b00000000000000000100111000010010;
assign LUT_1[34945] = 32'b11111111111111111110001010001110;
assign LUT_1[34946] = 32'b00000000000000000000100110100011;
assign LUT_1[34947] = 32'b11111111111111111001111000011111;
assign LUT_1[34948] = 32'b00000000000000001100110001101001;
assign LUT_1[34949] = 32'b00000000000000000110000011100101;
assign LUT_1[34950] = 32'b00000000000000001000011111111010;
assign LUT_1[34951] = 32'b00000000000000000001110001110110;
assign LUT_1[34952] = 32'b00000000000000000100000110000111;
assign LUT_1[34953] = 32'b11111111111111111101011000000011;
assign LUT_1[34954] = 32'b11111111111111111111110100011000;
assign LUT_1[34955] = 32'b11111111111111111001000110010100;
assign LUT_1[34956] = 32'b00000000000000001011111111011110;
assign LUT_1[34957] = 32'b00000000000000000101010001011010;
assign LUT_1[34958] = 32'b00000000000000000111101101101111;
assign LUT_1[34959] = 32'b00000000000000000000111111101011;
assign LUT_1[34960] = 32'b00000000000000000110110011110100;
assign LUT_1[34961] = 32'b00000000000000000000000101110000;
assign LUT_1[34962] = 32'b00000000000000000010100010000101;
assign LUT_1[34963] = 32'b11111111111111111011110100000001;
assign LUT_1[34964] = 32'b00000000000000001110101101001011;
assign LUT_1[34965] = 32'b00000000000000000111111111000111;
assign LUT_1[34966] = 32'b00000000000000001010011011011100;
assign LUT_1[34967] = 32'b00000000000000000011101101011000;
assign LUT_1[34968] = 32'b00000000000000000110000001101001;
assign LUT_1[34969] = 32'b11111111111111111111010011100101;
assign LUT_1[34970] = 32'b00000000000000000001101111111010;
assign LUT_1[34971] = 32'b11111111111111111011000001110110;
assign LUT_1[34972] = 32'b00000000000000001101111011000000;
assign LUT_1[34973] = 32'b00000000000000000111001100111100;
assign LUT_1[34974] = 32'b00000000000000001001101001010001;
assign LUT_1[34975] = 32'b00000000000000000010111011001101;
assign LUT_1[34976] = 32'b00000000000000000101110011010001;
assign LUT_1[34977] = 32'b11111111111111111111000101001101;
assign LUT_1[34978] = 32'b00000000000000000001100001100010;
assign LUT_1[34979] = 32'b11111111111111111010110011011110;
assign LUT_1[34980] = 32'b00000000000000001101101100101000;
assign LUT_1[34981] = 32'b00000000000000000110111110100100;
assign LUT_1[34982] = 32'b00000000000000001001011010111001;
assign LUT_1[34983] = 32'b00000000000000000010101100110101;
assign LUT_1[34984] = 32'b00000000000000000101000001000110;
assign LUT_1[34985] = 32'b11111111111111111110010011000010;
assign LUT_1[34986] = 32'b00000000000000000000101111010111;
assign LUT_1[34987] = 32'b11111111111111111010000001010011;
assign LUT_1[34988] = 32'b00000000000000001100111010011101;
assign LUT_1[34989] = 32'b00000000000000000110001100011001;
assign LUT_1[34990] = 32'b00000000000000001000101000101110;
assign LUT_1[34991] = 32'b00000000000000000001111010101010;
assign LUT_1[34992] = 32'b00000000000000000111101110110011;
assign LUT_1[34993] = 32'b00000000000000000001000000101111;
assign LUT_1[34994] = 32'b00000000000000000011011101000100;
assign LUT_1[34995] = 32'b11111111111111111100101111000000;
assign LUT_1[34996] = 32'b00000000000000001111101000001010;
assign LUT_1[34997] = 32'b00000000000000001000111010000110;
assign LUT_1[34998] = 32'b00000000000000001011010110011011;
assign LUT_1[34999] = 32'b00000000000000000100101000010111;
assign LUT_1[35000] = 32'b00000000000000000110111100101000;
assign LUT_1[35001] = 32'b00000000000000000000001110100100;
assign LUT_1[35002] = 32'b00000000000000000010101010111001;
assign LUT_1[35003] = 32'b11111111111111111011111100110101;
assign LUT_1[35004] = 32'b00000000000000001110110101111111;
assign LUT_1[35005] = 32'b00000000000000001000000111111011;
assign LUT_1[35006] = 32'b00000000000000001010100100010000;
assign LUT_1[35007] = 32'b00000000000000000011110110001100;
assign LUT_1[35008] = 32'b00000000000000000110110101111010;
assign LUT_1[35009] = 32'b00000000000000000000000111110110;
assign LUT_1[35010] = 32'b00000000000000000010100100001011;
assign LUT_1[35011] = 32'b11111111111111111011110110000111;
assign LUT_1[35012] = 32'b00000000000000001110101111010001;
assign LUT_1[35013] = 32'b00000000000000001000000001001101;
assign LUT_1[35014] = 32'b00000000000000001010011101100010;
assign LUT_1[35015] = 32'b00000000000000000011101111011110;
assign LUT_1[35016] = 32'b00000000000000000110000011101111;
assign LUT_1[35017] = 32'b11111111111111111111010101101011;
assign LUT_1[35018] = 32'b00000000000000000001110010000000;
assign LUT_1[35019] = 32'b11111111111111111011000011111100;
assign LUT_1[35020] = 32'b00000000000000001101111101000110;
assign LUT_1[35021] = 32'b00000000000000000111001111000010;
assign LUT_1[35022] = 32'b00000000000000001001101011010111;
assign LUT_1[35023] = 32'b00000000000000000010111101010011;
assign LUT_1[35024] = 32'b00000000000000001000110001011100;
assign LUT_1[35025] = 32'b00000000000000000010000011011000;
assign LUT_1[35026] = 32'b00000000000000000100011111101101;
assign LUT_1[35027] = 32'b11111111111111111101110001101001;
assign LUT_1[35028] = 32'b00000000000000010000101010110011;
assign LUT_1[35029] = 32'b00000000000000001001111100101111;
assign LUT_1[35030] = 32'b00000000000000001100011001000100;
assign LUT_1[35031] = 32'b00000000000000000101101011000000;
assign LUT_1[35032] = 32'b00000000000000000111111111010001;
assign LUT_1[35033] = 32'b00000000000000000001010001001101;
assign LUT_1[35034] = 32'b00000000000000000011101101100010;
assign LUT_1[35035] = 32'b11111111111111111100111111011110;
assign LUT_1[35036] = 32'b00000000000000001111111000101000;
assign LUT_1[35037] = 32'b00000000000000001001001010100100;
assign LUT_1[35038] = 32'b00000000000000001011100110111001;
assign LUT_1[35039] = 32'b00000000000000000100111000110101;
assign LUT_1[35040] = 32'b00000000000000000111110000111001;
assign LUT_1[35041] = 32'b00000000000000000001000010110101;
assign LUT_1[35042] = 32'b00000000000000000011011111001010;
assign LUT_1[35043] = 32'b11111111111111111100110001000110;
assign LUT_1[35044] = 32'b00000000000000001111101010010000;
assign LUT_1[35045] = 32'b00000000000000001000111100001100;
assign LUT_1[35046] = 32'b00000000000000001011011000100001;
assign LUT_1[35047] = 32'b00000000000000000100101010011101;
assign LUT_1[35048] = 32'b00000000000000000110111110101110;
assign LUT_1[35049] = 32'b00000000000000000000010000101010;
assign LUT_1[35050] = 32'b00000000000000000010101100111111;
assign LUT_1[35051] = 32'b11111111111111111011111110111011;
assign LUT_1[35052] = 32'b00000000000000001110111000000101;
assign LUT_1[35053] = 32'b00000000000000001000001010000001;
assign LUT_1[35054] = 32'b00000000000000001010100110010110;
assign LUT_1[35055] = 32'b00000000000000000011111000010010;
assign LUT_1[35056] = 32'b00000000000000001001101100011011;
assign LUT_1[35057] = 32'b00000000000000000010111110010111;
assign LUT_1[35058] = 32'b00000000000000000101011010101100;
assign LUT_1[35059] = 32'b11111111111111111110101100101000;
assign LUT_1[35060] = 32'b00000000000000010001100101110010;
assign LUT_1[35061] = 32'b00000000000000001010110111101110;
assign LUT_1[35062] = 32'b00000000000000001101010100000011;
assign LUT_1[35063] = 32'b00000000000000000110100101111111;
assign LUT_1[35064] = 32'b00000000000000001000111010010000;
assign LUT_1[35065] = 32'b00000000000000000010001100001100;
assign LUT_1[35066] = 32'b00000000000000000100101000100001;
assign LUT_1[35067] = 32'b11111111111111111101111010011101;
assign LUT_1[35068] = 32'b00000000000000010000110011100111;
assign LUT_1[35069] = 32'b00000000000000001010000101100011;
assign LUT_1[35070] = 32'b00000000000000001100100001111000;
assign LUT_1[35071] = 32'b00000000000000000101110011110100;
assign LUT_1[35072] = 32'b11111111111111111111101100011011;
assign LUT_1[35073] = 32'b11111111111111111000111110010111;
assign LUT_1[35074] = 32'b11111111111111111011011010101100;
assign LUT_1[35075] = 32'b11111111111111110100101100101000;
assign LUT_1[35076] = 32'b00000000000000000111100101110010;
assign LUT_1[35077] = 32'b00000000000000000000110111101110;
assign LUT_1[35078] = 32'b00000000000000000011010100000011;
assign LUT_1[35079] = 32'b11111111111111111100100101111111;
assign LUT_1[35080] = 32'b11111111111111111110111010010000;
assign LUT_1[35081] = 32'b11111111111111111000001100001100;
assign LUT_1[35082] = 32'b11111111111111111010101000100001;
assign LUT_1[35083] = 32'b11111111111111110011111010011101;
assign LUT_1[35084] = 32'b00000000000000000110110011100111;
assign LUT_1[35085] = 32'b00000000000000000000000101100011;
assign LUT_1[35086] = 32'b00000000000000000010100001111000;
assign LUT_1[35087] = 32'b11111111111111111011110011110100;
assign LUT_1[35088] = 32'b00000000000000000001100111111101;
assign LUT_1[35089] = 32'b11111111111111111010111001111001;
assign LUT_1[35090] = 32'b11111111111111111101010110001110;
assign LUT_1[35091] = 32'b11111111111111110110101000001010;
assign LUT_1[35092] = 32'b00000000000000001001100001010100;
assign LUT_1[35093] = 32'b00000000000000000010110011010000;
assign LUT_1[35094] = 32'b00000000000000000101001111100101;
assign LUT_1[35095] = 32'b11111111111111111110100001100001;
assign LUT_1[35096] = 32'b00000000000000000000110101110010;
assign LUT_1[35097] = 32'b11111111111111111010000111101110;
assign LUT_1[35098] = 32'b11111111111111111100100100000011;
assign LUT_1[35099] = 32'b11111111111111110101110101111111;
assign LUT_1[35100] = 32'b00000000000000001000101111001001;
assign LUT_1[35101] = 32'b00000000000000000010000001000101;
assign LUT_1[35102] = 32'b00000000000000000100011101011010;
assign LUT_1[35103] = 32'b11111111111111111101101111010110;
assign LUT_1[35104] = 32'b00000000000000000000100111011010;
assign LUT_1[35105] = 32'b11111111111111111001111001010110;
assign LUT_1[35106] = 32'b11111111111111111100010101101011;
assign LUT_1[35107] = 32'b11111111111111110101100111100111;
assign LUT_1[35108] = 32'b00000000000000001000100000110001;
assign LUT_1[35109] = 32'b00000000000000000001110010101101;
assign LUT_1[35110] = 32'b00000000000000000100001111000010;
assign LUT_1[35111] = 32'b11111111111111111101100000111110;
assign LUT_1[35112] = 32'b11111111111111111111110101001111;
assign LUT_1[35113] = 32'b11111111111111111001000111001011;
assign LUT_1[35114] = 32'b11111111111111111011100011100000;
assign LUT_1[35115] = 32'b11111111111111110100110101011100;
assign LUT_1[35116] = 32'b00000000000000000111101110100110;
assign LUT_1[35117] = 32'b00000000000000000001000000100010;
assign LUT_1[35118] = 32'b00000000000000000011011100110111;
assign LUT_1[35119] = 32'b11111111111111111100101110110011;
assign LUT_1[35120] = 32'b00000000000000000010100010111100;
assign LUT_1[35121] = 32'b11111111111111111011110100111000;
assign LUT_1[35122] = 32'b11111111111111111110010001001101;
assign LUT_1[35123] = 32'b11111111111111110111100011001001;
assign LUT_1[35124] = 32'b00000000000000001010011100010011;
assign LUT_1[35125] = 32'b00000000000000000011101110001111;
assign LUT_1[35126] = 32'b00000000000000000110001010100100;
assign LUT_1[35127] = 32'b11111111111111111111011100100000;
assign LUT_1[35128] = 32'b00000000000000000001110000110001;
assign LUT_1[35129] = 32'b11111111111111111011000010101101;
assign LUT_1[35130] = 32'b11111111111111111101011111000010;
assign LUT_1[35131] = 32'b11111111111111110110110000111110;
assign LUT_1[35132] = 32'b00000000000000001001101010001000;
assign LUT_1[35133] = 32'b00000000000000000010111100000100;
assign LUT_1[35134] = 32'b00000000000000000101011000011001;
assign LUT_1[35135] = 32'b11111111111111111110101010010101;
assign LUT_1[35136] = 32'b00000000000000000001101010000011;
assign LUT_1[35137] = 32'b11111111111111111010111011111111;
assign LUT_1[35138] = 32'b11111111111111111101011000010100;
assign LUT_1[35139] = 32'b11111111111111110110101010010000;
assign LUT_1[35140] = 32'b00000000000000001001100011011010;
assign LUT_1[35141] = 32'b00000000000000000010110101010110;
assign LUT_1[35142] = 32'b00000000000000000101010001101011;
assign LUT_1[35143] = 32'b11111111111111111110100011100111;
assign LUT_1[35144] = 32'b00000000000000000000110111111000;
assign LUT_1[35145] = 32'b11111111111111111010001001110100;
assign LUT_1[35146] = 32'b11111111111111111100100110001001;
assign LUT_1[35147] = 32'b11111111111111110101111000000101;
assign LUT_1[35148] = 32'b00000000000000001000110001001111;
assign LUT_1[35149] = 32'b00000000000000000010000011001011;
assign LUT_1[35150] = 32'b00000000000000000100011111100000;
assign LUT_1[35151] = 32'b11111111111111111101110001011100;
assign LUT_1[35152] = 32'b00000000000000000011100101100101;
assign LUT_1[35153] = 32'b11111111111111111100110111100001;
assign LUT_1[35154] = 32'b11111111111111111111010011110110;
assign LUT_1[35155] = 32'b11111111111111111000100101110010;
assign LUT_1[35156] = 32'b00000000000000001011011110111100;
assign LUT_1[35157] = 32'b00000000000000000100110000111000;
assign LUT_1[35158] = 32'b00000000000000000111001101001101;
assign LUT_1[35159] = 32'b00000000000000000000011111001001;
assign LUT_1[35160] = 32'b00000000000000000010110011011010;
assign LUT_1[35161] = 32'b11111111111111111100000101010110;
assign LUT_1[35162] = 32'b11111111111111111110100001101011;
assign LUT_1[35163] = 32'b11111111111111110111110011100111;
assign LUT_1[35164] = 32'b00000000000000001010101100110001;
assign LUT_1[35165] = 32'b00000000000000000011111110101101;
assign LUT_1[35166] = 32'b00000000000000000110011011000010;
assign LUT_1[35167] = 32'b11111111111111111111101100111110;
assign LUT_1[35168] = 32'b00000000000000000010100101000010;
assign LUT_1[35169] = 32'b11111111111111111011110110111110;
assign LUT_1[35170] = 32'b11111111111111111110010011010011;
assign LUT_1[35171] = 32'b11111111111111110111100101001111;
assign LUT_1[35172] = 32'b00000000000000001010011110011001;
assign LUT_1[35173] = 32'b00000000000000000011110000010101;
assign LUT_1[35174] = 32'b00000000000000000110001100101010;
assign LUT_1[35175] = 32'b11111111111111111111011110100110;
assign LUT_1[35176] = 32'b00000000000000000001110010110111;
assign LUT_1[35177] = 32'b11111111111111111011000100110011;
assign LUT_1[35178] = 32'b11111111111111111101100001001000;
assign LUT_1[35179] = 32'b11111111111111110110110011000100;
assign LUT_1[35180] = 32'b00000000000000001001101100001110;
assign LUT_1[35181] = 32'b00000000000000000010111110001010;
assign LUT_1[35182] = 32'b00000000000000000101011010011111;
assign LUT_1[35183] = 32'b11111111111111111110101100011011;
assign LUT_1[35184] = 32'b00000000000000000100100000100100;
assign LUT_1[35185] = 32'b11111111111111111101110010100000;
assign LUT_1[35186] = 32'b00000000000000000000001110110101;
assign LUT_1[35187] = 32'b11111111111111111001100000110001;
assign LUT_1[35188] = 32'b00000000000000001100011001111011;
assign LUT_1[35189] = 32'b00000000000000000101101011110111;
assign LUT_1[35190] = 32'b00000000000000001000001000001100;
assign LUT_1[35191] = 32'b00000000000000000001011010001000;
assign LUT_1[35192] = 32'b00000000000000000011101110011001;
assign LUT_1[35193] = 32'b11111111111111111101000000010101;
assign LUT_1[35194] = 32'b11111111111111111111011100101010;
assign LUT_1[35195] = 32'b11111111111111111000101110100110;
assign LUT_1[35196] = 32'b00000000000000001011100111110000;
assign LUT_1[35197] = 32'b00000000000000000100111001101100;
assign LUT_1[35198] = 32'b00000000000000000111010110000001;
assign LUT_1[35199] = 32'b00000000000000000000100111111101;
assign LUT_1[35200] = 32'b00000000000000000010101100011110;
assign LUT_1[35201] = 32'b11111111111111111011111110011010;
assign LUT_1[35202] = 32'b11111111111111111110011010101111;
assign LUT_1[35203] = 32'b11111111111111110111101100101011;
assign LUT_1[35204] = 32'b00000000000000001010100101110101;
assign LUT_1[35205] = 32'b00000000000000000011110111110001;
assign LUT_1[35206] = 32'b00000000000000000110010100000110;
assign LUT_1[35207] = 32'b11111111111111111111100110000010;
assign LUT_1[35208] = 32'b00000000000000000001111010010011;
assign LUT_1[35209] = 32'b11111111111111111011001100001111;
assign LUT_1[35210] = 32'b11111111111111111101101000100100;
assign LUT_1[35211] = 32'b11111111111111110110111010100000;
assign LUT_1[35212] = 32'b00000000000000001001110011101010;
assign LUT_1[35213] = 32'b00000000000000000011000101100110;
assign LUT_1[35214] = 32'b00000000000000000101100001111011;
assign LUT_1[35215] = 32'b11111111111111111110110011110111;
assign LUT_1[35216] = 32'b00000000000000000100101000000000;
assign LUT_1[35217] = 32'b11111111111111111101111001111100;
assign LUT_1[35218] = 32'b00000000000000000000010110010001;
assign LUT_1[35219] = 32'b11111111111111111001101000001101;
assign LUT_1[35220] = 32'b00000000000000001100100001010111;
assign LUT_1[35221] = 32'b00000000000000000101110011010011;
assign LUT_1[35222] = 32'b00000000000000001000001111101000;
assign LUT_1[35223] = 32'b00000000000000000001100001100100;
assign LUT_1[35224] = 32'b00000000000000000011110101110101;
assign LUT_1[35225] = 32'b11111111111111111101000111110001;
assign LUT_1[35226] = 32'b11111111111111111111100100000110;
assign LUT_1[35227] = 32'b11111111111111111000110110000010;
assign LUT_1[35228] = 32'b00000000000000001011101111001100;
assign LUT_1[35229] = 32'b00000000000000000101000001001000;
assign LUT_1[35230] = 32'b00000000000000000111011101011101;
assign LUT_1[35231] = 32'b00000000000000000000101111011001;
assign LUT_1[35232] = 32'b00000000000000000011100111011101;
assign LUT_1[35233] = 32'b11111111111111111100111001011001;
assign LUT_1[35234] = 32'b11111111111111111111010101101110;
assign LUT_1[35235] = 32'b11111111111111111000100111101010;
assign LUT_1[35236] = 32'b00000000000000001011100000110100;
assign LUT_1[35237] = 32'b00000000000000000100110010110000;
assign LUT_1[35238] = 32'b00000000000000000111001111000101;
assign LUT_1[35239] = 32'b00000000000000000000100001000001;
assign LUT_1[35240] = 32'b00000000000000000010110101010010;
assign LUT_1[35241] = 32'b11111111111111111100000111001110;
assign LUT_1[35242] = 32'b11111111111111111110100011100011;
assign LUT_1[35243] = 32'b11111111111111110111110101011111;
assign LUT_1[35244] = 32'b00000000000000001010101110101001;
assign LUT_1[35245] = 32'b00000000000000000100000000100101;
assign LUT_1[35246] = 32'b00000000000000000110011100111010;
assign LUT_1[35247] = 32'b11111111111111111111101110110110;
assign LUT_1[35248] = 32'b00000000000000000101100010111111;
assign LUT_1[35249] = 32'b11111111111111111110110100111011;
assign LUT_1[35250] = 32'b00000000000000000001010001010000;
assign LUT_1[35251] = 32'b11111111111111111010100011001100;
assign LUT_1[35252] = 32'b00000000000000001101011100010110;
assign LUT_1[35253] = 32'b00000000000000000110101110010010;
assign LUT_1[35254] = 32'b00000000000000001001001010100111;
assign LUT_1[35255] = 32'b00000000000000000010011100100011;
assign LUT_1[35256] = 32'b00000000000000000100110000110100;
assign LUT_1[35257] = 32'b11111111111111111110000010110000;
assign LUT_1[35258] = 32'b00000000000000000000011111000101;
assign LUT_1[35259] = 32'b11111111111111111001110001000001;
assign LUT_1[35260] = 32'b00000000000000001100101010001011;
assign LUT_1[35261] = 32'b00000000000000000101111100000111;
assign LUT_1[35262] = 32'b00000000000000001000011000011100;
assign LUT_1[35263] = 32'b00000000000000000001101010011000;
assign LUT_1[35264] = 32'b00000000000000000100101010000110;
assign LUT_1[35265] = 32'b11111111111111111101111100000010;
assign LUT_1[35266] = 32'b00000000000000000000011000010111;
assign LUT_1[35267] = 32'b11111111111111111001101010010011;
assign LUT_1[35268] = 32'b00000000000000001100100011011101;
assign LUT_1[35269] = 32'b00000000000000000101110101011001;
assign LUT_1[35270] = 32'b00000000000000001000010001101110;
assign LUT_1[35271] = 32'b00000000000000000001100011101010;
assign LUT_1[35272] = 32'b00000000000000000011110111111011;
assign LUT_1[35273] = 32'b11111111111111111101001001110111;
assign LUT_1[35274] = 32'b11111111111111111111100110001100;
assign LUT_1[35275] = 32'b11111111111111111000111000001000;
assign LUT_1[35276] = 32'b00000000000000001011110001010010;
assign LUT_1[35277] = 32'b00000000000000000101000011001110;
assign LUT_1[35278] = 32'b00000000000000000111011111100011;
assign LUT_1[35279] = 32'b00000000000000000000110001011111;
assign LUT_1[35280] = 32'b00000000000000000110100101101000;
assign LUT_1[35281] = 32'b11111111111111111111110111100100;
assign LUT_1[35282] = 32'b00000000000000000010010011111001;
assign LUT_1[35283] = 32'b11111111111111111011100101110101;
assign LUT_1[35284] = 32'b00000000000000001110011110111111;
assign LUT_1[35285] = 32'b00000000000000000111110000111011;
assign LUT_1[35286] = 32'b00000000000000001010001101010000;
assign LUT_1[35287] = 32'b00000000000000000011011111001100;
assign LUT_1[35288] = 32'b00000000000000000101110011011101;
assign LUT_1[35289] = 32'b11111111111111111111000101011001;
assign LUT_1[35290] = 32'b00000000000000000001100001101110;
assign LUT_1[35291] = 32'b11111111111111111010110011101010;
assign LUT_1[35292] = 32'b00000000000000001101101100110100;
assign LUT_1[35293] = 32'b00000000000000000110111110110000;
assign LUT_1[35294] = 32'b00000000000000001001011011000101;
assign LUT_1[35295] = 32'b00000000000000000010101101000001;
assign LUT_1[35296] = 32'b00000000000000000101100101000101;
assign LUT_1[35297] = 32'b11111111111111111110110111000001;
assign LUT_1[35298] = 32'b00000000000000000001010011010110;
assign LUT_1[35299] = 32'b11111111111111111010100101010010;
assign LUT_1[35300] = 32'b00000000000000001101011110011100;
assign LUT_1[35301] = 32'b00000000000000000110110000011000;
assign LUT_1[35302] = 32'b00000000000000001001001100101101;
assign LUT_1[35303] = 32'b00000000000000000010011110101001;
assign LUT_1[35304] = 32'b00000000000000000100110010111010;
assign LUT_1[35305] = 32'b11111111111111111110000100110110;
assign LUT_1[35306] = 32'b00000000000000000000100001001011;
assign LUT_1[35307] = 32'b11111111111111111001110011000111;
assign LUT_1[35308] = 32'b00000000000000001100101100010001;
assign LUT_1[35309] = 32'b00000000000000000101111110001101;
assign LUT_1[35310] = 32'b00000000000000001000011010100010;
assign LUT_1[35311] = 32'b00000000000000000001101100011110;
assign LUT_1[35312] = 32'b00000000000000000111100000100111;
assign LUT_1[35313] = 32'b00000000000000000000110010100011;
assign LUT_1[35314] = 32'b00000000000000000011001110111000;
assign LUT_1[35315] = 32'b11111111111111111100100000110100;
assign LUT_1[35316] = 32'b00000000000000001111011001111110;
assign LUT_1[35317] = 32'b00000000000000001000101011111010;
assign LUT_1[35318] = 32'b00000000000000001011001000001111;
assign LUT_1[35319] = 32'b00000000000000000100011010001011;
assign LUT_1[35320] = 32'b00000000000000000110101110011100;
assign LUT_1[35321] = 32'b00000000000000000000000000011000;
assign LUT_1[35322] = 32'b00000000000000000010011100101101;
assign LUT_1[35323] = 32'b11111111111111111011101110101001;
assign LUT_1[35324] = 32'b00000000000000001110100111110011;
assign LUT_1[35325] = 32'b00000000000000000111111001101111;
assign LUT_1[35326] = 32'b00000000000000001010010110000100;
assign LUT_1[35327] = 32'b00000000000000000011101000000000;
assign LUT_1[35328] = 32'b11111111111111111011100110101100;
assign LUT_1[35329] = 32'b11111111111111110100111000101000;
assign LUT_1[35330] = 32'b11111111111111110111010100111101;
assign LUT_1[35331] = 32'b11111111111111110000100110111001;
assign LUT_1[35332] = 32'b00000000000000000011100000000011;
assign LUT_1[35333] = 32'b11111111111111111100110001111111;
assign LUT_1[35334] = 32'b11111111111111111111001110010100;
assign LUT_1[35335] = 32'b11111111111111111000100000010000;
assign LUT_1[35336] = 32'b11111111111111111010110100100001;
assign LUT_1[35337] = 32'b11111111111111110100000110011101;
assign LUT_1[35338] = 32'b11111111111111110110100010110010;
assign LUT_1[35339] = 32'b11111111111111101111110100101110;
assign LUT_1[35340] = 32'b00000000000000000010101101111000;
assign LUT_1[35341] = 32'b11111111111111111011111111110100;
assign LUT_1[35342] = 32'b11111111111111111110011100001001;
assign LUT_1[35343] = 32'b11111111111111110111101110000101;
assign LUT_1[35344] = 32'b11111111111111111101100010001110;
assign LUT_1[35345] = 32'b11111111111111110110110100001010;
assign LUT_1[35346] = 32'b11111111111111111001010000011111;
assign LUT_1[35347] = 32'b11111111111111110010100010011011;
assign LUT_1[35348] = 32'b00000000000000000101011011100101;
assign LUT_1[35349] = 32'b11111111111111111110101101100001;
assign LUT_1[35350] = 32'b00000000000000000001001001110110;
assign LUT_1[35351] = 32'b11111111111111111010011011110010;
assign LUT_1[35352] = 32'b11111111111111111100110000000011;
assign LUT_1[35353] = 32'b11111111111111110110000001111111;
assign LUT_1[35354] = 32'b11111111111111111000011110010100;
assign LUT_1[35355] = 32'b11111111111111110001110000010000;
assign LUT_1[35356] = 32'b00000000000000000100101001011010;
assign LUT_1[35357] = 32'b11111111111111111101111011010110;
assign LUT_1[35358] = 32'b00000000000000000000010111101011;
assign LUT_1[35359] = 32'b11111111111111111001101001100111;
assign LUT_1[35360] = 32'b11111111111111111100100001101011;
assign LUT_1[35361] = 32'b11111111111111110101110011100111;
assign LUT_1[35362] = 32'b11111111111111111000001111111100;
assign LUT_1[35363] = 32'b11111111111111110001100001111000;
assign LUT_1[35364] = 32'b00000000000000000100011011000010;
assign LUT_1[35365] = 32'b11111111111111111101101100111110;
assign LUT_1[35366] = 32'b00000000000000000000001001010011;
assign LUT_1[35367] = 32'b11111111111111111001011011001111;
assign LUT_1[35368] = 32'b11111111111111111011101111100000;
assign LUT_1[35369] = 32'b11111111111111110101000001011100;
assign LUT_1[35370] = 32'b11111111111111110111011101110001;
assign LUT_1[35371] = 32'b11111111111111110000101111101101;
assign LUT_1[35372] = 32'b00000000000000000011101000110111;
assign LUT_1[35373] = 32'b11111111111111111100111010110011;
assign LUT_1[35374] = 32'b11111111111111111111010111001000;
assign LUT_1[35375] = 32'b11111111111111111000101001000100;
assign LUT_1[35376] = 32'b11111111111111111110011101001101;
assign LUT_1[35377] = 32'b11111111111111110111101111001001;
assign LUT_1[35378] = 32'b11111111111111111010001011011110;
assign LUT_1[35379] = 32'b11111111111111110011011101011010;
assign LUT_1[35380] = 32'b00000000000000000110010110100100;
assign LUT_1[35381] = 32'b11111111111111111111101000100000;
assign LUT_1[35382] = 32'b00000000000000000010000100110101;
assign LUT_1[35383] = 32'b11111111111111111011010110110001;
assign LUT_1[35384] = 32'b11111111111111111101101011000010;
assign LUT_1[35385] = 32'b11111111111111110110111100111110;
assign LUT_1[35386] = 32'b11111111111111111001011001010011;
assign LUT_1[35387] = 32'b11111111111111110010101011001111;
assign LUT_1[35388] = 32'b00000000000000000101100100011001;
assign LUT_1[35389] = 32'b11111111111111111110110110010101;
assign LUT_1[35390] = 32'b00000000000000000001010010101010;
assign LUT_1[35391] = 32'b11111111111111111010100100100110;
assign LUT_1[35392] = 32'b11111111111111111101100100010100;
assign LUT_1[35393] = 32'b11111111111111110110110110010000;
assign LUT_1[35394] = 32'b11111111111111111001010010100101;
assign LUT_1[35395] = 32'b11111111111111110010100100100001;
assign LUT_1[35396] = 32'b00000000000000000101011101101011;
assign LUT_1[35397] = 32'b11111111111111111110101111100111;
assign LUT_1[35398] = 32'b00000000000000000001001011111100;
assign LUT_1[35399] = 32'b11111111111111111010011101111000;
assign LUT_1[35400] = 32'b11111111111111111100110010001001;
assign LUT_1[35401] = 32'b11111111111111110110000100000101;
assign LUT_1[35402] = 32'b11111111111111111000100000011010;
assign LUT_1[35403] = 32'b11111111111111110001110010010110;
assign LUT_1[35404] = 32'b00000000000000000100101011100000;
assign LUT_1[35405] = 32'b11111111111111111101111101011100;
assign LUT_1[35406] = 32'b00000000000000000000011001110001;
assign LUT_1[35407] = 32'b11111111111111111001101011101101;
assign LUT_1[35408] = 32'b11111111111111111111011111110110;
assign LUT_1[35409] = 32'b11111111111111111000110001110010;
assign LUT_1[35410] = 32'b11111111111111111011001110000111;
assign LUT_1[35411] = 32'b11111111111111110100100000000011;
assign LUT_1[35412] = 32'b00000000000000000111011001001101;
assign LUT_1[35413] = 32'b00000000000000000000101011001001;
assign LUT_1[35414] = 32'b00000000000000000011000111011110;
assign LUT_1[35415] = 32'b11111111111111111100011001011010;
assign LUT_1[35416] = 32'b11111111111111111110101101101011;
assign LUT_1[35417] = 32'b11111111111111110111111111100111;
assign LUT_1[35418] = 32'b11111111111111111010011011111100;
assign LUT_1[35419] = 32'b11111111111111110011101101111000;
assign LUT_1[35420] = 32'b00000000000000000110100111000010;
assign LUT_1[35421] = 32'b11111111111111111111111000111110;
assign LUT_1[35422] = 32'b00000000000000000010010101010011;
assign LUT_1[35423] = 32'b11111111111111111011100111001111;
assign LUT_1[35424] = 32'b11111111111111111110011111010011;
assign LUT_1[35425] = 32'b11111111111111110111110001001111;
assign LUT_1[35426] = 32'b11111111111111111010001101100100;
assign LUT_1[35427] = 32'b11111111111111110011011111100000;
assign LUT_1[35428] = 32'b00000000000000000110011000101010;
assign LUT_1[35429] = 32'b11111111111111111111101010100110;
assign LUT_1[35430] = 32'b00000000000000000010000110111011;
assign LUT_1[35431] = 32'b11111111111111111011011000110111;
assign LUT_1[35432] = 32'b11111111111111111101101101001000;
assign LUT_1[35433] = 32'b11111111111111110110111111000100;
assign LUT_1[35434] = 32'b11111111111111111001011011011001;
assign LUT_1[35435] = 32'b11111111111111110010101101010101;
assign LUT_1[35436] = 32'b00000000000000000101100110011111;
assign LUT_1[35437] = 32'b11111111111111111110111000011011;
assign LUT_1[35438] = 32'b00000000000000000001010100110000;
assign LUT_1[35439] = 32'b11111111111111111010100110101100;
assign LUT_1[35440] = 32'b00000000000000000000011010110101;
assign LUT_1[35441] = 32'b11111111111111111001101100110001;
assign LUT_1[35442] = 32'b11111111111111111100001001000110;
assign LUT_1[35443] = 32'b11111111111111110101011011000010;
assign LUT_1[35444] = 32'b00000000000000001000010100001100;
assign LUT_1[35445] = 32'b00000000000000000001100110001000;
assign LUT_1[35446] = 32'b00000000000000000100000010011101;
assign LUT_1[35447] = 32'b11111111111111111101010100011001;
assign LUT_1[35448] = 32'b11111111111111111111101000101010;
assign LUT_1[35449] = 32'b11111111111111111000111010100110;
assign LUT_1[35450] = 32'b11111111111111111011010110111011;
assign LUT_1[35451] = 32'b11111111111111110100101000110111;
assign LUT_1[35452] = 32'b00000000000000000111100010000001;
assign LUT_1[35453] = 32'b00000000000000000000110011111101;
assign LUT_1[35454] = 32'b00000000000000000011010000010010;
assign LUT_1[35455] = 32'b11111111111111111100100010001110;
assign LUT_1[35456] = 32'b11111111111111111110100110101111;
assign LUT_1[35457] = 32'b11111111111111110111111000101011;
assign LUT_1[35458] = 32'b11111111111111111010010101000000;
assign LUT_1[35459] = 32'b11111111111111110011100110111100;
assign LUT_1[35460] = 32'b00000000000000000110100000000110;
assign LUT_1[35461] = 32'b11111111111111111111110010000010;
assign LUT_1[35462] = 32'b00000000000000000010001110010111;
assign LUT_1[35463] = 32'b11111111111111111011100000010011;
assign LUT_1[35464] = 32'b11111111111111111101110100100100;
assign LUT_1[35465] = 32'b11111111111111110111000110100000;
assign LUT_1[35466] = 32'b11111111111111111001100010110101;
assign LUT_1[35467] = 32'b11111111111111110010110100110001;
assign LUT_1[35468] = 32'b00000000000000000101101101111011;
assign LUT_1[35469] = 32'b11111111111111111110111111110111;
assign LUT_1[35470] = 32'b00000000000000000001011100001100;
assign LUT_1[35471] = 32'b11111111111111111010101110001000;
assign LUT_1[35472] = 32'b00000000000000000000100010010001;
assign LUT_1[35473] = 32'b11111111111111111001110100001101;
assign LUT_1[35474] = 32'b11111111111111111100010000100010;
assign LUT_1[35475] = 32'b11111111111111110101100010011110;
assign LUT_1[35476] = 32'b00000000000000001000011011101000;
assign LUT_1[35477] = 32'b00000000000000000001101101100100;
assign LUT_1[35478] = 32'b00000000000000000100001001111001;
assign LUT_1[35479] = 32'b11111111111111111101011011110101;
assign LUT_1[35480] = 32'b11111111111111111111110000000110;
assign LUT_1[35481] = 32'b11111111111111111001000010000010;
assign LUT_1[35482] = 32'b11111111111111111011011110010111;
assign LUT_1[35483] = 32'b11111111111111110100110000010011;
assign LUT_1[35484] = 32'b00000000000000000111101001011101;
assign LUT_1[35485] = 32'b00000000000000000000111011011001;
assign LUT_1[35486] = 32'b00000000000000000011010111101110;
assign LUT_1[35487] = 32'b11111111111111111100101001101010;
assign LUT_1[35488] = 32'b11111111111111111111100001101110;
assign LUT_1[35489] = 32'b11111111111111111000110011101010;
assign LUT_1[35490] = 32'b11111111111111111011001111111111;
assign LUT_1[35491] = 32'b11111111111111110100100001111011;
assign LUT_1[35492] = 32'b00000000000000000111011011000101;
assign LUT_1[35493] = 32'b00000000000000000000101101000001;
assign LUT_1[35494] = 32'b00000000000000000011001001010110;
assign LUT_1[35495] = 32'b11111111111111111100011011010010;
assign LUT_1[35496] = 32'b11111111111111111110101111100011;
assign LUT_1[35497] = 32'b11111111111111111000000001011111;
assign LUT_1[35498] = 32'b11111111111111111010011101110100;
assign LUT_1[35499] = 32'b11111111111111110011101111110000;
assign LUT_1[35500] = 32'b00000000000000000110101000111010;
assign LUT_1[35501] = 32'b11111111111111111111111010110110;
assign LUT_1[35502] = 32'b00000000000000000010010111001011;
assign LUT_1[35503] = 32'b11111111111111111011101001000111;
assign LUT_1[35504] = 32'b00000000000000000001011101010000;
assign LUT_1[35505] = 32'b11111111111111111010101111001100;
assign LUT_1[35506] = 32'b11111111111111111101001011100001;
assign LUT_1[35507] = 32'b11111111111111110110011101011101;
assign LUT_1[35508] = 32'b00000000000000001001010110100111;
assign LUT_1[35509] = 32'b00000000000000000010101000100011;
assign LUT_1[35510] = 32'b00000000000000000101000100111000;
assign LUT_1[35511] = 32'b11111111111111111110010110110100;
assign LUT_1[35512] = 32'b00000000000000000000101011000101;
assign LUT_1[35513] = 32'b11111111111111111001111101000001;
assign LUT_1[35514] = 32'b11111111111111111100011001010110;
assign LUT_1[35515] = 32'b11111111111111110101101011010010;
assign LUT_1[35516] = 32'b00000000000000001000100100011100;
assign LUT_1[35517] = 32'b00000000000000000001110110011000;
assign LUT_1[35518] = 32'b00000000000000000100010010101101;
assign LUT_1[35519] = 32'b11111111111111111101100100101001;
assign LUT_1[35520] = 32'b00000000000000000000100100010111;
assign LUT_1[35521] = 32'b11111111111111111001110110010011;
assign LUT_1[35522] = 32'b11111111111111111100010010101000;
assign LUT_1[35523] = 32'b11111111111111110101100100100100;
assign LUT_1[35524] = 32'b00000000000000001000011101101110;
assign LUT_1[35525] = 32'b00000000000000000001101111101010;
assign LUT_1[35526] = 32'b00000000000000000100001011111111;
assign LUT_1[35527] = 32'b11111111111111111101011101111011;
assign LUT_1[35528] = 32'b11111111111111111111110010001100;
assign LUT_1[35529] = 32'b11111111111111111001000100001000;
assign LUT_1[35530] = 32'b11111111111111111011100000011101;
assign LUT_1[35531] = 32'b11111111111111110100110010011001;
assign LUT_1[35532] = 32'b00000000000000000111101011100011;
assign LUT_1[35533] = 32'b00000000000000000000111101011111;
assign LUT_1[35534] = 32'b00000000000000000011011001110100;
assign LUT_1[35535] = 32'b11111111111111111100101011110000;
assign LUT_1[35536] = 32'b00000000000000000010011111111001;
assign LUT_1[35537] = 32'b11111111111111111011110001110101;
assign LUT_1[35538] = 32'b11111111111111111110001110001010;
assign LUT_1[35539] = 32'b11111111111111110111100000000110;
assign LUT_1[35540] = 32'b00000000000000001010011001010000;
assign LUT_1[35541] = 32'b00000000000000000011101011001100;
assign LUT_1[35542] = 32'b00000000000000000110000111100001;
assign LUT_1[35543] = 32'b11111111111111111111011001011101;
assign LUT_1[35544] = 32'b00000000000000000001101101101110;
assign LUT_1[35545] = 32'b11111111111111111010111111101010;
assign LUT_1[35546] = 32'b11111111111111111101011011111111;
assign LUT_1[35547] = 32'b11111111111111110110101101111011;
assign LUT_1[35548] = 32'b00000000000000001001100111000101;
assign LUT_1[35549] = 32'b00000000000000000010111001000001;
assign LUT_1[35550] = 32'b00000000000000000101010101010110;
assign LUT_1[35551] = 32'b11111111111111111110100111010010;
assign LUT_1[35552] = 32'b00000000000000000001011111010110;
assign LUT_1[35553] = 32'b11111111111111111010110001010010;
assign LUT_1[35554] = 32'b11111111111111111101001101100111;
assign LUT_1[35555] = 32'b11111111111111110110011111100011;
assign LUT_1[35556] = 32'b00000000000000001001011000101101;
assign LUT_1[35557] = 32'b00000000000000000010101010101001;
assign LUT_1[35558] = 32'b00000000000000000101000110111110;
assign LUT_1[35559] = 32'b11111111111111111110011000111010;
assign LUT_1[35560] = 32'b00000000000000000000101101001011;
assign LUT_1[35561] = 32'b11111111111111111001111111000111;
assign LUT_1[35562] = 32'b11111111111111111100011011011100;
assign LUT_1[35563] = 32'b11111111111111110101101101011000;
assign LUT_1[35564] = 32'b00000000000000001000100110100010;
assign LUT_1[35565] = 32'b00000000000000000001111000011110;
assign LUT_1[35566] = 32'b00000000000000000100010100110011;
assign LUT_1[35567] = 32'b11111111111111111101100110101111;
assign LUT_1[35568] = 32'b00000000000000000011011010111000;
assign LUT_1[35569] = 32'b11111111111111111100101100110100;
assign LUT_1[35570] = 32'b11111111111111111111001001001001;
assign LUT_1[35571] = 32'b11111111111111111000011011000101;
assign LUT_1[35572] = 32'b00000000000000001011010100001111;
assign LUT_1[35573] = 32'b00000000000000000100100110001011;
assign LUT_1[35574] = 32'b00000000000000000111000010100000;
assign LUT_1[35575] = 32'b00000000000000000000010100011100;
assign LUT_1[35576] = 32'b00000000000000000010101000101101;
assign LUT_1[35577] = 32'b11111111111111111011111010101001;
assign LUT_1[35578] = 32'b11111111111111111110010110111110;
assign LUT_1[35579] = 32'b11111111111111110111101000111010;
assign LUT_1[35580] = 32'b00000000000000001010100010000100;
assign LUT_1[35581] = 32'b00000000000000000011110100000000;
assign LUT_1[35582] = 32'b00000000000000000110010000010101;
assign LUT_1[35583] = 32'b11111111111111111111100010010001;
assign LUT_1[35584] = 32'b11111111111111111001011010111000;
assign LUT_1[35585] = 32'b11111111111111110010101100110100;
assign LUT_1[35586] = 32'b11111111111111110101001001001001;
assign LUT_1[35587] = 32'b11111111111111101110011011000101;
assign LUT_1[35588] = 32'b00000000000000000001010100001111;
assign LUT_1[35589] = 32'b11111111111111111010100110001011;
assign LUT_1[35590] = 32'b11111111111111111101000010100000;
assign LUT_1[35591] = 32'b11111111111111110110010100011100;
assign LUT_1[35592] = 32'b11111111111111111000101000101101;
assign LUT_1[35593] = 32'b11111111111111110001111010101001;
assign LUT_1[35594] = 32'b11111111111111110100010110111110;
assign LUT_1[35595] = 32'b11111111111111101101101000111010;
assign LUT_1[35596] = 32'b00000000000000000000100010000100;
assign LUT_1[35597] = 32'b11111111111111111001110100000000;
assign LUT_1[35598] = 32'b11111111111111111100010000010101;
assign LUT_1[35599] = 32'b11111111111111110101100010010001;
assign LUT_1[35600] = 32'b11111111111111111011010110011010;
assign LUT_1[35601] = 32'b11111111111111110100101000010110;
assign LUT_1[35602] = 32'b11111111111111110111000100101011;
assign LUT_1[35603] = 32'b11111111111111110000010110100111;
assign LUT_1[35604] = 32'b00000000000000000011001111110001;
assign LUT_1[35605] = 32'b11111111111111111100100001101101;
assign LUT_1[35606] = 32'b11111111111111111110111110000010;
assign LUT_1[35607] = 32'b11111111111111111000001111111110;
assign LUT_1[35608] = 32'b11111111111111111010100100001111;
assign LUT_1[35609] = 32'b11111111111111110011110110001011;
assign LUT_1[35610] = 32'b11111111111111110110010010100000;
assign LUT_1[35611] = 32'b11111111111111101111100100011100;
assign LUT_1[35612] = 32'b00000000000000000010011101100110;
assign LUT_1[35613] = 32'b11111111111111111011101111100010;
assign LUT_1[35614] = 32'b11111111111111111110001011110111;
assign LUT_1[35615] = 32'b11111111111111110111011101110011;
assign LUT_1[35616] = 32'b11111111111111111010010101110111;
assign LUT_1[35617] = 32'b11111111111111110011100111110011;
assign LUT_1[35618] = 32'b11111111111111110110000100001000;
assign LUT_1[35619] = 32'b11111111111111101111010110000100;
assign LUT_1[35620] = 32'b00000000000000000010001111001110;
assign LUT_1[35621] = 32'b11111111111111111011100001001010;
assign LUT_1[35622] = 32'b11111111111111111101111101011111;
assign LUT_1[35623] = 32'b11111111111111110111001111011011;
assign LUT_1[35624] = 32'b11111111111111111001100011101100;
assign LUT_1[35625] = 32'b11111111111111110010110101101000;
assign LUT_1[35626] = 32'b11111111111111110101010001111101;
assign LUT_1[35627] = 32'b11111111111111101110100011111001;
assign LUT_1[35628] = 32'b00000000000000000001011101000011;
assign LUT_1[35629] = 32'b11111111111111111010101110111111;
assign LUT_1[35630] = 32'b11111111111111111101001011010100;
assign LUT_1[35631] = 32'b11111111111111110110011101010000;
assign LUT_1[35632] = 32'b11111111111111111100010001011001;
assign LUT_1[35633] = 32'b11111111111111110101100011010101;
assign LUT_1[35634] = 32'b11111111111111110111111111101010;
assign LUT_1[35635] = 32'b11111111111111110001010001100110;
assign LUT_1[35636] = 32'b00000000000000000100001010110000;
assign LUT_1[35637] = 32'b11111111111111111101011100101100;
assign LUT_1[35638] = 32'b11111111111111111111111001000001;
assign LUT_1[35639] = 32'b11111111111111111001001010111101;
assign LUT_1[35640] = 32'b11111111111111111011011111001110;
assign LUT_1[35641] = 32'b11111111111111110100110001001010;
assign LUT_1[35642] = 32'b11111111111111110111001101011111;
assign LUT_1[35643] = 32'b11111111111111110000011111011011;
assign LUT_1[35644] = 32'b00000000000000000011011000100101;
assign LUT_1[35645] = 32'b11111111111111111100101010100001;
assign LUT_1[35646] = 32'b11111111111111111111000110110110;
assign LUT_1[35647] = 32'b11111111111111111000011000110010;
assign LUT_1[35648] = 32'b11111111111111111011011000100000;
assign LUT_1[35649] = 32'b11111111111111110100101010011100;
assign LUT_1[35650] = 32'b11111111111111110111000110110001;
assign LUT_1[35651] = 32'b11111111111111110000011000101101;
assign LUT_1[35652] = 32'b00000000000000000011010001110111;
assign LUT_1[35653] = 32'b11111111111111111100100011110011;
assign LUT_1[35654] = 32'b11111111111111111111000000001000;
assign LUT_1[35655] = 32'b11111111111111111000010010000100;
assign LUT_1[35656] = 32'b11111111111111111010100110010101;
assign LUT_1[35657] = 32'b11111111111111110011111000010001;
assign LUT_1[35658] = 32'b11111111111111110110010100100110;
assign LUT_1[35659] = 32'b11111111111111101111100110100010;
assign LUT_1[35660] = 32'b00000000000000000010011111101100;
assign LUT_1[35661] = 32'b11111111111111111011110001101000;
assign LUT_1[35662] = 32'b11111111111111111110001101111101;
assign LUT_1[35663] = 32'b11111111111111110111011111111001;
assign LUT_1[35664] = 32'b11111111111111111101010100000010;
assign LUT_1[35665] = 32'b11111111111111110110100101111110;
assign LUT_1[35666] = 32'b11111111111111111001000010010011;
assign LUT_1[35667] = 32'b11111111111111110010010100001111;
assign LUT_1[35668] = 32'b00000000000000000101001101011001;
assign LUT_1[35669] = 32'b11111111111111111110011111010101;
assign LUT_1[35670] = 32'b00000000000000000000111011101010;
assign LUT_1[35671] = 32'b11111111111111111010001101100110;
assign LUT_1[35672] = 32'b11111111111111111100100001110111;
assign LUT_1[35673] = 32'b11111111111111110101110011110011;
assign LUT_1[35674] = 32'b11111111111111111000010000001000;
assign LUT_1[35675] = 32'b11111111111111110001100010000100;
assign LUT_1[35676] = 32'b00000000000000000100011011001110;
assign LUT_1[35677] = 32'b11111111111111111101101101001010;
assign LUT_1[35678] = 32'b00000000000000000000001001011111;
assign LUT_1[35679] = 32'b11111111111111111001011011011011;
assign LUT_1[35680] = 32'b11111111111111111100010011011111;
assign LUT_1[35681] = 32'b11111111111111110101100101011011;
assign LUT_1[35682] = 32'b11111111111111111000000001110000;
assign LUT_1[35683] = 32'b11111111111111110001010011101100;
assign LUT_1[35684] = 32'b00000000000000000100001100110110;
assign LUT_1[35685] = 32'b11111111111111111101011110110010;
assign LUT_1[35686] = 32'b11111111111111111111111011000111;
assign LUT_1[35687] = 32'b11111111111111111001001101000011;
assign LUT_1[35688] = 32'b11111111111111111011100001010100;
assign LUT_1[35689] = 32'b11111111111111110100110011010000;
assign LUT_1[35690] = 32'b11111111111111110111001111100101;
assign LUT_1[35691] = 32'b11111111111111110000100001100001;
assign LUT_1[35692] = 32'b00000000000000000011011010101011;
assign LUT_1[35693] = 32'b11111111111111111100101100100111;
assign LUT_1[35694] = 32'b11111111111111111111001000111100;
assign LUT_1[35695] = 32'b11111111111111111000011010111000;
assign LUT_1[35696] = 32'b11111111111111111110001111000001;
assign LUT_1[35697] = 32'b11111111111111110111100000111101;
assign LUT_1[35698] = 32'b11111111111111111001111101010010;
assign LUT_1[35699] = 32'b11111111111111110011001111001110;
assign LUT_1[35700] = 32'b00000000000000000110001000011000;
assign LUT_1[35701] = 32'b11111111111111111111011010010100;
assign LUT_1[35702] = 32'b00000000000000000001110110101001;
assign LUT_1[35703] = 32'b11111111111111111011001000100101;
assign LUT_1[35704] = 32'b11111111111111111101011100110110;
assign LUT_1[35705] = 32'b11111111111111110110101110110010;
assign LUT_1[35706] = 32'b11111111111111111001001011000111;
assign LUT_1[35707] = 32'b11111111111111110010011101000011;
assign LUT_1[35708] = 32'b00000000000000000101010110001101;
assign LUT_1[35709] = 32'b11111111111111111110101000001001;
assign LUT_1[35710] = 32'b00000000000000000001000100011110;
assign LUT_1[35711] = 32'b11111111111111111010010110011010;
assign LUT_1[35712] = 32'b11111111111111111100011010111011;
assign LUT_1[35713] = 32'b11111111111111110101101100110111;
assign LUT_1[35714] = 32'b11111111111111111000001001001100;
assign LUT_1[35715] = 32'b11111111111111110001011011001000;
assign LUT_1[35716] = 32'b00000000000000000100010100010010;
assign LUT_1[35717] = 32'b11111111111111111101100110001110;
assign LUT_1[35718] = 32'b00000000000000000000000010100011;
assign LUT_1[35719] = 32'b11111111111111111001010100011111;
assign LUT_1[35720] = 32'b11111111111111111011101000110000;
assign LUT_1[35721] = 32'b11111111111111110100111010101100;
assign LUT_1[35722] = 32'b11111111111111110111010111000001;
assign LUT_1[35723] = 32'b11111111111111110000101000111101;
assign LUT_1[35724] = 32'b00000000000000000011100010000111;
assign LUT_1[35725] = 32'b11111111111111111100110100000011;
assign LUT_1[35726] = 32'b11111111111111111111010000011000;
assign LUT_1[35727] = 32'b11111111111111111000100010010100;
assign LUT_1[35728] = 32'b11111111111111111110010110011101;
assign LUT_1[35729] = 32'b11111111111111110111101000011001;
assign LUT_1[35730] = 32'b11111111111111111010000100101110;
assign LUT_1[35731] = 32'b11111111111111110011010110101010;
assign LUT_1[35732] = 32'b00000000000000000110001111110100;
assign LUT_1[35733] = 32'b11111111111111111111100001110000;
assign LUT_1[35734] = 32'b00000000000000000001111110000101;
assign LUT_1[35735] = 32'b11111111111111111011010000000001;
assign LUT_1[35736] = 32'b11111111111111111101100100010010;
assign LUT_1[35737] = 32'b11111111111111110110110110001110;
assign LUT_1[35738] = 32'b11111111111111111001010010100011;
assign LUT_1[35739] = 32'b11111111111111110010100100011111;
assign LUT_1[35740] = 32'b00000000000000000101011101101001;
assign LUT_1[35741] = 32'b11111111111111111110101111100101;
assign LUT_1[35742] = 32'b00000000000000000001001011111010;
assign LUT_1[35743] = 32'b11111111111111111010011101110110;
assign LUT_1[35744] = 32'b11111111111111111101010101111010;
assign LUT_1[35745] = 32'b11111111111111110110100111110110;
assign LUT_1[35746] = 32'b11111111111111111001000100001011;
assign LUT_1[35747] = 32'b11111111111111110010010110000111;
assign LUT_1[35748] = 32'b00000000000000000101001111010001;
assign LUT_1[35749] = 32'b11111111111111111110100001001101;
assign LUT_1[35750] = 32'b00000000000000000000111101100010;
assign LUT_1[35751] = 32'b11111111111111111010001111011110;
assign LUT_1[35752] = 32'b11111111111111111100100011101111;
assign LUT_1[35753] = 32'b11111111111111110101110101101011;
assign LUT_1[35754] = 32'b11111111111111111000010010000000;
assign LUT_1[35755] = 32'b11111111111111110001100011111100;
assign LUT_1[35756] = 32'b00000000000000000100011101000110;
assign LUT_1[35757] = 32'b11111111111111111101101111000010;
assign LUT_1[35758] = 32'b00000000000000000000001011010111;
assign LUT_1[35759] = 32'b11111111111111111001011101010011;
assign LUT_1[35760] = 32'b11111111111111111111010001011100;
assign LUT_1[35761] = 32'b11111111111111111000100011011000;
assign LUT_1[35762] = 32'b11111111111111111010111111101101;
assign LUT_1[35763] = 32'b11111111111111110100010001101001;
assign LUT_1[35764] = 32'b00000000000000000111001010110011;
assign LUT_1[35765] = 32'b00000000000000000000011100101111;
assign LUT_1[35766] = 32'b00000000000000000010111001000100;
assign LUT_1[35767] = 32'b11111111111111111100001011000000;
assign LUT_1[35768] = 32'b11111111111111111110011111010001;
assign LUT_1[35769] = 32'b11111111111111110111110001001101;
assign LUT_1[35770] = 32'b11111111111111111010001101100010;
assign LUT_1[35771] = 32'b11111111111111110011011111011110;
assign LUT_1[35772] = 32'b00000000000000000110011000101000;
assign LUT_1[35773] = 32'b11111111111111111111101010100100;
assign LUT_1[35774] = 32'b00000000000000000010000110111001;
assign LUT_1[35775] = 32'b11111111111111111011011000110101;
assign LUT_1[35776] = 32'b11111111111111111110011000100011;
assign LUT_1[35777] = 32'b11111111111111110111101010011111;
assign LUT_1[35778] = 32'b11111111111111111010000110110100;
assign LUT_1[35779] = 32'b11111111111111110011011000110000;
assign LUT_1[35780] = 32'b00000000000000000110010001111010;
assign LUT_1[35781] = 32'b11111111111111111111100011110110;
assign LUT_1[35782] = 32'b00000000000000000010000000001011;
assign LUT_1[35783] = 32'b11111111111111111011010010000111;
assign LUT_1[35784] = 32'b11111111111111111101100110011000;
assign LUT_1[35785] = 32'b11111111111111110110111000010100;
assign LUT_1[35786] = 32'b11111111111111111001010100101001;
assign LUT_1[35787] = 32'b11111111111111110010100110100101;
assign LUT_1[35788] = 32'b00000000000000000101011111101111;
assign LUT_1[35789] = 32'b11111111111111111110110001101011;
assign LUT_1[35790] = 32'b00000000000000000001001110000000;
assign LUT_1[35791] = 32'b11111111111111111010011111111100;
assign LUT_1[35792] = 32'b00000000000000000000010100000101;
assign LUT_1[35793] = 32'b11111111111111111001100110000001;
assign LUT_1[35794] = 32'b11111111111111111100000010010110;
assign LUT_1[35795] = 32'b11111111111111110101010100010010;
assign LUT_1[35796] = 32'b00000000000000001000001101011100;
assign LUT_1[35797] = 32'b00000000000000000001011111011000;
assign LUT_1[35798] = 32'b00000000000000000011111011101101;
assign LUT_1[35799] = 32'b11111111111111111101001101101001;
assign LUT_1[35800] = 32'b11111111111111111111100001111010;
assign LUT_1[35801] = 32'b11111111111111111000110011110110;
assign LUT_1[35802] = 32'b11111111111111111011010000001011;
assign LUT_1[35803] = 32'b11111111111111110100100010000111;
assign LUT_1[35804] = 32'b00000000000000000111011011010001;
assign LUT_1[35805] = 32'b00000000000000000000101101001101;
assign LUT_1[35806] = 32'b00000000000000000011001001100010;
assign LUT_1[35807] = 32'b11111111111111111100011011011110;
assign LUT_1[35808] = 32'b11111111111111111111010011100010;
assign LUT_1[35809] = 32'b11111111111111111000100101011110;
assign LUT_1[35810] = 32'b11111111111111111011000001110011;
assign LUT_1[35811] = 32'b11111111111111110100010011101111;
assign LUT_1[35812] = 32'b00000000000000000111001100111001;
assign LUT_1[35813] = 32'b00000000000000000000011110110101;
assign LUT_1[35814] = 32'b00000000000000000010111011001010;
assign LUT_1[35815] = 32'b11111111111111111100001101000110;
assign LUT_1[35816] = 32'b11111111111111111110100001010111;
assign LUT_1[35817] = 32'b11111111111111110111110011010011;
assign LUT_1[35818] = 32'b11111111111111111010001111101000;
assign LUT_1[35819] = 32'b11111111111111110011100001100100;
assign LUT_1[35820] = 32'b00000000000000000110011010101110;
assign LUT_1[35821] = 32'b11111111111111111111101100101010;
assign LUT_1[35822] = 32'b00000000000000000010001000111111;
assign LUT_1[35823] = 32'b11111111111111111011011010111011;
assign LUT_1[35824] = 32'b00000000000000000001001111000100;
assign LUT_1[35825] = 32'b11111111111111111010100001000000;
assign LUT_1[35826] = 32'b11111111111111111100111101010101;
assign LUT_1[35827] = 32'b11111111111111110110001111010001;
assign LUT_1[35828] = 32'b00000000000000001001001000011011;
assign LUT_1[35829] = 32'b00000000000000000010011010010111;
assign LUT_1[35830] = 32'b00000000000000000100110110101100;
assign LUT_1[35831] = 32'b11111111111111111110001000101000;
assign LUT_1[35832] = 32'b00000000000000000000011100111001;
assign LUT_1[35833] = 32'b11111111111111111001101110110101;
assign LUT_1[35834] = 32'b11111111111111111100001011001010;
assign LUT_1[35835] = 32'b11111111111111110101011101000110;
assign LUT_1[35836] = 32'b00000000000000001000010110010000;
assign LUT_1[35837] = 32'b00000000000000000001101000001100;
assign LUT_1[35838] = 32'b00000000000000000100000100100001;
assign LUT_1[35839] = 32'b11111111111111111101010110011101;
assign LUT_1[35840] = 32'b00000000000000001000001110111111;
assign LUT_1[35841] = 32'b00000000000000000001100000111011;
assign LUT_1[35842] = 32'b00000000000000000011111101010000;
assign LUT_1[35843] = 32'b11111111111111111101001111001100;
assign LUT_1[35844] = 32'b00000000000000010000001000010110;
assign LUT_1[35845] = 32'b00000000000000001001011010010010;
assign LUT_1[35846] = 32'b00000000000000001011110110100111;
assign LUT_1[35847] = 32'b00000000000000000101001000100011;
assign LUT_1[35848] = 32'b00000000000000000111011100110100;
assign LUT_1[35849] = 32'b00000000000000000000101110110000;
assign LUT_1[35850] = 32'b00000000000000000011001011000101;
assign LUT_1[35851] = 32'b11111111111111111100011101000001;
assign LUT_1[35852] = 32'b00000000000000001111010110001011;
assign LUT_1[35853] = 32'b00000000000000001000101000000111;
assign LUT_1[35854] = 32'b00000000000000001011000100011100;
assign LUT_1[35855] = 32'b00000000000000000100010110011000;
assign LUT_1[35856] = 32'b00000000000000001010001010100001;
assign LUT_1[35857] = 32'b00000000000000000011011100011101;
assign LUT_1[35858] = 32'b00000000000000000101111000110010;
assign LUT_1[35859] = 32'b11111111111111111111001010101110;
assign LUT_1[35860] = 32'b00000000000000010010000011111000;
assign LUT_1[35861] = 32'b00000000000000001011010101110100;
assign LUT_1[35862] = 32'b00000000000000001101110010001001;
assign LUT_1[35863] = 32'b00000000000000000111000100000101;
assign LUT_1[35864] = 32'b00000000000000001001011000010110;
assign LUT_1[35865] = 32'b00000000000000000010101010010010;
assign LUT_1[35866] = 32'b00000000000000000101000110100111;
assign LUT_1[35867] = 32'b11111111111111111110011000100011;
assign LUT_1[35868] = 32'b00000000000000010001010001101101;
assign LUT_1[35869] = 32'b00000000000000001010100011101001;
assign LUT_1[35870] = 32'b00000000000000001100111111111110;
assign LUT_1[35871] = 32'b00000000000000000110010001111010;
assign LUT_1[35872] = 32'b00000000000000001001001001111110;
assign LUT_1[35873] = 32'b00000000000000000010011011111010;
assign LUT_1[35874] = 32'b00000000000000000100111000001111;
assign LUT_1[35875] = 32'b11111111111111111110001010001011;
assign LUT_1[35876] = 32'b00000000000000010001000011010101;
assign LUT_1[35877] = 32'b00000000000000001010010101010001;
assign LUT_1[35878] = 32'b00000000000000001100110001100110;
assign LUT_1[35879] = 32'b00000000000000000110000011100010;
assign LUT_1[35880] = 32'b00000000000000001000010111110011;
assign LUT_1[35881] = 32'b00000000000000000001101001101111;
assign LUT_1[35882] = 32'b00000000000000000100000110000100;
assign LUT_1[35883] = 32'b11111111111111111101011000000000;
assign LUT_1[35884] = 32'b00000000000000010000010001001010;
assign LUT_1[35885] = 32'b00000000000000001001100011000110;
assign LUT_1[35886] = 32'b00000000000000001011111111011011;
assign LUT_1[35887] = 32'b00000000000000000101010001010111;
assign LUT_1[35888] = 32'b00000000000000001011000101100000;
assign LUT_1[35889] = 32'b00000000000000000100010111011100;
assign LUT_1[35890] = 32'b00000000000000000110110011110001;
assign LUT_1[35891] = 32'b00000000000000000000000101101101;
assign LUT_1[35892] = 32'b00000000000000010010111110110111;
assign LUT_1[35893] = 32'b00000000000000001100010000110011;
assign LUT_1[35894] = 32'b00000000000000001110101101001000;
assign LUT_1[35895] = 32'b00000000000000000111111111000100;
assign LUT_1[35896] = 32'b00000000000000001010010011010101;
assign LUT_1[35897] = 32'b00000000000000000011100101010001;
assign LUT_1[35898] = 32'b00000000000000000110000001100110;
assign LUT_1[35899] = 32'b11111111111111111111010011100010;
assign LUT_1[35900] = 32'b00000000000000010010001100101100;
assign LUT_1[35901] = 32'b00000000000000001011011110101000;
assign LUT_1[35902] = 32'b00000000000000001101111010111101;
assign LUT_1[35903] = 32'b00000000000000000111001100111001;
assign LUT_1[35904] = 32'b00000000000000001010001100100111;
assign LUT_1[35905] = 32'b00000000000000000011011110100011;
assign LUT_1[35906] = 32'b00000000000000000101111010111000;
assign LUT_1[35907] = 32'b11111111111111111111001100110100;
assign LUT_1[35908] = 32'b00000000000000010010000101111110;
assign LUT_1[35909] = 32'b00000000000000001011010111111010;
assign LUT_1[35910] = 32'b00000000000000001101110100001111;
assign LUT_1[35911] = 32'b00000000000000000111000110001011;
assign LUT_1[35912] = 32'b00000000000000001001011010011100;
assign LUT_1[35913] = 32'b00000000000000000010101100011000;
assign LUT_1[35914] = 32'b00000000000000000101001000101101;
assign LUT_1[35915] = 32'b11111111111111111110011010101001;
assign LUT_1[35916] = 32'b00000000000000010001010011110011;
assign LUT_1[35917] = 32'b00000000000000001010100101101111;
assign LUT_1[35918] = 32'b00000000000000001101000010000100;
assign LUT_1[35919] = 32'b00000000000000000110010100000000;
assign LUT_1[35920] = 32'b00000000000000001100001000001001;
assign LUT_1[35921] = 32'b00000000000000000101011010000101;
assign LUT_1[35922] = 32'b00000000000000000111110110011010;
assign LUT_1[35923] = 32'b00000000000000000001001000010110;
assign LUT_1[35924] = 32'b00000000000000010100000001100000;
assign LUT_1[35925] = 32'b00000000000000001101010011011100;
assign LUT_1[35926] = 32'b00000000000000001111101111110001;
assign LUT_1[35927] = 32'b00000000000000001001000001101101;
assign LUT_1[35928] = 32'b00000000000000001011010101111110;
assign LUT_1[35929] = 32'b00000000000000000100100111111010;
assign LUT_1[35930] = 32'b00000000000000000111000100001111;
assign LUT_1[35931] = 32'b00000000000000000000010110001011;
assign LUT_1[35932] = 32'b00000000000000010011001111010101;
assign LUT_1[35933] = 32'b00000000000000001100100001010001;
assign LUT_1[35934] = 32'b00000000000000001110111101100110;
assign LUT_1[35935] = 32'b00000000000000001000001111100010;
assign LUT_1[35936] = 32'b00000000000000001011000111100110;
assign LUT_1[35937] = 32'b00000000000000000100011001100010;
assign LUT_1[35938] = 32'b00000000000000000110110101110111;
assign LUT_1[35939] = 32'b00000000000000000000000111110011;
assign LUT_1[35940] = 32'b00000000000000010011000000111101;
assign LUT_1[35941] = 32'b00000000000000001100010010111001;
assign LUT_1[35942] = 32'b00000000000000001110101111001110;
assign LUT_1[35943] = 32'b00000000000000001000000001001010;
assign LUT_1[35944] = 32'b00000000000000001010010101011011;
assign LUT_1[35945] = 32'b00000000000000000011100111010111;
assign LUT_1[35946] = 32'b00000000000000000110000011101100;
assign LUT_1[35947] = 32'b11111111111111111111010101101000;
assign LUT_1[35948] = 32'b00000000000000010010001110110010;
assign LUT_1[35949] = 32'b00000000000000001011100000101110;
assign LUT_1[35950] = 32'b00000000000000001101111101000011;
assign LUT_1[35951] = 32'b00000000000000000111001110111111;
assign LUT_1[35952] = 32'b00000000000000001101000011001000;
assign LUT_1[35953] = 32'b00000000000000000110010101000100;
assign LUT_1[35954] = 32'b00000000000000001000110001011001;
assign LUT_1[35955] = 32'b00000000000000000010000011010101;
assign LUT_1[35956] = 32'b00000000000000010100111100011111;
assign LUT_1[35957] = 32'b00000000000000001110001110011011;
assign LUT_1[35958] = 32'b00000000000000010000101010110000;
assign LUT_1[35959] = 32'b00000000000000001001111100101100;
assign LUT_1[35960] = 32'b00000000000000001100010000111101;
assign LUT_1[35961] = 32'b00000000000000000101100010111001;
assign LUT_1[35962] = 32'b00000000000000000111111111001110;
assign LUT_1[35963] = 32'b00000000000000000001010001001010;
assign LUT_1[35964] = 32'b00000000000000010100001010010100;
assign LUT_1[35965] = 32'b00000000000000001101011100010000;
assign LUT_1[35966] = 32'b00000000000000001111111000100101;
assign LUT_1[35967] = 32'b00000000000000001001001010100001;
assign LUT_1[35968] = 32'b00000000000000001011001111000010;
assign LUT_1[35969] = 32'b00000000000000000100100000111110;
assign LUT_1[35970] = 32'b00000000000000000110111101010011;
assign LUT_1[35971] = 32'b00000000000000000000001111001111;
assign LUT_1[35972] = 32'b00000000000000010011001000011001;
assign LUT_1[35973] = 32'b00000000000000001100011010010101;
assign LUT_1[35974] = 32'b00000000000000001110110110101010;
assign LUT_1[35975] = 32'b00000000000000001000001000100110;
assign LUT_1[35976] = 32'b00000000000000001010011100110111;
assign LUT_1[35977] = 32'b00000000000000000011101110110011;
assign LUT_1[35978] = 32'b00000000000000000110001011001000;
assign LUT_1[35979] = 32'b11111111111111111111011101000100;
assign LUT_1[35980] = 32'b00000000000000010010010110001110;
assign LUT_1[35981] = 32'b00000000000000001011101000001010;
assign LUT_1[35982] = 32'b00000000000000001110000100011111;
assign LUT_1[35983] = 32'b00000000000000000111010110011011;
assign LUT_1[35984] = 32'b00000000000000001101001010100100;
assign LUT_1[35985] = 32'b00000000000000000110011100100000;
assign LUT_1[35986] = 32'b00000000000000001000111000110101;
assign LUT_1[35987] = 32'b00000000000000000010001010110001;
assign LUT_1[35988] = 32'b00000000000000010101000011111011;
assign LUT_1[35989] = 32'b00000000000000001110010101110111;
assign LUT_1[35990] = 32'b00000000000000010000110010001100;
assign LUT_1[35991] = 32'b00000000000000001010000100001000;
assign LUT_1[35992] = 32'b00000000000000001100011000011001;
assign LUT_1[35993] = 32'b00000000000000000101101010010101;
assign LUT_1[35994] = 32'b00000000000000001000000110101010;
assign LUT_1[35995] = 32'b00000000000000000001011000100110;
assign LUT_1[35996] = 32'b00000000000000010100010001110000;
assign LUT_1[35997] = 32'b00000000000000001101100011101100;
assign LUT_1[35998] = 32'b00000000000000010000000000000001;
assign LUT_1[35999] = 32'b00000000000000001001010001111101;
assign LUT_1[36000] = 32'b00000000000000001100001010000001;
assign LUT_1[36001] = 32'b00000000000000000101011011111101;
assign LUT_1[36002] = 32'b00000000000000000111111000010010;
assign LUT_1[36003] = 32'b00000000000000000001001010001110;
assign LUT_1[36004] = 32'b00000000000000010100000011011000;
assign LUT_1[36005] = 32'b00000000000000001101010101010100;
assign LUT_1[36006] = 32'b00000000000000001111110001101001;
assign LUT_1[36007] = 32'b00000000000000001001000011100101;
assign LUT_1[36008] = 32'b00000000000000001011010111110110;
assign LUT_1[36009] = 32'b00000000000000000100101001110010;
assign LUT_1[36010] = 32'b00000000000000000111000110000111;
assign LUT_1[36011] = 32'b00000000000000000000011000000011;
assign LUT_1[36012] = 32'b00000000000000010011010001001101;
assign LUT_1[36013] = 32'b00000000000000001100100011001001;
assign LUT_1[36014] = 32'b00000000000000001110111111011110;
assign LUT_1[36015] = 32'b00000000000000001000010001011010;
assign LUT_1[36016] = 32'b00000000000000001110000101100011;
assign LUT_1[36017] = 32'b00000000000000000111010111011111;
assign LUT_1[36018] = 32'b00000000000000001001110011110100;
assign LUT_1[36019] = 32'b00000000000000000011000101110000;
assign LUT_1[36020] = 32'b00000000000000010101111110111010;
assign LUT_1[36021] = 32'b00000000000000001111010000110110;
assign LUT_1[36022] = 32'b00000000000000010001101101001011;
assign LUT_1[36023] = 32'b00000000000000001010111111000111;
assign LUT_1[36024] = 32'b00000000000000001101010011011000;
assign LUT_1[36025] = 32'b00000000000000000110100101010100;
assign LUT_1[36026] = 32'b00000000000000001001000001101001;
assign LUT_1[36027] = 32'b00000000000000000010010011100101;
assign LUT_1[36028] = 32'b00000000000000010101001100101111;
assign LUT_1[36029] = 32'b00000000000000001110011110101011;
assign LUT_1[36030] = 32'b00000000000000010000111011000000;
assign LUT_1[36031] = 32'b00000000000000001010001100111100;
assign LUT_1[36032] = 32'b00000000000000001101001100101010;
assign LUT_1[36033] = 32'b00000000000000000110011110100110;
assign LUT_1[36034] = 32'b00000000000000001000111010111011;
assign LUT_1[36035] = 32'b00000000000000000010001100110111;
assign LUT_1[36036] = 32'b00000000000000010101000110000001;
assign LUT_1[36037] = 32'b00000000000000001110010111111101;
assign LUT_1[36038] = 32'b00000000000000010000110100010010;
assign LUT_1[36039] = 32'b00000000000000001010000110001110;
assign LUT_1[36040] = 32'b00000000000000001100011010011111;
assign LUT_1[36041] = 32'b00000000000000000101101100011011;
assign LUT_1[36042] = 32'b00000000000000001000001000110000;
assign LUT_1[36043] = 32'b00000000000000000001011010101100;
assign LUT_1[36044] = 32'b00000000000000010100010011110110;
assign LUT_1[36045] = 32'b00000000000000001101100101110010;
assign LUT_1[36046] = 32'b00000000000000010000000010000111;
assign LUT_1[36047] = 32'b00000000000000001001010100000011;
assign LUT_1[36048] = 32'b00000000000000001111001000001100;
assign LUT_1[36049] = 32'b00000000000000001000011010001000;
assign LUT_1[36050] = 32'b00000000000000001010110110011101;
assign LUT_1[36051] = 32'b00000000000000000100001000011001;
assign LUT_1[36052] = 32'b00000000000000010111000001100011;
assign LUT_1[36053] = 32'b00000000000000010000010011011111;
assign LUT_1[36054] = 32'b00000000000000010010101111110100;
assign LUT_1[36055] = 32'b00000000000000001100000001110000;
assign LUT_1[36056] = 32'b00000000000000001110010110000001;
assign LUT_1[36057] = 32'b00000000000000000111100111111101;
assign LUT_1[36058] = 32'b00000000000000001010000100010010;
assign LUT_1[36059] = 32'b00000000000000000011010110001110;
assign LUT_1[36060] = 32'b00000000000000010110001111011000;
assign LUT_1[36061] = 32'b00000000000000001111100001010100;
assign LUT_1[36062] = 32'b00000000000000010001111101101001;
assign LUT_1[36063] = 32'b00000000000000001011001111100101;
assign LUT_1[36064] = 32'b00000000000000001110000111101001;
assign LUT_1[36065] = 32'b00000000000000000111011001100101;
assign LUT_1[36066] = 32'b00000000000000001001110101111010;
assign LUT_1[36067] = 32'b00000000000000000011000111110110;
assign LUT_1[36068] = 32'b00000000000000010110000001000000;
assign LUT_1[36069] = 32'b00000000000000001111010010111100;
assign LUT_1[36070] = 32'b00000000000000010001101111010001;
assign LUT_1[36071] = 32'b00000000000000001011000001001101;
assign LUT_1[36072] = 32'b00000000000000001101010101011110;
assign LUT_1[36073] = 32'b00000000000000000110100111011010;
assign LUT_1[36074] = 32'b00000000000000001001000011101111;
assign LUT_1[36075] = 32'b00000000000000000010010101101011;
assign LUT_1[36076] = 32'b00000000000000010101001110110101;
assign LUT_1[36077] = 32'b00000000000000001110100000110001;
assign LUT_1[36078] = 32'b00000000000000010000111101000110;
assign LUT_1[36079] = 32'b00000000000000001010001111000010;
assign LUT_1[36080] = 32'b00000000000000010000000011001011;
assign LUT_1[36081] = 32'b00000000000000001001010101000111;
assign LUT_1[36082] = 32'b00000000000000001011110001011100;
assign LUT_1[36083] = 32'b00000000000000000101000011011000;
assign LUT_1[36084] = 32'b00000000000000010111111100100010;
assign LUT_1[36085] = 32'b00000000000000010001001110011110;
assign LUT_1[36086] = 32'b00000000000000010011101010110011;
assign LUT_1[36087] = 32'b00000000000000001100111100101111;
assign LUT_1[36088] = 32'b00000000000000001111010001000000;
assign LUT_1[36089] = 32'b00000000000000001000100010111100;
assign LUT_1[36090] = 32'b00000000000000001010111111010001;
assign LUT_1[36091] = 32'b00000000000000000100010001001101;
assign LUT_1[36092] = 32'b00000000000000010111001010010111;
assign LUT_1[36093] = 32'b00000000000000010000011100010011;
assign LUT_1[36094] = 32'b00000000000000010010111000101000;
assign LUT_1[36095] = 32'b00000000000000001100001010100100;
assign LUT_1[36096] = 32'b00000000000000000110000011001011;
assign LUT_1[36097] = 32'b11111111111111111111010101000111;
assign LUT_1[36098] = 32'b00000000000000000001110001011100;
assign LUT_1[36099] = 32'b11111111111111111011000011011000;
assign LUT_1[36100] = 32'b00000000000000001101111100100010;
assign LUT_1[36101] = 32'b00000000000000000111001110011110;
assign LUT_1[36102] = 32'b00000000000000001001101010110011;
assign LUT_1[36103] = 32'b00000000000000000010111100101111;
assign LUT_1[36104] = 32'b00000000000000000101010001000000;
assign LUT_1[36105] = 32'b11111111111111111110100010111100;
assign LUT_1[36106] = 32'b00000000000000000000111111010001;
assign LUT_1[36107] = 32'b11111111111111111010010001001101;
assign LUT_1[36108] = 32'b00000000000000001101001010010111;
assign LUT_1[36109] = 32'b00000000000000000110011100010011;
assign LUT_1[36110] = 32'b00000000000000001000111000101000;
assign LUT_1[36111] = 32'b00000000000000000010001010100100;
assign LUT_1[36112] = 32'b00000000000000000111111110101101;
assign LUT_1[36113] = 32'b00000000000000000001010000101001;
assign LUT_1[36114] = 32'b00000000000000000011101100111110;
assign LUT_1[36115] = 32'b11111111111111111100111110111010;
assign LUT_1[36116] = 32'b00000000000000001111111000000100;
assign LUT_1[36117] = 32'b00000000000000001001001010000000;
assign LUT_1[36118] = 32'b00000000000000001011100110010101;
assign LUT_1[36119] = 32'b00000000000000000100111000010001;
assign LUT_1[36120] = 32'b00000000000000000111001100100010;
assign LUT_1[36121] = 32'b00000000000000000000011110011110;
assign LUT_1[36122] = 32'b00000000000000000010111010110011;
assign LUT_1[36123] = 32'b11111111111111111100001100101111;
assign LUT_1[36124] = 32'b00000000000000001111000101111001;
assign LUT_1[36125] = 32'b00000000000000001000010111110101;
assign LUT_1[36126] = 32'b00000000000000001010110100001010;
assign LUT_1[36127] = 32'b00000000000000000100000110000110;
assign LUT_1[36128] = 32'b00000000000000000110111110001010;
assign LUT_1[36129] = 32'b00000000000000000000010000000110;
assign LUT_1[36130] = 32'b00000000000000000010101100011011;
assign LUT_1[36131] = 32'b11111111111111111011111110010111;
assign LUT_1[36132] = 32'b00000000000000001110110111100001;
assign LUT_1[36133] = 32'b00000000000000001000001001011101;
assign LUT_1[36134] = 32'b00000000000000001010100101110010;
assign LUT_1[36135] = 32'b00000000000000000011110111101110;
assign LUT_1[36136] = 32'b00000000000000000110001011111111;
assign LUT_1[36137] = 32'b11111111111111111111011101111011;
assign LUT_1[36138] = 32'b00000000000000000001111010010000;
assign LUT_1[36139] = 32'b11111111111111111011001100001100;
assign LUT_1[36140] = 32'b00000000000000001110000101010110;
assign LUT_1[36141] = 32'b00000000000000000111010111010010;
assign LUT_1[36142] = 32'b00000000000000001001110011100111;
assign LUT_1[36143] = 32'b00000000000000000011000101100011;
assign LUT_1[36144] = 32'b00000000000000001000111001101100;
assign LUT_1[36145] = 32'b00000000000000000010001011101000;
assign LUT_1[36146] = 32'b00000000000000000100100111111101;
assign LUT_1[36147] = 32'b11111111111111111101111001111001;
assign LUT_1[36148] = 32'b00000000000000010000110011000011;
assign LUT_1[36149] = 32'b00000000000000001010000100111111;
assign LUT_1[36150] = 32'b00000000000000001100100001010100;
assign LUT_1[36151] = 32'b00000000000000000101110011010000;
assign LUT_1[36152] = 32'b00000000000000001000000111100001;
assign LUT_1[36153] = 32'b00000000000000000001011001011101;
assign LUT_1[36154] = 32'b00000000000000000011110101110010;
assign LUT_1[36155] = 32'b11111111111111111101000111101110;
assign LUT_1[36156] = 32'b00000000000000010000000000111000;
assign LUT_1[36157] = 32'b00000000000000001001010010110100;
assign LUT_1[36158] = 32'b00000000000000001011101111001001;
assign LUT_1[36159] = 32'b00000000000000000101000001000101;
assign LUT_1[36160] = 32'b00000000000000001000000000110011;
assign LUT_1[36161] = 32'b00000000000000000001010010101111;
assign LUT_1[36162] = 32'b00000000000000000011101111000100;
assign LUT_1[36163] = 32'b11111111111111111101000001000000;
assign LUT_1[36164] = 32'b00000000000000001111111010001010;
assign LUT_1[36165] = 32'b00000000000000001001001100000110;
assign LUT_1[36166] = 32'b00000000000000001011101000011011;
assign LUT_1[36167] = 32'b00000000000000000100111010010111;
assign LUT_1[36168] = 32'b00000000000000000111001110101000;
assign LUT_1[36169] = 32'b00000000000000000000100000100100;
assign LUT_1[36170] = 32'b00000000000000000010111100111001;
assign LUT_1[36171] = 32'b11111111111111111100001110110101;
assign LUT_1[36172] = 32'b00000000000000001111000111111111;
assign LUT_1[36173] = 32'b00000000000000001000011001111011;
assign LUT_1[36174] = 32'b00000000000000001010110110010000;
assign LUT_1[36175] = 32'b00000000000000000100001000001100;
assign LUT_1[36176] = 32'b00000000000000001001111100010101;
assign LUT_1[36177] = 32'b00000000000000000011001110010001;
assign LUT_1[36178] = 32'b00000000000000000101101010100110;
assign LUT_1[36179] = 32'b11111111111111111110111100100010;
assign LUT_1[36180] = 32'b00000000000000010001110101101100;
assign LUT_1[36181] = 32'b00000000000000001011000111101000;
assign LUT_1[36182] = 32'b00000000000000001101100011111101;
assign LUT_1[36183] = 32'b00000000000000000110110101111001;
assign LUT_1[36184] = 32'b00000000000000001001001010001010;
assign LUT_1[36185] = 32'b00000000000000000010011100000110;
assign LUT_1[36186] = 32'b00000000000000000100111000011011;
assign LUT_1[36187] = 32'b11111111111111111110001010010111;
assign LUT_1[36188] = 32'b00000000000000010001000011100001;
assign LUT_1[36189] = 32'b00000000000000001010010101011101;
assign LUT_1[36190] = 32'b00000000000000001100110001110010;
assign LUT_1[36191] = 32'b00000000000000000110000011101110;
assign LUT_1[36192] = 32'b00000000000000001000111011110010;
assign LUT_1[36193] = 32'b00000000000000000010001101101110;
assign LUT_1[36194] = 32'b00000000000000000100101010000011;
assign LUT_1[36195] = 32'b11111111111111111101111011111111;
assign LUT_1[36196] = 32'b00000000000000010000110101001001;
assign LUT_1[36197] = 32'b00000000000000001010000111000101;
assign LUT_1[36198] = 32'b00000000000000001100100011011010;
assign LUT_1[36199] = 32'b00000000000000000101110101010110;
assign LUT_1[36200] = 32'b00000000000000001000001001100111;
assign LUT_1[36201] = 32'b00000000000000000001011011100011;
assign LUT_1[36202] = 32'b00000000000000000011110111111000;
assign LUT_1[36203] = 32'b11111111111111111101001001110100;
assign LUT_1[36204] = 32'b00000000000000010000000010111110;
assign LUT_1[36205] = 32'b00000000000000001001010100111010;
assign LUT_1[36206] = 32'b00000000000000001011110001001111;
assign LUT_1[36207] = 32'b00000000000000000101000011001011;
assign LUT_1[36208] = 32'b00000000000000001010110111010100;
assign LUT_1[36209] = 32'b00000000000000000100001001010000;
assign LUT_1[36210] = 32'b00000000000000000110100101100101;
assign LUT_1[36211] = 32'b11111111111111111111110111100001;
assign LUT_1[36212] = 32'b00000000000000010010110000101011;
assign LUT_1[36213] = 32'b00000000000000001100000010100111;
assign LUT_1[36214] = 32'b00000000000000001110011110111100;
assign LUT_1[36215] = 32'b00000000000000000111110000111000;
assign LUT_1[36216] = 32'b00000000000000001010000101001001;
assign LUT_1[36217] = 32'b00000000000000000011010111000101;
assign LUT_1[36218] = 32'b00000000000000000101110011011010;
assign LUT_1[36219] = 32'b11111111111111111111000101010110;
assign LUT_1[36220] = 32'b00000000000000010001111110100000;
assign LUT_1[36221] = 32'b00000000000000001011010000011100;
assign LUT_1[36222] = 32'b00000000000000001101101100110001;
assign LUT_1[36223] = 32'b00000000000000000110111110101101;
assign LUT_1[36224] = 32'b00000000000000001001000011001110;
assign LUT_1[36225] = 32'b00000000000000000010010101001010;
assign LUT_1[36226] = 32'b00000000000000000100110001011111;
assign LUT_1[36227] = 32'b11111111111111111110000011011011;
assign LUT_1[36228] = 32'b00000000000000010000111100100101;
assign LUT_1[36229] = 32'b00000000000000001010001110100001;
assign LUT_1[36230] = 32'b00000000000000001100101010110110;
assign LUT_1[36231] = 32'b00000000000000000101111100110010;
assign LUT_1[36232] = 32'b00000000000000001000010001000011;
assign LUT_1[36233] = 32'b00000000000000000001100010111111;
assign LUT_1[36234] = 32'b00000000000000000011111111010100;
assign LUT_1[36235] = 32'b11111111111111111101010001010000;
assign LUT_1[36236] = 32'b00000000000000010000001010011010;
assign LUT_1[36237] = 32'b00000000000000001001011100010110;
assign LUT_1[36238] = 32'b00000000000000001011111000101011;
assign LUT_1[36239] = 32'b00000000000000000101001010100111;
assign LUT_1[36240] = 32'b00000000000000001010111110110000;
assign LUT_1[36241] = 32'b00000000000000000100010000101100;
assign LUT_1[36242] = 32'b00000000000000000110101101000001;
assign LUT_1[36243] = 32'b11111111111111111111111110111101;
assign LUT_1[36244] = 32'b00000000000000010010111000000111;
assign LUT_1[36245] = 32'b00000000000000001100001010000011;
assign LUT_1[36246] = 32'b00000000000000001110100110011000;
assign LUT_1[36247] = 32'b00000000000000000111111000010100;
assign LUT_1[36248] = 32'b00000000000000001010001100100101;
assign LUT_1[36249] = 32'b00000000000000000011011110100001;
assign LUT_1[36250] = 32'b00000000000000000101111010110110;
assign LUT_1[36251] = 32'b11111111111111111111001100110010;
assign LUT_1[36252] = 32'b00000000000000010010000101111100;
assign LUT_1[36253] = 32'b00000000000000001011010111111000;
assign LUT_1[36254] = 32'b00000000000000001101110100001101;
assign LUT_1[36255] = 32'b00000000000000000111000110001001;
assign LUT_1[36256] = 32'b00000000000000001001111110001101;
assign LUT_1[36257] = 32'b00000000000000000011010000001001;
assign LUT_1[36258] = 32'b00000000000000000101101100011110;
assign LUT_1[36259] = 32'b11111111111111111110111110011010;
assign LUT_1[36260] = 32'b00000000000000010001110111100100;
assign LUT_1[36261] = 32'b00000000000000001011001001100000;
assign LUT_1[36262] = 32'b00000000000000001101100101110101;
assign LUT_1[36263] = 32'b00000000000000000110110111110001;
assign LUT_1[36264] = 32'b00000000000000001001001100000010;
assign LUT_1[36265] = 32'b00000000000000000010011101111110;
assign LUT_1[36266] = 32'b00000000000000000100111010010011;
assign LUT_1[36267] = 32'b11111111111111111110001100001111;
assign LUT_1[36268] = 32'b00000000000000010001000101011001;
assign LUT_1[36269] = 32'b00000000000000001010010111010101;
assign LUT_1[36270] = 32'b00000000000000001100110011101010;
assign LUT_1[36271] = 32'b00000000000000000110000101100110;
assign LUT_1[36272] = 32'b00000000000000001011111001101111;
assign LUT_1[36273] = 32'b00000000000000000101001011101011;
assign LUT_1[36274] = 32'b00000000000000000111101000000000;
assign LUT_1[36275] = 32'b00000000000000000000111001111100;
assign LUT_1[36276] = 32'b00000000000000010011110011000110;
assign LUT_1[36277] = 32'b00000000000000001101000101000010;
assign LUT_1[36278] = 32'b00000000000000001111100001010111;
assign LUT_1[36279] = 32'b00000000000000001000110011010011;
assign LUT_1[36280] = 32'b00000000000000001011000111100100;
assign LUT_1[36281] = 32'b00000000000000000100011001100000;
assign LUT_1[36282] = 32'b00000000000000000110110101110101;
assign LUT_1[36283] = 32'b00000000000000000000000111110001;
assign LUT_1[36284] = 32'b00000000000000010011000000111011;
assign LUT_1[36285] = 32'b00000000000000001100010010110111;
assign LUT_1[36286] = 32'b00000000000000001110101111001100;
assign LUT_1[36287] = 32'b00000000000000001000000001001000;
assign LUT_1[36288] = 32'b00000000000000001011000000110110;
assign LUT_1[36289] = 32'b00000000000000000100010010110010;
assign LUT_1[36290] = 32'b00000000000000000110101111000111;
assign LUT_1[36291] = 32'b00000000000000000000000001000011;
assign LUT_1[36292] = 32'b00000000000000010010111010001101;
assign LUT_1[36293] = 32'b00000000000000001100001100001001;
assign LUT_1[36294] = 32'b00000000000000001110101000011110;
assign LUT_1[36295] = 32'b00000000000000000111111010011010;
assign LUT_1[36296] = 32'b00000000000000001010001110101011;
assign LUT_1[36297] = 32'b00000000000000000011100000100111;
assign LUT_1[36298] = 32'b00000000000000000101111100111100;
assign LUT_1[36299] = 32'b11111111111111111111001110111000;
assign LUT_1[36300] = 32'b00000000000000010010001000000010;
assign LUT_1[36301] = 32'b00000000000000001011011001111110;
assign LUT_1[36302] = 32'b00000000000000001101110110010011;
assign LUT_1[36303] = 32'b00000000000000000111001000001111;
assign LUT_1[36304] = 32'b00000000000000001100111100011000;
assign LUT_1[36305] = 32'b00000000000000000110001110010100;
assign LUT_1[36306] = 32'b00000000000000001000101010101001;
assign LUT_1[36307] = 32'b00000000000000000001111100100101;
assign LUT_1[36308] = 32'b00000000000000010100110101101111;
assign LUT_1[36309] = 32'b00000000000000001110000111101011;
assign LUT_1[36310] = 32'b00000000000000010000100100000000;
assign LUT_1[36311] = 32'b00000000000000001001110101111100;
assign LUT_1[36312] = 32'b00000000000000001100001010001101;
assign LUT_1[36313] = 32'b00000000000000000101011100001001;
assign LUT_1[36314] = 32'b00000000000000000111111000011110;
assign LUT_1[36315] = 32'b00000000000000000001001010011010;
assign LUT_1[36316] = 32'b00000000000000010100000011100100;
assign LUT_1[36317] = 32'b00000000000000001101010101100000;
assign LUT_1[36318] = 32'b00000000000000001111110001110101;
assign LUT_1[36319] = 32'b00000000000000001001000011110001;
assign LUT_1[36320] = 32'b00000000000000001011111011110101;
assign LUT_1[36321] = 32'b00000000000000000101001101110001;
assign LUT_1[36322] = 32'b00000000000000000111101010000110;
assign LUT_1[36323] = 32'b00000000000000000000111100000010;
assign LUT_1[36324] = 32'b00000000000000010011110101001100;
assign LUT_1[36325] = 32'b00000000000000001101000111001000;
assign LUT_1[36326] = 32'b00000000000000001111100011011101;
assign LUT_1[36327] = 32'b00000000000000001000110101011001;
assign LUT_1[36328] = 32'b00000000000000001011001001101010;
assign LUT_1[36329] = 32'b00000000000000000100011011100110;
assign LUT_1[36330] = 32'b00000000000000000110110111111011;
assign LUT_1[36331] = 32'b00000000000000000000001001110111;
assign LUT_1[36332] = 32'b00000000000000010011000011000001;
assign LUT_1[36333] = 32'b00000000000000001100010100111101;
assign LUT_1[36334] = 32'b00000000000000001110110001010010;
assign LUT_1[36335] = 32'b00000000000000001000000011001110;
assign LUT_1[36336] = 32'b00000000000000001101110111010111;
assign LUT_1[36337] = 32'b00000000000000000111001001010011;
assign LUT_1[36338] = 32'b00000000000000001001100101101000;
assign LUT_1[36339] = 32'b00000000000000000010110111100100;
assign LUT_1[36340] = 32'b00000000000000010101110000101110;
assign LUT_1[36341] = 32'b00000000000000001111000010101010;
assign LUT_1[36342] = 32'b00000000000000010001011110111111;
assign LUT_1[36343] = 32'b00000000000000001010110000111011;
assign LUT_1[36344] = 32'b00000000000000001101000101001100;
assign LUT_1[36345] = 32'b00000000000000000110010111001000;
assign LUT_1[36346] = 32'b00000000000000001000110011011101;
assign LUT_1[36347] = 32'b00000000000000000010000101011001;
assign LUT_1[36348] = 32'b00000000000000010100111110100011;
assign LUT_1[36349] = 32'b00000000000000001110010000011111;
assign LUT_1[36350] = 32'b00000000000000010000101100110100;
assign LUT_1[36351] = 32'b00000000000000001001111110110000;
assign LUT_1[36352] = 32'b00000000000000000001111101011100;
assign LUT_1[36353] = 32'b11111111111111111011001111011000;
assign LUT_1[36354] = 32'b11111111111111111101101011101101;
assign LUT_1[36355] = 32'b11111111111111110110111101101001;
assign LUT_1[36356] = 32'b00000000000000001001110110110011;
assign LUT_1[36357] = 32'b00000000000000000011001000101111;
assign LUT_1[36358] = 32'b00000000000000000101100101000100;
assign LUT_1[36359] = 32'b11111111111111111110110111000000;
assign LUT_1[36360] = 32'b00000000000000000001001011010001;
assign LUT_1[36361] = 32'b11111111111111111010011101001101;
assign LUT_1[36362] = 32'b11111111111111111100111001100010;
assign LUT_1[36363] = 32'b11111111111111110110001011011110;
assign LUT_1[36364] = 32'b00000000000000001001000100101000;
assign LUT_1[36365] = 32'b00000000000000000010010110100100;
assign LUT_1[36366] = 32'b00000000000000000100110010111001;
assign LUT_1[36367] = 32'b11111111111111111110000100110101;
assign LUT_1[36368] = 32'b00000000000000000011111000111110;
assign LUT_1[36369] = 32'b11111111111111111101001010111010;
assign LUT_1[36370] = 32'b11111111111111111111100111001111;
assign LUT_1[36371] = 32'b11111111111111111000111001001011;
assign LUT_1[36372] = 32'b00000000000000001011110010010101;
assign LUT_1[36373] = 32'b00000000000000000101000100010001;
assign LUT_1[36374] = 32'b00000000000000000111100000100110;
assign LUT_1[36375] = 32'b00000000000000000000110010100010;
assign LUT_1[36376] = 32'b00000000000000000011000110110011;
assign LUT_1[36377] = 32'b11111111111111111100011000101111;
assign LUT_1[36378] = 32'b11111111111111111110110101000100;
assign LUT_1[36379] = 32'b11111111111111111000000111000000;
assign LUT_1[36380] = 32'b00000000000000001011000000001010;
assign LUT_1[36381] = 32'b00000000000000000100010010000110;
assign LUT_1[36382] = 32'b00000000000000000110101110011011;
assign LUT_1[36383] = 32'b00000000000000000000000000010111;
assign LUT_1[36384] = 32'b00000000000000000010111000011011;
assign LUT_1[36385] = 32'b11111111111111111100001010010111;
assign LUT_1[36386] = 32'b11111111111111111110100110101100;
assign LUT_1[36387] = 32'b11111111111111110111111000101000;
assign LUT_1[36388] = 32'b00000000000000001010110001110010;
assign LUT_1[36389] = 32'b00000000000000000100000011101110;
assign LUT_1[36390] = 32'b00000000000000000110100000000011;
assign LUT_1[36391] = 32'b11111111111111111111110001111111;
assign LUT_1[36392] = 32'b00000000000000000010000110010000;
assign LUT_1[36393] = 32'b11111111111111111011011000001100;
assign LUT_1[36394] = 32'b11111111111111111101110100100001;
assign LUT_1[36395] = 32'b11111111111111110111000110011101;
assign LUT_1[36396] = 32'b00000000000000001001111111100111;
assign LUT_1[36397] = 32'b00000000000000000011010001100011;
assign LUT_1[36398] = 32'b00000000000000000101101101111000;
assign LUT_1[36399] = 32'b11111111111111111110111111110100;
assign LUT_1[36400] = 32'b00000000000000000100110011111101;
assign LUT_1[36401] = 32'b11111111111111111110000101111001;
assign LUT_1[36402] = 32'b00000000000000000000100010001110;
assign LUT_1[36403] = 32'b11111111111111111001110100001010;
assign LUT_1[36404] = 32'b00000000000000001100101101010100;
assign LUT_1[36405] = 32'b00000000000000000101111111010000;
assign LUT_1[36406] = 32'b00000000000000001000011011100101;
assign LUT_1[36407] = 32'b00000000000000000001101101100001;
assign LUT_1[36408] = 32'b00000000000000000100000001110010;
assign LUT_1[36409] = 32'b11111111111111111101010011101110;
assign LUT_1[36410] = 32'b11111111111111111111110000000011;
assign LUT_1[36411] = 32'b11111111111111111001000001111111;
assign LUT_1[36412] = 32'b00000000000000001011111011001001;
assign LUT_1[36413] = 32'b00000000000000000101001101000101;
assign LUT_1[36414] = 32'b00000000000000000111101001011010;
assign LUT_1[36415] = 32'b00000000000000000000111011010110;
assign LUT_1[36416] = 32'b00000000000000000011111011000100;
assign LUT_1[36417] = 32'b11111111111111111101001101000000;
assign LUT_1[36418] = 32'b11111111111111111111101001010101;
assign LUT_1[36419] = 32'b11111111111111111000111011010001;
assign LUT_1[36420] = 32'b00000000000000001011110100011011;
assign LUT_1[36421] = 32'b00000000000000000101000110010111;
assign LUT_1[36422] = 32'b00000000000000000111100010101100;
assign LUT_1[36423] = 32'b00000000000000000000110100101000;
assign LUT_1[36424] = 32'b00000000000000000011001000111001;
assign LUT_1[36425] = 32'b11111111111111111100011010110101;
assign LUT_1[36426] = 32'b11111111111111111110110111001010;
assign LUT_1[36427] = 32'b11111111111111111000001001000110;
assign LUT_1[36428] = 32'b00000000000000001011000010010000;
assign LUT_1[36429] = 32'b00000000000000000100010100001100;
assign LUT_1[36430] = 32'b00000000000000000110110000100001;
assign LUT_1[36431] = 32'b00000000000000000000000010011101;
assign LUT_1[36432] = 32'b00000000000000000101110110100110;
assign LUT_1[36433] = 32'b11111111111111111111001000100010;
assign LUT_1[36434] = 32'b00000000000000000001100100110111;
assign LUT_1[36435] = 32'b11111111111111111010110110110011;
assign LUT_1[36436] = 32'b00000000000000001101101111111101;
assign LUT_1[36437] = 32'b00000000000000000111000001111001;
assign LUT_1[36438] = 32'b00000000000000001001011110001110;
assign LUT_1[36439] = 32'b00000000000000000010110000001010;
assign LUT_1[36440] = 32'b00000000000000000101000100011011;
assign LUT_1[36441] = 32'b11111111111111111110010110010111;
assign LUT_1[36442] = 32'b00000000000000000000110010101100;
assign LUT_1[36443] = 32'b11111111111111111010000100101000;
assign LUT_1[36444] = 32'b00000000000000001100111101110010;
assign LUT_1[36445] = 32'b00000000000000000110001111101110;
assign LUT_1[36446] = 32'b00000000000000001000101100000011;
assign LUT_1[36447] = 32'b00000000000000000001111101111111;
assign LUT_1[36448] = 32'b00000000000000000100110110000011;
assign LUT_1[36449] = 32'b11111111111111111110000111111111;
assign LUT_1[36450] = 32'b00000000000000000000100100010100;
assign LUT_1[36451] = 32'b11111111111111111001110110010000;
assign LUT_1[36452] = 32'b00000000000000001100101111011010;
assign LUT_1[36453] = 32'b00000000000000000110000001010110;
assign LUT_1[36454] = 32'b00000000000000001000011101101011;
assign LUT_1[36455] = 32'b00000000000000000001101111100111;
assign LUT_1[36456] = 32'b00000000000000000100000011111000;
assign LUT_1[36457] = 32'b11111111111111111101010101110100;
assign LUT_1[36458] = 32'b11111111111111111111110010001001;
assign LUT_1[36459] = 32'b11111111111111111001000100000101;
assign LUT_1[36460] = 32'b00000000000000001011111101001111;
assign LUT_1[36461] = 32'b00000000000000000101001111001011;
assign LUT_1[36462] = 32'b00000000000000000111101011100000;
assign LUT_1[36463] = 32'b00000000000000000000111101011100;
assign LUT_1[36464] = 32'b00000000000000000110110001100101;
assign LUT_1[36465] = 32'b00000000000000000000000011100001;
assign LUT_1[36466] = 32'b00000000000000000010011111110110;
assign LUT_1[36467] = 32'b11111111111111111011110001110010;
assign LUT_1[36468] = 32'b00000000000000001110101010111100;
assign LUT_1[36469] = 32'b00000000000000000111111100111000;
assign LUT_1[36470] = 32'b00000000000000001010011001001101;
assign LUT_1[36471] = 32'b00000000000000000011101011001001;
assign LUT_1[36472] = 32'b00000000000000000101111111011010;
assign LUT_1[36473] = 32'b11111111111111111111010001010110;
assign LUT_1[36474] = 32'b00000000000000000001101101101011;
assign LUT_1[36475] = 32'b11111111111111111010111111100111;
assign LUT_1[36476] = 32'b00000000000000001101111000110001;
assign LUT_1[36477] = 32'b00000000000000000111001010101101;
assign LUT_1[36478] = 32'b00000000000000001001100111000010;
assign LUT_1[36479] = 32'b00000000000000000010111000111110;
assign LUT_1[36480] = 32'b00000000000000000100111101011111;
assign LUT_1[36481] = 32'b11111111111111111110001111011011;
assign LUT_1[36482] = 32'b00000000000000000000101011110000;
assign LUT_1[36483] = 32'b11111111111111111001111101101100;
assign LUT_1[36484] = 32'b00000000000000001100110110110110;
assign LUT_1[36485] = 32'b00000000000000000110001000110010;
assign LUT_1[36486] = 32'b00000000000000001000100101000111;
assign LUT_1[36487] = 32'b00000000000000000001110111000011;
assign LUT_1[36488] = 32'b00000000000000000100001011010100;
assign LUT_1[36489] = 32'b11111111111111111101011101010000;
assign LUT_1[36490] = 32'b11111111111111111111111001100101;
assign LUT_1[36491] = 32'b11111111111111111001001011100001;
assign LUT_1[36492] = 32'b00000000000000001100000100101011;
assign LUT_1[36493] = 32'b00000000000000000101010110100111;
assign LUT_1[36494] = 32'b00000000000000000111110010111100;
assign LUT_1[36495] = 32'b00000000000000000001000100111000;
assign LUT_1[36496] = 32'b00000000000000000110111001000001;
assign LUT_1[36497] = 32'b00000000000000000000001010111101;
assign LUT_1[36498] = 32'b00000000000000000010100111010010;
assign LUT_1[36499] = 32'b11111111111111111011111001001110;
assign LUT_1[36500] = 32'b00000000000000001110110010011000;
assign LUT_1[36501] = 32'b00000000000000001000000100010100;
assign LUT_1[36502] = 32'b00000000000000001010100000101001;
assign LUT_1[36503] = 32'b00000000000000000011110010100101;
assign LUT_1[36504] = 32'b00000000000000000110000110110110;
assign LUT_1[36505] = 32'b11111111111111111111011000110010;
assign LUT_1[36506] = 32'b00000000000000000001110101000111;
assign LUT_1[36507] = 32'b11111111111111111011000111000011;
assign LUT_1[36508] = 32'b00000000000000001110000000001101;
assign LUT_1[36509] = 32'b00000000000000000111010010001001;
assign LUT_1[36510] = 32'b00000000000000001001101110011110;
assign LUT_1[36511] = 32'b00000000000000000011000000011010;
assign LUT_1[36512] = 32'b00000000000000000101111000011110;
assign LUT_1[36513] = 32'b11111111111111111111001010011010;
assign LUT_1[36514] = 32'b00000000000000000001100110101111;
assign LUT_1[36515] = 32'b11111111111111111010111000101011;
assign LUT_1[36516] = 32'b00000000000000001101110001110101;
assign LUT_1[36517] = 32'b00000000000000000111000011110001;
assign LUT_1[36518] = 32'b00000000000000001001100000000110;
assign LUT_1[36519] = 32'b00000000000000000010110010000010;
assign LUT_1[36520] = 32'b00000000000000000101000110010011;
assign LUT_1[36521] = 32'b11111111111111111110011000001111;
assign LUT_1[36522] = 32'b00000000000000000000110100100100;
assign LUT_1[36523] = 32'b11111111111111111010000110100000;
assign LUT_1[36524] = 32'b00000000000000001100111111101010;
assign LUT_1[36525] = 32'b00000000000000000110010001100110;
assign LUT_1[36526] = 32'b00000000000000001000101101111011;
assign LUT_1[36527] = 32'b00000000000000000001111111110111;
assign LUT_1[36528] = 32'b00000000000000000111110100000000;
assign LUT_1[36529] = 32'b00000000000000000001000101111100;
assign LUT_1[36530] = 32'b00000000000000000011100010010001;
assign LUT_1[36531] = 32'b11111111111111111100110100001101;
assign LUT_1[36532] = 32'b00000000000000001111101101010111;
assign LUT_1[36533] = 32'b00000000000000001000111111010011;
assign LUT_1[36534] = 32'b00000000000000001011011011101000;
assign LUT_1[36535] = 32'b00000000000000000100101101100100;
assign LUT_1[36536] = 32'b00000000000000000111000001110101;
assign LUT_1[36537] = 32'b00000000000000000000010011110001;
assign LUT_1[36538] = 32'b00000000000000000010110000000110;
assign LUT_1[36539] = 32'b11111111111111111100000010000010;
assign LUT_1[36540] = 32'b00000000000000001110111011001100;
assign LUT_1[36541] = 32'b00000000000000001000001101001000;
assign LUT_1[36542] = 32'b00000000000000001010101001011101;
assign LUT_1[36543] = 32'b00000000000000000011111011011001;
assign LUT_1[36544] = 32'b00000000000000000110111011000111;
assign LUT_1[36545] = 32'b00000000000000000000001101000011;
assign LUT_1[36546] = 32'b00000000000000000010101001011000;
assign LUT_1[36547] = 32'b11111111111111111011111011010100;
assign LUT_1[36548] = 32'b00000000000000001110110100011110;
assign LUT_1[36549] = 32'b00000000000000001000000110011010;
assign LUT_1[36550] = 32'b00000000000000001010100010101111;
assign LUT_1[36551] = 32'b00000000000000000011110100101011;
assign LUT_1[36552] = 32'b00000000000000000110001000111100;
assign LUT_1[36553] = 32'b11111111111111111111011010111000;
assign LUT_1[36554] = 32'b00000000000000000001110111001101;
assign LUT_1[36555] = 32'b11111111111111111011001001001001;
assign LUT_1[36556] = 32'b00000000000000001110000010010011;
assign LUT_1[36557] = 32'b00000000000000000111010100001111;
assign LUT_1[36558] = 32'b00000000000000001001110000100100;
assign LUT_1[36559] = 32'b00000000000000000011000010100000;
assign LUT_1[36560] = 32'b00000000000000001000110110101001;
assign LUT_1[36561] = 32'b00000000000000000010001000100101;
assign LUT_1[36562] = 32'b00000000000000000100100100111010;
assign LUT_1[36563] = 32'b11111111111111111101110110110110;
assign LUT_1[36564] = 32'b00000000000000010000110000000000;
assign LUT_1[36565] = 32'b00000000000000001010000001111100;
assign LUT_1[36566] = 32'b00000000000000001100011110010001;
assign LUT_1[36567] = 32'b00000000000000000101110000001101;
assign LUT_1[36568] = 32'b00000000000000001000000100011110;
assign LUT_1[36569] = 32'b00000000000000000001010110011010;
assign LUT_1[36570] = 32'b00000000000000000011110010101111;
assign LUT_1[36571] = 32'b11111111111111111101000100101011;
assign LUT_1[36572] = 32'b00000000000000001111111101110101;
assign LUT_1[36573] = 32'b00000000000000001001001111110001;
assign LUT_1[36574] = 32'b00000000000000001011101100000110;
assign LUT_1[36575] = 32'b00000000000000000100111110000010;
assign LUT_1[36576] = 32'b00000000000000000111110110000110;
assign LUT_1[36577] = 32'b00000000000000000001001000000010;
assign LUT_1[36578] = 32'b00000000000000000011100100010111;
assign LUT_1[36579] = 32'b11111111111111111100110110010011;
assign LUT_1[36580] = 32'b00000000000000001111101111011101;
assign LUT_1[36581] = 32'b00000000000000001001000001011001;
assign LUT_1[36582] = 32'b00000000000000001011011101101110;
assign LUT_1[36583] = 32'b00000000000000000100101111101010;
assign LUT_1[36584] = 32'b00000000000000000111000011111011;
assign LUT_1[36585] = 32'b00000000000000000000010101110111;
assign LUT_1[36586] = 32'b00000000000000000010110010001100;
assign LUT_1[36587] = 32'b11111111111111111100000100001000;
assign LUT_1[36588] = 32'b00000000000000001110111101010010;
assign LUT_1[36589] = 32'b00000000000000001000001111001110;
assign LUT_1[36590] = 32'b00000000000000001010101011100011;
assign LUT_1[36591] = 32'b00000000000000000011111101011111;
assign LUT_1[36592] = 32'b00000000000000001001110001101000;
assign LUT_1[36593] = 32'b00000000000000000011000011100100;
assign LUT_1[36594] = 32'b00000000000000000101011111111001;
assign LUT_1[36595] = 32'b11111111111111111110110001110101;
assign LUT_1[36596] = 32'b00000000000000010001101010111111;
assign LUT_1[36597] = 32'b00000000000000001010111100111011;
assign LUT_1[36598] = 32'b00000000000000001101011001010000;
assign LUT_1[36599] = 32'b00000000000000000110101011001100;
assign LUT_1[36600] = 32'b00000000000000001000111111011101;
assign LUT_1[36601] = 32'b00000000000000000010010001011001;
assign LUT_1[36602] = 32'b00000000000000000100101101101110;
assign LUT_1[36603] = 32'b11111111111111111101111111101010;
assign LUT_1[36604] = 32'b00000000000000010000111000110100;
assign LUT_1[36605] = 32'b00000000000000001010001010110000;
assign LUT_1[36606] = 32'b00000000000000001100100111000101;
assign LUT_1[36607] = 32'b00000000000000000101111001000001;
assign LUT_1[36608] = 32'b11111111111111111111110001101000;
assign LUT_1[36609] = 32'b11111111111111111001000011100100;
assign LUT_1[36610] = 32'b11111111111111111011011111111001;
assign LUT_1[36611] = 32'b11111111111111110100110001110101;
assign LUT_1[36612] = 32'b00000000000000000111101010111111;
assign LUT_1[36613] = 32'b00000000000000000000111100111011;
assign LUT_1[36614] = 32'b00000000000000000011011001010000;
assign LUT_1[36615] = 32'b11111111111111111100101011001100;
assign LUT_1[36616] = 32'b11111111111111111110111111011101;
assign LUT_1[36617] = 32'b11111111111111111000010001011001;
assign LUT_1[36618] = 32'b11111111111111111010101101101110;
assign LUT_1[36619] = 32'b11111111111111110011111111101010;
assign LUT_1[36620] = 32'b00000000000000000110111000110100;
assign LUT_1[36621] = 32'b00000000000000000000001010110000;
assign LUT_1[36622] = 32'b00000000000000000010100111000101;
assign LUT_1[36623] = 32'b11111111111111111011111001000001;
assign LUT_1[36624] = 32'b00000000000000000001101101001010;
assign LUT_1[36625] = 32'b11111111111111111010111111000110;
assign LUT_1[36626] = 32'b11111111111111111101011011011011;
assign LUT_1[36627] = 32'b11111111111111110110101101010111;
assign LUT_1[36628] = 32'b00000000000000001001100110100001;
assign LUT_1[36629] = 32'b00000000000000000010111000011101;
assign LUT_1[36630] = 32'b00000000000000000101010100110010;
assign LUT_1[36631] = 32'b11111111111111111110100110101110;
assign LUT_1[36632] = 32'b00000000000000000000111010111111;
assign LUT_1[36633] = 32'b11111111111111111010001100111011;
assign LUT_1[36634] = 32'b11111111111111111100101001010000;
assign LUT_1[36635] = 32'b11111111111111110101111011001100;
assign LUT_1[36636] = 32'b00000000000000001000110100010110;
assign LUT_1[36637] = 32'b00000000000000000010000110010010;
assign LUT_1[36638] = 32'b00000000000000000100100010100111;
assign LUT_1[36639] = 32'b11111111111111111101110100100011;
assign LUT_1[36640] = 32'b00000000000000000000101100100111;
assign LUT_1[36641] = 32'b11111111111111111001111110100011;
assign LUT_1[36642] = 32'b11111111111111111100011010111000;
assign LUT_1[36643] = 32'b11111111111111110101101100110100;
assign LUT_1[36644] = 32'b00000000000000001000100101111110;
assign LUT_1[36645] = 32'b00000000000000000001110111111010;
assign LUT_1[36646] = 32'b00000000000000000100010100001111;
assign LUT_1[36647] = 32'b11111111111111111101100110001011;
assign LUT_1[36648] = 32'b11111111111111111111111010011100;
assign LUT_1[36649] = 32'b11111111111111111001001100011000;
assign LUT_1[36650] = 32'b11111111111111111011101000101101;
assign LUT_1[36651] = 32'b11111111111111110100111010101001;
assign LUT_1[36652] = 32'b00000000000000000111110011110011;
assign LUT_1[36653] = 32'b00000000000000000001000101101111;
assign LUT_1[36654] = 32'b00000000000000000011100010000100;
assign LUT_1[36655] = 32'b11111111111111111100110100000000;
assign LUT_1[36656] = 32'b00000000000000000010101000001001;
assign LUT_1[36657] = 32'b11111111111111111011111010000101;
assign LUT_1[36658] = 32'b11111111111111111110010110011010;
assign LUT_1[36659] = 32'b11111111111111110111101000010110;
assign LUT_1[36660] = 32'b00000000000000001010100001100000;
assign LUT_1[36661] = 32'b00000000000000000011110011011100;
assign LUT_1[36662] = 32'b00000000000000000110001111110001;
assign LUT_1[36663] = 32'b11111111111111111111100001101101;
assign LUT_1[36664] = 32'b00000000000000000001110101111110;
assign LUT_1[36665] = 32'b11111111111111111011000111111010;
assign LUT_1[36666] = 32'b11111111111111111101100100001111;
assign LUT_1[36667] = 32'b11111111111111110110110110001011;
assign LUT_1[36668] = 32'b00000000000000001001101111010101;
assign LUT_1[36669] = 32'b00000000000000000011000001010001;
assign LUT_1[36670] = 32'b00000000000000000101011101100110;
assign LUT_1[36671] = 32'b11111111111111111110101111100010;
assign LUT_1[36672] = 32'b00000000000000000001101111010000;
assign LUT_1[36673] = 32'b11111111111111111011000001001100;
assign LUT_1[36674] = 32'b11111111111111111101011101100001;
assign LUT_1[36675] = 32'b11111111111111110110101111011101;
assign LUT_1[36676] = 32'b00000000000000001001101000100111;
assign LUT_1[36677] = 32'b00000000000000000010111010100011;
assign LUT_1[36678] = 32'b00000000000000000101010110111000;
assign LUT_1[36679] = 32'b11111111111111111110101000110100;
assign LUT_1[36680] = 32'b00000000000000000000111101000101;
assign LUT_1[36681] = 32'b11111111111111111010001111000001;
assign LUT_1[36682] = 32'b11111111111111111100101011010110;
assign LUT_1[36683] = 32'b11111111111111110101111101010010;
assign LUT_1[36684] = 32'b00000000000000001000110110011100;
assign LUT_1[36685] = 32'b00000000000000000010001000011000;
assign LUT_1[36686] = 32'b00000000000000000100100100101101;
assign LUT_1[36687] = 32'b11111111111111111101110110101001;
assign LUT_1[36688] = 32'b00000000000000000011101010110010;
assign LUT_1[36689] = 32'b11111111111111111100111100101110;
assign LUT_1[36690] = 32'b11111111111111111111011001000011;
assign LUT_1[36691] = 32'b11111111111111111000101010111111;
assign LUT_1[36692] = 32'b00000000000000001011100100001001;
assign LUT_1[36693] = 32'b00000000000000000100110110000101;
assign LUT_1[36694] = 32'b00000000000000000111010010011010;
assign LUT_1[36695] = 32'b00000000000000000000100100010110;
assign LUT_1[36696] = 32'b00000000000000000010111000100111;
assign LUT_1[36697] = 32'b11111111111111111100001010100011;
assign LUT_1[36698] = 32'b11111111111111111110100110111000;
assign LUT_1[36699] = 32'b11111111111111110111111000110100;
assign LUT_1[36700] = 32'b00000000000000001010110001111110;
assign LUT_1[36701] = 32'b00000000000000000100000011111010;
assign LUT_1[36702] = 32'b00000000000000000110100000001111;
assign LUT_1[36703] = 32'b11111111111111111111110010001011;
assign LUT_1[36704] = 32'b00000000000000000010101010001111;
assign LUT_1[36705] = 32'b11111111111111111011111100001011;
assign LUT_1[36706] = 32'b11111111111111111110011000100000;
assign LUT_1[36707] = 32'b11111111111111110111101010011100;
assign LUT_1[36708] = 32'b00000000000000001010100011100110;
assign LUT_1[36709] = 32'b00000000000000000011110101100010;
assign LUT_1[36710] = 32'b00000000000000000110010001110111;
assign LUT_1[36711] = 32'b11111111111111111111100011110011;
assign LUT_1[36712] = 32'b00000000000000000001111000000100;
assign LUT_1[36713] = 32'b11111111111111111011001010000000;
assign LUT_1[36714] = 32'b11111111111111111101100110010101;
assign LUT_1[36715] = 32'b11111111111111110110111000010001;
assign LUT_1[36716] = 32'b00000000000000001001110001011011;
assign LUT_1[36717] = 32'b00000000000000000011000011010111;
assign LUT_1[36718] = 32'b00000000000000000101011111101100;
assign LUT_1[36719] = 32'b11111111111111111110110001101000;
assign LUT_1[36720] = 32'b00000000000000000100100101110001;
assign LUT_1[36721] = 32'b11111111111111111101110111101101;
assign LUT_1[36722] = 32'b00000000000000000000010100000010;
assign LUT_1[36723] = 32'b11111111111111111001100101111110;
assign LUT_1[36724] = 32'b00000000000000001100011111001000;
assign LUT_1[36725] = 32'b00000000000000000101110001000100;
assign LUT_1[36726] = 32'b00000000000000001000001101011001;
assign LUT_1[36727] = 32'b00000000000000000001011111010101;
assign LUT_1[36728] = 32'b00000000000000000011110011100110;
assign LUT_1[36729] = 32'b11111111111111111101000101100010;
assign LUT_1[36730] = 32'b11111111111111111111100001110111;
assign LUT_1[36731] = 32'b11111111111111111000110011110011;
assign LUT_1[36732] = 32'b00000000000000001011101100111101;
assign LUT_1[36733] = 32'b00000000000000000100111110111001;
assign LUT_1[36734] = 32'b00000000000000000111011011001110;
assign LUT_1[36735] = 32'b00000000000000000000101101001010;
assign LUT_1[36736] = 32'b00000000000000000010110001101011;
assign LUT_1[36737] = 32'b11111111111111111100000011100111;
assign LUT_1[36738] = 32'b11111111111111111110011111111100;
assign LUT_1[36739] = 32'b11111111111111110111110001111000;
assign LUT_1[36740] = 32'b00000000000000001010101011000010;
assign LUT_1[36741] = 32'b00000000000000000011111100111110;
assign LUT_1[36742] = 32'b00000000000000000110011001010011;
assign LUT_1[36743] = 32'b11111111111111111111101011001111;
assign LUT_1[36744] = 32'b00000000000000000001111111100000;
assign LUT_1[36745] = 32'b11111111111111111011010001011100;
assign LUT_1[36746] = 32'b11111111111111111101101101110001;
assign LUT_1[36747] = 32'b11111111111111110110111111101101;
assign LUT_1[36748] = 32'b00000000000000001001111000110111;
assign LUT_1[36749] = 32'b00000000000000000011001010110011;
assign LUT_1[36750] = 32'b00000000000000000101100111001000;
assign LUT_1[36751] = 32'b11111111111111111110111001000100;
assign LUT_1[36752] = 32'b00000000000000000100101101001101;
assign LUT_1[36753] = 32'b11111111111111111101111111001001;
assign LUT_1[36754] = 32'b00000000000000000000011011011110;
assign LUT_1[36755] = 32'b11111111111111111001101101011010;
assign LUT_1[36756] = 32'b00000000000000001100100110100100;
assign LUT_1[36757] = 32'b00000000000000000101111000100000;
assign LUT_1[36758] = 32'b00000000000000001000010100110101;
assign LUT_1[36759] = 32'b00000000000000000001100110110001;
assign LUT_1[36760] = 32'b00000000000000000011111011000010;
assign LUT_1[36761] = 32'b11111111111111111101001100111110;
assign LUT_1[36762] = 32'b11111111111111111111101001010011;
assign LUT_1[36763] = 32'b11111111111111111000111011001111;
assign LUT_1[36764] = 32'b00000000000000001011110100011001;
assign LUT_1[36765] = 32'b00000000000000000101000110010101;
assign LUT_1[36766] = 32'b00000000000000000111100010101010;
assign LUT_1[36767] = 32'b00000000000000000000110100100110;
assign LUT_1[36768] = 32'b00000000000000000011101100101010;
assign LUT_1[36769] = 32'b11111111111111111100111110100110;
assign LUT_1[36770] = 32'b11111111111111111111011010111011;
assign LUT_1[36771] = 32'b11111111111111111000101100110111;
assign LUT_1[36772] = 32'b00000000000000001011100110000001;
assign LUT_1[36773] = 32'b00000000000000000100110111111101;
assign LUT_1[36774] = 32'b00000000000000000111010100010010;
assign LUT_1[36775] = 32'b00000000000000000000100110001110;
assign LUT_1[36776] = 32'b00000000000000000010111010011111;
assign LUT_1[36777] = 32'b11111111111111111100001100011011;
assign LUT_1[36778] = 32'b11111111111111111110101000110000;
assign LUT_1[36779] = 32'b11111111111111110111111010101100;
assign LUT_1[36780] = 32'b00000000000000001010110011110110;
assign LUT_1[36781] = 32'b00000000000000000100000101110010;
assign LUT_1[36782] = 32'b00000000000000000110100010000111;
assign LUT_1[36783] = 32'b11111111111111111111110100000011;
assign LUT_1[36784] = 32'b00000000000000000101101000001100;
assign LUT_1[36785] = 32'b11111111111111111110111010001000;
assign LUT_1[36786] = 32'b00000000000000000001010110011101;
assign LUT_1[36787] = 32'b11111111111111111010101000011001;
assign LUT_1[36788] = 32'b00000000000000001101100001100011;
assign LUT_1[36789] = 32'b00000000000000000110110011011111;
assign LUT_1[36790] = 32'b00000000000000001001001111110100;
assign LUT_1[36791] = 32'b00000000000000000010100001110000;
assign LUT_1[36792] = 32'b00000000000000000100110110000001;
assign LUT_1[36793] = 32'b11111111111111111110000111111101;
assign LUT_1[36794] = 32'b00000000000000000000100100010010;
assign LUT_1[36795] = 32'b11111111111111111001110110001110;
assign LUT_1[36796] = 32'b00000000000000001100101111011000;
assign LUT_1[36797] = 32'b00000000000000000110000001010100;
assign LUT_1[36798] = 32'b00000000000000001000011101101001;
assign LUT_1[36799] = 32'b00000000000000000001101111100101;
assign LUT_1[36800] = 32'b00000000000000000100101111010011;
assign LUT_1[36801] = 32'b11111111111111111110000001001111;
assign LUT_1[36802] = 32'b00000000000000000000011101100100;
assign LUT_1[36803] = 32'b11111111111111111001101111100000;
assign LUT_1[36804] = 32'b00000000000000001100101000101010;
assign LUT_1[36805] = 32'b00000000000000000101111010100110;
assign LUT_1[36806] = 32'b00000000000000001000010110111011;
assign LUT_1[36807] = 32'b00000000000000000001101000110111;
assign LUT_1[36808] = 32'b00000000000000000011111101001000;
assign LUT_1[36809] = 32'b11111111111111111101001111000100;
assign LUT_1[36810] = 32'b11111111111111111111101011011001;
assign LUT_1[36811] = 32'b11111111111111111000111101010101;
assign LUT_1[36812] = 32'b00000000000000001011110110011111;
assign LUT_1[36813] = 32'b00000000000000000101001000011011;
assign LUT_1[36814] = 32'b00000000000000000111100100110000;
assign LUT_1[36815] = 32'b00000000000000000000110110101100;
assign LUT_1[36816] = 32'b00000000000000000110101010110101;
assign LUT_1[36817] = 32'b11111111111111111111111100110001;
assign LUT_1[36818] = 32'b00000000000000000010011001000110;
assign LUT_1[36819] = 32'b11111111111111111011101011000010;
assign LUT_1[36820] = 32'b00000000000000001110100100001100;
assign LUT_1[36821] = 32'b00000000000000000111110110001000;
assign LUT_1[36822] = 32'b00000000000000001010010010011101;
assign LUT_1[36823] = 32'b00000000000000000011100100011001;
assign LUT_1[36824] = 32'b00000000000000000101111000101010;
assign LUT_1[36825] = 32'b11111111111111111111001010100110;
assign LUT_1[36826] = 32'b00000000000000000001100110111011;
assign LUT_1[36827] = 32'b11111111111111111010111000110111;
assign LUT_1[36828] = 32'b00000000000000001101110010000001;
assign LUT_1[36829] = 32'b00000000000000000111000011111101;
assign LUT_1[36830] = 32'b00000000000000001001100000010010;
assign LUT_1[36831] = 32'b00000000000000000010110010001110;
assign LUT_1[36832] = 32'b00000000000000000101101010010010;
assign LUT_1[36833] = 32'b11111111111111111110111100001110;
assign LUT_1[36834] = 32'b00000000000000000001011000100011;
assign LUT_1[36835] = 32'b11111111111111111010101010011111;
assign LUT_1[36836] = 32'b00000000000000001101100011101001;
assign LUT_1[36837] = 32'b00000000000000000110110101100101;
assign LUT_1[36838] = 32'b00000000000000001001010001111010;
assign LUT_1[36839] = 32'b00000000000000000010100011110110;
assign LUT_1[36840] = 32'b00000000000000000100111000000111;
assign LUT_1[36841] = 32'b11111111111111111110001010000011;
assign LUT_1[36842] = 32'b00000000000000000000100110011000;
assign LUT_1[36843] = 32'b11111111111111111001111000010100;
assign LUT_1[36844] = 32'b00000000000000001100110001011110;
assign LUT_1[36845] = 32'b00000000000000000110000011011010;
assign LUT_1[36846] = 32'b00000000000000001000011111101111;
assign LUT_1[36847] = 32'b00000000000000000001110001101011;
assign LUT_1[36848] = 32'b00000000000000000111100101110100;
assign LUT_1[36849] = 32'b00000000000000000000110111110000;
assign LUT_1[36850] = 32'b00000000000000000011010100000101;
assign LUT_1[36851] = 32'b11111111111111111100100110000001;
assign LUT_1[36852] = 32'b00000000000000001111011111001011;
assign LUT_1[36853] = 32'b00000000000000001000110001000111;
assign LUT_1[36854] = 32'b00000000000000001011001101011100;
assign LUT_1[36855] = 32'b00000000000000000100011111011000;
assign LUT_1[36856] = 32'b00000000000000000110110011101001;
assign LUT_1[36857] = 32'b00000000000000000000000101100101;
assign LUT_1[36858] = 32'b00000000000000000010100001111010;
assign LUT_1[36859] = 32'b11111111111111111011110011110110;
assign LUT_1[36860] = 32'b00000000000000001110101101000000;
assign LUT_1[36861] = 32'b00000000000000000111111110111100;
assign LUT_1[36862] = 32'b00000000000000001010011011010001;
assign LUT_1[36863] = 32'b00000000000000000011101101001101;
assign LUT_1[36864] = 32'b00000000000000000000101011011010;
assign LUT_1[36865] = 32'b11111111111111111001111101010110;
assign LUT_1[36866] = 32'b11111111111111111100011001101011;
assign LUT_1[36867] = 32'b11111111111111110101101011100111;
assign LUT_1[36868] = 32'b00000000000000001000100100110001;
assign LUT_1[36869] = 32'b00000000000000000001110110101101;
assign LUT_1[36870] = 32'b00000000000000000100010011000010;
assign LUT_1[36871] = 32'b11111111111111111101100100111110;
assign LUT_1[36872] = 32'b11111111111111111111111001001111;
assign LUT_1[36873] = 32'b11111111111111111001001011001011;
assign LUT_1[36874] = 32'b11111111111111111011100111100000;
assign LUT_1[36875] = 32'b11111111111111110100111001011100;
assign LUT_1[36876] = 32'b00000000000000000111110010100110;
assign LUT_1[36877] = 32'b00000000000000000001000100100010;
assign LUT_1[36878] = 32'b00000000000000000011100000110111;
assign LUT_1[36879] = 32'b11111111111111111100110010110011;
assign LUT_1[36880] = 32'b00000000000000000010100110111100;
assign LUT_1[36881] = 32'b11111111111111111011111000111000;
assign LUT_1[36882] = 32'b11111111111111111110010101001101;
assign LUT_1[36883] = 32'b11111111111111110111100111001001;
assign LUT_1[36884] = 32'b00000000000000001010100000010011;
assign LUT_1[36885] = 32'b00000000000000000011110010001111;
assign LUT_1[36886] = 32'b00000000000000000110001110100100;
assign LUT_1[36887] = 32'b11111111111111111111100000100000;
assign LUT_1[36888] = 32'b00000000000000000001110100110001;
assign LUT_1[36889] = 32'b11111111111111111011000110101101;
assign LUT_1[36890] = 32'b11111111111111111101100011000010;
assign LUT_1[36891] = 32'b11111111111111110110110100111110;
assign LUT_1[36892] = 32'b00000000000000001001101110001000;
assign LUT_1[36893] = 32'b00000000000000000011000000000100;
assign LUT_1[36894] = 32'b00000000000000000101011100011001;
assign LUT_1[36895] = 32'b11111111111111111110101110010101;
assign LUT_1[36896] = 32'b00000000000000000001100110011001;
assign LUT_1[36897] = 32'b11111111111111111010111000010101;
assign LUT_1[36898] = 32'b11111111111111111101010100101010;
assign LUT_1[36899] = 32'b11111111111111110110100110100110;
assign LUT_1[36900] = 32'b00000000000000001001011111110000;
assign LUT_1[36901] = 32'b00000000000000000010110001101100;
assign LUT_1[36902] = 32'b00000000000000000101001110000001;
assign LUT_1[36903] = 32'b11111111111111111110011111111101;
assign LUT_1[36904] = 32'b00000000000000000000110100001110;
assign LUT_1[36905] = 32'b11111111111111111010000110001010;
assign LUT_1[36906] = 32'b11111111111111111100100010011111;
assign LUT_1[36907] = 32'b11111111111111110101110100011011;
assign LUT_1[36908] = 32'b00000000000000001000101101100101;
assign LUT_1[36909] = 32'b00000000000000000001111111100001;
assign LUT_1[36910] = 32'b00000000000000000100011011110110;
assign LUT_1[36911] = 32'b11111111111111111101101101110010;
assign LUT_1[36912] = 32'b00000000000000000011100001111011;
assign LUT_1[36913] = 32'b11111111111111111100110011110111;
assign LUT_1[36914] = 32'b11111111111111111111010000001100;
assign LUT_1[36915] = 32'b11111111111111111000100010001000;
assign LUT_1[36916] = 32'b00000000000000001011011011010010;
assign LUT_1[36917] = 32'b00000000000000000100101101001110;
assign LUT_1[36918] = 32'b00000000000000000111001001100011;
assign LUT_1[36919] = 32'b00000000000000000000011011011111;
assign LUT_1[36920] = 32'b00000000000000000010101111110000;
assign LUT_1[36921] = 32'b11111111111111111100000001101100;
assign LUT_1[36922] = 32'b11111111111111111110011110000001;
assign LUT_1[36923] = 32'b11111111111111110111101111111101;
assign LUT_1[36924] = 32'b00000000000000001010101001000111;
assign LUT_1[36925] = 32'b00000000000000000011111011000011;
assign LUT_1[36926] = 32'b00000000000000000110010111011000;
assign LUT_1[36927] = 32'b11111111111111111111101001010100;
assign LUT_1[36928] = 32'b00000000000000000010101001000010;
assign LUT_1[36929] = 32'b11111111111111111011111010111110;
assign LUT_1[36930] = 32'b11111111111111111110010111010011;
assign LUT_1[36931] = 32'b11111111111111110111101001001111;
assign LUT_1[36932] = 32'b00000000000000001010100010011001;
assign LUT_1[36933] = 32'b00000000000000000011110100010101;
assign LUT_1[36934] = 32'b00000000000000000110010000101010;
assign LUT_1[36935] = 32'b11111111111111111111100010100110;
assign LUT_1[36936] = 32'b00000000000000000001110110110111;
assign LUT_1[36937] = 32'b11111111111111111011001000110011;
assign LUT_1[36938] = 32'b11111111111111111101100101001000;
assign LUT_1[36939] = 32'b11111111111111110110110111000100;
assign LUT_1[36940] = 32'b00000000000000001001110000001110;
assign LUT_1[36941] = 32'b00000000000000000011000010001010;
assign LUT_1[36942] = 32'b00000000000000000101011110011111;
assign LUT_1[36943] = 32'b11111111111111111110110000011011;
assign LUT_1[36944] = 32'b00000000000000000100100100100100;
assign LUT_1[36945] = 32'b11111111111111111101110110100000;
assign LUT_1[36946] = 32'b00000000000000000000010010110101;
assign LUT_1[36947] = 32'b11111111111111111001100100110001;
assign LUT_1[36948] = 32'b00000000000000001100011101111011;
assign LUT_1[36949] = 32'b00000000000000000101101111110111;
assign LUT_1[36950] = 32'b00000000000000001000001100001100;
assign LUT_1[36951] = 32'b00000000000000000001011110001000;
assign LUT_1[36952] = 32'b00000000000000000011110010011001;
assign LUT_1[36953] = 32'b11111111111111111101000100010101;
assign LUT_1[36954] = 32'b11111111111111111111100000101010;
assign LUT_1[36955] = 32'b11111111111111111000110010100110;
assign LUT_1[36956] = 32'b00000000000000001011101011110000;
assign LUT_1[36957] = 32'b00000000000000000100111101101100;
assign LUT_1[36958] = 32'b00000000000000000111011010000001;
assign LUT_1[36959] = 32'b00000000000000000000101011111101;
assign LUT_1[36960] = 32'b00000000000000000011100100000001;
assign LUT_1[36961] = 32'b11111111111111111100110101111101;
assign LUT_1[36962] = 32'b11111111111111111111010010010010;
assign LUT_1[36963] = 32'b11111111111111111000100100001110;
assign LUT_1[36964] = 32'b00000000000000001011011101011000;
assign LUT_1[36965] = 32'b00000000000000000100101111010100;
assign LUT_1[36966] = 32'b00000000000000000111001011101001;
assign LUT_1[36967] = 32'b00000000000000000000011101100101;
assign LUT_1[36968] = 32'b00000000000000000010110001110110;
assign LUT_1[36969] = 32'b11111111111111111100000011110010;
assign LUT_1[36970] = 32'b11111111111111111110100000000111;
assign LUT_1[36971] = 32'b11111111111111110111110010000011;
assign LUT_1[36972] = 32'b00000000000000001010101011001101;
assign LUT_1[36973] = 32'b00000000000000000011111101001001;
assign LUT_1[36974] = 32'b00000000000000000110011001011110;
assign LUT_1[36975] = 32'b11111111111111111111101011011010;
assign LUT_1[36976] = 32'b00000000000000000101011111100011;
assign LUT_1[36977] = 32'b11111111111111111110110001011111;
assign LUT_1[36978] = 32'b00000000000000000001001101110100;
assign LUT_1[36979] = 32'b11111111111111111010011111110000;
assign LUT_1[36980] = 32'b00000000000000001101011000111010;
assign LUT_1[36981] = 32'b00000000000000000110101010110110;
assign LUT_1[36982] = 32'b00000000000000001001000111001011;
assign LUT_1[36983] = 32'b00000000000000000010011001000111;
assign LUT_1[36984] = 32'b00000000000000000100101101011000;
assign LUT_1[36985] = 32'b11111111111111111101111111010100;
assign LUT_1[36986] = 32'b00000000000000000000011011101001;
assign LUT_1[36987] = 32'b11111111111111111001101101100101;
assign LUT_1[36988] = 32'b00000000000000001100100110101111;
assign LUT_1[36989] = 32'b00000000000000000101111000101011;
assign LUT_1[36990] = 32'b00000000000000001000010101000000;
assign LUT_1[36991] = 32'b00000000000000000001100110111100;
assign LUT_1[36992] = 32'b00000000000000000011101011011101;
assign LUT_1[36993] = 32'b11111111111111111100111101011001;
assign LUT_1[36994] = 32'b11111111111111111111011001101110;
assign LUT_1[36995] = 32'b11111111111111111000101011101010;
assign LUT_1[36996] = 32'b00000000000000001011100100110100;
assign LUT_1[36997] = 32'b00000000000000000100110110110000;
assign LUT_1[36998] = 32'b00000000000000000111010011000101;
assign LUT_1[36999] = 32'b00000000000000000000100101000001;
assign LUT_1[37000] = 32'b00000000000000000010111001010010;
assign LUT_1[37001] = 32'b11111111111111111100001011001110;
assign LUT_1[37002] = 32'b11111111111111111110100111100011;
assign LUT_1[37003] = 32'b11111111111111110111111001011111;
assign LUT_1[37004] = 32'b00000000000000001010110010101001;
assign LUT_1[37005] = 32'b00000000000000000100000100100101;
assign LUT_1[37006] = 32'b00000000000000000110100000111010;
assign LUT_1[37007] = 32'b11111111111111111111110010110110;
assign LUT_1[37008] = 32'b00000000000000000101100110111111;
assign LUT_1[37009] = 32'b11111111111111111110111000111011;
assign LUT_1[37010] = 32'b00000000000000000001010101010000;
assign LUT_1[37011] = 32'b11111111111111111010100111001100;
assign LUT_1[37012] = 32'b00000000000000001101100000010110;
assign LUT_1[37013] = 32'b00000000000000000110110010010010;
assign LUT_1[37014] = 32'b00000000000000001001001110100111;
assign LUT_1[37015] = 32'b00000000000000000010100000100011;
assign LUT_1[37016] = 32'b00000000000000000100110100110100;
assign LUT_1[37017] = 32'b11111111111111111110000110110000;
assign LUT_1[37018] = 32'b00000000000000000000100011000101;
assign LUT_1[37019] = 32'b11111111111111111001110101000001;
assign LUT_1[37020] = 32'b00000000000000001100101110001011;
assign LUT_1[37021] = 32'b00000000000000000110000000000111;
assign LUT_1[37022] = 32'b00000000000000001000011100011100;
assign LUT_1[37023] = 32'b00000000000000000001101110011000;
assign LUT_1[37024] = 32'b00000000000000000100100110011100;
assign LUT_1[37025] = 32'b11111111111111111101111000011000;
assign LUT_1[37026] = 32'b00000000000000000000010100101101;
assign LUT_1[37027] = 32'b11111111111111111001100110101001;
assign LUT_1[37028] = 32'b00000000000000001100011111110011;
assign LUT_1[37029] = 32'b00000000000000000101110001101111;
assign LUT_1[37030] = 32'b00000000000000001000001110000100;
assign LUT_1[37031] = 32'b00000000000000000001100000000000;
assign LUT_1[37032] = 32'b00000000000000000011110100010001;
assign LUT_1[37033] = 32'b11111111111111111101000110001101;
assign LUT_1[37034] = 32'b11111111111111111111100010100010;
assign LUT_1[37035] = 32'b11111111111111111000110100011110;
assign LUT_1[37036] = 32'b00000000000000001011101101101000;
assign LUT_1[37037] = 32'b00000000000000000100111111100100;
assign LUT_1[37038] = 32'b00000000000000000111011011111001;
assign LUT_1[37039] = 32'b00000000000000000000101101110101;
assign LUT_1[37040] = 32'b00000000000000000110100001111110;
assign LUT_1[37041] = 32'b11111111111111111111110011111010;
assign LUT_1[37042] = 32'b00000000000000000010010000001111;
assign LUT_1[37043] = 32'b11111111111111111011100010001011;
assign LUT_1[37044] = 32'b00000000000000001110011011010101;
assign LUT_1[37045] = 32'b00000000000000000111101101010001;
assign LUT_1[37046] = 32'b00000000000000001010001001100110;
assign LUT_1[37047] = 32'b00000000000000000011011011100010;
assign LUT_1[37048] = 32'b00000000000000000101101111110011;
assign LUT_1[37049] = 32'b11111111111111111111000001101111;
assign LUT_1[37050] = 32'b00000000000000000001011110000100;
assign LUT_1[37051] = 32'b11111111111111111010110000000000;
assign LUT_1[37052] = 32'b00000000000000001101101001001010;
assign LUT_1[37053] = 32'b00000000000000000110111011000110;
assign LUT_1[37054] = 32'b00000000000000001001010111011011;
assign LUT_1[37055] = 32'b00000000000000000010101001010111;
assign LUT_1[37056] = 32'b00000000000000000101101001000101;
assign LUT_1[37057] = 32'b11111111111111111110111011000001;
assign LUT_1[37058] = 32'b00000000000000000001010111010110;
assign LUT_1[37059] = 32'b11111111111111111010101001010010;
assign LUT_1[37060] = 32'b00000000000000001101100010011100;
assign LUT_1[37061] = 32'b00000000000000000110110100011000;
assign LUT_1[37062] = 32'b00000000000000001001010000101101;
assign LUT_1[37063] = 32'b00000000000000000010100010101001;
assign LUT_1[37064] = 32'b00000000000000000100110110111010;
assign LUT_1[37065] = 32'b11111111111111111110001000110110;
assign LUT_1[37066] = 32'b00000000000000000000100101001011;
assign LUT_1[37067] = 32'b11111111111111111001110111000111;
assign LUT_1[37068] = 32'b00000000000000001100110000010001;
assign LUT_1[37069] = 32'b00000000000000000110000010001101;
assign LUT_1[37070] = 32'b00000000000000001000011110100010;
assign LUT_1[37071] = 32'b00000000000000000001110000011110;
assign LUT_1[37072] = 32'b00000000000000000111100100100111;
assign LUT_1[37073] = 32'b00000000000000000000110110100011;
assign LUT_1[37074] = 32'b00000000000000000011010010111000;
assign LUT_1[37075] = 32'b11111111111111111100100100110100;
assign LUT_1[37076] = 32'b00000000000000001111011101111110;
assign LUT_1[37077] = 32'b00000000000000001000101111111010;
assign LUT_1[37078] = 32'b00000000000000001011001100001111;
assign LUT_1[37079] = 32'b00000000000000000100011110001011;
assign LUT_1[37080] = 32'b00000000000000000110110010011100;
assign LUT_1[37081] = 32'b00000000000000000000000100011000;
assign LUT_1[37082] = 32'b00000000000000000010100000101101;
assign LUT_1[37083] = 32'b11111111111111111011110010101001;
assign LUT_1[37084] = 32'b00000000000000001110101011110011;
assign LUT_1[37085] = 32'b00000000000000000111111101101111;
assign LUT_1[37086] = 32'b00000000000000001010011010000100;
assign LUT_1[37087] = 32'b00000000000000000011101100000000;
assign LUT_1[37088] = 32'b00000000000000000110100100000100;
assign LUT_1[37089] = 32'b11111111111111111111110110000000;
assign LUT_1[37090] = 32'b00000000000000000010010010010101;
assign LUT_1[37091] = 32'b11111111111111111011100100010001;
assign LUT_1[37092] = 32'b00000000000000001110011101011011;
assign LUT_1[37093] = 32'b00000000000000000111101111010111;
assign LUT_1[37094] = 32'b00000000000000001010001011101100;
assign LUT_1[37095] = 32'b00000000000000000011011101101000;
assign LUT_1[37096] = 32'b00000000000000000101110001111001;
assign LUT_1[37097] = 32'b11111111111111111111000011110101;
assign LUT_1[37098] = 32'b00000000000000000001100000001010;
assign LUT_1[37099] = 32'b11111111111111111010110010000110;
assign LUT_1[37100] = 32'b00000000000000001101101011010000;
assign LUT_1[37101] = 32'b00000000000000000110111101001100;
assign LUT_1[37102] = 32'b00000000000000001001011001100001;
assign LUT_1[37103] = 32'b00000000000000000010101011011101;
assign LUT_1[37104] = 32'b00000000000000001000011111100110;
assign LUT_1[37105] = 32'b00000000000000000001110001100010;
assign LUT_1[37106] = 32'b00000000000000000100001101110111;
assign LUT_1[37107] = 32'b11111111111111111101011111110011;
assign LUT_1[37108] = 32'b00000000000000010000011000111101;
assign LUT_1[37109] = 32'b00000000000000001001101010111001;
assign LUT_1[37110] = 32'b00000000000000001100000111001110;
assign LUT_1[37111] = 32'b00000000000000000101011001001010;
assign LUT_1[37112] = 32'b00000000000000000111101101011011;
assign LUT_1[37113] = 32'b00000000000000000000111111010111;
assign LUT_1[37114] = 32'b00000000000000000011011011101100;
assign LUT_1[37115] = 32'b11111111111111111100101101101000;
assign LUT_1[37116] = 32'b00000000000000001111100110110010;
assign LUT_1[37117] = 32'b00000000000000001000111000101110;
assign LUT_1[37118] = 32'b00000000000000001011010101000011;
assign LUT_1[37119] = 32'b00000000000000000100100110111111;
assign LUT_1[37120] = 32'b11111111111111111110011111100110;
assign LUT_1[37121] = 32'b11111111111111110111110001100010;
assign LUT_1[37122] = 32'b11111111111111111010001101110111;
assign LUT_1[37123] = 32'b11111111111111110011011111110011;
assign LUT_1[37124] = 32'b00000000000000000110011000111101;
assign LUT_1[37125] = 32'b11111111111111111111101010111001;
assign LUT_1[37126] = 32'b00000000000000000010000111001110;
assign LUT_1[37127] = 32'b11111111111111111011011001001010;
assign LUT_1[37128] = 32'b11111111111111111101101101011011;
assign LUT_1[37129] = 32'b11111111111111110110111111010111;
assign LUT_1[37130] = 32'b11111111111111111001011011101100;
assign LUT_1[37131] = 32'b11111111111111110010101101101000;
assign LUT_1[37132] = 32'b00000000000000000101100110110010;
assign LUT_1[37133] = 32'b11111111111111111110111000101110;
assign LUT_1[37134] = 32'b00000000000000000001010101000011;
assign LUT_1[37135] = 32'b11111111111111111010100110111111;
assign LUT_1[37136] = 32'b00000000000000000000011011001000;
assign LUT_1[37137] = 32'b11111111111111111001101101000100;
assign LUT_1[37138] = 32'b11111111111111111100001001011001;
assign LUT_1[37139] = 32'b11111111111111110101011011010101;
assign LUT_1[37140] = 32'b00000000000000001000010100011111;
assign LUT_1[37141] = 32'b00000000000000000001100110011011;
assign LUT_1[37142] = 32'b00000000000000000100000010110000;
assign LUT_1[37143] = 32'b11111111111111111101010100101100;
assign LUT_1[37144] = 32'b11111111111111111111101000111101;
assign LUT_1[37145] = 32'b11111111111111111000111010111001;
assign LUT_1[37146] = 32'b11111111111111111011010111001110;
assign LUT_1[37147] = 32'b11111111111111110100101001001010;
assign LUT_1[37148] = 32'b00000000000000000111100010010100;
assign LUT_1[37149] = 32'b00000000000000000000110100010000;
assign LUT_1[37150] = 32'b00000000000000000011010000100101;
assign LUT_1[37151] = 32'b11111111111111111100100010100001;
assign LUT_1[37152] = 32'b11111111111111111111011010100101;
assign LUT_1[37153] = 32'b11111111111111111000101100100001;
assign LUT_1[37154] = 32'b11111111111111111011001000110110;
assign LUT_1[37155] = 32'b11111111111111110100011010110010;
assign LUT_1[37156] = 32'b00000000000000000111010011111100;
assign LUT_1[37157] = 32'b00000000000000000000100101111000;
assign LUT_1[37158] = 32'b00000000000000000011000010001101;
assign LUT_1[37159] = 32'b11111111111111111100010100001001;
assign LUT_1[37160] = 32'b11111111111111111110101000011010;
assign LUT_1[37161] = 32'b11111111111111110111111010010110;
assign LUT_1[37162] = 32'b11111111111111111010010110101011;
assign LUT_1[37163] = 32'b11111111111111110011101000100111;
assign LUT_1[37164] = 32'b00000000000000000110100001110001;
assign LUT_1[37165] = 32'b11111111111111111111110011101101;
assign LUT_1[37166] = 32'b00000000000000000010010000000010;
assign LUT_1[37167] = 32'b11111111111111111011100001111110;
assign LUT_1[37168] = 32'b00000000000000000001010110000111;
assign LUT_1[37169] = 32'b11111111111111111010101000000011;
assign LUT_1[37170] = 32'b11111111111111111101000100011000;
assign LUT_1[37171] = 32'b11111111111111110110010110010100;
assign LUT_1[37172] = 32'b00000000000000001001001111011110;
assign LUT_1[37173] = 32'b00000000000000000010100001011010;
assign LUT_1[37174] = 32'b00000000000000000100111101101111;
assign LUT_1[37175] = 32'b11111111111111111110001111101011;
assign LUT_1[37176] = 32'b00000000000000000000100011111100;
assign LUT_1[37177] = 32'b11111111111111111001110101111000;
assign LUT_1[37178] = 32'b11111111111111111100010010001101;
assign LUT_1[37179] = 32'b11111111111111110101100100001001;
assign LUT_1[37180] = 32'b00000000000000001000011101010011;
assign LUT_1[37181] = 32'b00000000000000000001101111001111;
assign LUT_1[37182] = 32'b00000000000000000100001011100100;
assign LUT_1[37183] = 32'b11111111111111111101011101100000;
assign LUT_1[37184] = 32'b00000000000000000000011101001110;
assign LUT_1[37185] = 32'b11111111111111111001101111001010;
assign LUT_1[37186] = 32'b11111111111111111100001011011111;
assign LUT_1[37187] = 32'b11111111111111110101011101011011;
assign LUT_1[37188] = 32'b00000000000000001000010110100101;
assign LUT_1[37189] = 32'b00000000000000000001101000100001;
assign LUT_1[37190] = 32'b00000000000000000100000100110110;
assign LUT_1[37191] = 32'b11111111111111111101010110110010;
assign LUT_1[37192] = 32'b11111111111111111111101011000011;
assign LUT_1[37193] = 32'b11111111111111111000111100111111;
assign LUT_1[37194] = 32'b11111111111111111011011001010100;
assign LUT_1[37195] = 32'b11111111111111110100101011010000;
assign LUT_1[37196] = 32'b00000000000000000111100100011010;
assign LUT_1[37197] = 32'b00000000000000000000110110010110;
assign LUT_1[37198] = 32'b00000000000000000011010010101011;
assign LUT_1[37199] = 32'b11111111111111111100100100100111;
assign LUT_1[37200] = 32'b00000000000000000010011000110000;
assign LUT_1[37201] = 32'b11111111111111111011101010101100;
assign LUT_1[37202] = 32'b11111111111111111110000111000001;
assign LUT_1[37203] = 32'b11111111111111110111011000111101;
assign LUT_1[37204] = 32'b00000000000000001010010010000111;
assign LUT_1[37205] = 32'b00000000000000000011100100000011;
assign LUT_1[37206] = 32'b00000000000000000110000000011000;
assign LUT_1[37207] = 32'b11111111111111111111010010010100;
assign LUT_1[37208] = 32'b00000000000000000001100110100101;
assign LUT_1[37209] = 32'b11111111111111111010111000100001;
assign LUT_1[37210] = 32'b11111111111111111101010100110110;
assign LUT_1[37211] = 32'b11111111111111110110100110110010;
assign LUT_1[37212] = 32'b00000000000000001001011111111100;
assign LUT_1[37213] = 32'b00000000000000000010110001111000;
assign LUT_1[37214] = 32'b00000000000000000101001110001101;
assign LUT_1[37215] = 32'b11111111111111111110100000001001;
assign LUT_1[37216] = 32'b00000000000000000001011000001101;
assign LUT_1[37217] = 32'b11111111111111111010101010001001;
assign LUT_1[37218] = 32'b11111111111111111101000110011110;
assign LUT_1[37219] = 32'b11111111111111110110011000011010;
assign LUT_1[37220] = 32'b00000000000000001001010001100100;
assign LUT_1[37221] = 32'b00000000000000000010100011100000;
assign LUT_1[37222] = 32'b00000000000000000100111111110101;
assign LUT_1[37223] = 32'b11111111111111111110010001110001;
assign LUT_1[37224] = 32'b00000000000000000000100110000010;
assign LUT_1[37225] = 32'b11111111111111111001110111111110;
assign LUT_1[37226] = 32'b11111111111111111100010100010011;
assign LUT_1[37227] = 32'b11111111111111110101100110001111;
assign LUT_1[37228] = 32'b00000000000000001000011111011001;
assign LUT_1[37229] = 32'b00000000000000000001110001010101;
assign LUT_1[37230] = 32'b00000000000000000100001101101010;
assign LUT_1[37231] = 32'b11111111111111111101011111100110;
assign LUT_1[37232] = 32'b00000000000000000011010011101111;
assign LUT_1[37233] = 32'b11111111111111111100100101101011;
assign LUT_1[37234] = 32'b11111111111111111111000010000000;
assign LUT_1[37235] = 32'b11111111111111111000010011111100;
assign LUT_1[37236] = 32'b00000000000000001011001101000110;
assign LUT_1[37237] = 32'b00000000000000000100011111000010;
assign LUT_1[37238] = 32'b00000000000000000110111011010111;
assign LUT_1[37239] = 32'b00000000000000000000001101010011;
assign LUT_1[37240] = 32'b00000000000000000010100001100100;
assign LUT_1[37241] = 32'b11111111111111111011110011100000;
assign LUT_1[37242] = 32'b11111111111111111110001111110101;
assign LUT_1[37243] = 32'b11111111111111110111100001110001;
assign LUT_1[37244] = 32'b00000000000000001010011010111011;
assign LUT_1[37245] = 32'b00000000000000000011101100110111;
assign LUT_1[37246] = 32'b00000000000000000110001001001100;
assign LUT_1[37247] = 32'b11111111111111111111011011001000;
assign LUT_1[37248] = 32'b00000000000000000001011111101001;
assign LUT_1[37249] = 32'b11111111111111111010110001100101;
assign LUT_1[37250] = 32'b11111111111111111101001101111010;
assign LUT_1[37251] = 32'b11111111111111110110011111110110;
assign LUT_1[37252] = 32'b00000000000000001001011001000000;
assign LUT_1[37253] = 32'b00000000000000000010101010111100;
assign LUT_1[37254] = 32'b00000000000000000101000111010001;
assign LUT_1[37255] = 32'b11111111111111111110011001001101;
assign LUT_1[37256] = 32'b00000000000000000000101101011110;
assign LUT_1[37257] = 32'b11111111111111111001111111011010;
assign LUT_1[37258] = 32'b11111111111111111100011011101111;
assign LUT_1[37259] = 32'b11111111111111110101101101101011;
assign LUT_1[37260] = 32'b00000000000000001000100110110101;
assign LUT_1[37261] = 32'b00000000000000000001111000110001;
assign LUT_1[37262] = 32'b00000000000000000100010101000110;
assign LUT_1[37263] = 32'b11111111111111111101100111000010;
assign LUT_1[37264] = 32'b00000000000000000011011011001011;
assign LUT_1[37265] = 32'b11111111111111111100101101000111;
assign LUT_1[37266] = 32'b11111111111111111111001001011100;
assign LUT_1[37267] = 32'b11111111111111111000011011011000;
assign LUT_1[37268] = 32'b00000000000000001011010100100010;
assign LUT_1[37269] = 32'b00000000000000000100100110011110;
assign LUT_1[37270] = 32'b00000000000000000111000010110011;
assign LUT_1[37271] = 32'b00000000000000000000010100101111;
assign LUT_1[37272] = 32'b00000000000000000010101001000000;
assign LUT_1[37273] = 32'b11111111111111111011111010111100;
assign LUT_1[37274] = 32'b11111111111111111110010111010001;
assign LUT_1[37275] = 32'b11111111111111110111101001001101;
assign LUT_1[37276] = 32'b00000000000000001010100010010111;
assign LUT_1[37277] = 32'b00000000000000000011110100010011;
assign LUT_1[37278] = 32'b00000000000000000110010000101000;
assign LUT_1[37279] = 32'b11111111111111111111100010100100;
assign LUT_1[37280] = 32'b00000000000000000010011010101000;
assign LUT_1[37281] = 32'b11111111111111111011101100100100;
assign LUT_1[37282] = 32'b11111111111111111110001000111001;
assign LUT_1[37283] = 32'b11111111111111110111011010110101;
assign LUT_1[37284] = 32'b00000000000000001010010011111111;
assign LUT_1[37285] = 32'b00000000000000000011100101111011;
assign LUT_1[37286] = 32'b00000000000000000110000010010000;
assign LUT_1[37287] = 32'b11111111111111111111010100001100;
assign LUT_1[37288] = 32'b00000000000000000001101000011101;
assign LUT_1[37289] = 32'b11111111111111111010111010011001;
assign LUT_1[37290] = 32'b11111111111111111101010110101110;
assign LUT_1[37291] = 32'b11111111111111110110101000101010;
assign LUT_1[37292] = 32'b00000000000000001001100001110100;
assign LUT_1[37293] = 32'b00000000000000000010110011110000;
assign LUT_1[37294] = 32'b00000000000000000101010000000101;
assign LUT_1[37295] = 32'b11111111111111111110100010000001;
assign LUT_1[37296] = 32'b00000000000000000100010110001010;
assign LUT_1[37297] = 32'b11111111111111111101101000000110;
assign LUT_1[37298] = 32'b00000000000000000000000100011011;
assign LUT_1[37299] = 32'b11111111111111111001010110010111;
assign LUT_1[37300] = 32'b00000000000000001100001111100001;
assign LUT_1[37301] = 32'b00000000000000000101100001011101;
assign LUT_1[37302] = 32'b00000000000000000111111101110010;
assign LUT_1[37303] = 32'b00000000000000000001001111101110;
assign LUT_1[37304] = 32'b00000000000000000011100011111111;
assign LUT_1[37305] = 32'b11111111111111111100110101111011;
assign LUT_1[37306] = 32'b11111111111111111111010010010000;
assign LUT_1[37307] = 32'b11111111111111111000100100001100;
assign LUT_1[37308] = 32'b00000000000000001011011101010110;
assign LUT_1[37309] = 32'b00000000000000000100101111010010;
assign LUT_1[37310] = 32'b00000000000000000111001011100111;
assign LUT_1[37311] = 32'b00000000000000000000011101100011;
assign LUT_1[37312] = 32'b00000000000000000011011101010001;
assign LUT_1[37313] = 32'b11111111111111111100101111001101;
assign LUT_1[37314] = 32'b11111111111111111111001011100010;
assign LUT_1[37315] = 32'b11111111111111111000011101011110;
assign LUT_1[37316] = 32'b00000000000000001011010110101000;
assign LUT_1[37317] = 32'b00000000000000000100101000100100;
assign LUT_1[37318] = 32'b00000000000000000111000100111001;
assign LUT_1[37319] = 32'b00000000000000000000010110110101;
assign LUT_1[37320] = 32'b00000000000000000010101011000110;
assign LUT_1[37321] = 32'b11111111111111111011111101000010;
assign LUT_1[37322] = 32'b11111111111111111110011001010111;
assign LUT_1[37323] = 32'b11111111111111110111101011010011;
assign LUT_1[37324] = 32'b00000000000000001010100100011101;
assign LUT_1[37325] = 32'b00000000000000000011110110011001;
assign LUT_1[37326] = 32'b00000000000000000110010010101110;
assign LUT_1[37327] = 32'b11111111111111111111100100101010;
assign LUT_1[37328] = 32'b00000000000000000101011000110011;
assign LUT_1[37329] = 32'b11111111111111111110101010101111;
assign LUT_1[37330] = 32'b00000000000000000001000111000100;
assign LUT_1[37331] = 32'b11111111111111111010011001000000;
assign LUT_1[37332] = 32'b00000000000000001101010010001010;
assign LUT_1[37333] = 32'b00000000000000000110100100000110;
assign LUT_1[37334] = 32'b00000000000000001001000000011011;
assign LUT_1[37335] = 32'b00000000000000000010010010010111;
assign LUT_1[37336] = 32'b00000000000000000100100110101000;
assign LUT_1[37337] = 32'b11111111111111111101111000100100;
assign LUT_1[37338] = 32'b00000000000000000000010100111001;
assign LUT_1[37339] = 32'b11111111111111111001100110110101;
assign LUT_1[37340] = 32'b00000000000000001100011111111111;
assign LUT_1[37341] = 32'b00000000000000000101110001111011;
assign LUT_1[37342] = 32'b00000000000000001000001110010000;
assign LUT_1[37343] = 32'b00000000000000000001100000001100;
assign LUT_1[37344] = 32'b00000000000000000100011000010000;
assign LUT_1[37345] = 32'b11111111111111111101101010001100;
assign LUT_1[37346] = 32'b00000000000000000000000110100001;
assign LUT_1[37347] = 32'b11111111111111111001011000011101;
assign LUT_1[37348] = 32'b00000000000000001100010001100111;
assign LUT_1[37349] = 32'b00000000000000000101100011100011;
assign LUT_1[37350] = 32'b00000000000000000111111111111000;
assign LUT_1[37351] = 32'b00000000000000000001010001110100;
assign LUT_1[37352] = 32'b00000000000000000011100110000101;
assign LUT_1[37353] = 32'b11111111111111111100111000000001;
assign LUT_1[37354] = 32'b11111111111111111111010100010110;
assign LUT_1[37355] = 32'b11111111111111111000100110010010;
assign LUT_1[37356] = 32'b00000000000000001011011111011100;
assign LUT_1[37357] = 32'b00000000000000000100110001011000;
assign LUT_1[37358] = 32'b00000000000000000111001101101101;
assign LUT_1[37359] = 32'b00000000000000000000011111101001;
assign LUT_1[37360] = 32'b00000000000000000110010011110010;
assign LUT_1[37361] = 32'b11111111111111111111100101101110;
assign LUT_1[37362] = 32'b00000000000000000010000010000011;
assign LUT_1[37363] = 32'b11111111111111111011010011111111;
assign LUT_1[37364] = 32'b00000000000000001110001101001001;
assign LUT_1[37365] = 32'b00000000000000000111011111000101;
assign LUT_1[37366] = 32'b00000000000000001001111011011010;
assign LUT_1[37367] = 32'b00000000000000000011001101010110;
assign LUT_1[37368] = 32'b00000000000000000101100001100111;
assign LUT_1[37369] = 32'b11111111111111111110110011100011;
assign LUT_1[37370] = 32'b00000000000000000001001111111000;
assign LUT_1[37371] = 32'b11111111111111111010100001110100;
assign LUT_1[37372] = 32'b00000000000000001101011010111110;
assign LUT_1[37373] = 32'b00000000000000000110101100111010;
assign LUT_1[37374] = 32'b00000000000000001001001001001111;
assign LUT_1[37375] = 32'b00000000000000000010011011001011;
assign LUT_1[37376] = 32'b11111111111111111010011001110111;
assign LUT_1[37377] = 32'b11111111111111110011101011110011;
assign LUT_1[37378] = 32'b11111111111111110110001000001000;
assign LUT_1[37379] = 32'b11111111111111101111011010000100;
assign LUT_1[37380] = 32'b00000000000000000010010011001110;
assign LUT_1[37381] = 32'b11111111111111111011100101001010;
assign LUT_1[37382] = 32'b11111111111111111110000001011111;
assign LUT_1[37383] = 32'b11111111111111110111010011011011;
assign LUT_1[37384] = 32'b11111111111111111001100111101100;
assign LUT_1[37385] = 32'b11111111111111110010111001101000;
assign LUT_1[37386] = 32'b11111111111111110101010101111101;
assign LUT_1[37387] = 32'b11111111111111101110100111111001;
assign LUT_1[37388] = 32'b00000000000000000001100001000011;
assign LUT_1[37389] = 32'b11111111111111111010110010111111;
assign LUT_1[37390] = 32'b11111111111111111101001111010100;
assign LUT_1[37391] = 32'b11111111111111110110100001010000;
assign LUT_1[37392] = 32'b11111111111111111100010101011001;
assign LUT_1[37393] = 32'b11111111111111110101100111010101;
assign LUT_1[37394] = 32'b11111111111111111000000011101010;
assign LUT_1[37395] = 32'b11111111111111110001010101100110;
assign LUT_1[37396] = 32'b00000000000000000100001110110000;
assign LUT_1[37397] = 32'b11111111111111111101100000101100;
assign LUT_1[37398] = 32'b11111111111111111111111101000001;
assign LUT_1[37399] = 32'b11111111111111111001001110111101;
assign LUT_1[37400] = 32'b11111111111111111011100011001110;
assign LUT_1[37401] = 32'b11111111111111110100110101001010;
assign LUT_1[37402] = 32'b11111111111111110111010001011111;
assign LUT_1[37403] = 32'b11111111111111110000100011011011;
assign LUT_1[37404] = 32'b00000000000000000011011100100101;
assign LUT_1[37405] = 32'b11111111111111111100101110100001;
assign LUT_1[37406] = 32'b11111111111111111111001010110110;
assign LUT_1[37407] = 32'b11111111111111111000011100110010;
assign LUT_1[37408] = 32'b11111111111111111011010100110110;
assign LUT_1[37409] = 32'b11111111111111110100100110110010;
assign LUT_1[37410] = 32'b11111111111111110111000011000111;
assign LUT_1[37411] = 32'b11111111111111110000010101000011;
assign LUT_1[37412] = 32'b00000000000000000011001110001101;
assign LUT_1[37413] = 32'b11111111111111111100100000001001;
assign LUT_1[37414] = 32'b11111111111111111110111100011110;
assign LUT_1[37415] = 32'b11111111111111111000001110011010;
assign LUT_1[37416] = 32'b11111111111111111010100010101011;
assign LUT_1[37417] = 32'b11111111111111110011110100100111;
assign LUT_1[37418] = 32'b11111111111111110110010000111100;
assign LUT_1[37419] = 32'b11111111111111101111100010111000;
assign LUT_1[37420] = 32'b00000000000000000010011100000010;
assign LUT_1[37421] = 32'b11111111111111111011101101111110;
assign LUT_1[37422] = 32'b11111111111111111110001010010011;
assign LUT_1[37423] = 32'b11111111111111110111011100001111;
assign LUT_1[37424] = 32'b11111111111111111101010000011000;
assign LUT_1[37425] = 32'b11111111111111110110100010010100;
assign LUT_1[37426] = 32'b11111111111111111000111110101001;
assign LUT_1[37427] = 32'b11111111111111110010010000100101;
assign LUT_1[37428] = 32'b00000000000000000101001001101111;
assign LUT_1[37429] = 32'b11111111111111111110011011101011;
assign LUT_1[37430] = 32'b00000000000000000000111000000000;
assign LUT_1[37431] = 32'b11111111111111111010001001111100;
assign LUT_1[37432] = 32'b11111111111111111100011110001101;
assign LUT_1[37433] = 32'b11111111111111110101110000001001;
assign LUT_1[37434] = 32'b11111111111111111000001100011110;
assign LUT_1[37435] = 32'b11111111111111110001011110011010;
assign LUT_1[37436] = 32'b00000000000000000100010111100100;
assign LUT_1[37437] = 32'b11111111111111111101101001100000;
assign LUT_1[37438] = 32'b00000000000000000000000101110101;
assign LUT_1[37439] = 32'b11111111111111111001010111110001;
assign LUT_1[37440] = 32'b11111111111111111100010111011111;
assign LUT_1[37441] = 32'b11111111111111110101101001011011;
assign LUT_1[37442] = 32'b11111111111111111000000101110000;
assign LUT_1[37443] = 32'b11111111111111110001010111101100;
assign LUT_1[37444] = 32'b00000000000000000100010000110110;
assign LUT_1[37445] = 32'b11111111111111111101100010110010;
assign LUT_1[37446] = 32'b11111111111111111111111111000111;
assign LUT_1[37447] = 32'b11111111111111111001010001000011;
assign LUT_1[37448] = 32'b11111111111111111011100101010100;
assign LUT_1[37449] = 32'b11111111111111110100110111010000;
assign LUT_1[37450] = 32'b11111111111111110111010011100101;
assign LUT_1[37451] = 32'b11111111111111110000100101100001;
assign LUT_1[37452] = 32'b00000000000000000011011110101011;
assign LUT_1[37453] = 32'b11111111111111111100110000100111;
assign LUT_1[37454] = 32'b11111111111111111111001100111100;
assign LUT_1[37455] = 32'b11111111111111111000011110111000;
assign LUT_1[37456] = 32'b11111111111111111110010011000001;
assign LUT_1[37457] = 32'b11111111111111110111100100111101;
assign LUT_1[37458] = 32'b11111111111111111010000001010010;
assign LUT_1[37459] = 32'b11111111111111110011010011001110;
assign LUT_1[37460] = 32'b00000000000000000110001100011000;
assign LUT_1[37461] = 32'b11111111111111111111011110010100;
assign LUT_1[37462] = 32'b00000000000000000001111010101001;
assign LUT_1[37463] = 32'b11111111111111111011001100100101;
assign LUT_1[37464] = 32'b11111111111111111101100000110110;
assign LUT_1[37465] = 32'b11111111111111110110110010110010;
assign LUT_1[37466] = 32'b11111111111111111001001111000111;
assign LUT_1[37467] = 32'b11111111111111110010100001000011;
assign LUT_1[37468] = 32'b00000000000000000101011010001101;
assign LUT_1[37469] = 32'b11111111111111111110101100001001;
assign LUT_1[37470] = 32'b00000000000000000001001000011110;
assign LUT_1[37471] = 32'b11111111111111111010011010011010;
assign LUT_1[37472] = 32'b11111111111111111101010010011110;
assign LUT_1[37473] = 32'b11111111111111110110100100011010;
assign LUT_1[37474] = 32'b11111111111111111001000000101111;
assign LUT_1[37475] = 32'b11111111111111110010010010101011;
assign LUT_1[37476] = 32'b00000000000000000101001011110101;
assign LUT_1[37477] = 32'b11111111111111111110011101110001;
assign LUT_1[37478] = 32'b00000000000000000000111010000110;
assign LUT_1[37479] = 32'b11111111111111111010001100000010;
assign LUT_1[37480] = 32'b11111111111111111100100000010011;
assign LUT_1[37481] = 32'b11111111111111110101110010001111;
assign LUT_1[37482] = 32'b11111111111111111000001110100100;
assign LUT_1[37483] = 32'b11111111111111110001100000100000;
assign LUT_1[37484] = 32'b00000000000000000100011001101010;
assign LUT_1[37485] = 32'b11111111111111111101101011100110;
assign LUT_1[37486] = 32'b00000000000000000000000111111011;
assign LUT_1[37487] = 32'b11111111111111111001011001110111;
assign LUT_1[37488] = 32'b11111111111111111111001110000000;
assign LUT_1[37489] = 32'b11111111111111111000011111111100;
assign LUT_1[37490] = 32'b11111111111111111010111100010001;
assign LUT_1[37491] = 32'b11111111111111110100001110001101;
assign LUT_1[37492] = 32'b00000000000000000111000111010111;
assign LUT_1[37493] = 32'b00000000000000000000011001010011;
assign LUT_1[37494] = 32'b00000000000000000010110101101000;
assign LUT_1[37495] = 32'b11111111111111111100000111100100;
assign LUT_1[37496] = 32'b11111111111111111110011011110101;
assign LUT_1[37497] = 32'b11111111111111110111101101110001;
assign LUT_1[37498] = 32'b11111111111111111010001010000110;
assign LUT_1[37499] = 32'b11111111111111110011011100000010;
assign LUT_1[37500] = 32'b00000000000000000110010101001100;
assign LUT_1[37501] = 32'b11111111111111111111100111001000;
assign LUT_1[37502] = 32'b00000000000000000010000011011101;
assign LUT_1[37503] = 32'b11111111111111111011010101011001;
assign LUT_1[37504] = 32'b11111111111111111101011001111010;
assign LUT_1[37505] = 32'b11111111111111110110101011110110;
assign LUT_1[37506] = 32'b11111111111111111001001000001011;
assign LUT_1[37507] = 32'b11111111111111110010011010000111;
assign LUT_1[37508] = 32'b00000000000000000101010011010001;
assign LUT_1[37509] = 32'b11111111111111111110100101001101;
assign LUT_1[37510] = 32'b00000000000000000001000001100010;
assign LUT_1[37511] = 32'b11111111111111111010010011011110;
assign LUT_1[37512] = 32'b11111111111111111100100111101111;
assign LUT_1[37513] = 32'b11111111111111110101111001101011;
assign LUT_1[37514] = 32'b11111111111111111000010110000000;
assign LUT_1[37515] = 32'b11111111111111110001100111111100;
assign LUT_1[37516] = 32'b00000000000000000100100001000110;
assign LUT_1[37517] = 32'b11111111111111111101110011000010;
assign LUT_1[37518] = 32'b00000000000000000000001111010111;
assign LUT_1[37519] = 32'b11111111111111111001100001010011;
assign LUT_1[37520] = 32'b11111111111111111111010101011100;
assign LUT_1[37521] = 32'b11111111111111111000100111011000;
assign LUT_1[37522] = 32'b11111111111111111011000011101101;
assign LUT_1[37523] = 32'b11111111111111110100010101101001;
assign LUT_1[37524] = 32'b00000000000000000111001110110011;
assign LUT_1[37525] = 32'b00000000000000000000100000101111;
assign LUT_1[37526] = 32'b00000000000000000010111101000100;
assign LUT_1[37527] = 32'b11111111111111111100001111000000;
assign LUT_1[37528] = 32'b11111111111111111110100011010001;
assign LUT_1[37529] = 32'b11111111111111110111110101001101;
assign LUT_1[37530] = 32'b11111111111111111010010001100010;
assign LUT_1[37531] = 32'b11111111111111110011100011011110;
assign LUT_1[37532] = 32'b00000000000000000110011100101000;
assign LUT_1[37533] = 32'b11111111111111111111101110100100;
assign LUT_1[37534] = 32'b00000000000000000010001010111001;
assign LUT_1[37535] = 32'b11111111111111111011011100110101;
assign LUT_1[37536] = 32'b11111111111111111110010100111001;
assign LUT_1[37537] = 32'b11111111111111110111100110110101;
assign LUT_1[37538] = 32'b11111111111111111010000011001010;
assign LUT_1[37539] = 32'b11111111111111110011010101000110;
assign LUT_1[37540] = 32'b00000000000000000110001110010000;
assign LUT_1[37541] = 32'b11111111111111111111100000001100;
assign LUT_1[37542] = 32'b00000000000000000001111100100001;
assign LUT_1[37543] = 32'b11111111111111111011001110011101;
assign LUT_1[37544] = 32'b11111111111111111101100010101110;
assign LUT_1[37545] = 32'b11111111111111110110110100101010;
assign LUT_1[37546] = 32'b11111111111111111001010000111111;
assign LUT_1[37547] = 32'b11111111111111110010100010111011;
assign LUT_1[37548] = 32'b00000000000000000101011100000101;
assign LUT_1[37549] = 32'b11111111111111111110101110000001;
assign LUT_1[37550] = 32'b00000000000000000001001010010110;
assign LUT_1[37551] = 32'b11111111111111111010011100010010;
assign LUT_1[37552] = 32'b00000000000000000000010000011011;
assign LUT_1[37553] = 32'b11111111111111111001100010010111;
assign LUT_1[37554] = 32'b11111111111111111011111110101100;
assign LUT_1[37555] = 32'b11111111111111110101010000101000;
assign LUT_1[37556] = 32'b00000000000000001000001001110010;
assign LUT_1[37557] = 32'b00000000000000000001011011101110;
assign LUT_1[37558] = 32'b00000000000000000011111000000011;
assign LUT_1[37559] = 32'b11111111111111111101001001111111;
assign LUT_1[37560] = 32'b11111111111111111111011110010000;
assign LUT_1[37561] = 32'b11111111111111111000110000001100;
assign LUT_1[37562] = 32'b11111111111111111011001100100001;
assign LUT_1[37563] = 32'b11111111111111110100011110011101;
assign LUT_1[37564] = 32'b00000000000000000111010111100111;
assign LUT_1[37565] = 32'b00000000000000000000101001100011;
assign LUT_1[37566] = 32'b00000000000000000011000101111000;
assign LUT_1[37567] = 32'b11111111111111111100010111110100;
assign LUT_1[37568] = 32'b11111111111111111111010111100010;
assign LUT_1[37569] = 32'b11111111111111111000101001011110;
assign LUT_1[37570] = 32'b11111111111111111011000101110011;
assign LUT_1[37571] = 32'b11111111111111110100010111101111;
assign LUT_1[37572] = 32'b00000000000000000111010000111001;
assign LUT_1[37573] = 32'b00000000000000000000100010110101;
assign LUT_1[37574] = 32'b00000000000000000010111111001010;
assign LUT_1[37575] = 32'b11111111111111111100010001000110;
assign LUT_1[37576] = 32'b11111111111111111110100101010111;
assign LUT_1[37577] = 32'b11111111111111110111110111010011;
assign LUT_1[37578] = 32'b11111111111111111010010011101000;
assign LUT_1[37579] = 32'b11111111111111110011100101100100;
assign LUT_1[37580] = 32'b00000000000000000110011110101110;
assign LUT_1[37581] = 32'b11111111111111111111110000101010;
assign LUT_1[37582] = 32'b00000000000000000010001100111111;
assign LUT_1[37583] = 32'b11111111111111111011011110111011;
assign LUT_1[37584] = 32'b00000000000000000001010011000100;
assign LUT_1[37585] = 32'b11111111111111111010100101000000;
assign LUT_1[37586] = 32'b11111111111111111101000001010101;
assign LUT_1[37587] = 32'b11111111111111110110010011010001;
assign LUT_1[37588] = 32'b00000000000000001001001100011011;
assign LUT_1[37589] = 32'b00000000000000000010011110010111;
assign LUT_1[37590] = 32'b00000000000000000100111010101100;
assign LUT_1[37591] = 32'b11111111111111111110001100101000;
assign LUT_1[37592] = 32'b00000000000000000000100000111001;
assign LUT_1[37593] = 32'b11111111111111111001110010110101;
assign LUT_1[37594] = 32'b11111111111111111100001111001010;
assign LUT_1[37595] = 32'b11111111111111110101100001000110;
assign LUT_1[37596] = 32'b00000000000000001000011010010000;
assign LUT_1[37597] = 32'b00000000000000000001101100001100;
assign LUT_1[37598] = 32'b00000000000000000100001000100001;
assign LUT_1[37599] = 32'b11111111111111111101011010011101;
assign LUT_1[37600] = 32'b00000000000000000000010010100001;
assign LUT_1[37601] = 32'b11111111111111111001100100011101;
assign LUT_1[37602] = 32'b11111111111111111100000000110010;
assign LUT_1[37603] = 32'b11111111111111110101010010101110;
assign LUT_1[37604] = 32'b00000000000000001000001011111000;
assign LUT_1[37605] = 32'b00000000000000000001011101110100;
assign LUT_1[37606] = 32'b00000000000000000011111010001001;
assign LUT_1[37607] = 32'b11111111111111111101001100000101;
assign LUT_1[37608] = 32'b11111111111111111111100000010110;
assign LUT_1[37609] = 32'b11111111111111111000110010010010;
assign LUT_1[37610] = 32'b11111111111111111011001110100111;
assign LUT_1[37611] = 32'b11111111111111110100100000100011;
assign LUT_1[37612] = 32'b00000000000000000111011001101101;
assign LUT_1[37613] = 32'b00000000000000000000101011101001;
assign LUT_1[37614] = 32'b00000000000000000011000111111110;
assign LUT_1[37615] = 32'b11111111111111111100011001111010;
assign LUT_1[37616] = 32'b00000000000000000010001110000011;
assign LUT_1[37617] = 32'b11111111111111111011011111111111;
assign LUT_1[37618] = 32'b11111111111111111101111100010100;
assign LUT_1[37619] = 32'b11111111111111110111001110010000;
assign LUT_1[37620] = 32'b00000000000000001010000111011010;
assign LUT_1[37621] = 32'b00000000000000000011011001010110;
assign LUT_1[37622] = 32'b00000000000000000101110101101011;
assign LUT_1[37623] = 32'b11111111111111111111000111100111;
assign LUT_1[37624] = 32'b00000000000000000001011011111000;
assign LUT_1[37625] = 32'b11111111111111111010101101110100;
assign LUT_1[37626] = 32'b11111111111111111101001010001001;
assign LUT_1[37627] = 32'b11111111111111110110011100000101;
assign LUT_1[37628] = 32'b00000000000000001001010101001111;
assign LUT_1[37629] = 32'b00000000000000000010100111001011;
assign LUT_1[37630] = 32'b00000000000000000101000011100000;
assign LUT_1[37631] = 32'b11111111111111111110010101011100;
assign LUT_1[37632] = 32'b11111111111111111000001110000011;
assign LUT_1[37633] = 32'b11111111111111110001011111111111;
assign LUT_1[37634] = 32'b11111111111111110011111100010100;
assign LUT_1[37635] = 32'b11111111111111101101001110010000;
assign LUT_1[37636] = 32'b00000000000000000000000111011010;
assign LUT_1[37637] = 32'b11111111111111111001011001010110;
assign LUT_1[37638] = 32'b11111111111111111011110101101011;
assign LUT_1[37639] = 32'b11111111111111110101000111100111;
assign LUT_1[37640] = 32'b11111111111111110111011011111000;
assign LUT_1[37641] = 32'b11111111111111110000101101110100;
assign LUT_1[37642] = 32'b11111111111111110011001010001001;
assign LUT_1[37643] = 32'b11111111111111101100011100000101;
assign LUT_1[37644] = 32'b11111111111111111111010101001111;
assign LUT_1[37645] = 32'b11111111111111111000100111001011;
assign LUT_1[37646] = 32'b11111111111111111011000011100000;
assign LUT_1[37647] = 32'b11111111111111110100010101011100;
assign LUT_1[37648] = 32'b11111111111111111010001001100101;
assign LUT_1[37649] = 32'b11111111111111110011011011100001;
assign LUT_1[37650] = 32'b11111111111111110101110111110110;
assign LUT_1[37651] = 32'b11111111111111101111001001110010;
assign LUT_1[37652] = 32'b00000000000000000010000010111100;
assign LUT_1[37653] = 32'b11111111111111111011010100111000;
assign LUT_1[37654] = 32'b11111111111111111101110001001101;
assign LUT_1[37655] = 32'b11111111111111110111000011001001;
assign LUT_1[37656] = 32'b11111111111111111001010111011010;
assign LUT_1[37657] = 32'b11111111111111110010101001010110;
assign LUT_1[37658] = 32'b11111111111111110101000101101011;
assign LUT_1[37659] = 32'b11111111111111101110010111100111;
assign LUT_1[37660] = 32'b00000000000000000001010000110001;
assign LUT_1[37661] = 32'b11111111111111111010100010101101;
assign LUT_1[37662] = 32'b11111111111111111100111111000010;
assign LUT_1[37663] = 32'b11111111111111110110010000111110;
assign LUT_1[37664] = 32'b11111111111111111001001001000010;
assign LUT_1[37665] = 32'b11111111111111110010011010111110;
assign LUT_1[37666] = 32'b11111111111111110100110111010011;
assign LUT_1[37667] = 32'b11111111111111101110001001001111;
assign LUT_1[37668] = 32'b00000000000000000001000010011001;
assign LUT_1[37669] = 32'b11111111111111111010010100010101;
assign LUT_1[37670] = 32'b11111111111111111100110000101010;
assign LUT_1[37671] = 32'b11111111111111110110000010100110;
assign LUT_1[37672] = 32'b11111111111111111000010110110111;
assign LUT_1[37673] = 32'b11111111111111110001101000110011;
assign LUT_1[37674] = 32'b11111111111111110100000101001000;
assign LUT_1[37675] = 32'b11111111111111101101010111000100;
assign LUT_1[37676] = 32'b00000000000000000000010000001110;
assign LUT_1[37677] = 32'b11111111111111111001100010001010;
assign LUT_1[37678] = 32'b11111111111111111011111110011111;
assign LUT_1[37679] = 32'b11111111111111110101010000011011;
assign LUT_1[37680] = 32'b11111111111111111011000100100100;
assign LUT_1[37681] = 32'b11111111111111110100010110100000;
assign LUT_1[37682] = 32'b11111111111111110110110010110101;
assign LUT_1[37683] = 32'b11111111111111110000000100110001;
assign LUT_1[37684] = 32'b00000000000000000010111101111011;
assign LUT_1[37685] = 32'b11111111111111111100001111110111;
assign LUT_1[37686] = 32'b11111111111111111110101100001100;
assign LUT_1[37687] = 32'b11111111111111110111111110001000;
assign LUT_1[37688] = 32'b11111111111111111010010010011001;
assign LUT_1[37689] = 32'b11111111111111110011100100010101;
assign LUT_1[37690] = 32'b11111111111111110110000000101010;
assign LUT_1[37691] = 32'b11111111111111101111010010100110;
assign LUT_1[37692] = 32'b00000000000000000010001011110000;
assign LUT_1[37693] = 32'b11111111111111111011011101101100;
assign LUT_1[37694] = 32'b11111111111111111101111010000001;
assign LUT_1[37695] = 32'b11111111111111110111001011111101;
assign LUT_1[37696] = 32'b11111111111111111010001011101011;
assign LUT_1[37697] = 32'b11111111111111110011011101100111;
assign LUT_1[37698] = 32'b11111111111111110101111001111100;
assign LUT_1[37699] = 32'b11111111111111101111001011111000;
assign LUT_1[37700] = 32'b00000000000000000010000101000010;
assign LUT_1[37701] = 32'b11111111111111111011010110111110;
assign LUT_1[37702] = 32'b11111111111111111101110011010011;
assign LUT_1[37703] = 32'b11111111111111110111000101001111;
assign LUT_1[37704] = 32'b11111111111111111001011001100000;
assign LUT_1[37705] = 32'b11111111111111110010101011011100;
assign LUT_1[37706] = 32'b11111111111111110101000111110001;
assign LUT_1[37707] = 32'b11111111111111101110011001101101;
assign LUT_1[37708] = 32'b00000000000000000001010010110111;
assign LUT_1[37709] = 32'b11111111111111111010100100110011;
assign LUT_1[37710] = 32'b11111111111111111101000001001000;
assign LUT_1[37711] = 32'b11111111111111110110010011000100;
assign LUT_1[37712] = 32'b11111111111111111100000111001101;
assign LUT_1[37713] = 32'b11111111111111110101011001001001;
assign LUT_1[37714] = 32'b11111111111111110111110101011110;
assign LUT_1[37715] = 32'b11111111111111110001000111011010;
assign LUT_1[37716] = 32'b00000000000000000100000000100100;
assign LUT_1[37717] = 32'b11111111111111111101010010100000;
assign LUT_1[37718] = 32'b11111111111111111111101110110101;
assign LUT_1[37719] = 32'b11111111111111111001000000110001;
assign LUT_1[37720] = 32'b11111111111111111011010101000010;
assign LUT_1[37721] = 32'b11111111111111110100100110111110;
assign LUT_1[37722] = 32'b11111111111111110111000011010011;
assign LUT_1[37723] = 32'b11111111111111110000010101001111;
assign LUT_1[37724] = 32'b00000000000000000011001110011001;
assign LUT_1[37725] = 32'b11111111111111111100100000010101;
assign LUT_1[37726] = 32'b11111111111111111110111100101010;
assign LUT_1[37727] = 32'b11111111111111111000001110100110;
assign LUT_1[37728] = 32'b11111111111111111011000110101010;
assign LUT_1[37729] = 32'b11111111111111110100011000100110;
assign LUT_1[37730] = 32'b11111111111111110110110100111011;
assign LUT_1[37731] = 32'b11111111111111110000000110110111;
assign LUT_1[37732] = 32'b00000000000000000011000000000001;
assign LUT_1[37733] = 32'b11111111111111111100010001111101;
assign LUT_1[37734] = 32'b11111111111111111110101110010010;
assign LUT_1[37735] = 32'b11111111111111111000000000001110;
assign LUT_1[37736] = 32'b11111111111111111010010100011111;
assign LUT_1[37737] = 32'b11111111111111110011100110011011;
assign LUT_1[37738] = 32'b11111111111111110110000010110000;
assign LUT_1[37739] = 32'b11111111111111101111010100101100;
assign LUT_1[37740] = 32'b00000000000000000010001101110110;
assign LUT_1[37741] = 32'b11111111111111111011011111110010;
assign LUT_1[37742] = 32'b11111111111111111101111100000111;
assign LUT_1[37743] = 32'b11111111111111110111001110000011;
assign LUT_1[37744] = 32'b11111111111111111101000010001100;
assign LUT_1[37745] = 32'b11111111111111110110010100001000;
assign LUT_1[37746] = 32'b11111111111111111000110000011101;
assign LUT_1[37747] = 32'b11111111111111110010000010011001;
assign LUT_1[37748] = 32'b00000000000000000100111011100011;
assign LUT_1[37749] = 32'b11111111111111111110001101011111;
assign LUT_1[37750] = 32'b00000000000000000000101001110100;
assign LUT_1[37751] = 32'b11111111111111111001111011110000;
assign LUT_1[37752] = 32'b11111111111111111100010000000001;
assign LUT_1[37753] = 32'b11111111111111110101100001111101;
assign LUT_1[37754] = 32'b11111111111111110111111110010010;
assign LUT_1[37755] = 32'b11111111111111110001010000001110;
assign LUT_1[37756] = 32'b00000000000000000100001001011000;
assign LUT_1[37757] = 32'b11111111111111111101011011010100;
assign LUT_1[37758] = 32'b11111111111111111111110111101001;
assign LUT_1[37759] = 32'b11111111111111111001001001100101;
assign LUT_1[37760] = 32'b11111111111111111011001110000110;
assign LUT_1[37761] = 32'b11111111111111110100100000000010;
assign LUT_1[37762] = 32'b11111111111111110110111100010111;
assign LUT_1[37763] = 32'b11111111111111110000001110010011;
assign LUT_1[37764] = 32'b00000000000000000011000111011101;
assign LUT_1[37765] = 32'b11111111111111111100011001011001;
assign LUT_1[37766] = 32'b11111111111111111110110101101110;
assign LUT_1[37767] = 32'b11111111111111111000000111101010;
assign LUT_1[37768] = 32'b11111111111111111010011011111011;
assign LUT_1[37769] = 32'b11111111111111110011101101110111;
assign LUT_1[37770] = 32'b11111111111111110110001010001100;
assign LUT_1[37771] = 32'b11111111111111101111011100001000;
assign LUT_1[37772] = 32'b00000000000000000010010101010010;
assign LUT_1[37773] = 32'b11111111111111111011100111001110;
assign LUT_1[37774] = 32'b11111111111111111110000011100011;
assign LUT_1[37775] = 32'b11111111111111110111010101011111;
assign LUT_1[37776] = 32'b11111111111111111101001001101000;
assign LUT_1[37777] = 32'b11111111111111110110011011100100;
assign LUT_1[37778] = 32'b11111111111111111000110111111001;
assign LUT_1[37779] = 32'b11111111111111110010001001110101;
assign LUT_1[37780] = 32'b00000000000000000101000010111111;
assign LUT_1[37781] = 32'b11111111111111111110010100111011;
assign LUT_1[37782] = 32'b00000000000000000000110001010000;
assign LUT_1[37783] = 32'b11111111111111111010000011001100;
assign LUT_1[37784] = 32'b11111111111111111100010111011101;
assign LUT_1[37785] = 32'b11111111111111110101101001011001;
assign LUT_1[37786] = 32'b11111111111111111000000101101110;
assign LUT_1[37787] = 32'b11111111111111110001010111101010;
assign LUT_1[37788] = 32'b00000000000000000100010000110100;
assign LUT_1[37789] = 32'b11111111111111111101100010110000;
assign LUT_1[37790] = 32'b11111111111111111111111111000101;
assign LUT_1[37791] = 32'b11111111111111111001010001000001;
assign LUT_1[37792] = 32'b11111111111111111100001001000101;
assign LUT_1[37793] = 32'b11111111111111110101011011000001;
assign LUT_1[37794] = 32'b11111111111111110111110111010110;
assign LUT_1[37795] = 32'b11111111111111110001001001010010;
assign LUT_1[37796] = 32'b00000000000000000100000010011100;
assign LUT_1[37797] = 32'b11111111111111111101010100011000;
assign LUT_1[37798] = 32'b11111111111111111111110000101101;
assign LUT_1[37799] = 32'b11111111111111111001000010101001;
assign LUT_1[37800] = 32'b11111111111111111011010110111010;
assign LUT_1[37801] = 32'b11111111111111110100101000110110;
assign LUT_1[37802] = 32'b11111111111111110111000101001011;
assign LUT_1[37803] = 32'b11111111111111110000010111000111;
assign LUT_1[37804] = 32'b00000000000000000011010000010001;
assign LUT_1[37805] = 32'b11111111111111111100100010001101;
assign LUT_1[37806] = 32'b11111111111111111110111110100010;
assign LUT_1[37807] = 32'b11111111111111111000010000011110;
assign LUT_1[37808] = 32'b11111111111111111110000100100111;
assign LUT_1[37809] = 32'b11111111111111110111010110100011;
assign LUT_1[37810] = 32'b11111111111111111001110010111000;
assign LUT_1[37811] = 32'b11111111111111110011000100110100;
assign LUT_1[37812] = 32'b00000000000000000101111101111110;
assign LUT_1[37813] = 32'b11111111111111111111001111111010;
assign LUT_1[37814] = 32'b00000000000000000001101100001111;
assign LUT_1[37815] = 32'b11111111111111111010111110001011;
assign LUT_1[37816] = 32'b11111111111111111101010010011100;
assign LUT_1[37817] = 32'b11111111111111110110100100011000;
assign LUT_1[37818] = 32'b11111111111111111001000000101101;
assign LUT_1[37819] = 32'b11111111111111110010010010101001;
assign LUT_1[37820] = 32'b00000000000000000101001011110011;
assign LUT_1[37821] = 32'b11111111111111111110011101101111;
assign LUT_1[37822] = 32'b00000000000000000000111010000100;
assign LUT_1[37823] = 32'b11111111111111111010001100000000;
assign LUT_1[37824] = 32'b11111111111111111101001011101110;
assign LUT_1[37825] = 32'b11111111111111110110011101101010;
assign LUT_1[37826] = 32'b11111111111111111000111001111111;
assign LUT_1[37827] = 32'b11111111111111110010001011111011;
assign LUT_1[37828] = 32'b00000000000000000101000101000101;
assign LUT_1[37829] = 32'b11111111111111111110010111000001;
assign LUT_1[37830] = 32'b00000000000000000000110011010110;
assign LUT_1[37831] = 32'b11111111111111111010000101010010;
assign LUT_1[37832] = 32'b11111111111111111100011001100011;
assign LUT_1[37833] = 32'b11111111111111110101101011011111;
assign LUT_1[37834] = 32'b11111111111111111000000111110100;
assign LUT_1[37835] = 32'b11111111111111110001011001110000;
assign LUT_1[37836] = 32'b00000000000000000100010010111010;
assign LUT_1[37837] = 32'b11111111111111111101100100110110;
assign LUT_1[37838] = 32'b00000000000000000000000001001011;
assign LUT_1[37839] = 32'b11111111111111111001010011000111;
assign LUT_1[37840] = 32'b11111111111111111111000111010000;
assign LUT_1[37841] = 32'b11111111111111111000011001001100;
assign LUT_1[37842] = 32'b11111111111111111010110101100001;
assign LUT_1[37843] = 32'b11111111111111110100000111011101;
assign LUT_1[37844] = 32'b00000000000000000111000000100111;
assign LUT_1[37845] = 32'b00000000000000000000010010100011;
assign LUT_1[37846] = 32'b00000000000000000010101110111000;
assign LUT_1[37847] = 32'b11111111111111111100000000110100;
assign LUT_1[37848] = 32'b11111111111111111110010101000101;
assign LUT_1[37849] = 32'b11111111111111110111100111000001;
assign LUT_1[37850] = 32'b11111111111111111010000011010110;
assign LUT_1[37851] = 32'b11111111111111110011010101010010;
assign LUT_1[37852] = 32'b00000000000000000110001110011100;
assign LUT_1[37853] = 32'b11111111111111111111100000011000;
assign LUT_1[37854] = 32'b00000000000000000001111100101101;
assign LUT_1[37855] = 32'b11111111111111111011001110101001;
assign LUT_1[37856] = 32'b11111111111111111110000110101101;
assign LUT_1[37857] = 32'b11111111111111110111011000101001;
assign LUT_1[37858] = 32'b11111111111111111001110100111110;
assign LUT_1[37859] = 32'b11111111111111110011000110111010;
assign LUT_1[37860] = 32'b00000000000000000110000000000100;
assign LUT_1[37861] = 32'b11111111111111111111010010000000;
assign LUT_1[37862] = 32'b00000000000000000001101110010101;
assign LUT_1[37863] = 32'b11111111111111111011000000010001;
assign LUT_1[37864] = 32'b11111111111111111101010100100010;
assign LUT_1[37865] = 32'b11111111111111110110100110011110;
assign LUT_1[37866] = 32'b11111111111111111001000010110011;
assign LUT_1[37867] = 32'b11111111111111110010010100101111;
assign LUT_1[37868] = 32'b00000000000000000101001101111001;
assign LUT_1[37869] = 32'b11111111111111111110011111110101;
assign LUT_1[37870] = 32'b00000000000000000000111100001010;
assign LUT_1[37871] = 32'b11111111111111111010001110000110;
assign LUT_1[37872] = 32'b00000000000000000000000010001111;
assign LUT_1[37873] = 32'b11111111111111111001010100001011;
assign LUT_1[37874] = 32'b11111111111111111011110000100000;
assign LUT_1[37875] = 32'b11111111111111110101000010011100;
assign LUT_1[37876] = 32'b00000000000000000111111011100110;
assign LUT_1[37877] = 32'b00000000000000000001001101100010;
assign LUT_1[37878] = 32'b00000000000000000011101001110111;
assign LUT_1[37879] = 32'b11111111111111111100111011110011;
assign LUT_1[37880] = 32'b11111111111111111111010000000100;
assign LUT_1[37881] = 32'b11111111111111111000100010000000;
assign LUT_1[37882] = 32'b11111111111111111010111110010101;
assign LUT_1[37883] = 32'b11111111111111110100010000010001;
assign LUT_1[37884] = 32'b00000000000000000111001001011011;
assign LUT_1[37885] = 32'b00000000000000000000011011010111;
assign LUT_1[37886] = 32'b00000000000000000010110111101100;
assign LUT_1[37887] = 32'b11111111111111111100001001101000;
assign LUT_1[37888] = 32'b00000000000000000111000010001010;
assign LUT_1[37889] = 32'b00000000000000000000010100000110;
assign LUT_1[37890] = 32'b00000000000000000010110000011011;
assign LUT_1[37891] = 32'b11111111111111111100000010010111;
assign LUT_1[37892] = 32'b00000000000000001110111011100001;
assign LUT_1[37893] = 32'b00000000000000001000001101011101;
assign LUT_1[37894] = 32'b00000000000000001010101001110010;
assign LUT_1[37895] = 32'b00000000000000000011111011101110;
assign LUT_1[37896] = 32'b00000000000000000110001111111111;
assign LUT_1[37897] = 32'b11111111111111111111100001111011;
assign LUT_1[37898] = 32'b00000000000000000001111110010000;
assign LUT_1[37899] = 32'b11111111111111111011010000001100;
assign LUT_1[37900] = 32'b00000000000000001110001001010110;
assign LUT_1[37901] = 32'b00000000000000000111011011010010;
assign LUT_1[37902] = 32'b00000000000000001001110111100111;
assign LUT_1[37903] = 32'b00000000000000000011001001100011;
assign LUT_1[37904] = 32'b00000000000000001000111101101100;
assign LUT_1[37905] = 32'b00000000000000000010001111101000;
assign LUT_1[37906] = 32'b00000000000000000100101011111101;
assign LUT_1[37907] = 32'b11111111111111111101111101111001;
assign LUT_1[37908] = 32'b00000000000000010000110111000011;
assign LUT_1[37909] = 32'b00000000000000001010001000111111;
assign LUT_1[37910] = 32'b00000000000000001100100101010100;
assign LUT_1[37911] = 32'b00000000000000000101110111010000;
assign LUT_1[37912] = 32'b00000000000000001000001011100001;
assign LUT_1[37913] = 32'b00000000000000000001011101011101;
assign LUT_1[37914] = 32'b00000000000000000011111001110010;
assign LUT_1[37915] = 32'b11111111111111111101001011101110;
assign LUT_1[37916] = 32'b00000000000000010000000100111000;
assign LUT_1[37917] = 32'b00000000000000001001010110110100;
assign LUT_1[37918] = 32'b00000000000000001011110011001001;
assign LUT_1[37919] = 32'b00000000000000000101000101000101;
assign LUT_1[37920] = 32'b00000000000000000111111101001001;
assign LUT_1[37921] = 32'b00000000000000000001001111000101;
assign LUT_1[37922] = 32'b00000000000000000011101011011010;
assign LUT_1[37923] = 32'b11111111111111111100111101010110;
assign LUT_1[37924] = 32'b00000000000000001111110110100000;
assign LUT_1[37925] = 32'b00000000000000001001001000011100;
assign LUT_1[37926] = 32'b00000000000000001011100100110001;
assign LUT_1[37927] = 32'b00000000000000000100110110101101;
assign LUT_1[37928] = 32'b00000000000000000111001010111110;
assign LUT_1[37929] = 32'b00000000000000000000011100111010;
assign LUT_1[37930] = 32'b00000000000000000010111001001111;
assign LUT_1[37931] = 32'b11111111111111111100001011001011;
assign LUT_1[37932] = 32'b00000000000000001111000100010101;
assign LUT_1[37933] = 32'b00000000000000001000010110010001;
assign LUT_1[37934] = 32'b00000000000000001010110010100110;
assign LUT_1[37935] = 32'b00000000000000000100000100100010;
assign LUT_1[37936] = 32'b00000000000000001001111000101011;
assign LUT_1[37937] = 32'b00000000000000000011001010100111;
assign LUT_1[37938] = 32'b00000000000000000101100110111100;
assign LUT_1[37939] = 32'b11111111111111111110111000111000;
assign LUT_1[37940] = 32'b00000000000000010001110010000010;
assign LUT_1[37941] = 32'b00000000000000001011000011111110;
assign LUT_1[37942] = 32'b00000000000000001101100000010011;
assign LUT_1[37943] = 32'b00000000000000000110110010001111;
assign LUT_1[37944] = 32'b00000000000000001001000110100000;
assign LUT_1[37945] = 32'b00000000000000000010011000011100;
assign LUT_1[37946] = 32'b00000000000000000100110100110001;
assign LUT_1[37947] = 32'b11111111111111111110000110101101;
assign LUT_1[37948] = 32'b00000000000000010000111111110111;
assign LUT_1[37949] = 32'b00000000000000001010010001110011;
assign LUT_1[37950] = 32'b00000000000000001100101110001000;
assign LUT_1[37951] = 32'b00000000000000000110000000000100;
assign LUT_1[37952] = 32'b00000000000000001000111111110010;
assign LUT_1[37953] = 32'b00000000000000000010010001101110;
assign LUT_1[37954] = 32'b00000000000000000100101110000011;
assign LUT_1[37955] = 32'b11111111111111111101111111111111;
assign LUT_1[37956] = 32'b00000000000000010000111001001001;
assign LUT_1[37957] = 32'b00000000000000001010001011000101;
assign LUT_1[37958] = 32'b00000000000000001100100111011010;
assign LUT_1[37959] = 32'b00000000000000000101111001010110;
assign LUT_1[37960] = 32'b00000000000000001000001101100111;
assign LUT_1[37961] = 32'b00000000000000000001011111100011;
assign LUT_1[37962] = 32'b00000000000000000011111011111000;
assign LUT_1[37963] = 32'b11111111111111111101001101110100;
assign LUT_1[37964] = 32'b00000000000000010000000110111110;
assign LUT_1[37965] = 32'b00000000000000001001011000111010;
assign LUT_1[37966] = 32'b00000000000000001011110101001111;
assign LUT_1[37967] = 32'b00000000000000000101000111001011;
assign LUT_1[37968] = 32'b00000000000000001010111011010100;
assign LUT_1[37969] = 32'b00000000000000000100001101010000;
assign LUT_1[37970] = 32'b00000000000000000110101001100101;
assign LUT_1[37971] = 32'b11111111111111111111111011100001;
assign LUT_1[37972] = 32'b00000000000000010010110100101011;
assign LUT_1[37973] = 32'b00000000000000001100000110100111;
assign LUT_1[37974] = 32'b00000000000000001110100010111100;
assign LUT_1[37975] = 32'b00000000000000000111110100111000;
assign LUT_1[37976] = 32'b00000000000000001010001001001001;
assign LUT_1[37977] = 32'b00000000000000000011011011000101;
assign LUT_1[37978] = 32'b00000000000000000101110111011010;
assign LUT_1[37979] = 32'b11111111111111111111001001010110;
assign LUT_1[37980] = 32'b00000000000000010010000010100000;
assign LUT_1[37981] = 32'b00000000000000001011010100011100;
assign LUT_1[37982] = 32'b00000000000000001101110000110001;
assign LUT_1[37983] = 32'b00000000000000000111000010101101;
assign LUT_1[37984] = 32'b00000000000000001001111010110001;
assign LUT_1[37985] = 32'b00000000000000000011001100101101;
assign LUT_1[37986] = 32'b00000000000000000101101001000010;
assign LUT_1[37987] = 32'b11111111111111111110111010111110;
assign LUT_1[37988] = 32'b00000000000000010001110100001000;
assign LUT_1[37989] = 32'b00000000000000001011000110000100;
assign LUT_1[37990] = 32'b00000000000000001101100010011001;
assign LUT_1[37991] = 32'b00000000000000000110110100010101;
assign LUT_1[37992] = 32'b00000000000000001001001000100110;
assign LUT_1[37993] = 32'b00000000000000000010011010100010;
assign LUT_1[37994] = 32'b00000000000000000100110110110111;
assign LUT_1[37995] = 32'b11111111111111111110001000110011;
assign LUT_1[37996] = 32'b00000000000000010001000001111101;
assign LUT_1[37997] = 32'b00000000000000001010010011111001;
assign LUT_1[37998] = 32'b00000000000000001100110000001110;
assign LUT_1[37999] = 32'b00000000000000000110000010001010;
assign LUT_1[38000] = 32'b00000000000000001011110110010011;
assign LUT_1[38001] = 32'b00000000000000000101001000001111;
assign LUT_1[38002] = 32'b00000000000000000111100100100100;
assign LUT_1[38003] = 32'b00000000000000000000110110100000;
assign LUT_1[38004] = 32'b00000000000000010011101111101010;
assign LUT_1[38005] = 32'b00000000000000001101000001100110;
assign LUT_1[38006] = 32'b00000000000000001111011101111011;
assign LUT_1[38007] = 32'b00000000000000001000101111110111;
assign LUT_1[38008] = 32'b00000000000000001011000100001000;
assign LUT_1[38009] = 32'b00000000000000000100010110000100;
assign LUT_1[38010] = 32'b00000000000000000110110010011001;
assign LUT_1[38011] = 32'b00000000000000000000000100010101;
assign LUT_1[38012] = 32'b00000000000000010010111101011111;
assign LUT_1[38013] = 32'b00000000000000001100001111011011;
assign LUT_1[38014] = 32'b00000000000000001110101011110000;
assign LUT_1[38015] = 32'b00000000000000000111111101101100;
assign LUT_1[38016] = 32'b00000000000000001010000010001101;
assign LUT_1[38017] = 32'b00000000000000000011010100001001;
assign LUT_1[38018] = 32'b00000000000000000101110000011110;
assign LUT_1[38019] = 32'b11111111111111111111000010011010;
assign LUT_1[38020] = 32'b00000000000000010001111011100100;
assign LUT_1[38021] = 32'b00000000000000001011001101100000;
assign LUT_1[38022] = 32'b00000000000000001101101001110101;
assign LUT_1[38023] = 32'b00000000000000000110111011110001;
assign LUT_1[38024] = 32'b00000000000000001001010000000010;
assign LUT_1[38025] = 32'b00000000000000000010100001111110;
assign LUT_1[38026] = 32'b00000000000000000100111110010011;
assign LUT_1[38027] = 32'b11111111111111111110010000001111;
assign LUT_1[38028] = 32'b00000000000000010001001001011001;
assign LUT_1[38029] = 32'b00000000000000001010011011010101;
assign LUT_1[38030] = 32'b00000000000000001100110111101010;
assign LUT_1[38031] = 32'b00000000000000000110001001100110;
assign LUT_1[38032] = 32'b00000000000000001011111101101111;
assign LUT_1[38033] = 32'b00000000000000000101001111101011;
assign LUT_1[38034] = 32'b00000000000000000111101100000000;
assign LUT_1[38035] = 32'b00000000000000000000111101111100;
assign LUT_1[38036] = 32'b00000000000000010011110111000110;
assign LUT_1[38037] = 32'b00000000000000001101001001000010;
assign LUT_1[38038] = 32'b00000000000000001111100101010111;
assign LUT_1[38039] = 32'b00000000000000001000110111010011;
assign LUT_1[38040] = 32'b00000000000000001011001011100100;
assign LUT_1[38041] = 32'b00000000000000000100011101100000;
assign LUT_1[38042] = 32'b00000000000000000110111001110101;
assign LUT_1[38043] = 32'b00000000000000000000001011110001;
assign LUT_1[38044] = 32'b00000000000000010011000100111011;
assign LUT_1[38045] = 32'b00000000000000001100010110110111;
assign LUT_1[38046] = 32'b00000000000000001110110011001100;
assign LUT_1[38047] = 32'b00000000000000001000000101001000;
assign LUT_1[38048] = 32'b00000000000000001010111101001100;
assign LUT_1[38049] = 32'b00000000000000000100001111001000;
assign LUT_1[38050] = 32'b00000000000000000110101011011101;
assign LUT_1[38051] = 32'b11111111111111111111111101011001;
assign LUT_1[38052] = 32'b00000000000000010010110110100011;
assign LUT_1[38053] = 32'b00000000000000001100001000011111;
assign LUT_1[38054] = 32'b00000000000000001110100100110100;
assign LUT_1[38055] = 32'b00000000000000000111110110110000;
assign LUT_1[38056] = 32'b00000000000000001010001011000001;
assign LUT_1[38057] = 32'b00000000000000000011011100111101;
assign LUT_1[38058] = 32'b00000000000000000101111001010010;
assign LUT_1[38059] = 32'b11111111111111111111001011001110;
assign LUT_1[38060] = 32'b00000000000000010010000100011000;
assign LUT_1[38061] = 32'b00000000000000001011010110010100;
assign LUT_1[38062] = 32'b00000000000000001101110010101001;
assign LUT_1[38063] = 32'b00000000000000000111000100100101;
assign LUT_1[38064] = 32'b00000000000000001100111000101110;
assign LUT_1[38065] = 32'b00000000000000000110001010101010;
assign LUT_1[38066] = 32'b00000000000000001000100110111111;
assign LUT_1[38067] = 32'b00000000000000000001111000111011;
assign LUT_1[38068] = 32'b00000000000000010100110010000101;
assign LUT_1[38069] = 32'b00000000000000001110000100000001;
assign LUT_1[38070] = 32'b00000000000000010000100000010110;
assign LUT_1[38071] = 32'b00000000000000001001110010010010;
assign LUT_1[38072] = 32'b00000000000000001100000110100011;
assign LUT_1[38073] = 32'b00000000000000000101011000011111;
assign LUT_1[38074] = 32'b00000000000000000111110100110100;
assign LUT_1[38075] = 32'b00000000000000000001000110110000;
assign LUT_1[38076] = 32'b00000000000000010011111111111010;
assign LUT_1[38077] = 32'b00000000000000001101010001110110;
assign LUT_1[38078] = 32'b00000000000000001111101110001011;
assign LUT_1[38079] = 32'b00000000000000001001000000000111;
assign LUT_1[38080] = 32'b00000000000000001011111111110101;
assign LUT_1[38081] = 32'b00000000000000000101010001110001;
assign LUT_1[38082] = 32'b00000000000000000111101110000110;
assign LUT_1[38083] = 32'b00000000000000000001000000000010;
assign LUT_1[38084] = 32'b00000000000000010011111001001100;
assign LUT_1[38085] = 32'b00000000000000001101001011001000;
assign LUT_1[38086] = 32'b00000000000000001111100111011101;
assign LUT_1[38087] = 32'b00000000000000001000111001011001;
assign LUT_1[38088] = 32'b00000000000000001011001101101010;
assign LUT_1[38089] = 32'b00000000000000000100011111100110;
assign LUT_1[38090] = 32'b00000000000000000110111011111011;
assign LUT_1[38091] = 32'b00000000000000000000001101110111;
assign LUT_1[38092] = 32'b00000000000000010011000111000001;
assign LUT_1[38093] = 32'b00000000000000001100011000111101;
assign LUT_1[38094] = 32'b00000000000000001110110101010010;
assign LUT_1[38095] = 32'b00000000000000001000000111001110;
assign LUT_1[38096] = 32'b00000000000000001101111011010111;
assign LUT_1[38097] = 32'b00000000000000000111001101010011;
assign LUT_1[38098] = 32'b00000000000000001001101001101000;
assign LUT_1[38099] = 32'b00000000000000000010111011100100;
assign LUT_1[38100] = 32'b00000000000000010101110100101110;
assign LUT_1[38101] = 32'b00000000000000001111000110101010;
assign LUT_1[38102] = 32'b00000000000000010001100010111111;
assign LUT_1[38103] = 32'b00000000000000001010110100111011;
assign LUT_1[38104] = 32'b00000000000000001101001001001100;
assign LUT_1[38105] = 32'b00000000000000000110011011001000;
assign LUT_1[38106] = 32'b00000000000000001000110111011101;
assign LUT_1[38107] = 32'b00000000000000000010001001011001;
assign LUT_1[38108] = 32'b00000000000000010101000010100011;
assign LUT_1[38109] = 32'b00000000000000001110010100011111;
assign LUT_1[38110] = 32'b00000000000000010000110000110100;
assign LUT_1[38111] = 32'b00000000000000001010000010110000;
assign LUT_1[38112] = 32'b00000000000000001100111010110100;
assign LUT_1[38113] = 32'b00000000000000000110001100110000;
assign LUT_1[38114] = 32'b00000000000000001000101001000101;
assign LUT_1[38115] = 32'b00000000000000000001111011000001;
assign LUT_1[38116] = 32'b00000000000000010100110100001011;
assign LUT_1[38117] = 32'b00000000000000001110000110000111;
assign LUT_1[38118] = 32'b00000000000000010000100010011100;
assign LUT_1[38119] = 32'b00000000000000001001110100011000;
assign LUT_1[38120] = 32'b00000000000000001100001000101001;
assign LUT_1[38121] = 32'b00000000000000000101011010100101;
assign LUT_1[38122] = 32'b00000000000000000111110110111010;
assign LUT_1[38123] = 32'b00000000000000000001001000110110;
assign LUT_1[38124] = 32'b00000000000000010100000010000000;
assign LUT_1[38125] = 32'b00000000000000001101010011111100;
assign LUT_1[38126] = 32'b00000000000000001111110000010001;
assign LUT_1[38127] = 32'b00000000000000001001000010001101;
assign LUT_1[38128] = 32'b00000000000000001110110110010110;
assign LUT_1[38129] = 32'b00000000000000001000001000010010;
assign LUT_1[38130] = 32'b00000000000000001010100100100111;
assign LUT_1[38131] = 32'b00000000000000000011110110100011;
assign LUT_1[38132] = 32'b00000000000000010110101111101101;
assign LUT_1[38133] = 32'b00000000000000010000000001101001;
assign LUT_1[38134] = 32'b00000000000000010010011101111110;
assign LUT_1[38135] = 32'b00000000000000001011101111111010;
assign LUT_1[38136] = 32'b00000000000000001110000100001011;
assign LUT_1[38137] = 32'b00000000000000000111010110000111;
assign LUT_1[38138] = 32'b00000000000000001001110010011100;
assign LUT_1[38139] = 32'b00000000000000000011000100011000;
assign LUT_1[38140] = 32'b00000000000000010101111101100010;
assign LUT_1[38141] = 32'b00000000000000001111001111011110;
assign LUT_1[38142] = 32'b00000000000000010001101011110011;
assign LUT_1[38143] = 32'b00000000000000001010111101101111;
assign LUT_1[38144] = 32'b00000000000000000100110110010110;
assign LUT_1[38145] = 32'b11111111111111111110001000010010;
assign LUT_1[38146] = 32'b00000000000000000000100100100111;
assign LUT_1[38147] = 32'b11111111111111111001110110100011;
assign LUT_1[38148] = 32'b00000000000000001100101111101101;
assign LUT_1[38149] = 32'b00000000000000000110000001101001;
assign LUT_1[38150] = 32'b00000000000000001000011101111110;
assign LUT_1[38151] = 32'b00000000000000000001101111111010;
assign LUT_1[38152] = 32'b00000000000000000100000100001011;
assign LUT_1[38153] = 32'b11111111111111111101010110000111;
assign LUT_1[38154] = 32'b11111111111111111111110010011100;
assign LUT_1[38155] = 32'b11111111111111111001000100011000;
assign LUT_1[38156] = 32'b00000000000000001011111101100010;
assign LUT_1[38157] = 32'b00000000000000000101001111011110;
assign LUT_1[38158] = 32'b00000000000000000111101011110011;
assign LUT_1[38159] = 32'b00000000000000000000111101101111;
assign LUT_1[38160] = 32'b00000000000000000110110001111000;
assign LUT_1[38161] = 32'b00000000000000000000000011110100;
assign LUT_1[38162] = 32'b00000000000000000010100000001001;
assign LUT_1[38163] = 32'b11111111111111111011110010000101;
assign LUT_1[38164] = 32'b00000000000000001110101011001111;
assign LUT_1[38165] = 32'b00000000000000000111111101001011;
assign LUT_1[38166] = 32'b00000000000000001010011001100000;
assign LUT_1[38167] = 32'b00000000000000000011101011011100;
assign LUT_1[38168] = 32'b00000000000000000101111111101101;
assign LUT_1[38169] = 32'b11111111111111111111010001101001;
assign LUT_1[38170] = 32'b00000000000000000001101101111110;
assign LUT_1[38171] = 32'b11111111111111111010111111111010;
assign LUT_1[38172] = 32'b00000000000000001101111001000100;
assign LUT_1[38173] = 32'b00000000000000000111001011000000;
assign LUT_1[38174] = 32'b00000000000000001001100111010101;
assign LUT_1[38175] = 32'b00000000000000000010111001010001;
assign LUT_1[38176] = 32'b00000000000000000101110001010101;
assign LUT_1[38177] = 32'b11111111111111111111000011010001;
assign LUT_1[38178] = 32'b00000000000000000001011111100110;
assign LUT_1[38179] = 32'b11111111111111111010110001100010;
assign LUT_1[38180] = 32'b00000000000000001101101010101100;
assign LUT_1[38181] = 32'b00000000000000000110111100101000;
assign LUT_1[38182] = 32'b00000000000000001001011000111101;
assign LUT_1[38183] = 32'b00000000000000000010101010111001;
assign LUT_1[38184] = 32'b00000000000000000100111111001010;
assign LUT_1[38185] = 32'b11111111111111111110010001000110;
assign LUT_1[38186] = 32'b00000000000000000000101101011011;
assign LUT_1[38187] = 32'b11111111111111111001111111010111;
assign LUT_1[38188] = 32'b00000000000000001100111000100001;
assign LUT_1[38189] = 32'b00000000000000000110001010011101;
assign LUT_1[38190] = 32'b00000000000000001000100110110010;
assign LUT_1[38191] = 32'b00000000000000000001111000101110;
assign LUT_1[38192] = 32'b00000000000000000111101100110111;
assign LUT_1[38193] = 32'b00000000000000000000111110110011;
assign LUT_1[38194] = 32'b00000000000000000011011011001000;
assign LUT_1[38195] = 32'b11111111111111111100101101000100;
assign LUT_1[38196] = 32'b00000000000000001111100110001110;
assign LUT_1[38197] = 32'b00000000000000001000111000001010;
assign LUT_1[38198] = 32'b00000000000000001011010100011111;
assign LUT_1[38199] = 32'b00000000000000000100100110011011;
assign LUT_1[38200] = 32'b00000000000000000110111010101100;
assign LUT_1[38201] = 32'b00000000000000000000001100101000;
assign LUT_1[38202] = 32'b00000000000000000010101000111101;
assign LUT_1[38203] = 32'b11111111111111111011111010111001;
assign LUT_1[38204] = 32'b00000000000000001110110100000011;
assign LUT_1[38205] = 32'b00000000000000001000000101111111;
assign LUT_1[38206] = 32'b00000000000000001010100010010100;
assign LUT_1[38207] = 32'b00000000000000000011110100010000;
assign LUT_1[38208] = 32'b00000000000000000110110011111110;
assign LUT_1[38209] = 32'b00000000000000000000000101111010;
assign LUT_1[38210] = 32'b00000000000000000010100010001111;
assign LUT_1[38211] = 32'b11111111111111111011110100001011;
assign LUT_1[38212] = 32'b00000000000000001110101101010101;
assign LUT_1[38213] = 32'b00000000000000000111111111010001;
assign LUT_1[38214] = 32'b00000000000000001010011011100110;
assign LUT_1[38215] = 32'b00000000000000000011101101100010;
assign LUT_1[38216] = 32'b00000000000000000110000001110011;
assign LUT_1[38217] = 32'b11111111111111111111010011101111;
assign LUT_1[38218] = 32'b00000000000000000001110000000100;
assign LUT_1[38219] = 32'b11111111111111111011000010000000;
assign LUT_1[38220] = 32'b00000000000000001101111011001010;
assign LUT_1[38221] = 32'b00000000000000000111001101000110;
assign LUT_1[38222] = 32'b00000000000000001001101001011011;
assign LUT_1[38223] = 32'b00000000000000000010111011010111;
assign LUT_1[38224] = 32'b00000000000000001000101111100000;
assign LUT_1[38225] = 32'b00000000000000000010000001011100;
assign LUT_1[38226] = 32'b00000000000000000100011101110001;
assign LUT_1[38227] = 32'b11111111111111111101101111101101;
assign LUT_1[38228] = 32'b00000000000000010000101000110111;
assign LUT_1[38229] = 32'b00000000000000001001111010110011;
assign LUT_1[38230] = 32'b00000000000000001100010111001000;
assign LUT_1[38231] = 32'b00000000000000000101101001000100;
assign LUT_1[38232] = 32'b00000000000000000111111101010101;
assign LUT_1[38233] = 32'b00000000000000000001001111010001;
assign LUT_1[38234] = 32'b00000000000000000011101011100110;
assign LUT_1[38235] = 32'b11111111111111111100111101100010;
assign LUT_1[38236] = 32'b00000000000000001111110110101100;
assign LUT_1[38237] = 32'b00000000000000001001001000101000;
assign LUT_1[38238] = 32'b00000000000000001011100100111101;
assign LUT_1[38239] = 32'b00000000000000000100110110111001;
assign LUT_1[38240] = 32'b00000000000000000111101110111101;
assign LUT_1[38241] = 32'b00000000000000000001000000111001;
assign LUT_1[38242] = 32'b00000000000000000011011101001110;
assign LUT_1[38243] = 32'b11111111111111111100101111001010;
assign LUT_1[38244] = 32'b00000000000000001111101000010100;
assign LUT_1[38245] = 32'b00000000000000001000111010010000;
assign LUT_1[38246] = 32'b00000000000000001011010110100101;
assign LUT_1[38247] = 32'b00000000000000000100101000100001;
assign LUT_1[38248] = 32'b00000000000000000110111100110010;
assign LUT_1[38249] = 32'b00000000000000000000001110101110;
assign LUT_1[38250] = 32'b00000000000000000010101011000011;
assign LUT_1[38251] = 32'b11111111111111111011111100111111;
assign LUT_1[38252] = 32'b00000000000000001110110110001001;
assign LUT_1[38253] = 32'b00000000000000001000001000000101;
assign LUT_1[38254] = 32'b00000000000000001010100100011010;
assign LUT_1[38255] = 32'b00000000000000000011110110010110;
assign LUT_1[38256] = 32'b00000000000000001001101010011111;
assign LUT_1[38257] = 32'b00000000000000000010111100011011;
assign LUT_1[38258] = 32'b00000000000000000101011000110000;
assign LUT_1[38259] = 32'b11111111111111111110101010101100;
assign LUT_1[38260] = 32'b00000000000000010001100011110110;
assign LUT_1[38261] = 32'b00000000000000001010110101110010;
assign LUT_1[38262] = 32'b00000000000000001101010010000111;
assign LUT_1[38263] = 32'b00000000000000000110100100000011;
assign LUT_1[38264] = 32'b00000000000000001000111000010100;
assign LUT_1[38265] = 32'b00000000000000000010001010010000;
assign LUT_1[38266] = 32'b00000000000000000100100110100101;
assign LUT_1[38267] = 32'b11111111111111111101111000100001;
assign LUT_1[38268] = 32'b00000000000000010000110001101011;
assign LUT_1[38269] = 32'b00000000000000001010000011100111;
assign LUT_1[38270] = 32'b00000000000000001100011111111100;
assign LUT_1[38271] = 32'b00000000000000000101110001111000;
assign LUT_1[38272] = 32'b00000000000000000111110110011001;
assign LUT_1[38273] = 32'b00000000000000000001001000010101;
assign LUT_1[38274] = 32'b00000000000000000011100100101010;
assign LUT_1[38275] = 32'b11111111111111111100110110100110;
assign LUT_1[38276] = 32'b00000000000000001111101111110000;
assign LUT_1[38277] = 32'b00000000000000001001000001101100;
assign LUT_1[38278] = 32'b00000000000000001011011110000001;
assign LUT_1[38279] = 32'b00000000000000000100101111111101;
assign LUT_1[38280] = 32'b00000000000000000111000100001110;
assign LUT_1[38281] = 32'b00000000000000000000010110001010;
assign LUT_1[38282] = 32'b00000000000000000010110010011111;
assign LUT_1[38283] = 32'b11111111111111111100000100011011;
assign LUT_1[38284] = 32'b00000000000000001110111101100101;
assign LUT_1[38285] = 32'b00000000000000001000001111100001;
assign LUT_1[38286] = 32'b00000000000000001010101011110110;
assign LUT_1[38287] = 32'b00000000000000000011111101110010;
assign LUT_1[38288] = 32'b00000000000000001001110001111011;
assign LUT_1[38289] = 32'b00000000000000000011000011110111;
assign LUT_1[38290] = 32'b00000000000000000101100000001100;
assign LUT_1[38291] = 32'b11111111111111111110110010001000;
assign LUT_1[38292] = 32'b00000000000000010001101011010010;
assign LUT_1[38293] = 32'b00000000000000001010111101001110;
assign LUT_1[38294] = 32'b00000000000000001101011001100011;
assign LUT_1[38295] = 32'b00000000000000000110101011011111;
assign LUT_1[38296] = 32'b00000000000000001000111111110000;
assign LUT_1[38297] = 32'b00000000000000000010010001101100;
assign LUT_1[38298] = 32'b00000000000000000100101110000001;
assign LUT_1[38299] = 32'b11111111111111111101111111111101;
assign LUT_1[38300] = 32'b00000000000000010000111001000111;
assign LUT_1[38301] = 32'b00000000000000001010001011000011;
assign LUT_1[38302] = 32'b00000000000000001100100111011000;
assign LUT_1[38303] = 32'b00000000000000000101111001010100;
assign LUT_1[38304] = 32'b00000000000000001000110001011000;
assign LUT_1[38305] = 32'b00000000000000000010000011010100;
assign LUT_1[38306] = 32'b00000000000000000100011111101001;
assign LUT_1[38307] = 32'b11111111111111111101110001100101;
assign LUT_1[38308] = 32'b00000000000000010000101010101111;
assign LUT_1[38309] = 32'b00000000000000001001111100101011;
assign LUT_1[38310] = 32'b00000000000000001100011001000000;
assign LUT_1[38311] = 32'b00000000000000000101101010111100;
assign LUT_1[38312] = 32'b00000000000000000111111111001101;
assign LUT_1[38313] = 32'b00000000000000000001010001001001;
assign LUT_1[38314] = 32'b00000000000000000011101101011110;
assign LUT_1[38315] = 32'b11111111111111111100111111011010;
assign LUT_1[38316] = 32'b00000000000000001111111000100100;
assign LUT_1[38317] = 32'b00000000000000001001001010100000;
assign LUT_1[38318] = 32'b00000000000000001011100110110101;
assign LUT_1[38319] = 32'b00000000000000000100111000110001;
assign LUT_1[38320] = 32'b00000000000000001010101100111010;
assign LUT_1[38321] = 32'b00000000000000000011111110110110;
assign LUT_1[38322] = 32'b00000000000000000110011011001011;
assign LUT_1[38323] = 32'b11111111111111111111101101000111;
assign LUT_1[38324] = 32'b00000000000000010010100110010001;
assign LUT_1[38325] = 32'b00000000000000001011111000001101;
assign LUT_1[38326] = 32'b00000000000000001110010100100010;
assign LUT_1[38327] = 32'b00000000000000000111100110011110;
assign LUT_1[38328] = 32'b00000000000000001001111010101111;
assign LUT_1[38329] = 32'b00000000000000000011001100101011;
assign LUT_1[38330] = 32'b00000000000000000101101001000000;
assign LUT_1[38331] = 32'b11111111111111111110111010111100;
assign LUT_1[38332] = 32'b00000000000000010001110100000110;
assign LUT_1[38333] = 32'b00000000000000001011000110000010;
assign LUT_1[38334] = 32'b00000000000000001101100010010111;
assign LUT_1[38335] = 32'b00000000000000000110110100010011;
assign LUT_1[38336] = 32'b00000000000000001001110100000001;
assign LUT_1[38337] = 32'b00000000000000000011000101111101;
assign LUT_1[38338] = 32'b00000000000000000101100010010010;
assign LUT_1[38339] = 32'b11111111111111111110110100001110;
assign LUT_1[38340] = 32'b00000000000000010001101101011000;
assign LUT_1[38341] = 32'b00000000000000001010111111010100;
assign LUT_1[38342] = 32'b00000000000000001101011011101001;
assign LUT_1[38343] = 32'b00000000000000000110101101100101;
assign LUT_1[38344] = 32'b00000000000000001001000001110110;
assign LUT_1[38345] = 32'b00000000000000000010010011110010;
assign LUT_1[38346] = 32'b00000000000000000100110000000111;
assign LUT_1[38347] = 32'b11111111111111111110000010000011;
assign LUT_1[38348] = 32'b00000000000000010000111011001101;
assign LUT_1[38349] = 32'b00000000000000001010001101001001;
assign LUT_1[38350] = 32'b00000000000000001100101001011110;
assign LUT_1[38351] = 32'b00000000000000000101111011011010;
assign LUT_1[38352] = 32'b00000000000000001011101111100011;
assign LUT_1[38353] = 32'b00000000000000000101000001011111;
assign LUT_1[38354] = 32'b00000000000000000111011101110100;
assign LUT_1[38355] = 32'b00000000000000000000101111110000;
assign LUT_1[38356] = 32'b00000000000000010011101000111010;
assign LUT_1[38357] = 32'b00000000000000001100111010110110;
assign LUT_1[38358] = 32'b00000000000000001111010111001011;
assign LUT_1[38359] = 32'b00000000000000001000101001000111;
assign LUT_1[38360] = 32'b00000000000000001010111101011000;
assign LUT_1[38361] = 32'b00000000000000000100001111010100;
assign LUT_1[38362] = 32'b00000000000000000110101011101001;
assign LUT_1[38363] = 32'b11111111111111111111111101100101;
assign LUT_1[38364] = 32'b00000000000000010010110110101111;
assign LUT_1[38365] = 32'b00000000000000001100001000101011;
assign LUT_1[38366] = 32'b00000000000000001110100101000000;
assign LUT_1[38367] = 32'b00000000000000000111110110111100;
assign LUT_1[38368] = 32'b00000000000000001010101111000000;
assign LUT_1[38369] = 32'b00000000000000000100000000111100;
assign LUT_1[38370] = 32'b00000000000000000110011101010001;
assign LUT_1[38371] = 32'b11111111111111111111101111001101;
assign LUT_1[38372] = 32'b00000000000000010010101000010111;
assign LUT_1[38373] = 32'b00000000000000001011111010010011;
assign LUT_1[38374] = 32'b00000000000000001110010110101000;
assign LUT_1[38375] = 32'b00000000000000000111101000100100;
assign LUT_1[38376] = 32'b00000000000000001001111100110101;
assign LUT_1[38377] = 32'b00000000000000000011001110110001;
assign LUT_1[38378] = 32'b00000000000000000101101011000110;
assign LUT_1[38379] = 32'b11111111111111111110111101000010;
assign LUT_1[38380] = 32'b00000000000000010001110110001100;
assign LUT_1[38381] = 32'b00000000000000001011001000001000;
assign LUT_1[38382] = 32'b00000000000000001101100100011101;
assign LUT_1[38383] = 32'b00000000000000000110110110011001;
assign LUT_1[38384] = 32'b00000000000000001100101010100010;
assign LUT_1[38385] = 32'b00000000000000000101111100011110;
assign LUT_1[38386] = 32'b00000000000000001000011000110011;
assign LUT_1[38387] = 32'b00000000000000000001101010101111;
assign LUT_1[38388] = 32'b00000000000000010100100011111001;
assign LUT_1[38389] = 32'b00000000000000001101110101110101;
assign LUT_1[38390] = 32'b00000000000000010000010010001010;
assign LUT_1[38391] = 32'b00000000000000001001100100000110;
assign LUT_1[38392] = 32'b00000000000000001011111000010111;
assign LUT_1[38393] = 32'b00000000000000000101001010010011;
assign LUT_1[38394] = 32'b00000000000000000111100110101000;
assign LUT_1[38395] = 32'b00000000000000000000111000100100;
assign LUT_1[38396] = 32'b00000000000000010011110001101110;
assign LUT_1[38397] = 32'b00000000000000001101000011101010;
assign LUT_1[38398] = 32'b00000000000000001111011111111111;
assign LUT_1[38399] = 32'b00000000000000001000110001111011;
assign LUT_1[38400] = 32'b00000000000000000000110000100111;
assign LUT_1[38401] = 32'b11111111111111111010000010100011;
assign LUT_1[38402] = 32'b11111111111111111100011110111000;
assign LUT_1[38403] = 32'b11111111111111110101110000110100;
assign LUT_1[38404] = 32'b00000000000000001000101001111110;
assign LUT_1[38405] = 32'b00000000000000000001111011111010;
assign LUT_1[38406] = 32'b00000000000000000100011000001111;
assign LUT_1[38407] = 32'b11111111111111111101101010001011;
assign LUT_1[38408] = 32'b11111111111111111111111110011100;
assign LUT_1[38409] = 32'b11111111111111111001010000011000;
assign LUT_1[38410] = 32'b11111111111111111011101100101101;
assign LUT_1[38411] = 32'b11111111111111110100111110101001;
assign LUT_1[38412] = 32'b00000000000000000111110111110011;
assign LUT_1[38413] = 32'b00000000000000000001001001101111;
assign LUT_1[38414] = 32'b00000000000000000011100110000100;
assign LUT_1[38415] = 32'b11111111111111111100111000000000;
assign LUT_1[38416] = 32'b00000000000000000010101100001001;
assign LUT_1[38417] = 32'b11111111111111111011111110000101;
assign LUT_1[38418] = 32'b11111111111111111110011010011010;
assign LUT_1[38419] = 32'b11111111111111110111101100010110;
assign LUT_1[38420] = 32'b00000000000000001010100101100000;
assign LUT_1[38421] = 32'b00000000000000000011110111011100;
assign LUT_1[38422] = 32'b00000000000000000110010011110001;
assign LUT_1[38423] = 32'b11111111111111111111100101101101;
assign LUT_1[38424] = 32'b00000000000000000001111001111110;
assign LUT_1[38425] = 32'b11111111111111111011001011111010;
assign LUT_1[38426] = 32'b11111111111111111101101000001111;
assign LUT_1[38427] = 32'b11111111111111110110111010001011;
assign LUT_1[38428] = 32'b00000000000000001001110011010101;
assign LUT_1[38429] = 32'b00000000000000000011000101010001;
assign LUT_1[38430] = 32'b00000000000000000101100001100110;
assign LUT_1[38431] = 32'b11111111111111111110110011100010;
assign LUT_1[38432] = 32'b00000000000000000001101011100110;
assign LUT_1[38433] = 32'b11111111111111111010111101100010;
assign LUT_1[38434] = 32'b11111111111111111101011001110111;
assign LUT_1[38435] = 32'b11111111111111110110101011110011;
assign LUT_1[38436] = 32'b00000000000000001001100100111101;
assign LUT_1[38437] = 32'b00000000000000000010110110111001;
assign LUT_1[38438] = 32'b00000000000000000101010011001110;
assign LUT_1[38439] = 32'b11111111111111111110100101001010;
assign LUT_1[38440] = 32'b00000000000000000000111001011011;
assign LUT_1[38441] = 32'b11111111111111111010001011010111;
assign LUT_1[38442] = 32'b11111111111111111100100111101100;
assign LUT_1[38443] = 32'b11111111111111110101111001101000;
assign LUT_1[38444] = 32'b00000000000000001000110010110010;
assign LUT_1[38445] = 32'b00000000000000000010000100101110;
assign LUT_1[38446] = 32'b00000000000000000100100001000011;
assign LUT_1[38447] = 32'b11111111111111111101110010111111;
assign LUT_1[38448] = 32'b00000000000000000011100111001000;
assign LUT_1[38449] = 32'b11111111111111111100111001000100;
assign LUT_1[38450] = 32'b11111111111111111111010101011001;
assign LUT_1[38451] = 32'b11111111111111111000100111010101;
assign LUT_1[38452] = 32'b00000000000000001011100000011111;
assign LUT_1[38453] = 32'b00000000000000000100110010011011;
assign LUT_1[38454] = 32'b00000000000000000111001110110000;
assign LUT_1[38455] = 32'b00000000000000000000100000101100;
assign LUT_1[38456] = 32'b00000000000000000010110100111101;
assign LUT_1[38457] = 32'b11111111111111111100000110111001;
assign LUT_1[38458] = 32'b11111111111111111110100011001110;
assign LUT_1[38459] = 32'b11111111111111110111110101001010;
assign LUT_1[38460] = 32'b00000000000000001010101110010100;
assign LUT_1[38461] = 32'b00000000000000000100000000010000;
assign LUT_1[38462] = 32'b00000000000000000110011100100101;
assign LUT_1[38463] = 32'b11111111111111111111101110100001;
assign LUT_1[38464] = 32'b00000000000000000010101110001111;
assign LUT_1[38465] = 32'b11111111111111111100000000001011;
assign LUT_1[38466] = 32'b11111111111111111110011100100000;
assign LUT_1[38467] = 32'b11111111111111110111101110011100;
assign LUT_1[38468] = 32'b00000000000000001010100111100110;
assign LUT_1[38469] = 32'b00000000000000000011111001100010;
assign LUT_1[38470] = 32'b00000000000000000110010101110111;
assign LUT_1[38471] = 32'b11111111111111111111100111110011;
assign LUT_1[38472] = 32'b00000000000000000001111100000100;
assign LUT_1[38473] = 32'b11111111111111111011001110000000;
assign LUT_1[38474] = 32'b11111111111111111101101010010101;
assign LUT_1[38475] = 32'b11111111111111110110111100010001;
assign LUT_1[38476] = 32'b00000000000000001001110101011011;
assign LUT_1[38477] = 32'b00000000000000000011000111010111;
assign LUT_1[38478] = 32'b00000000000000000101100011101100;
assign LUT_1[38479] = 32'b11111111111111111110110101101000;
assign LUT_1[38480] = 32'b00000000000000000100101001110001;
assign LUT_1[38481] = 32'b11111111111111111101111011101101;
assign LUT_1[38482] = 32'b00000000000000000000011000000010;
assign LUT_1[38483] = 32'b11111111111111111001101001111110;
assign LUT_1[38484] = 32'b00000000000000001100100011001000;
assign LUT_1[38485] = 32'b00000000000000000101110101000100;
assign LUT_1[38486] = 32'b00000000000000001000010001011001;
assign LUT_1[38487] = 32'b00000000000000000001100011010101;
assign LUT_1[38488] = 32'b00000000000000000011110111100110;
assign LUT_1[38489] = 32'b11111111111111111101001001100010;
assign LUT_1[38490] = 32'b11111111111111111111100101110111;
assign LUT_1[38491] = 32'b11111111111111111000110111110011;
assign LUT_1[38492] = 32'b00000000000000001011110000111101;
assign LUT_1[38493] = 32'b00000000000000000101000010111001;
assign LUT_1[38494] = 32'b00000000000000000111011111001110;
assign LUT_1[38495] = 32'b00000000000000000000110001001010;
assign LUT_1[38496] = 32'b00000000000000000011101001001110;
assign LUT_1[38497] = 32'b11111111111111111100111011001010;
assign LUT_1[38498] = 32'b11111111111111111111010111011111;
assign LUT_1[38499] = 32'b11111111111111111000101001011011;
assign LUT_1[38500] = 32'b00000000000000001011100010100101;
assign LUT_1[38501] = 32'b00000000000000000100110100100001;
assign LUT_1[38502] = 32'b00000000000000000111010000110110;
assign LUT_1[38503] = 32'b00000000000000000000100010110010;
assign LUT_1[38504] = 32'b00000000000000000010110111000011;
assign LUT_1[38505] = 32'b11111111111111111100001000111111;
assign LUT_1[38506] = 32'b11111111111111111110100101010100;
assign LUT_1[38507] = 32'b11111111111111110111110111010000;
assign LUT_1[38508] = 32'b00000000000000001010110000011010;
assign LUT_1[38509] = 32'b00000000000000000100000010010110;
assign LUT_1[38510] = 32'b00000000000000000110011110101011;
assign LUT_1[38511] = 32'b11111111111111111111110000100111;
assign LUT_1[38512] = 32'b00000000000000000101100100110000;
assign LUT_1[38513] = 32'b11111111111111111110110110101100;
assign LUT_1[38514] = 32'b00000000000000000001010011000001;
assign LUT_1[38515] = 32'b11111111111111111010100100111101;
assign LUT_1[38516] = 32'b00000000000000001101011110000111;
assign LUT_1[38517] = 32'b00000000000000000110110000000011;
assign LUT_1[38518] = 32'b00000000000000001001001100011000;
assign LUT_1[38519] = 32'b00000000000000000010011110010100;
assign LUT_1[38520] = 32'b00000000000000000100110010100101;
assign LUT_1[38521] = 32'b11111111111111111110000100100001;
assign LUT_1[38522] = 32'b00000000000000000000100000110110;
assign LUT_1[38523] = 32'b11111111111111111001110010110010;
assign LUT_1[38524] = 32'b00000000000000001100101011111100;
assign LUT_1[38525] = 32'b00000000000000000101111101111000;
assign LUT_1[38526] = 32'b00000000000000001000011010001101;
assign LUT_1[38527] = 32'b00000000000000000001101100001001;
assign LUT_1[38528] = 32'b00000000000000000011110000101010;
assign LUT_1[38529] = 32'b11111111111111111101000010100110;
assign LUT_1[38530] = 32'b11111111111111111111011110111011;
assign LUT_1[38531] = 32'b11111111111111111000110000110111;
assign LUT_1[38532] = 32'b00000000000000001011101010000001;
assign LUT_1[38533] = 32'b00000000000000000100111011111101;
assign LUT_1[38534] = 32'b00000000000000000111011000010010;
assign LUT_1[38535] = 32'b00000000000000000000101010001110;
assign LUT_1[38536] = 32'b00000000000000000010111110011111;
assign LUT_1[38537] = 32'b11111111111111111100010000011011;
assign LUT_1[38538] = 32'b11111111111111111110101100110000;
assign LUT_1[38539] = 32'b11111111111111110111111110101100;
assign LUT_1[38540] = 32'b00000000000000001010110111110110;
assign LUT_1[38541] = 32'b00000000000000000100001001110010;
assign LUT_1[38542] = 32'b00000000000000000110100110000111;
assign LUT_1[38543] = 32'b11111111111111111111111000000011;
assign LUT_1[38544] = 32'b00000000000000000101101100001100;
assign LUT_1[38545] = 32'b11111111111111111110111110001000;
assign LUT_1[38546] = 32'b00000000000000000001011010011101;
assign LUT_1[38547] = 32'b11111111111111111010101100011001;
assign LUT_1[38548] = 32'b00000000000000001101100101100011;
assign LUT_1[38549] = 32'b00000000000000000110110111011111;
assign LUT_1[38550] = 32'b00000000000000001001010011110100;
assign LUT_1[38551] = 32'b00000000000000000010100101110000;
assign LUT_1[38552] = 32'b00000000000000000100111010000001;
assign LUT_1[38553] = 32'b11111111111111111110001011111101;
assign LUT_1[38554] = 32'b00000000000000000000101000010010;
assign LUT_1[38555] = 32'b11111111111111111001111010001110;
assign LUT_1[38556] = 32'b00000000000000001100110011011000;
assign LUT_1[38557] = 32'b00000000000000000110000101010100;
assign LUT_1[38558] = 32'b00000000000000001000100001101001;
assign LUT_1[38559] = 32'b00000000000000000001110011100101;
assign LUT_1[38560] = 32'b00000000000000000100101011101001;
assign LUT_1[38561] = 32'b11111111111111111101111101100101;
assign LUT_1[38562] = 32'b00000000000000000000011001111010;
assign LUT_1[38563] = 32'b11111111111111111001101011110110;
assign LUT_1[38564] = 32'b00000000000000001100100101000000;
assign LUT_1[38565] = 32'b00000000000000000101110110111100;
assign LUT_1[38566] = 32'b00000000000000001000010011010001;
assign LUT_1[38567] = 32'b00000000000000000001100101001101;
assign LUT_1[38568] = 32'b00000000000000000011111001011110;
assign LUT_1[38569] = 32'b11111111111111111101001011011010;
assign LUT_1[38570] = 32'b11111111111111111111100111101111;
assign LUT_1[38571] = 32'b11111111111111111000111001101011;
assign LUT_1[38572] = 32'b00000000000000001011110010110101;
assign LUT_1[38573] = 32'b00000000000000000101000100110001;
assign LUT_1[38574] = 32'b00000000000000000111100001000110;
assign LUT_1[38575] = 32'b00000000000000000000110011000010;
assign LUT_1[38576] = 32'b00000000000000000110100111001011;
assign LUT_1[38577] = 32'b11111111111111111111111001000111;
assign LUT_1[38578] = 32'b00000000000000000010010101011100;
assign LUT_1[38579] = 32'b11111111111111111011100111011000;
assign LUT_1[38580] = 32'b00000000000000001110100000100010;
assign LUT_1[38581] = 32'b00000000000000000111110010011110;
assign LUT_1[38582] = 32'b00000000000000001010001110110011;
assign LUT_1[38583] = 32'b00000000000000000011100000101111;
assign LUT_1[38584] = 32'b00000000000000000101110101000000;
assign LUT_1[38585] = 32'b11111111111111111111000110111100;
assign LUT_1[38586] = 32'b00000000000000000001100011010001;
assign LUT_1[38587] = 32'b11111111111111111010110101001101;
assign LUT_1[38588] = 32'b00000000000000001101101110010111;
assign LUT_1[38589] = 32'b00000000000000000111000000010011;
assign LUT_1[38590] = 32'b00000000000000001001011100101000;
assign LUT_1[38591] = 32'b00000000000000000010101110100100;
assign LUT_1[38592] = 32'b00000000000000000101101110010010;
assign LUT_1[38593] = 32'b11111111111111111111000000001110;
assign LUT_1[38594] = 32'b00000000000000000001011100100011;
assign LUT_1[38595] = 32'b11111111111111111010101110011111;
assign LUT_1[38596] = 32'b00000000000000001101100111101001;
assign LUT_1[38597] = 32'b00000000000000000110111001100101;
assign LUT_1[38598] = 32'b00000000000000001001010101111010;
assign LUT_1[38599] = 32'b00000000000000000010100111110110;
assign LUT_1[38600] = 32'b00000000000000000100111100000111;
assign LUT_1[38601] = 32'b11111111111111111110001110000011;
assign LUT_1[38602] = 32'b00000000000000000000101010011000;
assign LUT_1[38603] = 32'b11111111111111111001111100010100;
assign LUT_1[38604] = 32'b00000000000000001100110101011110;
assign LUT_1[38605] = 32'b00000000000000000110000111011010;
assign LUT_1[38606] = 32'b00000000000000001000100011101111;
assign LUT_1[38607] = 32'b00000000000000000001110101101011;
assign LUT_1[38608] = 32'b00000000000000000111101001110100;
assign LUT_1[38609] = 32'b00000000000000000000111011110000;
assign LUT_1[38610] = 32'b00000000000000000011011000000101;
assign LUT_1[38611] = 32'b11111111111111111100101010000001;
assign LUT_1[38612] = 32'b00000000000000001111100011001011;
assign LUT_1[38613] = 32'b00000000000000001000110101000111;
assign LUT_1[38614] = 32'b00000000000000001011010001011100;
assign LUT_1[38615] = 32'b00000000000000000100100011011000;
assign LUT_1[38616] = 32'b00000000000000000110110111101001;
assign LUT_1[38617] = 32'b00000000000000000000001001100101;
assign LUT_1[38618] = 32'b00000000000000000010100101111010;
assign LUT_1[38619] = 32'b11111111111111111011110111110110;
assign LUT_1[38620] = 32'b00000000000000001110110001000000;
assign LUT_1[38621] = 32'b00000000000000001000000010111100;
assign LUT_1[38622] = 32'b00000000000000001010011111010001;
assign LUT_1[38623] = 32'b00000000000000000011110001001101;
assign LUT_1[38624] = 32'b00000000000000000110101001010001;
assign LUT_1[38625] = 32'b11111111111111111111111011001101;
assign LUT_1[38626] = 32'b00000000000000000010010111100010;
assign LUT_1[38627] = 32'b11111111111111111011101001011110;
assign LUT_1[38628] = 32'b00000000000000001110100010101000;
assign LUT_1[38629] = 32'b00000000000000000111110100100100;
assign LUT_1[38630] = 32'b00000000000000001010010000111001;
assign LUT_1[38631] = 32'b00000000000000000011100010110101;
assign LUT_1[38632] = 32'b00000000000000000101110111000110;
assign LUT_1[38633] = 32'b11111111111111111111001001000010;
assign LUT_1[38634] = 32'b00000000000000000001100101010111;
assign LUT_1[38635] = 32'b11111111111111111010110111010011;
assign LUT_1[38636] = 32'b00000000000000001101110000011101;
assign LUT_1[38637] = 32'b00000000000000000111000010011001;
assign LUT_1[38638] = 32'b00000000000000001001011110101110;
assign LUT_1[38639] = 32'b00000000000000000010110000101010;
assign LUT_1[38640] = 32'b00000000000000001000100100110011;
assign LUT_1[38641] = 32'b00000000000000000001110110101111;
assign LUT_1[38642] = 32'b00000000000000000100010011000100;
assign LUT_1[38643] = 32'b11111111111111111101100101000000;
assign LUT_1[38644] = 32'b00000000000000010000011110001010;
assign LUT_1[38645] = 32'b00000000000000001001110000000110;
assign LUT_1[38646] = 32'b00000000000000001100001100011011;
assign LUT_1[38647] = 32'b00000000000000000101011110010111;
assign LUT_1[38648] = 32'b00000000000000000111110010101000;
assign LUT_1[38649] = 32'b00000000000000000001000100100100;
assign LUT_1[38650] = 32'b00000000000000000011100000111001;
assign LUT_1[38651] = 32'b11111111111111111100110010110101;
assign LUT_1[38652] = 32'b00000000000000001111101011111111;
assign LUT_1[38653] = 32'b00000000000000001000111101111011;
assign LUT_1[38654] = 32'b00000000000000001011011010010000;
assign LUT_1[38655] = 32'b00000000000000000100101100001100;
assign LUT_1[38656] = 32'b11111111111111111110100100110011;
assign LUT_1[38657] = 32'b11111111111111110111110110101111;
assign LUT_1[38658] = 32'b11111111111111111010010011000100;
assign LUT_1[38659] = 32'b11111111111111110011100101000000;
assign LUT_1[38660] = 32'b00000000000000000110011110001010;
assign LUT_1[38661] = 32'b11111111111111111111110000000110;
assign LUT_1[38662] = 32'b00000000000000000010001100011011;
assign LUT_1[38663] = 32'b11111111111111111011011110010111;
assign LUT_1[38664] = 32'b11111111111111111101110010101000;
assign LUT_1[38665] = 32'b11111111111111110111000100100100;
assign LUT_1[38666] = 32'b11111111111111111001100000111001;
assign LUT_1[38667] = 32'b11111111111111110010110010110101;
assign LUT_1[38668] = 32'b00000000000000000101101011111111;
assign LUT_1[38669] = 32'b11111111111111111110111101111011;
assign LUT_1[38670] = 32'b00000000000000000001011010010000;
assign LUT_1[38671] = 32'b11111111111111111010101100001100;
assign LUT_1[38672] = 32'b00000000000000000000100000010101;
assign LUT_1[38673] = 32'b11111111111111111001110010010001;
assign LUT_1[38674] = 32'b11111111111111111100001110100110;
assign LUT_1[38675] = 32'b11111111111111110101100000100010;
assign LUT_1[38676] = 32'b00000000000000001000011001101100;
assign LUT_1[38677] = 32'b00000000000000000001101011101000;
assign LUT_1[38678] = 32'b00000000000000000100000111111101;
assign LUT_1[38679] = 32'b11111111111111111101011001111001;
assign LUT_1[38680] = 32'b11111111111111111111101110001010;
assign LUT_1[38681] = 32'b11111111111111111001000000000110;
assign LUT_1[38682] = 32'b11111111111111111011011100011011;
assign LUT_1[38683] = 32'b11111111111111110100101110010111;
assign LUT_1[38684] = 32'b00000000000000000111100111100001;
assign LUT_1[38685] = 32'b00000000000000000000111001011101;
assign LUT_1[38686] = 32'b00000000000000000011010101110010;
assign LUT_1[38687] = 32'b11111111111111111100100111101110;
assign LUT_1[38688] = 32'b11111111111111111111011111110010;
assign LUT_1[38689] = 32'b11111111111111111000110001101110;
assign LUT_1[38690] = 32'b11111111111111111011001110000011;
assign LUT_1[38691] = 32'b11111111111111110100011111111111;
assign LUT_1[38692] = 32'b00000000000000000111011001001001;
assign LUT_1[38693] = 32'b00000000000000000000101011000101;
assign LUT_1[38694] = 32'b00000000000000000011000111011010;
assign LUT_1[38695] = 32'b11111111111111111100011001010110;
assign LUT_1[38696] = 32'b11111111111111111110101101100111;
assign LUT_1[38697] = 32'b11111111111111110111111111100011;
assign LUT_1[38698] = 32'b11111111111111111010011011111000;
assign LUT_1[38699] = 32'b11111111111111110011101101110100;
assign LUT_1[38700] = 32'b00000000000000000110100110111110;
assign LUT_1[38701] = 32'b11111111111111111111111000111010;
assign LUT_1[38702] = 32'b00000000000000000010010101001111;
assign LUT_1[38703] = 32'b11111111111111111011100111001011;
assign LUT_1[38704] = 32'b00000000000000000001011011010100;
assign LUT_1[38705] = 32'b11111111111111111010101101010000;
assign LUT_1[38706] = 32'b11111111111111111101001001100101;
assign LUT_1[38707] = 32'b11111111111111110110011011100001;
assign LUT_1[38708] = 32'b00000000000000001001010100101011;
assign LUT_1[38709] = 32'b00000000000000000010100110100111;
assign LUT_1[38710] = 32'b00000000000000000101000010111100;
assign LUT_1[38711] = 32'b11111111111111111110010100111000;
assign LUT_1[38712] = 32'b00000000000000000000101001001001;
assign LUT_1[38713] = 32'b11111111111111111001111011000101;
assign LUT_1[38714] = 32'b11111111111111111100010111011010;
assign LUT_1[38715] = 32'b11111111111111110101101001010110;
assign LUT_1[38716] = 32'b00000000000000001000100010100000;
assign LUT_1[38717] = 32'b00000000000000000001110100011100;
assign LUT_1[38718] = 32'b00000000000000000100010000110001;
assign LUT_1[38719] = 32'b11111111111111111101100010101101;
assign LUT_1[38720] = 32'b00000000000000000000100010011011;
assign LUT_1[38721] = 32'b11111111111111111001110100010111;
assign LUT_1[38722] = 32'b11111111111111111100010000101100;
assign LUT_1[38723] = 32'b11111111111111110101100010101000;
assign LUT_1[38724] = 32'b00000000000000001000011011110010;
assign LUT_1[38725] = 32'b00000000000000000001101101101110;
assign LUT_1[38726] = 32'b00000000000000000100001010000011;
assign LUT_1[38727] = 32'b11111111111111111101011011111111;
assign LUT_1[38728] = 32'b11111111111111111111110000010000;
assign LUT_1[38729] = 32'b11111111111111111001000010001100;
assign LUT_1[38730] = 32'b11111111111111111011011110100001;
assign LUT_1[38731] = 32'b11111111111111110100110000011101;
assign LUT_1[38732] = 32'b00000000000000000111101001100111;
assign LUT_1[38733] = 32'b00000000000000000000111011100011;
assign LUT_1[38734] = 32'b00000000000000000011010111111000;
assign LUT_1[38735] = 32'b11111111111111111100101001110100;
assign LUT_1[38736] = 32'b00000000000000000010011101111101;
assign LUT_1[38737] = 32'b11111111111111111011101111111001;
assign LUT_1[38738] = 32'b11111111111111111110001100001110;
assign LUT_1[38739] = 32'b11111111111111110111011110001010;
assign LUT_1[38740] = 32'b00000000000000001010010111010100;
assign LUT_1[38741] = 32'b00000000000000000011101001010000;
assign LUT_1[38742] = 32'b00000000000000000110000101100101;
assign LUT_1[38743] = 32'b11111111111111111111010111100001;
assign LUT_1[38744] = 32'b00000000000000000001101011110010;
assign LUT_1[38745] = 32'b11111111111111111010111101101110;
assign LUT_1[38746] = 32'b11111111111111111101011010000011;
assign LUT_1[38747] = 32'b11111111111111110110101011111111;
assign LUT_1[38748] = 32'b00000000000000001001100101001001;
assign LUT_1[38749] = 32'b00000000000000000010110111000101;
assign LUT_1[38750] = 32'b00000000000000000101010011011010;
assign LUT_1[38751] = 32'b11111111111111111110100101010110;
assign LUT_1[38752] = 32'b00000000000000000001011101011010;
assign LUT_1[38753] = 32'b11111111111111111010101111010110;
assign LUT_1[38754] = 32'b11111111111111111101001011101011;
assign LUT_1[38755] = 32'b11111111111111110110011101100111;
assign LUT_1[38756] = 32'b00000000000000001001010110110001;
assign LUT_1[38757] = 32'b00000000000000000010101000101101;
assign LUT_1[38758] = 32'b00000000000000000101000101000010;
assign LUT_1[38759] = 32'b11111111111111111110010110111110;
assign LUT_1[38760] = 32'b00000000000000000000101011001111;
assign LUT_1[38761] = 32'b11111111111111111001111101001011;
assign LUT_1[38762] = 32'b11111111111111111100011001100000;
assign LUT_1[38763] = 32'b11111111111111110101101011011100;
assign LUT_1[38764] = 32'b00000000000000001000100100100110;
assign LUT_1[38765] = 32'b00000000000000000001110110100010;
assign LUT_1[38766] = 32'b00000000000000000100010010110111;
assign LUT_1[38767] = 32'b11111111111111111101100100110011;
assign LUT_1[38768] = 32'b00000000000000000011011000111100;
assign LUT_1[38769] = 32'b11111111111111111100101010111000;
assign LUT_1[38770] = 32'b11111111111111111111000111001101;
assign LUT_1[38771] = 32'b11111111111111111000011001001001;
assign LUT_1[38772] = 32'b00000000000000001011010010010011;
assign LUT_1[38773] = 32'b00000000000000000100100100001111;
assign LUT_1[38774] = 32'b00000000000000000111000000100100;
assign LUT_1[38775] = 32'b00000000000000000000010010100000;
assign LUT_1[38776] = 32'b00000000000000000010100110110001;
assign LUT_1[38777] = 32'b11111111111111111011111000101101;
assign LUT_1[38778] = 32'b11111111111111111110010101000010;
assign LUT_1[38779] = 32'b11111111111111110111100110111110;
assign LUT_1[38780] = 32'b00000000000000001010100000001000;
assign LUT_1[38781] = 32'b00000000000000000011110010000100;
assign LUT_1[38782] = 32'b00000000000000000110001110011001;
assign LUT_1[38783] = 32'b11111111111111111111100000010101;
assign LUT_1[38784] = 32'b00000000000000000001100100110110;
assign LUT_1[38785] = 32'b11111111111111111010110110110010;
assign LUT_1[38786] = 32'b11111111111111111101010011000111;
assign LUT_1[38787] = 32'b11111111111111110110100101000011;
assign LUT_1[38788] = 32'b00000000000000001001011110001101;
assign LUT_1[38789] = 32'b00000000000000000010110000001001;
assign LUT_1[38790] = 32'b00000000000000000101001100011110;
assign LUT_1[38791] = 32'b11111111111111111110011110011010;
assign LUT_1[38792] = 32'b00000000000000000000110010101011;
assign LUT_1[38793] = 32'b11111111111111111010000100100111;
assign LUT_1[38794] = 32'b11111111111111111100100000111100;
assign LUT_1[38795] = 32'b11111111111111110101110010111000;
assign LUT_1[38796] = 32'b00000000000000001000101100000010;
assign LUT_1[38797] = 32'b00000000000000000001111101111110;
assign LUT_1[38798] = 32'b00000000000000000100011010010011;
assign LUT_1[38799] = 32'b11111111111111111101101100001111;
assign LUT_1[38800] = 32'b00000000000000000011100000011000;
assign LUT_1[38801] = 32'b11111111111111111100110010010100;
assign LUT_1[38802] = 32'b11111111111111111111001110101001;
assign LUT_1[38803] = 32'b11111111111111111000100000100101;
assign LUT_1[38804] = 32'b00000000000000001011011001101111;
assign LUT_1[38805] = 32'b00000000000000000100101011101011;
assign LUT_1[38806] = 32'b00000000000000000111001000000000;
assign LUT_1[38807] = 32'b00000000000000000000011001111100;
assign LUT_1[38808] = 32'b00000000000000000010101110001101;
assign LUT_1[38809] = 32'b11111111111111111100000000001001;
assign LUT_1[38810] = 32'b11111111111111111110011100011110;
assign LUT_1[38811] = 32'b11111111111111110111101110011010;
assign LUT_1[38812] = 32'b00000000000000001010100111100100;
assign LUT_1[38813] = 32'b00000000000000000011111001100000;
assign LUT_1[38814] = 32'b00000000000000000110010101110101;
assign LUT_1[38815] = 32'b11111111111111111111100111110001;
assign LUT_1[38816] = 32'b00000000000000000010011111110101;
assign LUT_1[38817] = 32'b11111111111111111011110001110001;
assign LUT_1[38818] = 32'b11111111111111111110001110000110;
assign LUT_1[38819] = 32'b11111111111111110111100000000010;
assign LUT_1[38820] = 32'b00000000000000001010011001001100;
assign LUT_1[38821] = 32'b00000000000000000011101011001000;
assign LUT_1[38822] = 32'b00000000000000000110000111011101;
assign LUT_1[38823] = 32'b11111111111111111111011001011001;
assign LUT_1[38824] = 32'b00000000000000000001101101101010;
assign LUT_1[38825] = 32'b11111111111111111010111111100110;
assign LUT_1[38826] = 32'b11111111111111111101011011111011;
assign LUT_1[38827] = 32'b11111111111111110110101101110111;
assign LUT_1[38828] = 32'b00000000000000001001100111000001;
assign LUT_1[38829] = 32'b00000000000000000010111000111101;
assign LUT_1[38830] = 32'b00000000000000000101010101010010;
assign LUT_1[38831] = 32'b11111111111111111110100111001110;
assign LUT_1[38832] = 32'b00000000000000000100011011010111;
assign LUT_1[38833] = 32'b11111111111111111101101101010011;
assign LUT_1[38834] = 32'b00000000000000000000001001101000;
assign LUT_1[38835] = 32'b11111111111111111001011011100100;
assign LUT_1[38836] = 32'b00000000000000001100010100101110;
assign LUT_1[38837] = 32'b00000000000000000101100110101010;
assign LUT_1[38838] = 32'b00000000000000001000000010111111;
assign LUT_1[38839] = 32'b00000000000000000001010100111011;
assign LUT_1[38840] = 32'b00000000000000000011101001001100;
assign LUT_1[38841] = 32'b11111111111111111100111011001000;
assign LUT_1[38842] = 32'b11111111111111111111010111011101;
assign LUT_1[38843] = 32'b11111111111111111000101001011001;
assign LUT_1[38844] = 32'b00000000000000001011100010100011;
assign LUT_1[38845] = 32'b00000000000000000100110100011111;
assign LUT_1[38846] = 32'b00000000000000000111010000110100;
assign LUT_1[38847] = 32'b00000000000000000000100010110000;
assign LUT_1[38848] = 32'b00000000000000000011100010011110;
assign LUT_1[38849] = 32'b11111111111111111100110100011010;
assign LUT_1[38850] = 32'b11111111111111111111010000101111;
assign LUT_1[38851] = 32'b11111111111111111000100010101011;
assign LUT_1[38852] = 32'b00000000000000001011011011110101;
assign LUT_1[38853] = 32'b00000000000000000100101101110001;
assign LUT_1[38854] = 32'b00000000000000000111001010000110;
assign LUT_1[38855] = 32'b00000000000000000000011100000010;
assign LUT_1[38856] = 32'b00000000000000000010110000010011;
assign LUT_1[38857] = 32'b11111111111111111100000010001111;
assign LUT_1[38858] = 32'b11111111111111111110011110100100;
assign LUT_1[38859] = 32'b11111111111111110111110000100000;
assign LUT_1[38860] = 32'b00000000000000001010101001101010;
assign LUT_1[38861] = 32'b00000000000000000011111011100110;
assign LUT_1[38862] = 32'b00000000000000000110010111111011;
assign LUT_1[38863] = 32'b11111111111111111111101001110111;
assign LUT_1[38864] = 32'b00000000000000000101011110000000;
assign LUT_1[38865] = 32'b11111111111111111110101111111100;
assign LUT_1[38866] = 32'b00000000000000000001001100010001;
assign LUT_1[38867] = 32'b11111111111111111010011110001101;
assign LUT_1[38868] = 32'b00000000000000001101010111010111;
assign LUT_1[38869] = 32'b00000000000000000110101001010011;
assign LUT_1[38870] = 32'b00000000000000001001000101101000;
assign LUT_1[38871] = 32'b00000000000000000010010111100100;
assign LUT_1[38872] = 32'b00000000000000000100101011110101;
assign LUT_1[38873] = 32'b11111111111111111101111101110001;
assign LUT_1[38874] = 32'b00000000000000000000011010000110;
assign LUT_1[38875] = 32'b11111111111111111001101100000010;
assign LUT_1[38876] = 32'b00000000000000001100100101001100;
assign LUT_1[38877] = 32'b00000000000000000101110111001000;
assign LUT_1[38878] = 32'b00000000000000001000010011011101;
assign LUT_1[38879] = 32'b00000000000000000001100101011001;
assign LUT_1[38880] = 32'b00000000000000000100011101011101;
assign LUT_1[38881] = 32'b11111111111111111101101111011001;
assign LUT_1[38882] = 32'b00000000000000000000001011101110;
assign LUT_1[38883] = 32'b11111111111111111001011101101010;
assign LUT_1[38884] = 32'b00000000000000001100010110110100;
assign LUT_1[38885] = 32'b00000000000000000101101000110000;
assign LUT_1[38886] = 32'b00000000000000001000000101000101;
assign LUT_1[38887] = 32'b00000000000000000001010111000001;
assign LUT_1[38888] = 32'b00000000000000000011101011010010;
assign LUT_1[38889] = 32'b11111111111111111100111101001110;
assign LUT_1[38890] = 32'b11111111111111111111011001100011;
assign LUT_1[38891] = 32'b11111111111111111000101011011111;
assign LUT_1[38892] = 32'b00000000000000001011100100101001;
assign LUT_1[38893] = 32'b00000000000000000100110110100101;
assign LUT_1[38894] = 32'b00000000000000000111010010111010;
assign LUT_1[38895] = 32'b00000000000000000000100100110110;
assign LUT_1[38896] = 32'b00000000000000000110011000111111;
assign LUT_1[38897] = 32'b11111111111111111111101010111011;
assign LUT_1[38898] = 32'b00000000000000000010000111010000;
assign LUT_1[38899] = 32'b11111111111111111011011001001100;
assign LUT_1[38900] = 32'b00000000000000001110010010010110;
assign LUT_1[38901] = 32'b00000000000000000111100100010010;
assign LUT_1[38902] = 32'b00000000000000001010000000100111;
assign LUT_1[38903] = 32'b00000000000000000011010010100011;
assign LUT_1[38904] = 32'b00000000000000000101100110110100;
assign LUT_1[38905] = 32'b11111111111111111110111000110000;
assign LUT_1[38906] = 32'b00000000000000000001010101000101;
assign LUT_1[38907] = 32'b11111111111111111010100111000001;
assign LUT_1[38908] = 32'b00000000000000001101100000001011;
assign LUT_1[38909] = 32'b00000000000000000110110010000111;
assign LUT_1[38910] = 32'b00000000000000001001001110011100;
assign LUT_1[38911] = 32'b00000000000000000010100000011000;
assign LUT_1[38912] = 32'b00000000000000000001101101010101;
assign LUT_1[38913] = 32'b11111111111111111010111111010001;
assign LUT_1[38914] = 32'b11111111111111111101011011100110;
assign LUT_1[38915] = 32'b11111111111111110110101101100010;
assign LUT_1[38916] = 32'b00000000000000001001100110101100;
assign LUT_1[38917] = 32'b00000000000000000010111000101000;
assign LUT_1[38918] = 32'b00000000000000000101010100111101;
assign LUT_1[38919] = 32'b11111111111111111110100110111001;
assign LUT_1[38920] = 32'b00000000000000000000111011001010;
assign LUT_1[38921] = 32'b11111111111111111010001101000110;
assign LUT_1[38922] = 32'b11111111111111111100101001011011;
assign LUT_1[38923] = 32'b11111111111111110101111011010111;
assign LUT_1[38924] = 32'b00000000000000001000110100100001;
assign LUT_1[38925] = 32'b00000000000000000010000110011101;
assign LUT_1[38926] = 32'b00000000000000000100100010110010;
assign LUT_1[38927] = 32'b11111111111111111101110100101110;
assign LUT_1[38928] = 32'b00000000000000000011101000110111;
assign LUT_1[38929] = 32'b11111111111111111100111010110011;
assign LUT_1[38930] = 32'b11111111111111111111010111001000;
assign LUT_1[38931] = 32'b11111111111111111000101001000100;
assign LUT_1[38932] = 32'b00000000000000001011100010001110;
assign LUT_1[38933] = 32'b00000000000000000100110100001010;
assign LUT_1[38934] = 32'b00000000000000000111010000011111;
assign LUT_1[38935] = 32'b00000000000000000000100010011011;
assign LUT_1[38936] = 32'b00000000000000000010110110101100;
assign LUT_1[38937] = 32'b11111111111111111100001000101000;
assign LUT_1[38938] = 32'b11111111111111111110100100111101;
assign LUT_1[38939] = 32'b11111111111111110111110110111001;
assign LUT_1[38940] = 32'b00000000000000001010110000000011;
assign LUT_1[38941] = 32'b00000000000000000100000001111111;
assign LUT_1[38942] = 32'b00000000000000000110011110010100;
assign LUT_1[38943] = 32'b11111111111111111111110000010000;
assign LUT_1[38944] = 32'b00000000000000000010101000010100;
assign LUT_1[38945] = 32'b11111111111111111011111010010000;
assign LUT_1[38946] = 32'b11111111111111111110010110100101;
assign LUT_1[38947] = 32'b11111111111111110111101000100001;
assign LUT_1[38948] = 32'b00000000000000001010100001101011;
assign LUT_1[38949] = 32'b00000000000000000011110011100111;
assign LUT_1[38950] = 32'b00000000000000000110001111111100;
assign LUT_1[38951] = 32'b11111111111111111111100001111000;
assign LUT_1[38952] = 32'b00000000000000000001110110001001;
assign LUT_1[38953] = 32'b11111111111111111011001000000101;
assign LUT_1[38954] = 32'b11111111111111111101100100011010;
assign LUT_1[38955] = 32'b11111111111111110110110110010110;
assign LUT_1[38956] = 32'b00000000000000001001101111100000;
assign LUT_1[38957] = 32'b00000000000000000011000001011100;
assign LUT_1[38958] = 32'b00000000000000000101011101110001;
assign LUT_1[38959] = 32'b11111111111111111110101111101101;
assign LUT_1[38960] = 32'b00000000000000000100100011110110;
assign LUT_1[38961] = 32'b11111111111111111101110101110010;
assign LUT_1[38962] = 32'b00000000000000000000010010000111;
assign LUT_1[38963] = 32'b11111111111111111001100100000011;
assign LUT_1[38964] = 32'b00000000000000001100011101001101;
assign LUT_1[38965] = 32'b00000000000000000101101111001001;
assign LUT_1[38966] = 32'b00000000000000001000001011011110;
assign LUT_1[38967] = 32'b00000000000000000001011101011010;
assign LUT_1[38968] = 32'b00000000000000000011110001101011;
assign LUT_1[38969] = 32'b11111111111111111101000011100111;
assign LUT_1[38970] = 32'b11111111111111111111011111111100;
assign LUT_1[38971] = 32'b11111111111111111000110001111000;
assign LUT_1[38972] = 32'b00000000000000001011101011000010;
assign LUT_1[38973] = 32'b00000000000000000100111100111110;
assign LUT_1[38974] = 32'b00000000000000000111011001010011;
assign LUT_1[38975] = 32'b00000000000000000000101011001111;
assign LUT_1[38976] = 32'b00000000000000000011101010111101;
assign LUT_1[38977] = 32'b11111111111111111100111100111001;
assign LUT_1[38978] = 32'b11111111111111111111011001001110;
assign LUT_1[38979] = 32'b11111111111111111000101011001010;
assign LUT_1[38980] = 32'b00000000000000001011100100010100;
assign LUT_1[38981] = 32'b00000000000000000100110110010000;
assign LUT_1[38982] = 32'b00000000000000000111010010100101;
assign LUT_1[38983] = 32'b00000000000000000000100100100001;
assign LUT_1[38984] = 32'b00000000000000000010111000110010;
assign LUT_1[38985] = 32'b11111111111111111100001010101110;
assign LUT_1[38986] = 32'b11111111111111111110100111000011;
assign LUT_1[38987] = 32'b11111111111111110111111000111111;
assign LUT_1[38988] = 32'b00000000000000001010110010001001;
assign LUT_1[38989] = 32'b00000000000000000100000100000101;
assign LUT_1[38990] = 32'b00000000000000000110100000011010;
assign LUT_1[38991] = 32'b11111111111111111111110010010110;
assign LUT_1[38992] = 32'b00000000000000000101100110011111;
assign LUT_1[38993] = 32'b11111111111111111110111000011011;
assign LUT_1[38994] = 32'b00000000000000000001010100110000;
assign LUT_1[38995] = 32'b11111111111111111010100110101100;
assign LUT_1[38996] = 32'b00000000000000001101011111110110;
assign LUT_1[38997] = 32'b00000000000000000110110001110010;
assign LUT_1[38998] = 32'b00000000000000001001001110000111;
assign LUT_1[38999] = 32'b00000000000000000010100000000011;
assign LUT_1[39000] = 32'b00000000000000000100110100010100;
assign LUT_1[39001] = 32'b11111111111111111110000110010000;
assign LUT_1[39002] = 32'b00000000000000000000100010100101;
assign LUT_1[39003] = 32'b11111111111111111001110100100001;
assign LUT_1[39004] = 32'b00000000000000001100101101101011;
assign LUT_1[39005] = 32'b00000000000000000101111111100111;
assign LUT_1[39006] = 32'b00000000000000001000011011111100;
assign LUT_1[39007] = 32'b00000000000000000001101101111000;
assign LUT_1[39008] = 32'b00000000000000000100100101111100;
assign LUT_1[39009] = 32'b11111111111111111101110111111000;
assign LUT_1[39010] = 32'b00000000000000000000010100001101;
assign LUT_1[39011] = 32'b11111111111111111001100110001001;
assign LUT_1[39012] = 32'b00000000000000001100011111010011;
assign LUT_1[39013] = 32'b00000000000000000101110001001111;
assign LUT_1[39014] = 32'b00000000000000001000001101100100;
assign LUT_1[39015] = 32'b00000000000000000001011111100000;
assign LUT_1[39016] = 32'b00000000000000000011110011110001;
assign LUT_1[39017] = 32'b11111111111111111101000101101101;
assign LUT_1[39018] = 32'b11111111111111111111100010000010;
assign LUT_1[39019] = 32'b11111111111111111000110011111110;
assign LUT_1[39020] = 32'b00000000000000001011101101001000;
assign LUT_1[39021] = 32'b00000000000000000100111111000100;
assign LUT_1[39022] = 32'b00000000000000000111011011011001;
assign LUT_1[39023] = 32'b00000000000000000000101101010101;
assign LUT_1[39024] = 32'b00000000000000000110100001011110;
assign LUT_1[39025] = 32'b11111111111111111111110011011010;
assign LUT_1[39026] = 32'b00000000000000000010001111101111;
assign LUT_1[39027] = 32'b11111111111111111011100001101011;
assign LUT_1[39028] = 32'b00000000000000001110011010110101;
assign LUT_1[39029] = 32'b00000000000000000111101100110001;
assign LUT_1[39030] = 32'b00000000000000001010001001000110;
assign LUT_1[39031] = 32'b00000000000000000011011011000010;
assign LUT_1[39032] = 32'b00000000000000000101101111010011;
assign LUT_1[39033] = 32'b11111111111111111111000001001111;
assign LUT_1[39034] = 32'b00000000000000000001011101100100;
assign LUT_1[39035] = 32'b11111111111111111010101111100000;
assign LUT_1[39036] = 32'b00000000000000001101101000101010;
assign LUT_1[39037] = 32'b00000000000000000110111010100110;
assign LUT_1[39038] = 32'b00000000000000001001010110111011;
assign LUT_1[39039] = 32'b00000000000000000010101000110111;
assign LUT_1[39040] = 32'b00000000000000000100101101011000;
assign LUT_1[39041] = 32'b11111111111111111101111111010100;
assign LUT_1[39042] = 32'b00000000000000000000011011101001;
assign LUT_1[39043] = 32'b11111111111111111001101101100101;
assign LUT_1[39044] = 32'b00000000000000001100100110101111;
assign LUT_1[39045] = 32'b00000000000000000101111000101011;
assign LUT_1[39046] = 32'b00000000000000001000010101000000;
assign LUT_1[39047] = 32'b00000000000000000001100110111100;
assign LUT_1[39048] = 32'b00000000000000000011111011001101;
assign LUT_1[39049] = 32'b11111111111111111101001101001001;
assign LUT_1[39050] = 32'b11111111111111111111101001011110;
assign LUT_1[39051] = 32'b11111111111111111000111011011010;
assign LUT_1[39052] = 32'b00000000000000001011110100100100;
assign LUT_1[39053] = 32'b00000000000000000101000110100000;
assign LUT_1[39054] = 32'b00000000000000000111100010110101;
assign LUT_1[39055] = 32'b00000000000000000000110100110001;
assign LUT_1[39056] = 32'b00000000000000000110101000111010;
assign LUT_1[39057] = 32'b11111111111111111111111010110110;
assign LUT_1[39058] = 32'b00000000000000000010010111001011;
assign LUT_1[39059] = 32'b11111111111111111011101001000111;
assign LUT_1[39060] = 32'b00000000000000001110100010010001;
assign LUT_1[39061] = 32'b00000000000000000111110100001101;
assign LUT_1[39062] = 32'b00000000000000001010010000100010;
assign LUT_1[39063] = 32'b00000000000000000011100010011110;
assign LUT_1[39064] = 32'b00000000000000000101110110101111;
assign LUT_1[39065] = 32'b11111111111111111111001000101011;
assign LUT_1[39066] = 32'b00000000000000000001100101000000;
assign LUT_1[39067] = 32'b11111111111111111010110110111100;
assign LUT_1[39068] = 32'b00000000000000001101110000000110;
assign LUT_1[39069] = 32'b00000000000000000111000010000010;
assign LUT_1[39070] = 32'b00000000000000001001011110010111;
assign LUT_1[39071] = 32'b00000000000000000010110000010011;
assign LUT_1[39072] = 32'b00000000000000000101101000010111;
assign LUT_1[39073] = 32'b11111111111111111110111010010011;
assign LUT_1[39074] = 32'b00000000000000000001010110101000;
assign LUT_1[39075] = 32'b11111111111111111010101000100100;
assign LUT_1[39076] = 32'b00000000000000001101100001101110;
assign LUT_1[39077] = 32'b00000000000000000110110011101010;
assign LUT_1[39078] = 32'b00000000000000001001001111111111;
assign LUT_1[39079] = 32'b00000000000000000010100001111011;
assign LUT_1[39080] = 32'b00000000000000000100110110001100;
assign LUT_1[39081] = 32'b11111111111111111110001000001000;
assign LUT_1[39082] = 32'b00000000000000000000100100011101;
assign LUT_1[39083] = 32'b11111111111111111001110110011001;
assign LUT_1[39084] = 32'b00000000000000001100101111100011;
assign LUT_1[39085] = 32'b00000000000000000110000001011111;
assign LUT_1[39086] = 32'b00000000000000001000011101110100;
assign LUT_1[39087] = 32'b00000000000000000001101111110000;
assign LUT_1[39088] = 32'b00000000000000000111100011111001;
assign LUT_1[39089] = 32'b00000000000000000000110101110101;
assign LUT_1[39090] = 32'b00000000000000000011010010001010;
assign LUT_1[39091] = 32'b11111111111111111100100100000110;
assign LUT_1[39092] = 32'b00000000000000001111011101010000;
assign LUT_1[39093] = 32'b00000000000000001000101111001100;
assign LUT_1[39094] = 32'b00000000000000001011001011100001;
assign LUT_1[39095] = 32'b00000000000000000100011101011101;
assign LUT_1[39096] = 32'b00000000000000000110110001101110;
assign LUT_1[39097] = 32'b00000000000000000000000011101010;
assign LUT_1[39098] = 32'b00000000000000000010011111111111;
assign LUT_1[39099] = 32'b11111111111111111011110001111011;
assign LUT_1[39100] = 32'b00000000000000001110101011000101;
assign LUT_1[39101] = 32'b00000000000000000111111101000001;
assign LUT_1[39102] = 32'b00000000000000001010011001010110;
assign LUT_1[39103] = 32'b00000000000000000011101011010010;
assign LUT_1[39104] = 32'b00000000000000000110101011000000;
assign LUT_1[39105] = 32'b11111111111111111111111100111100;
assign LUT_1[39106] = 32'b00000000000000000010011001010001;
assign LUT_1[39107] = 32'b11111111111111111011101011001101;
assign LUT_1[39108] = 32'b00000000000000001110100100010111;
assign LUT_1[39109] = 32'b00000000000000000111110110010011;
assign LUT_1[39110] = 32'b00000000000000001010010010101000;
assign LUT_1[39111] = 32'b00000000000000000011100100100100;
assign LUT_1[39112] = 32'b00000000000000000101111000110101;
assign LUT_1[39113] = 32'b11111111111111111111001010110001;
assign LUT_1[39114] = 32'b00000000000000000001100111000110;
assign LUT_1[39115] = 32'b11111111111111111010111001000010;
assign LUT_1[39116] = 32'b00000000000000001101110010001100;
assign LUT_1[39117] = 32'b00000000000000000111000100001000;
assign LUT_1[39118] = 32'b00000000000000001001100000011101;
assign LUT_1[39119] = 32'b00000000000000000010110010011001;
assign LUT_1[39120] = 32'b00000000000000001000100110100010;
assign LUT_1[39121] = 32'b00000000000000000001111000011110;
assign LUT_1[39122] = 32'b00000000000000000100010100110011;
assign LUT_1[39123] = 32'b11111111111111111101100110101111;
assign LUT_1[39124] = 32'b00000000000000010000011111111001;
assign LUT_1[39125] = 32'b00000000000000001001110001110101;
assign LUT_1[39126] = 32'b00000000000000001100001110001010;
assign LUT_1[39127] = 32'b00000000000000000101100000000110;
assign LUT_1[39128] = 32'b00000000000000000111110100010111;
assign LUT_1[39129] = 32'b00000000000000000001000110010011;
assign LUT_1[39130] = 32'b00000000000000000011100010101000;
assign LUT_1[39131] = 32'b11111111111111111100110100100100;
assign LUT_1[39132] = 32'b00000000000000001111101101101110;
assign LUT_1[39133] = 32'b00000000000000001000111111101010;
assign LUT_1[39134] = 32'b00000000000000001011011011111111;
assign LUT_1[39135] = 32'b00000000000000000100101101111011;
assign LUT_1[39136] = 32'b00000000000000000111100101111111;
assign LUT_1[39137] = 32'b00000000000000000000110111111011;
assign LUT_1[39138] = 32'b00000000000000000011010100010000;
assign LUT_1[39139] = 32'b11111111111111111100100110001100;
assign LUT_1[39140] = 32'b00000000000000001111011111010110;
assign LUT_1[39141] = 32'b00000000000000001000110001010010;
assign LUT_1[39142] = 32'b00000000000000001011001101100111;
assign LUT_1[39143] = 32'b00000000000000000100011111100011;
assign LUT_1[39144] = 32'b00000000000000000110110011110100;
assign LUT_1[39145] = 32'b00000000000000000000000101110000;
assign LUT_1[39146] = 32'b00000000000000000010100010000101;
assign LUT_1[39147] = 32'b11111111111111111011110100000001;
assign LUT_1[39148] = 32'b00000000000000001110101101001011;
assign LUT_1[39149] = 32'b00000000000000000111111111000111;
assign LUT_1[39150] = 32'b00000000000000001010011011011100;
assign LUT_1[39151] = 32'b00000000000000000011101101011000;
assign LUT_1[39152] = 32'b00000000000000001001100001100001;
assign LUT_1[39153] = 32'b00000000000000000010110011011101;
assign LUT_1[39154] = 32'b00000000000000000101001111110010;
assign LUT_1[39155] = 32'b11111111111111111110100001101110;
assign LUT_1[39156] = 32'b00000000000000010001011010111000;
assign LUT_1[39157] = 32'b00000000000000001010101100110100;
assign LUT_1[39158] = 32'b00000000000000001101001001001001;
assign LUT_1[39159] = 32'b00000000000000000110011011000101;
assign LUT_1[39160] = 32'b00000000000000001000101111010110;
assign LUT_1[39161] = 32'b00000000000000000010000001010010;
assign LUT_1[39162] = 32'b00000000000000000100011101100111;
assign LUT_1[39163] = 32'b11111111111111111101101111100011;
assign LUT_1[39164] = 32'b00000000000000010000101000101101;
assign LUT_1[39165] = 32'b00000000000000001001111010101001;
assign LUT_1[39166] = 32'b00000000000000001100010110111110;
assign LUT_1[39167] = 32'b00000000000000000101101000111010;
assign LUT_1[39168] = 32'b11111111111111111111100001100001;
assign LUT_1[39169] = 32'b11111111111111111000110011011101;
assign LUT_1[39170] = 32'b11111111111111111011001111110010;
assign LUT_1[39171] = 32'b11111111111111110100100001101110;
assign LUT_1[39172] = 32'b00000000000000000111011010111000;
assign LUT_1[39173] = 32'b00000000000000000000101100110100;
assign LUT_1[39174] = 32'b00000000000000000011001001001001;
assign LUT_1[39175] = 32'b11111111111111111100011011000101;
assign LUT_1[39176] = 32'b11111111111111111110101111010110;
assign LUT_1[39177] = 32'b11111111111111111000000001010010;
assign LUT_1[39178] = 32'b11111111111111111010011101100111;
assign LUT_1[39179] = 32'b11111111111111110011101111100011;
assign LUT_1[39180] = 32'b00000000000000000110101000101101;
assign LUT_1[39181] = 32'b11111111111111111111111010101001;
assign LUT_1[39182] = 32'b00000000000000000010010110111110;
assign LUT_1[39183] = 32'b11111111111111111011101000111010;
assign LUT_1[39184] = 32'b00000000000000000001011101000011;
assign LUT_1[39185] = 32'b11111111111111111010101110111111;
assign LUT_1[39186] = 32'b11111111111111111101001011010100;
assign LUT_1[39187] = 32'b11111111111111110110011101010000;
assign LUT_1[39188] = 32'b00000000000000001001010110011010;
assign LUT_1[39189] = 32'b00000000000000000010101000010110;
assign LUT_1[39190] = 32'b00000000000000000101000100101011;
assign LUT_1[39191] = 32'b11111111111111111110010110100111;
assign LUT_1[39192] = 32'b00000000000000000000101010111000;
assign LUT_1[39193] = 32'b11111111111111111001111100110100;
assign LUT_1[39194] = 32'b11111111111111111100011001001001;
assign LUT_1[39195] = 32'b11111111111111110101101011000101;
assign LUT_1[39196] = 32'b00000000000000001000100100001111;
assign LUT_1[39197] = 32'b00000000000000000001110110001011;
assign LUT_1[39198] = 32'b00000000000000000100010010100000;
assign LUT_1[39199] = 32'b11111111111111111101100100011100;
assign LUT_1[39200] = 32'b00000000000000000000011100100000;
assign LUT_1[39201] = 32'b11111111111111111001101110011100;
assign LUT_1[39202] = 32'b11111111111111111100001010110001;
assign LUT_1[39203] = 32'b11111111111111110101011100101101;
assign LUT_1[39204] = 32'b00000000000000001000010101110111;
assign LUT_1[39205] = 32'b00000000000000000001100111110011;
assign LUT_1[39206] = 32'b00000000000000000100000100001000;
assign LUT_1[39207] = 32'b11111111111111111101010110000100;
assign LUT_1[39208] = 32'b11111111111111111111101010010101;
assign LUT_1[39209] = 32'b11111111111111111000111100010001;
assign LUT_1[39210] = 32'b11111111111111111011011000100110;
assign LUT_1[39211] = 32'b11111111111111110100101010100010;
assign LUT_1[39212] = 32'b00000000000000000111100011101100;
assign LUT_1[39213] = 32'b00000000000000000000110101101000;
assign LUT_1[39214] = 32'b00000000000000000011010001111101;
assign LUT_1[39215] = 32'b11111111111111111100100011111001;
assign LUT_1[39216] = 32'b00000000000000000010011000000010;
assign LUT_1[39217] = 32'b11111111111111111011101001111110;
assign LUT_1[39218] = 32'b11111111111111111110000110010011;
assign LUT_1[39219] = 32'b11111111111111110111011000001111;
assign LUT_1[39220] = 32'b00000000000000001010010001011001;
assign LUT_1[39221] = 32'b00000000000000000011100011010101;
assign LUT_1[39222] = 32'b00000000000000000101111111101010;
assign LUT_1[39223] = 32'b11111111111111111111010001100110;
assign LUT_1[39224] = 32'b00000000000000000001100101110111;
assign LUT_1[39225] = 32'b11111111111111111010110111110011;
assign LUT_1[39226] = 32'b11111111111111111101010100001000;
assign LUT_1[39227] = 32'b11111111111111110110100110000100;
assign LUT_1[39228] = 32'b00000000000000001001011111001110;
assign LUT_1[39229] = 32'b00000000000000000010110001001010;
assign LUT_1[39230] = 32'b00000000000000000101001101011111;
assign LUT_1[39231] = 32'b11111111111111111110011111011011;
assign LUT_1[39232] = 32'b00000000000000000001011111001001;
assign LUT_1[39233] = 32'b11111111111111111010110001000101;
assign LUT_1[39234] = 32'b11111111111111111101001101011010;
assign LUT_1[39235] = 32'b11111111111111110110011111010110;
assign LUT_1[39236] = 32'b00000000000000001001011000100000;
assign LUT_1[39237] = 32'b00000000000000000010101010011100;
assign LUT_1[39238] = 32'b00000000000000000101000110110001;
assign LUT_1[39239] = 32'b11111111111111111110011000101101;
assign LUT_1[39240] = 32'b00000000000000000000101100111110;
assign LUT_1[39241] = 32'b11111111111111111001111110111010;
assign LUT_1[39242] = 32'b11111111111111111100011011001111;
assign LUT_1[39243] = 32'b11111111111111110101101101001011;
assign LUT_1[39244] = 32'b00000000000000001000100110010101;
assign LUT_1[39245] = 32'b00000000000000000001111000010001;
assign LUT_1[39246] = 32'b00000000000000000100010100100110;
assign LUT_1[39247] = 32'b11111111111111111101100110100010;
assign LUT_1[39248] = 32'b00000000000000000011011010101011;
assign LUT_1[39249] = 32'b11111111111111111100101100100111;
assign LUT_1[39250] = 32'b11111111111111111111001000111100;
assign LUT_1[39251] = 32'b11111111111111111000011010111000;
assign LUT_1[39252] = 32'b00000000000000001011010100000010;
assign LUT_1[39253] = 32'b00000000000000000100100101111110;
assign LUT_1[39254] = 32'b00000000000000000111000010010011;
assign LUT_1[39255] = 32'b00000000000000000000010100001111;
assign LUT_1[39256] = 32'b00000000000000000010101000100000;
assign LUT_1[39257] = 32'b11111111111111111011111010011100;
assign LUT_1[39258] = 32'b11111111111111111110010110110001;
assign LUT_1[39259] = 32'b11111111111111110111101000101101;
assign LUT_1[39260] = 32'b00000000000000001010100001110111;
assign LUT_1[39261] = 32'b00000000000000000011110011110011;
assign LUT_1[39262] = 32'b00000000000000000110010000001000;
assign LUT_1[39263] = 32'b11111111111111111111100010000100;
assign LUT_1[39264] = 32'b00000000000000000010011010001000;
assign LUT_1[39265] = 32'b11111111111111111011101100000100;
assign LUT_1[39266] = 32'b11111111111111111110001000011001;
assign LUT_1[39267] = 32'b11111111111111110111011010010101;
assign LUT_1[39268] = 32'b00000000000000001010010011011111;
assign LUT_1[39269] = 32'b00000000000000000011100101011011;
assign LUT_1[39270] = 32'b00000000000000000110000001110000;
assign LUT_1[39271] = 32'b11111111111111111111010011101100;
assign LUT_1[39272] = 32'b00000000000000000001100111111101;
assign LUT_1[39273] = 32'b11111111111111111010111001111001;
assign LUT_1[39274] = 32'b11111111111111111101010110001110;
assign LUT_1[39275] = 32'b11111111111111110110101000001010;
assign LUT_1[39276] = 32'b00000000000000001001100001010100;
assign LUT_1[39277] = 32'b00000000000000000010110011010000;
assign LUT_1[39278] = 32'b00000000000000000101001111100101;
assign LUT_1[39279] = 32'b11111111111111111110100001100001;
assign LUT_1[39280] = 32'b00000000000000000100010101101010;
assign LUT_1[39281] = 32'b11111111111111111101100111100110;
assign LUT_1[39282] = 32'b00000000000000000000000011111011;
assign LUT_1[39283] = 32'b11111111111111111001010101110111;
assign LUT_1[39284] = 32'b00000000000000001100001111000001;
assign LUT_1[39285] = 32'b00000000000000000101100000111101;
assign LUT_1[39286] = 32'b00000000000000000111111101010010;
assign LUT_1[39287] = 32'b00000000000000000001001111001110;
assign LUT_1[39288] = 32'b00000000000000000011100011011111;
assign LUT_1[39289] = 32'b11111111111111111100110101011011;
assign LUT_1[39290] = 32'b11111111111111111111010001110000;
assign LUT_1[39291] = 32'b11111111111111111000100011101100;
assign LUT_1[39292] = 32'b00000000000000001011011100110110;
assign LUT_1[39293] = 32'b00000000000000000100101110110010;
assign LUT_1[39294] = 32'b00000000000000000111001011000111;
assign LUT_1[39295] = 32'b00000000000000000000011101000011;
assign LUT_1[39296] = 32'b00000000000000000010100001100100;
assign LUT_1[39297] = 32'b11111111111111111011110011100000;
assign LUT_1[39298] = 32'b11111111111111111110001111110101;
assign LUT_1[39299] = 32'b11111111111111110111100001110001;
assign LUT_1[39300] = 32'b00000000000000001010011010111011;
assign LUT_1[39301] = 32'b00000000000000000011101100110111;
assign LUT_1[39302] = 32'b00000000000000000110001001001100;
assign LUT_1[39303] = 32'b11111111111111111111011011001000;
assign LUT_1[39304] = 32'b00000000000000000001101111011001;
assign LUT_1[39305] = 32'b11111111111111111011000001010101;
assign LUT_1[39306] = 32'b11111111111111111101011101101010;
assign LUT_1[39307] = 32'b11111111111111110110101111100110;
assign LUT_1[39308] = 32'b00000000000000001001101000110000;
assign LUT_1[39309] = 32'b00000000000000000010111010101100;
assign LUT_1[39310] = 32'b00000000000000000101010111000001;
assign LUT_1[39311] = 32'b11111111111111111110101000111101;
assign LUT_1[39312] = 32'b00000000000000000100011101000110;
assign LUT_1[39313] = 32'b11111111111111111101101111000010;
assign LUT_1[39314] = 32'b00000000000000000000001011010111;
assign LUT_1[39315] = 32'b11111111111111111001011101010011;
assign LUT_1[39316] = 32'b00000000000000001100010110011101;
assign LUT_1[39317] = 32'b00000000000000000101101000011001;
assign LUT_1[39318] = 32'b00000000000000001000000100101110;
assign LUT_1[39319] = 32'b00000000000000000001010110101010;
assign LUT_1[39320] = 32'b00000000000000000011101010111011;
assign LUT_1[39321] = 32'b11111111111111111100111100110111;
assign LUT_1[39322] = 32'b11111111111111111111011001001100;
assign LUT_1[39323] = 32'b11111111111111111000101011001000;
assign LUT_1[39324] = 32'b00000000000000001011100100010010;
assign LUT_1[39325] = 32'b00000000000000000100110110001110;
assign LUT_1[39326] = 32'b00000000000000000111010010100011;
assign LUT_1[39327] = 32'b00000000000000000000100100011111;
assign LUT_1[39328] = 32'b00000000000000000011011100100011;
assign LUT_1[39329] = 32'b11111111111111111100101110011111;
assign LUT_1[39330] = 32'b11111111111111111111001010110100;
assign LUT_1[39331] = 32'b11111111111111111000011100110000;
assign LUT_1[39332] = 32'b00000000000000001011010101111010;
assign LUT_1[39333] = 32'b00000000000000000100100111110110;
assign LUT_1[39334] = 32'b00000000000000000111000100001011;
assign LUT_1[39335] = 32'b00000000000000000000010110000111;
assign LUT_1[39336] = 32'b00000000000000000010101010011000;
assign LUT_1[39337] = 32'b11111111111111111011111100010100;
assign LUT_1[39338] = 32'b11111111111111111110011000101001;
assign LUT_1[39339] = 32'b11111111111111110111101010100101;
assign LUT_1[39340] = 32'b00000000000000001010100011101111;
assign LUT_1[39341] = 32'b00000000000000000011110101101011;
assign LUT_1[39342] = 32'b00000000000000000110010010000000;
assign LUT_1[39343] = 32'b11111111111111111111100011111100;
assign LUT_1[39344] = 32'b00000000000000000101011000000101;
assign LUT_1[39345] = 32'b11111111111111111110101010000001;
assign LUT_1[39346] = 32'b00000000000000000001000110010110;
assign LUT_1[39347] = 32'b11111111111111111010011000010010;
assign LUT_1[39348] = 32'b00000000000000001101010001011100;
assign LUT_1[39349] = 32'b00000000000000000110100011011000;
assign LUT_1[39350] = 32'b00000000000000001000111111101101;
assign LUT_1[39351] = 32'b00000000000000000010010001101001;
assign LUT_1[39352] = 32'b00000000000000000100100101111010;
assign LUT_1[39353] = 32'b11111111111111111101110111110110;
assign LUT_1[39354] = 32'b00000000000000000000010100001011;
assign LUT_1[39355] = 32'b11111111111111111001100110000111;
assign LUT_1[39356] = 32'b00000000000000001100011111010001;
assign LUT_1[39357] = 32'b00000000000000000101110001001101;
assign LUT_1[39358] = 32'b00000000000000001000001101100010;
assign LUT_1[39359] = 32'b00000000000000000001011111011110;
assign LUT_1[39360] = 32'b00000000000000000100011111001100;
assign LUT_1[39361] = 32'b11111111111111111101110001001000;
assign LUT_1[39362] = 32'b00000000000000000000001101011101;
assign LUT_1[39363] = 32'b11111111111111111001011111011001;
assign LUT_1[39364] = 32'b00000000000000001100011000100011;
assign LUT_1[39365] = 32'b00000000000000000101101010011111;
assign LUT_1[39366] = 32'b00000000000000001000000110110100;
assign LUT_1[39367] = 32'b00000000000000000001011000110000;
assign LUT_1[39368] = 32'b00000000000000000011101101000001;
assign LUT_1[39369] = 32'b11111111111111111100111110111101;
assign LUT_1[39370] = 32'b11111111111111111111011011010010;
assign LUT_1[39371] = 32'b11111111111111111000101101001110;
assign LUT_1[39372] = 32'b00000000000000001011100110011000;
assign LUT_1[39373] = 32'b00000000000000000100111000010100;
assign LUT_1[39374] = 32'b00000000000000000111010100101001;
assign LUT_1[39375] = 32'b00000000000000000000100110100101;
assign LUT_1[39376] = 32'b00000000000000000110011010101110;
assign LUT_1[39377] = 32'b11111111111111111111101100101010;
assign LUT_1[39378] = 32'b00000000000000000010001000111111;
assign LUT_1[39379] = 32'b11111111111111111011011010111011;
assign LUT_1[39380] = 32'b00000000000000001110010100000101;
assign LUT_1[39381] = 32'b00000000000000000111100110000001;
assign LUT_1[39382] = 32'b00000000000000001010000010010110;
assign LUT_1[39383] = 32'b00000000000000000011010100010010;
assign LUT_1[39384] = 32'b00000000000000000101101000100011;
assign LUT_1[39385] = 32'b11111111111111111110111010011111;
assign LUT_1[39386] = 32'b00000000000000000001010110110100;
assign LUT_1[39387] = 32'b11111111111111111010101000110000;
assign LUT_1[39388] = 32'b00000000000000001101100001111010;
assign LUT_1[39389] = 32'b00000000000000000110110011110110;
assign LUT_1[39390] = 32'b00000000000000001001010000001011;
assign LUT_1[39391] = 32'b00000000000000000010100010000111;
assign LUT_1[39392] = 32'b00000000000000000101011010001011;
assign LUT_1[39393] = 32'b11111111111111111110101100000111;
assign LUT_1[39394] = 32'b00000000000000000001001000011100;
assign LUT_1[39395] = 32'b11111111111111111010011010011000;
assign LUT_1[39396] = 32'b00000000000000001101010011100010;
assign LUT_1[39397] = 32'b00000000000000000110100101011110;
assign LUT_1[39398] = 32'b00000000000000001001000001110011;
assign LUT_1[39399] = 32'b00000000000000000010010011101111;
assign LUT_1[39400] = 32'b00000000000000000100101000000000;
assign LUT_1[39401] = 32'b11111111111111111101111001111100;
assign LUT_1[39402] = 32'b00000000000000000000010110010001;
assign LUT_1[39403] = 32'b11111111111111111001101000001101;
assign LUT_1[39404] = 32'b00000000000000001100100001010111;
assign LUT_1[39405] = 32'b00000000000000000101110011010011;
assign LUT_1[39406] = 32'b00000000000000001000001111101000;
assign LUT_1[39407] = 32'b00000000000000000001100001100100;
assign LUT_1[39408] = 32'b00000000000000000111010101101101;
assign LUT_1[39409] = 32'b00000000000000000000100111101001;
assign LUT_1[39410] = 32'b00000000000000000011000011111110;
assign LUT_1[39411] = 32'b11111111111111111100010101111010;
assign LUT_1[39412] = 32'b00000000000000001111001111000100;
assign LUT_1[39413] = 32'b00000000000000001000100001000000;
assign LUT_1[39414] = 32'b00000000000000001010111101010101;
assign LUT_1[39415] = 32'b00000000000000000100001111010001;
assign LUT_1[39416] = 32'b00000000000000000110100011100010;
assign LUT_1[39417] = 32'b11111111111111111111110101011110;
assign LUT_1[39418] = 32'b00000000000000000010010001110011;
assign LUT_1[39419] = 32'b11111111111111111011100011101111;
assign LUT_1[39420] = 32'b00000000000000001110011100111001;
assign LUT_1[39421] = 32'b00000000000000000111101110110101;
assign LUT_1[39422] = 32'b00000000000000001010001011001010;
assign LUT_1[39423] = 32'b00000000000000000011011101000110;
assign LUT_1[39424] = 32'b11111111111111111011011011110010;
assign LUT_1[39425] = 32'b11111111111111110100101101101110;
assign LUT_1[39426] = 32'b11111111111111110111001010000011;
assign LUT_1[39427] = 32'b11111111111111110000011011111111;
assign LUT_1[39428] = 32'b00000000000000000011010101001001;
assign LUT_1[39429] = 32'b11111111111111111100100111000101;
assign LUT_1[39430] = 32'b11111111111111111111000011011010;
assign LUT_1[39431] = 32'b11111111111111111000010101010110;
assign LUT_1[39432] = 32'b11111111111111111010101001100111;
assign LUT_1[39433] = 32'b11111111111111110011111011100011;
assign LUT_1[39434] = 32'b11111111111111110110010111111000;
assign LUT_1[39435] = 32'b11111111111111101111101001110100;
assign LUT_1[39436] = 32'b00000000000000000010100010111110;
assign LUT_1[39437] = 32'b11111111111111111011110100111010;
assign LUT_1[39438] = 32'b11111111111111111110010001001111;
assign LUT_1[39439] = 32'b11111111111111110111100011001011;
assign LUT_1[39440] = 32'b11111111111111111101010111010100;
assign LUT_1[39441] = 32'b11111111111111110110101001010000;
assign LUT_1[39442] = 32'b11111111111111111001000101100101;
assign LUT_1[39443] = 32'b11111111111111110010010111100001;
assign LUT_1[39444] = 32'b00000000000000000101010000101011;
assign LUT_1[39445] = 32'b11111111111111111110100010100111;
assign LUT_1[39446] = 32'b00000000000000000000111110111100;
assign LUT_1[39447] = 32'b11111111111111111010010000111000;
assign LUT_1[39448] = 32'b11111111111111111100100101001001;
assign LUT_1[39449] = 32'b11111111111111110101110111000101;
assign LUT_1[39450] = 32'b11111111111111111000010011011010;
assign LUT_1[39451] = 32'b11111111111111110001100101010110;
assign LUT_1[39452] = 32'b00000000000000000100011110100000;
assign LUT_1[39453] = 32'b11111111111111111101110000011100;
assign LUT_1[39454] = 32'b00000000000000000000001100110001;
assign LUT_1[39455] = 32'b11111111111111111001011110101101;
assign LUT_1[39456] = 32'b11111111111111111100010110110001;
assign LUT_1[39457] = 32'b11111111111111110101101000101101;
assign LUT_1[39458] = 32'b11111111111111111000000101000010;
assign LUT_1[39459] = 32'b11111111111111110001010110111110;
assign LUT_1[39460] = 32'b00000000000000000100010000001000;
assign LUT_1[39461] = 32'b11111111111111111101100010000100;
assign LUT_1[39462] = 32'b11111111111111111111111110011001;
assign LUT_1[39463] = 32'b11111111111111111001010000010101;
assign LUT_1[39464] = 32'b11111111111111111011100100100110;
assign LUT_1[39465] = 32'b11111111111111110100110110100010;
assign LUT_1[39466] = 32'b11111111111111110111010010110111;
assign LUT_1[39467] = 32'b11111111111111110000100100110011;
assign LUT_1[39468] = 32'b00000000000000000011011101111101;
assign LUT_1[39469] = 32'b11111111111111111100101111111001;
assign LUT_1[39470] = 32'b11111111111111111111001100001110;
assign LUT_1[39471] = 32'b11111111111111111000011110001010;
assign LUT_1[39472] = 32'b11111111111111111110010010010011;
assign LUT_1[39473] = 32'b11111111111111110111100100001111;
assign LUT_1[39474] = 32'b11111111111111111010000000100100;
assign LUT_1[39475] = 32'b11111111111111110011010010100000;
assign LUT_1[39476] = 32'b00000000000000000110001011101010;
assign LUT_1[39477] = 32'b11111111111111111111011101100110;
assign LUT_1[39478] = 32'b00000000000000000001111001111011;
assign LUT_1[39479] = 32'b11111111111111111011001011110111;
assign LUT_1[39480] = 32'b11111111111111111101100000001000;
assign LUT_1[39481] = 32'b11111111111111110110110010000100;
assign LUT_1[39482] = 32'b11111111111111111001001110011001;
assign LUT_1[39483] = 32'b11111111111111110010100000010101;
assign LUT_1[39484] = 32'b00000000000000000101011001011111;
assign LUT_1[39485] = 32'b11111111111111111110101011011011;
assign LUT_1[39486] = 32'b00000000000000000001000111110000;
assign LUT_1[39487] = 32'b11111111111111111010011001101100;
assign LUT_1[39488] = 32'b11111111111111111101011001011010;
assign LUT_1[39489] = 32'b11111111111111110110101011010110;
assign LUT_1[39490] = 32'b11111111111111111001000111101011;
assign LUT_1[39491] = 32'b11111111111111110010011001100111;
assign LUT_1[39492] = 32'b00000000000000000101010010110001;
assign LUT_1[39493] = 32'b11111111111111111110100100101101;
assign LUT_1[39494] = 32'b00000000000000000001000001000010;
assign LUT_1[39495] = 32'b11111111111111111010010010111110;
assign LUT_1[39496] = 32'b11111111111111111100100111001111;
assign LUT_1[39497] = 32'b11111111111111110101111001001011;
assign LUT_1[39498] = 32'b11111111111111111000010101100000;
assign LUT_1[39499] = 32'b11111111111111110001100111011100;
assign LUT_1[39500] = 32'b00000000000000000100100000100110;
assign LUT_1[39501] = 32'b11111111111111111101110010100010;
assign LUT_1[39502] = 32'b00000000000000000000001110110111;
assign LUT_1[39503] = 32'b11111111111111111001100000110011;
assign LUT_1[39504] = 32'b11111111111111111111010100111100;
assign LUT_1[39505] = 32'b11111111111111111000100110111000;
assign LUT_1[39506] = 32'b11111111111111111011000011001101;
assign LUT_1[39507] = 32'b11111111111111110100010101001001;
assign LUT_1[39508] = 32'b00000000000000000111001110010011;
assign LUT_1[39509] = 32'b00000000000000000000100000001111;
assign LUT_1[39510] = 32'b00000000000000000010111100100100;
assign LUT_1[39511] = 32'b11111111111111111100001110100000;
assign LUT_1[39512] = 32'b11111111111111111110100010110001;
assign LUT_1[39513] = 32'b11111111111111110111110100101101;
assign LUT_1[39514] = 32'b11111111111111111010010001000010;
assign LUT_1[39515] = 32'b11111111111111110011100010111110;
assign LUT_1[39516] = 32'b00000000000000000110011100001000;
assign LUT_1[39517] = 32'b11111111111111111111101110000100;
assign LUT_1[39518] = 32'b00000000000000000010001010011001;
assign LUT_1[39519] = 32'b11111111111111111011011100010101;
assign LUT_1[39520] = 32'b11111111111111111110010100011001;
assign LUT_1[39521] = 32'b11111111111111110111100110010101;
assign LUT_1[39522] = 32'b11111111111111111010000010101010;
assign LUT_1[39523] = 32'b11111111111111110011010100100110;
assign LUT_1[39524] = 32'b00000000000000000110001101110000;
assign LUT_1[39525] = 32'b11111111111111111111011111101100;
assign LUT_1[39526] = 32'b00000000000000000001111100000001;
assign LUT_1[39527] = 32'b11111111111111111011001101111101;
assign LUT_1[39528] = 32'b11111111111111111101100010001110;
assign LUT_1[39529] = 32'b11111111111111110110110100001010;
assign LUT_1[39530] = 32'b11111111111111111001010000011111;
assign LUT_1[39531] = 32'b11111111111111110010100010011011;
assign LUT_1[39532] = 32'b00000000000000000101011011100101;
assign LUT_1[39533] = 32'b11111111111111111110101101100001;
assign LUT_1[39534] = 32'b00000000000000000001001001110110;
assign LUT_1[39535] = 32'b11111111111111111010011011110010;
assign LUT_1[39536] = 32'b00000000000000000000001111111011;
assign LUT_1[39537] = 32'b11111111111111111001100001110111;
assign LUT_1[39538] = 32'b11111111111111111011111110001100;
assign LUT_1[39539] = 32'b11111111111111110101010000001000;
assign LUT_1[39540] = 32'b00000000000000001000001001010010;
assign LUT_1[39541] = 32'b00000000000000000001011011001110;
assign LUT_1[39542] = 32'b00000000000000000011110111100011;
assign LUT_1[39543] = 32'b11111111111111111101001001011111;
assign LUT_1[39544] = 32'b11111111111111111111011101110000;
assign LUT_1[39545] = 32'b11111111111111111000101111101100;
assign LUT_1[39546] = 32'b11111111111111111011001100000001;
assign LUT_1[39547] = 32'b11111111111111110100011101111101;
assign LUT_1[39548] = 32'b00000000000000000111010111000111;
assign LUT_1[39549] = 32'b00000000000000000000101001000011;
assign LUT_1[39550] = 32'b00000000000000000011000101011000;
assign LUT_1[39551] = 32'b11111111111111111100010111010100;
assign LUT_1[39552] = 32'b11111111111111111110011011110101;
assign LUT_1[39553] = 32'b11111111111111110111101101110001;
assign LUT_1[39554] = 32'b11111111111111111010001010000110;
assign LUT_1[39555] = 32'b11111111111111110011011100000010;
assign LUT_1[39556] = 32'b00000000000000000110010101001100;
assign LUT_1[39557] = 32'b11111111111111111111100111001000;
assign LUT_1[39558] = 32'b00000000000000000010000011011101;
assign LUT_1[39559] = 32'b11111111111111111011010101011001;
assign LUT_1[39560] = 32'b11111111111111111101101001101010;
assign LUT_1[39561] = 32'b11111111111111110110111011100110;
assign LUT_1[39562] = 32'b11111111111111111001010111111011;
assign LUT_1[39563] = 32'b11111111111111110010101001110111;
assign LUT_1[39564] = 32'b00000000000000000101100011000001;
assign LUT_1[39565] = 32'b11111111111111111110110100111101;
assign LUT_1[39566] = 32'b00000000000000000001010001010010;
assign LUT_1[39567] = 32'b11111111111111111010100011001110;
assign LUT_1[39568] = 32'b00000000000000000000010111010111;
assign LUT_1[39569] = 32'b11111111111111111001101001010011;
assign LUT_1[39570] = 32'b11111111111111111100000101101000;
assign LUT_1[39571] = 32'b11111111111111110101010111100100;
assign LUT_1[39572] = 32'b00000000000000001000010000101110;
assign LUT_1[39573] = 32'b00000000000000000001100010101010;
assign LUT_1[39574] = 32'b00000000000000000011111110111111;
assign LUT_1[39575] = 32'b11111111111111111101010000111011;
assign LUT_1[39576] = 32'b11111111111111111111100101001100;
assign LUT_1[39577] = 32'b11111111111111111000110111001000;
assign LUT_1[39578] = 32'b11111111111111111011010011011101;
assign LUT_1[39579] = 32'b11111111111111110100100101011001;
assign LUT_1[39580] = 32'b00000000000000000111011110100011;
assign LUT_1[39581] = 32'b00000000000000000000110000011111;
assign LUT_1[39582] = 32'b00000000000000000011001100110100;
assign LUT_1[39583] = 32'b11111111111111111100011110110000;
assign LUT_1[39584] = 32'b11111111111111111111010110110100;
assign LUT_1[39585] = 32'b11111111111111111000101000110000;
assign LUT_1[39586] = 32'b11111111111111111011000101000101;
assign LUT_1[39587] = 32'b11111111111111110100010111000001;
assign LUT_1[39588] = 32'b00000000000000000111010000001011;
assign LUT_1[39589] = 32'b00000000000000000000100010000111;
assign LUT_1[39590] = 32'b00000000000000000010111110011100;
assign LUT_1[39591] = 32'b11111111111111111100010000011000;
assign LUT_1[39592] = 32'b11111111111111111110100100101001;
assign LUT_1[39593] = 32'b11111111111111110111110110100101;
assign LUT_1[39594] = 32'b11111111111111111010010010111010;
assign LUT_1[39595] = 32'b11111111111111110011100100110110;
assign LUT_1[39596] = 32'b00000000000000000110011110000000;
assign LUT_1[39597] = 32'b11111111111111111111101111111100;
assign LUT_1[39598] = 32'b00000000000000000010001100010001;
assign LUT_1[39599] = 32'b11111111111111111011011110001101;
assign LUT_1[39600] = 32'b00000000000000000001010010010110;
assign LUT_1[39601] = 32'b11111111111111111010100100010010;
assign LUT_1[39602] = 32'b11111111111111111101000000100111;
assign LUT_1[39603] = 32'b11111111111111110110010010100011;
assign LUT_1[39604] = 32'b00000000000000001001001011101101;
assign LUT_1[39605] = 32'b00000000000000000010011101101001;
assign LUT_1[39606] = 32'b00000000000000000100111001111110;
assign LUT_1[39607] = 32'b11111111111111111110001011111010;
assign LUT_1[39608] = 32'b00000000000000000000100000001011;
assign LUT_1[39609] = 32'b11111111111111111001110010000111;
assign LUT_1[39610] = 32'b11111111111111111100001110011100;
assign LUT_1[39611] = 32'b11111111111111110101100000011000;
assign LUT_1[39612] = 32'b00000000000000001000011001100010;
assign LUT_1[39613] = 32'b00000000000000000001101011011110;
assign LUT_1[39614] = 32'b00000000000000000100000111110011;
assign LUT_1[39615] = 32'b11111111111111111101011001101111;
assign LUT_1[39616] = 32'b00000000000000000000011001011101;
assign LUT_1[39617] = 32'b11111111111111111001101011011001;
assign LUT_1[39618] = 32'b11111111111111111100000111101110;
assign LUT_1[39619] = 32'b11111111111111110101011001101010;
assign LUT_1[39620] = 32'b00000000000000001000010010110100;
assign LUT_1[39621] = 32'b00000000000000000001100100110000;
assign LUT_1[39622] = 32'b00000000000000000100000001000101;
assign LUT_1[39623] = 32'b11111111111111111101010011000001;
assign LUT_1[39624] = 32'b11111111111111111111100111010010;
assign LUT_1[39625] = 32'b11111111111111111000111001001110;
assign LUT_1[39626] = 32'b11111111111111111011010101100011;
assign LUT_1[39627] = 32'b11111111111111110100100111011111;
assign LUT_1[39628] = 32'b00000000000000000111100000101001;
assign LUT_1[39629] = 32'b00000000000000000000110010100101;
assign LUT_1[39630] = 32'b00000000000000000011001110111010;
assign LUT_1[39631] = 32'b11111111111111111100100000110110;
assign LUT_1[39632] = 32'b00000000000000000010010100111111;
assign LUT_1[39633] = 32'b11111111111111111011100110111011;
assign LUT_1[39634] = 32'b11111111111111111110000011010000;
assign LUT_1[39635] = 32'b11111111111111110111010101001100;
assign LUT_1[39636] = 32'b00000000000000001010001110010110;
assign LUT_1[39637] = 32'b00000000000000000011100000010010;
assign LUT_1[39638] = 32'b00000000000000000101111100100111;
assign LUT_1[39639] = 32'b11111111111111111111001110100011;
assign LUT_1[39640] = 32'b00000000000000000001100010110100;
assign LUT_1[39641] = 32'b11111111111111111010110100110000;
assign LUT_1[39642] = 32'b11111111111111111101010001000101;
assign LUT_1[39643] = 32'b11111111111111110110100011000001;
assign LUT_1[39644] = 32'b00000000000000001001011100001011;
assign LUT_1[39645] = 32'b00000000000000000010101110000111;
assign LUT_1[39646] = 32'b00000000000000000101001010011100;
assign LUT_1[39647] = 32'b11111111111111111110011100011000;
assign LUT_1[39648] = 32'b00000000000000000001010100011100;
assign LUT_1[39649] = 32'b11111111111111111010100110011000;
assign LUT_1[39650] = 32'b11111111111111111101000010101101;
assign LUT_1[39651] = 32'b11111111111111110110010100101001;
assign LUT_1[39652] = 32'b00000000000000001001001101110011;
assign LUT_1[39653] = 32'b00000000000000000010011111101111;
assign LUT_1[39654] = 32'b00000000000000000100111100000100;
assign LUT_1[39655] = 32'b11111111111111111110001110000000;
assign LUT_1[39656] = 32'b00000000000000000000100010010001;
assign LUT_1[39657] = 32'b11111111111111111001110100001101;
assign LUT_1[39658] = 32'b11111111111111111100010000100010;
assign LUT_1[39659] = 32'b11111111111111110101100010011110;
assign LUT_1[39660] = 32'b00000000000000001000011011101000;
assign LUT_1[39661] = 32'b00000000000000000001101101100100;
assign LUT_1[39662] = 32'b00000000000000000100001001111001;
assign LUT_1[39663] = 32'b11111111111111111101011011110101;
assign LUT_1[39664] = 32'b00000000000000000011001111111110;
assign LUT_1[39665] = 32'b11111111111111111100100001111010;
assign LUT_1[39666] = 32'b11111111111111111110111110001111;
assign LUT_1[39667] = 32'b11111111111111111000010000001011;
assign LUT_1[39668] = 32'b00000000000000001011001001010101;
assign LUT_1[39669] = 32'b00000000000000000100011011010001;
assign LUT_1[39670] = 32'b00000000000000000110110111100110;
assign LUT_1[39671] = 32'b00000000000000000000001001100010;
assign LUT_1[39672] = 32'b00000000000000000010011101110011;
assign LUT_1[39673] = 32'b11111111111111111011101111101111;
assign LUT_1[39674] = 32'b11111111111111111110001100000100;
assign LUT_1[39675] = 32'b11111111111111110111011110000000;
assign LUT_1[39676] = 32'b00000000000000001010010111001010;
assign LUT_1[39677] = 32'b00000000000000000011101001000110;
assign LUT_1[39678] = 32'b00000000000000000110000101011011;
assign LUT_1[39679] = 32'b11111111111111111111010111010111;
assign LUT_1[39680] = 32'b11111111111111111001001111111110;
assign LUT_1[39681] = 32'b11111111111111110010100001111010;
assign LUT_1[39682] = 32'b11111111111111110100111110001111;
assign LUT_1[39683] = 32'b11111111111111101110010000001011;
assign LUT_1[39684] = 32'b00000000000000000001001001010101;
assign LUT_1[39685] = 32'b11111111111111111010011011010001;
assign LUT_1[39686] = 32'b11111111111111111100110111100110;
assign LUT_1[39687] = 32'b11111111111111110110001001100010;
assign LUT_1[39688] = 32'b11111111111111111000011101110011;
assign LUT_1[39689] = 32'b11111111111111110001101111101111;
assign LUT_1[39690] = 32'b11111111111111110100001100000100;
assign LUT_1[39691] = 32'b11111111111111101101011110000000;
assign LUT_1[39692] = 32'b00000000000000000000010111001010;
assign LUT_1[39693] = 32'b11111111111111111001101001000110;
assign LUT_1[39694] = 32'b11111111111111111100000101011011;
assign LUT_1[39695] = 32'b11111111111111110101010111010111;
assign LUT_1[39696] = 32'b11111111111111111011001011100000;
assign LUT_1[39697] = 32'b11111111111111110100011101011100;
assign LUT_1[39698] = 32'b11111111111111110110111001110001;
assign LUT_1[39699] = 32'b11111111111111110000001011101101;
assign LUT_1[39700] = 32'b00000000000000000011000100110111;
assign LUT_1[39701] = 32'b11111111111111111100010110110011;
assign LUT_1[39702] = 32'b11111111111111111110110011001000;
assign LUT_1[39703] = 32'b11111111111111111000000101000100;
assign LUT_1[39704] = 32'b11111111111111111010011001010101;
assign LUT_1[39705] = 32'b11111111111111110011101011010001;
assign LUT_1[39706] = 32'b11111111111111110110000111100110;
assign LUT_1[39707] = 32'b11111111111111101111011001100010;
assign LUT_1[39708] = 32'b00000000000000000010010010101100;
assign LUT_1[39709] = 32'b11111111111111111011100100101000;
assign LUT_1[39710] = 32'b11111111111111111110000000111101;
assign LUT_1[39711] = 32'b11111111111111110111010010111001;
assign LUT_1[39712] = 32'b11111111111111111010001010111101;
assign LUT_1[39713] = 32'b11111111111111110011011100111001;
assign LUT_1[39714] = 32'b11111111111111110101111001001110;
assign LUT_1[39715] = 32'b11111111111111101111001011001010;
assign LUT_1[39716] = 32'b00000000000000000010000100010100;
assign LUT_1[39717] = 32'b11111111111111111011010110010000;
assign LUT_1[39718] = 32'b11111111111111111101110010100101;
assign LUT_1[39719] = 32'b11111111111111110111000100100001;
assign LUT_1[39720] = 32'b11111111111111111001011000110010;
assign LUT_1[39721] = 32'b11111111111111110010101010101110;
assign LUT_1[39722] = 32'b11111111111111110101000111000011;
assign LUT_1[39723] = 32'b11111111111111101110011000111111;
assign LUT_1[39724] = 32'b00000000000000000001010010001001;
assign LUT_1[39725] = 32'b11111111111111111010100100000101;
assign LUT_1[39726] = 32'b11111111111111111101000000011010;
assign LUT_1[39727] = 32'b11111111111111110110010010010110;
assign LUT_1[39728] = 32'b11111111111111111100000110011111;
assign LUT_1[39729] = 32'b11111111111111110101011000011011;
assign LUT_1[39730] = 32'b11111111111111110111110100110000;
assign LUT_1[39731] = 32'b11111111111111110001000110101100;
assign LUT_1[39732] = 32'b00000000000000000011111111110110;
assign LUT_1[39733] = 32'b11111111111111111101010001110010;
assign LUT_1[39734] = 32'b11111111111111111111101110000111;
assign LUT_1[39735] = 32'b11111111111111111001000000000011;
assign LUT_1[39736] = 32'b11111111111111111011010100010100;
assign LUT_1[39737] = 32'b11111111111111110100100110010000;
assign LUT_1[39738] = 32'b11111111111111110111000010100101;
assign LUT_1[39739] = 32'b11111111111111110000010100100001;
assign LUT_1[39740] = 32'b00000000000000000011001101101011;
assign LUT_1[39741] = 32'b11111111111111111100011111100111;
assign LUT_1[39742] = 32'b11111111111111111110111011111100;
assign LUT_1[39743] = 32'b11111111111111111000001101111000;
assign LUT_1[39744] = 32'b11111111111111111011001101100110;
assign LUT_1[39745] = 32'b11111111111111110100011111100010;
assign LUT_1[39746] = 32'b11111111111111110110111011110111;
assign LUT_1[39747] = 32'b11111111111111110000001101110011;
assign LUT_1[39748] = 32'b00000000000000000011000110111101;
assign LUT_1[39749] = 32'b11111111111111111100011000111001;
assign LUT_1[39750] = 32'b11111111111111111110110101001110;
assign LUT_1[39751] = 32'b11111111111111111000000111001010;
assign LUT_1[39752] = 32'b11111111111111111010011011011011;
assign LUT_1[39753] = 32'b11111111111111110011101101010111;
assign LUT_1[39754] = 32'b11111111111111110110001001101100;
assign LUT_1[39755] = 32'b11111111111111101111011011101000;
assign LUT_1[39756] = 32'b00000000000000000010010100110010;
assign LUT_1[39757] = 32'b11111111111111111011100110101110;
assign LUT_1[39758] = 32'b11111111111111111110000011000011;
assign LUT_1[39759] = 32'b11111111111111110111010100111111;
assign LUT_1[39760] = 32'b11111111111111111101001001001000;
assign LUT_1[39761] = 32'b11111111111111110110011011000100;
assign LUT_1[39762] = 32'b11111111111111111000110111011001;
assign LUT_1[39763] = 32'b11111111111111110010001001010101;
assign LUT_1[39764] = 32'b00000000000000000101000010011111;
assign LUT_1[39765] = 32'b11111111111111111110010100011011;
assign LUT_1[39766] = 32'b00000000000000000000110000110000;
assign LUT_1[39767] = 32'b11111111111111111010000010101100;
assign LUT_1[39768] = 32'b11111111111111111100010110111101;
assign LUT_1[39769] = 32'b11111111111111110101101000111001;
assign LUT_1[39770] = 32'b11111111111111111000000101001110;
assign LUT_1[39771] = 32'b11111111111111110001010111001010;
assign LUT_1[39772] = 32'b00000000000000000100010000010100;
assign LUT_1[39773] = 32'b11111111111111111101100010010000;
assign LUT_1[39774] = 32'b11111111111111111111111110100101;
assign LUT_1[39775] = 32'b11111111111111111001010000100001;
assign LUT_1[39776] = 32'b11111111111111111100001000100101;
assign LUT_1[39777] = 32'b11111111111111110101011010100001;
assign LUT_1[39778] = 32'b11111111111111110111110110110110;
assign LUT_1[39779] = 32'b11111111111111110001001000110010;
assign LUT_1[39780] = 32'b00000000000000000100000001111100;
assign LUT_1[39781] = 32'b11111111111111111101010011111000;
assign LUT_1[39782] = 32'b11111111111111111111110000001101;
assign LUT_1[39783] = 32'b11111111111111111001000010001001;
assign LUT_1[39784] = 32'b11111111111111111011010110011010;
assign LUT_1[39785] = 32'b11111111111111110100101000010110;
assign LUT_1[39786] = 32'b11111111111111110111000100101011;
assign LUT_1[39787] = 32'b11111111111111110000010110100111;
assign LUT_1[39788] = 32'b00000000000000000011001111110001;
assign LUT_1[39789] = 32'b11111111111111111100100001101101;
assign LUT_1[39790] = 32'b11111111111111111110111110000010;
assign LUT_1[39791] = 32'b11111111111111111000001111111110;
assign LUT_1[39792] = 32'b11111111111111111110000100000111;
assign LUT_1[39793] = 32'b11111111111111110111010110000011;
assign LUT_1[39794] = 32'b11111111111111111001110010011000;
assign LUT_1[39795] = 32'b11111111111111110011000100010100;
assign LUT_1[39796] = 32'b00000000000000000101111101011110;
assign LUT_1[39797] = 32'b11111111111111111111001111011010;
assign LUT_1[39798] = 32'b00000000000000000001101011101111;
assign LUT_1[39799] = 32'b11111111111111111010111101101011;
assign LUT_1[39800] = 32'b11111111111111111101010001111100;
assign LUT_1[39801] = 32'b11111111111111110110100011111000;
assign LUT_1[39802] = 32'b11111111111111111001000000001101;
assign LUT_1[39803] = 32'b11111111111111110010010010001001;
assign LUT_1[39804] = 32'b00000000000000000101001011010011;
assign LUT_1[39805] = 32'b11111111111111111110011101001111;
assign LUT_1[39806] = 32'b00000000000000000000111001100100;
assign LUT_1[39807] = 32'b11111111111111111010001011100000;
assign LUT_1[39808] = 32'b11111111111111111100010000000001;
assign LUT_1[39809] = 32'b11111111111111110101100001111101;
assign LUT_1[39810] = 32'b11111111111111110111111110010010;
assign LUT_1[39811] = 32'b11111111111111110001010000001110;
assign LUT_1[39812] = 32'b00000000000000000100001001011000;
assign LUT_1[39813] = 32'b11111111111111111101011011010100;
assign LUT_1[39814] = 32'b11111111111111111111110111101001;
assign LUT_1[39815] = 32'b11111111111111111001001001100101;
assign LUT_1[39816] = 32'b11111111111111111011011101110110;
assign LUT_1[39817] = 32'b11111111111111110100101111110010;
assign LUT_1[39818] = 32'b11111111111111110111001100000111;
assign LUT_1[39819] = 32'b11111111111111110000011110000011;
assign LUT_1[39820] = 32'b00000000000000000011010111001101;
assign LUT_1[39821] = 32'b11111111111111111100101001001001;
assign LUT_1[39822] = 32'b11111111111111111111000101011110;
assign LUT_1[39823] = 32'b11111111111111111000010111011010;
assign LUT_1[39824] = 32'b11111111111111111110001011100011;
assign LUT_1[39825] = 32'b11111111111111110111011101011111;
assign LUT_1[39826] = 32'b11111111111111111001111001110100;
assign LUT_1[39827] = 32'b11111111111111110011001011110000;
assign LUT_1[39828] = 32'b00000000000000000110000100111010;
assign LUT_1[39829] = 32'b11111111111111111111010110110110;
assign LUT_1[39830] = 32'b00000000000000000001110011001011;
assign LUT_1[39831] = 32'b11111111111111111011000101000111;
assign LUT_1[39832] = 32'b11111111111111111101011001011000;
assign LUT_1[39833] = 32'b11111111111111110110101011010100;
assign LUT_1[39834] = 32'b11111111111111111001000111101001;
assign LUT_1[39835] = 32'b11111111111111110010011001100101;
assign LUT_1[39836] = 32'b00000000000000000101010010101111;
assign LUT_1[39837] = 32'b11111111111111111110100100101011;
assign LUT_1[39838] = 32'b00000000000000000001000001000000;
assign LUT_1[39839] = 32'b11111111111111111010010010111100;
assign LUT_1[39840] = 32'b11111111111111111101001011000000;
assign LUT_1[39841] = 32'b11111111111111110110011100111100;
assign LUT_1[39842] = 32'b11111111111111111000111001010001;
assign LUT_1[39843] = 32'b11111111111111110010001011001101;
assign LUT_1[39844] = 32'b00000000000000000101000100010111;
assign LUT_1[39845] = 32'b11111111111111111110010110010011;
assign LUT_1[39846] = 32'b00000000000000000000110010101000;
assign LUT_1[39847] = 32'b11111111111111111010000100100100;
assign LUT_1[39848] = 32'b11111111111111111100011000110101;
assign LUT_1[39849] = 32'b11111111111111110101101010110001;
assign LUT_1[39850] = 32'b11111111111111111000000111000110;
assign LUT_1[39851] = 32'b11111111111111110001011001000010;
assign LUT_1[39852] = 32'b00000000000000000100010010001100;
assign LUT_1[39853] = 32'b11111111111111111101100100001000;
assign LUT_1[39854] = 32'b00000000000000000000000000011101;
assign LUT_1[39855] = 32'b11111111111111111001010010011001;
assign LUT_1[39856] = 32'b11111111111111111111000110100010;
assign LUT_1[39857] = 32'b11111111111111111000011000011110;
assign LUT_1[39858] = 32'b11111111111111111010110100110011;
assign LUT_1[39859] = 32'b11111111111111110100000110101111;
assign LUT_1[39860] = 32'b00000000000000000110111111111001;
assign LUT_1[39861] = 32'b00000000000000000000010001110101;
assign LUT_1[39862] = 32'b00000000000000000010101110001010;
assign LUT_1[39863] = 32'b11111111111111111100000000000110;
assign LUT_1[39864] = 32'b11111111111111111110010100010111;
assign LUT_1[39865] = 32'b11111111111111110111100110010011;
assign LUT_1[39866] = 32'b11111111111111111010000010101000;
assign LUT_1[39867] = 32'b11111111111111110011010100100100;
assign LUT_1[39868] = 32'b00000000000000000110001101101110;
assign LUT_1[39869] = 32'b11111111111111111111011111101010;
assign LUT_1[39870] = 32'b00000000000000000001111011111111;
assign LUT_1[39871] = 32'b11111111111111111011001101111011;
assign LUT_1[39872] = 32'b11111111111111111110001101101001;
assign LUT_1[39873] = 32'b11111111111111110111011111100101;
assign LUT_1[39874] = 32'b11111111111111111001111011111010;
assign LUT_1[39875] = 32'b11111111111111110011001101110110;
assign LUT_1[39876] = 32'b00000000000000000110000111000000;
assign LUT_1[39877] = 32'b11111111111111111111011000111100;
assign LUT_1[39878] = 32'b00000000000000000001110101010001;
assign LUT_1[39879] = 32'b11111111111111111011000111001101;
assign LUT_1[39880] = 32'b11111111111111111101011011011110;
assign LUT_1[39881] = 32'b11111111111111110110101101011010;
assign LUT_1[39882] = 32'b11111111111111111001001001101111;
assign LUT_1[39883] = 32'b11111111111111110010011011101011;
assign LUT_1[39884] = 32'b00000000000000000101010100110101;
assign LUT_1[39885] = 32'b11111111111111111110100110110001;
assign LUT_1[39886] = 32'b00000000000000000001000011000110;
assign LUT_1[39887] = 32'b11111111111111111010010101000010;
assign LUT_1[39888] = 32'b00000000000000000000001001001011;
assign LUT_1[39889] = 32'b11111111111111111001011011000111;
assign LUT_1[39890] = 32'b11111111111111111011110111011100;
assign LUT_1[39891] = 32'b11111111111111110101001001011000;
assign LUT_1[39892] = 32'b00000000000000001000000010100010;
assign LUT_1[39893] = 32'b00000000000000000001010100011110;
assign LUT_1[39894] = 32'b00000000000000000011110000110011;
assign LUT_1[39895] = 32'b11111111111111111101000010101111;
assign LUT_1[39896] = 32'b11111111111111111111010111000000;
assign LUT_1[39897] = 32'b11111111111111111000101000111100;
assign LUT_1[39898] = 32'b11111111111111111011000101010001;
assign LUT_1[39899] = 32'b11111111111111110100010111001101;
assign LUT_1[39900] = 32'b00000000000000000111010000010111;
assign LUT_1[39901] = 32'b00000000000000000000100010010011;
assign LUT_1[39902] = 32'b00000000000000000010111110101000;
assign LUT_1[39903] = 32'b11111111111111111100010000100100;
assign LUT_1[39904] = 32'b11111111111111111111001000101000;
assign LUT_1[39905] = 32'b11111111111111111000011010100100;
assign LUT_1[39906] = 32'b11111111111111111010110110111001;
assign LUT_1[39907] = 32'b11111111111111110100001000110101;
assign LUT_1[39908] = 32'b00000000000000000111000001111111;
assign LUT_1[39909] = 32'b00000000000000000000010011111011;
assign LUT_1[39910] = 32'b00000000000000000010110000010000;
assign LUT_1[39911] = 32'b11111111111111111100000010001100;
assign LUT_1[39912] = 32'b11111111111111111110010110011101;
assign LUT_1[39913] = 32'b11111111111111110111101000011001;
assign LUT_1[39914] = 32'b11111111111111111010000100101110;
assign LUT_1[39915] = 32'b11111111111111110011010110101010;
assign LUT_1[39916] = 32'b00000000000000000110001111110100;
assign LUT_1[39917] = 32'b11111111111111111111100001110000;
assign LUT_1[39918] = 32'b00000000000000000001111110000101;
assign LUT_1[39919] = 32'b11111111111111111011010000000001;
assign LUT_1[39920] = 32'b00000000000000000001000100001010;
assign LUT_1[39921] = 32'b11111111111111111010010110000110;
assign LUT_1[39922] = 32'b11111111111111111100110010011011;
assign LUT_1[39923] = 32'b11111111111111110110000100010111;
assign LUT_1[39924] = 32'b00000000000000001000111101100001;
assign LUT_1[39925] = 32'b00000000000000000010001111011101;
assign LUT_1[39926] = 32'b00000000000000000100101011110010;
assign LUT_1[39927] = 32'b11111111111111111101111101101110;
assign LUT_1[39928] = 32'b00000000000000000000010001111111;
assign LUT_1[39929] = 32'b11111111111111111001100011111011;
assign LUT_1[39930] = 32'b11111111111111111100000000010000;
assign LUT_1[39931] = 32'b11111111111111110101010010001100;
assign LUT_1[39932] = 32'b00000000000000001000001011010110;
assign LUT_1[39933] = 32'b00000000000000000001011101010010;
assign LUT_1[39934] = 32'b00000000000000000011111001100111;
assign LUT_1[39935] = 32'b11111111111111111101001011100011;
assign LUT_1[39936] = 32'b00000000000000001000000100000101;
assign LUT_1[39937] = 32'b00000000000000000001010110000001;
assign LUT_1[39938] = 32'b00000000000000000011110010010110;
assign LUT_1[39939] = 32'b11111111111111111101000100010010;
assign LUT_1[39940] = 32'b00000000000000001111111101011100;
assign LUT_1[39941] = 32'b00000000000000001001001111011000;
assign LUT_1[39942] = 32'b00000000000000001011101011101101;
assign LUT_1[39943] = 32'b00000000000000000100111101101001;
assign LUT_1[39944] = 32'b00000000000000000111010001111010;
assign LUT_1[39945] = 32'b00000000000000000000100011110110;
assign LUT_1[39946] = 32'b00000000000000000011000000001011;
assign LUT_1[39947] = 32'b11111111111111111100010010000111;
assign LUT_1[39948] = 32'b00000000000000001111001011010001;
assign LUT_1[39949] = 32'b00000000000000001000011101001101;
assign LUT_1[39950] = 32'b00000000000000001010111001100010;
assign LUT_1[39951] = 32'b00000000000000000100001011011110;
assign LUT_1[39952] = 32'b00000000000000001001111111100111;
assign LUT_1[39953] = 32'b00000000000000000011010001100011;
assign LUT_1[39954] = 32'b00000000000000000101101101111000;
assign LUT_1[39955] = 32'b11111111111111111110111111110100;
assign LUT_1[39956] = 32'b00000000000000010001111000111110;
assign LUT_1[39957] = 32'b00000000000000001011001010111010;
assign LUT_1[39958] = 32'b00000000000000001101100111001111;
assign LUT_1[39959] = 32'b00000000000000000110111001001011;
assign LUT_1[39960] = 32'b00000000000000001001001101011100;
assign LUT_1[39961] = 32'b00000000000000000010011111011000;
assign LUT_1[39962] = 32'b00000000000000000100111011101101;
assign LUT_1[39963] = 32'b11111111111111111110001101101001;
assign LUT_1[39964] = 32'b00000000000000010001000110110011;
assign LUT_1[39965] = 32'b00000000000000001010011000101111;
assign LUT_1[39966] = 32'b00000000000000001100110101000100;
assign LUT_1[39967] = 32'b00000000000000000110000111000000;
assign LUT_1[39968] = 32'b00000000000000001000111111000100;
assign LUT_1[39969] = 32'b00000000000000000010010001000000;
assign LUT_1[39970] = 32'b00000000000000000100101101010101;
assign LUT_1[39971] = 32'b11111111111111111101111111010001;
assign LUT_1[39972] = 32'b00000000000000010000111000011011;
assign LUT_1[39973] = 32'b00000000000000001010001010010111;
assign LUT_1[39974] = 32'b00000000000000001100100110101100;
assign LUT_1[39975] = 32'b00000000000000000101111000101000;
assign LUT_1[39976] = 32'b00000000000000001000001100111001;
assign LUT_1[39977] = 32'b00000000000000000001011110110101;
assign LUT_1[39978] = 32'b00000000000000000011111011001010;
assign LUT_1[39979] = 32'b11111111111111111101001101000110;
assign LUT_1[39980] = 32'b00000000000000010000000110010000;
assign LUT_1[39981] = 32'b00000000000000001001011000001100;
assign LUT_1[39982] = 32'b00000000000000001011110100100001;
assign LUT_1[39983] = 32'b00000000000000000101000110011101;
assign LUT_1[39984] = 32'b00000000000000001010111010100110;
assign LUT_1[39985] = 32'b00000000000000000100001100100010;
assign LUT_1[39986] = 32'b00000000000000000110101000110111;
assign LUT_1[39987] = 32'b11111111111111111111111010110011;
assign LUT_1[39988] = 32'b00000000000000010010110011111101;
assign LUT_1[39989] = 32'b00000000000000001100000101111001;
assign LUT_1[39990] = 32'b00000000000000001110100010001110;
assign LUT_1[39991] = 32'b00000000000000000111110100001010;
assign LUT_1[39992] = 32'b00000000000000001010001000011011;
assign LUT_1[39993] = 32'b00000000000000000011011010010111;
assign LUT_1[39994] = 32'b00000000000000000101110110101100;
assign LUT_1[39995] = 32'b11111111111111111111001000101000;
assign LUT_1[39996] = 32'b00000000000000010010000001110010;
assign LUT_1[39997] = 32'b00000000000000001011010011101110;
assign LUT_1[39998] = 32'b00000000000000001101110000000011;
assign LUT_1[39999] = 32'b00000000000000000111000001111111;
assign LUT_1[40000] = 32'b00000000000000001010000001101101;
assign LUT_1[40001] = 32'b00000000000000000011010011101001;
assign LUT_1[40002] = 32'b00000000000000000101101111111110;
assign LUT_1[40003] = 32'b11111111111111111111000001111010;
assign LUT_1[40004] = 32'b00000000000000010001111011000100;
assign LUT_1[40005] = 32'b00000000000000001011001101000000;
assign LUT_1[40006] = 32'b00000000000000001101101001010101;
assign LUT_1[40007] = 32'b00000000000000000110111011010001;
assign LUT_1[40008] = 32'b00000000000000001001001111100010;
assign LUT_1[40009] = 32'b00000000000000000010100001011110;
assign LUT_1[40010] = 32'b00000000000000000100111101110011;
assign LUT_1[40011] = 32'b11111111111111111110001111101111;
assign LUT_1[40012] = 32'b00000000000000010001001000111001;
assign LUT_1[40013] = 32'b00000000000000001010011010110101;
assign LUT_1[40014] = 32'b00000000000000001100110111001010;
assign LUT_1[40015] = 32'b00000000000000000110001001000110;
assign LUT_1[40016] = 32'b00000000000000001011111101001111;
assign LUT_1[40017] = 32'b00000000000000000101001111001011;
assign LUT_1[40018] = 32'b00000000000000000111101011100000;
assign LUT_1[40019] = 32'b00000000000000000000111101011100;
assign LUT_1[40020] = 32'b00000000000000010011110110100110;
assign LUT_1[40021] = 32'b00000000000000001101001000100010;
assign LUT_1[40022] = 32'b00000000000000001111100100110111;
assign LUT_1[40023] = 32'b00000000000000001000110110110011;
assign LUT_1[40024] = 32'b00000000000000001011001011000100;
assign LUT_1[40025] = 32'b00000000000000000100011101000000;
assign LUT_1[40026] = 32'b00000000000000000110111001010101;
assign LUT_1[40027] = 32'b00000000000000000000001011010001;
assign LUT_1[40028] = 32'b00000000000000010011000100011011;
assign LUT_1[40029] = 32'b00000000000000001100010110010111;
assign LUT_1[40030] = 32'b00000000000000001110110010101100;
assign LUT_1[40031] = 32'b00000000000000001000000100101000;
assign LUT_1[40032] = 32'b00000000000000001010111100101100;
assign LUT_1[40033] = 32'b00000000000000000100001110101000;
assign LUT_1[40034] = 32'b00000000000000000110101010111101;
assign LUT_1[40035] = 32'b11111111111111111111111100111001;
assign LUT_1[40036] = 32'b00000000000000010010110110000011;
assign LUT_1[40037] = 32'b00000000000000001100000111111111;
assign LUT_1[40038] = 32'b00000000000000001110100100010100;
assign LUT_1[40039] = 32'b00000000000000000111110110010000;
assign LUT_1[40040] = 32'b00000000000000001010001010100001;
assign LUT_1[40041] = 32'b00000000000000000011011100011101;
assign LUT_1[40042] = 32'b00000000000000000101111000110010;
assign LUT_1[40043] = 32'b11111111111111111111001010101110;
assign LUT_1[40044] = 32'b00000000000000010010000011111000;
assign LUT_1[40045] = 32'b00000000000000001011010101110100;
assign LUT_1[40046] = 32'b00000000000000001101110010001001;
assign LUT_1[40047] = 32'b00000000000000000111000100000101;
assign LUT_1[40048] = 32'b00000000000000001100111000001110;
assign LUT_1[40049] = 32'b00000000000000000110001010001010;
assign LUT_1[40050] = 32'b00000000000000001000100110011111;
assign LUT_1[40051] = 32'b00000000000000000001111000011011;
assign LUT_1[40052] = 32'b00000000000000010100110001100101;
assign LUT_1[40053] = 32'b00000000000000001110000011100001;
assign LUT_1[40054] = 32'b00000000000000010000011111110110;
assign LUT_1[40055] = 32'b00000000000000001001110001110010;
assign LUT_1[40056] = 32'b00000000000000001100000110000011;
assign LUT_1[40057] = 32'b00000000000000000101010111111111;
assign LUT_1[40058] = 32'b00000000000000000111110100010100;
assign LUT_1[40059] = 32'b00000000000000000001000110010000;
assign LUT_1[40060] = 32'b00000000000000010011111111011010;
assign LUT_1[40061] = 32'b00000000000000001101010001010110;
assign LUT_1[40062] = 32'b00000000000000001111101101101011;
assign LUT_1[40063] = 32'b00000000000000001000111111100111;
assign LUT_1[40064] = 32'b00000000000000001011000100001000;
assign LUT_1[40065] = 32'b00000000000000000100010110000100;
assign LUT_1[40066] = 32'b00000000000000000110110010011001;
assign LUT_1[40067] = 32'b00000000000000000000000100010101;
assign LUT_1[40068] = 32'b00000000000000010010111101011111;
assign LUT_1[40069] = 32'b00000000000000001100001111011011;
assign LUT_1[40070] = 32'b00000000000000001110101011110000;
assign LUT_1[40071] = 32'b00000000000000000111111101101100;
assign LUT_1[40072] = 32'b00000000000000001010010001111101;
assign LUT_1[40073] = 32'b00000000000000000011100011111001;
assign LUT_1[40074] = 32'b00000000000000000110000000001110;
assign LUT_1[40075] = 32'b11111111111111111111010010001010;
assign LUT_1[40076] = 32'b00000000000000010010001011010100;
assign LUT_1[40077] = 32'b00000000000000001011011101010000;
assign LUT_1[40078] = 32'b00000000000000001101111001100101;
assign LUT_1[40079] = 32'b00000000000000000111001011100001;
assign LUT_1[40080] = 32'b00000000000000001100111111101010;
assign LUT_1[40081] = 32'b00000000000000000110010001100110;
assign LUT_1[40082] = 32'b00000000000000001000101101111011;
assign LUT_1[40083] = 32'b00000000000000000001111111110111;
assign LUT_1[40084] = 32'b00000000000000010100111001000001;
assign LUT_1[40085] = 32'b00000000000000001110001010111101;
assign LUT_1[40086] = 32'b00000000000000010000100111010010;
assign LUT_1[40087] = 32'b00000000000000001001111001001110;
assign LUT_1[40088] = 32'b00000000000000001100001101011111;
assign LUT_1[40089] = 32'b00000000000000000101011111011011;
assign LUT_1[40090] = 32'b00000000000000000111111011110000;
assign LUT_1[40091] = 32'b00000000000000000001001101101100;
assign LUT_1[40092] = 32'b00000000000000010100000110110110;
assign LUT_1[40093] = 32'b00000000000000001101011000110010;
assign LUT_1[40094] = 32'b00000000000000001111110101000111;
assign LUT_1[40095] = 32'b00000000000000001001000111000011;
assign LUT_1[40096] = 32'b00000000000000001011111111000111;
assign LUT_1[40097] = 32'b00000000000000000101010001000011;
assign LUT_1[40098] = 32'b00000000000000000111101101011000;
assign LUT_1[40099] = 32'b00000000000000000000111111010100;
assign LUT_1[40100] = 32'b00000000000000010011111000011110;
assign LUT_1[40101] = 32'b00000000000000001101001010011010;
assign LUT_1[40102] = 32'b00000000000000001111100110101111;
assign LUT_1[40103] = 32'b00000000000000001000111000101011;
assign LUT_1[40104] = 32'b00000000000000001011001100111100;
assign LUT_1[40105] = 32'b00000000000000000100011110111000;
assign LUT_1[40106] = 32'b00000000000000000110111011001101;
assign LUT_1[40107] = 32'b00000000000000000000001101001001;
assign LUT_1[40108] = 32'b00000000000000010011000110010011;
assign LUT_1[40109] = 32'b00000000000000001100011000001111;
assign LUT_1[40110] = 32'b00000000000000001110110100100100;
assign LUT_1[40111] = 32'b00000000000000001000000110100000;
assign LUT_1[40112] = 32'b00000000000000001101111010101001;
assign LUT_1[40113] = 32'b00000000000000000111001100100101;
assign LUT_1[40114] = 32'b00000000000000001001101000111010;
assign LUT_1[40115] = 32'b00000000000000000010111010110110;
assign LUT_1[40116] = 32'b00000000000000010101110100000000;
assign LUT_1[40117] = 32'b00000000000000001111000101111100;
assign LUT_1[40118] = 32'b00000000000000010001100010010001;
assign LUT_1[40119] = 32'b00000000000000001010110100001101;
assign LUT_1[40120] = 32'b00000000000000001101001000011110;
assign LUT_1[40121] = 32'b00000000000000000110011010011010;
assign LUT_1[40122] = 32'b00000000000000001000110110101111;
assign LUT_1[40123] = 32'b00000000000000000010001000101011;
assign LUT_1[40124] = 32'b00000000000000010101000001110101;
assign LUT_1[40125] = 32'b00000000000000001110010011110001;
assign LUT_1[40126] = 32'b00000000000000010000110000000110;
assign LUT_1[40127] = 32'b00000000000000001010000010000010;
assign LUT_1[40128] = 32'b00000000000000001101000001110000;
assign LUT_1[40129] = 32'b00000000000000000110010011101100;
assign LUT_1[40130] = 32'b00000000000000001000110000000001;
assign LUT_1[40131] = 32'b00000000000000000010000001111101;
assign LUT_1[40132] = 32'b00000000000000010100111011000111;
assign LUT_1[40133] = 32'b00000000000000001110001101000011;
assign LUT_1[40134] = 32'b00000000000000010000101001011000;
assign LUT_1[40135] = 32'b00000000000000001001111011010100;
assign LUT_1[40136] = 32'b00000000000000001100001111100101;
assign LUT_1[40137] = 32'b00000000000000000101100001100001;
assign LUT_1[40138] = 32'b00000000000000000111111101110110;
assign LUT_1[40139] = 32'b00000000000000000001001111110010;
assign LUT_1[40140] = 32'b00000000000000010100001000111100;
assign LUT_1[40141] = 32'b00000000000000001101011010111000;
assign LUT_1[40142] = 32'b00000000000000001111110111001101;
assign LUT_1[40143] = 32'b00000000000000001001001001001001;
assign LUT_1[40144] = 32'b00000000000000001110111101010010;
assign LUT_1[40145] = 32'b00000000000000001000001111001110;
assign LUT_1[40146] = 32'b00000000000000001010101011100011;
assign LUT_1[40147] = 32'b00000000000000000011111101011111;
assign LUT_1[40148] = 32'b00000000000000010110110110101001;
assign LUT_1[40149] = 32'b00000000000000010000001000100101;
assign LUT_1[40150] = 32'b00000000000000010010100100111010;
assign LUT_1[40151] = 32'b00000000000000001011110110110110;
assign LUT_1[40152] = 32'b00000000000000001110001011000111;
assign LUT_1[40153] = 32'b00000000000000000111011101000011;
assign LUT_1[40154] = 32'b00000000000000001001111001011000;
assign LUT_1[40155] = 32'b00000000000000000011001011010100;
assign LUT_1[40156] = 32'b00000000000000010110000100011110;
assign LUT_1[40157] = 32'b00000000000000001111010110011010;
assign LUT_1[40158] = 32'b00000000000000010001110010101111;
assign LUT_1[40159] = 32'b00000000000000001011000100101011;
assign LUT_1[40160] = 32'b00000000000000001101111100101111;
assign LUT_1[40161] = 32'b00000000000000000111001110101011;
assign LUT_1[40162] = 32'b00000000000000001001101011000000;
assign LUT_1[40163] = 32'b00000000000000000010111100111100;
assign LUT_1[40164] = 32'b00000000000000010101110110000110;
assign LUT_1[40165] = 32'b00000000000000001111001000000010;
assign LUT_1[40166] = 32'b00000000000000010001100100010111;
assign LUT_1[40167] = 32'b00000000000000001010110110010011;
assign LUT_1[40168] = 32'b00000000000000001101001010100100;
assign LUT_1[40169] = 32'b00000000000000000110011100100000;
assign LUT_1[40170] = 32'b00000000000000001000111000110101;
assign LUT_1[40171] = 32'b00000000000000000010001010110001;
assign LUT_1[40172] = 32'b00000000000000010101000011111011;
assign LUT_1[40173] = 32'b00000000000000001110010101110111;
assign LUT_1[40174] = 32'b00000000000000010000110010001100;
assign LUT_1[40175] = 32'b00000000000000001010000100001000;
assign LUT_1[40176] = 32'b00000000000000001111111000010001;
assign LUT_1[40177] = 32'b00000000000000001001001010001101;
assign LUT_1[40178] = 32'b00000000000000001011100110100010;
assign LUT_1[40179] = 32'b00000000000000000100111000011110;
assign LUT_1[40180] = 32'b00000000000000010111110001101000;
assign LUT_1[40181] = 32'b00000000000000010001000011100100;
assign LUT_1[40182] = 32'b00000000000000010011011111111001;
assign LUT_1[40183] = 32'b00000000000000001100110001110101;
assign LUT_1[40184] = 32'b00000000000000001111000110000110;
assign LUT_1[40185] = 32'b00000000000000001000011000000010;
assign LUT_1[40186] = 32'b00000000000000001010110100010111;
assign LUT_1[40187] = 32'b00000000000000000100000110010011;
assign LUT_1[40188] = 32'b00000000000000010110111111011101;
assign LUT_1[40189] = 32'b00000000000000010000010001011001;
assign LUT_1[40190] = 32'b00000000000000010010101101101110;
assign LUT_1[40191] = 32'b00000000000000001011111111101010;
assign LUT_1[40192] = 32'b00000000000000000101111000010001;
assign LUT_1[40193] = 32'b11111111111111111111001010001101;
assign LUT_1[40194] = 32'b00000000000000000001100110100010;
assign LUT_1[40195] = 32'b11111111111111111010111000011110;
assign LUT_1[40196] = 32'b00000000000000001101110001101000;
assign LUT_1[40197] = 32'b00000000000000000111000011100100;
assign LUT_1[40198] = 32'b00000000000000001001011111111001;
assign LUT_1[40199] = 32'b00000000000000000010110001110101;
assign LUT_1[40200] = 32'b00000000000000000101000110000110;
assign LUT_1[40201] = 32'b11111111111111111110011000000010;
assign LUT_1[40202] = 32'b00000000000000000000110100010111;
assign LUT_1[40203] = 32'b11111111111111111010000110010011;
assign LUT_1[40204] = 32'b00000000000000001100111111011101;
assign LUT_1[40205] = 32'b00000000000000000110010001011001;
assign LUT_1[40206] = 32'b00000000000000001000101101101110;
assign LUT_1[40207] = 32'b00000000000000000001111111101010;
assign LUT_1[40208] = 32'b00000000000000000111110011110011;
assign LUT_1[40209] = 32'b00000000000000000001000101101111;
assign LUT_1[40210] = 32'b00000000000000000011100010000100;
assign LUT_1[40211] = 32'b11111111111111111100110100000000;
assign LUT_1[40212] = 32'b00000000000000001111101101001010;
assign LUT_1[40213] = 32'b00000000000000001000111111000110;
assign LUT_1[40214] = 32'b00000000000000001011011011011011;
assign LUT_1[40215] = 32'b00000000000000000100101101010111;
assign LUT_1[40216] = 32'b00000000000000000111000001101000;
assign LUT_1[40217] = 32'b00000000000000000000010011100100;
assign LUT_1[40218] = 32'b00000000000000000010101111111001;
assign LUT_1[40219] = 32'b11111111111111111100000001110101;
assign LUT_1[40220] = 32'b00000000000000001110111010111111;
assign LUT_1[40221] = 32'b00000000000000001000001100111011;
assign LUT_1[40222] = 32'b00000000000000001010101001010000;
assign LUT_1[40223] = 32'b00000000000000000011111011001100;
assign LUT_1[40224] = 32'b00000000000000000110110011010000;
assign LUT_1[40225] = 32'b00000000000000000000000101001100;
assign LUT_1[40226] = 32'b00000000000000000010100001100001;
assign LUT_1[40227] = 32'b11111111111111111011110011011101;
assign LUT_1[40228] = 32'b00000000000000001110101100100111;
assign LUT_1[40229] = 32'b00000000000000000111111110100011;
assign LUT_1[40230] = 32'b00000000000000001010011010111000;
assign LUT_1[40231] = 32'b00000000000000000011101100110100;
assign LUT_1[40232] = 32'b00000000000000000110000001000101;
assign LUT_1[40233] = 32'b11111111111111111111010011000001;
assign LUT_1[40234] = 32'b00000000000000000001101111010110;
assign LUT_1[40235] = 32'b11111111111111111011000001010010;
assign LUT_1[40236] = 32'b00000000000000001101111010011100;
assign LUT_1[40237] = 32'b00000000000000000111001100011000;
assign LUT_1[40238] = 32'b00000000000000001001101000101101;
assign LUT_1[40239] = 32'b00000000000000000010111010101001;
assign LUT_1[40240] = 32'b00000000000000001000101110110010;
assign LUT_1[40241] = 32'b00000000000000000010000000101110;
assign LUT_1[40242] = 32'b00000000000000000100011101000011;
assign LUT_1[40243] = 32'b11111111111111111101101110111111;
assign LUT_1[40244] = 32'b00000000000000010000101000001001;
assign LUT_1[40245] = 32'b00000000000000001001111010000101;
assign LUT_1[40246] = 32'b00000000000000001100010110011010;
assign LUT_1[40247] = 32'b00000000000000000101101000010110;
assign LUT_1[40248] = 32'b00000000000000000111111100100111;
assign LUT_1[40249] = 32'b00000000000000000001001110100011;
assign LUT_1[40250] = 32'b00000000000000000011101010111000;
assign LUT_1[40251] = 32'b11111111111111111100111100110100;
assign LUT_1[40252] = 32'b00000000000000001111110101111110;
assign LUT_1[40253] = 32'b00000000000000001001000111111010;
assign LUT_1[40254] = 32'b00000000000000001011100100001111;
assign LUT_1[40255] = 32'b00000000000000000100110110001011;
assign LUT_1[40256] = 32'b00000000000000000111110101111001;
assign LUT_1[40257] = 32'b00000000000000000001000111110101;
assign LUT_1[40258] = 32'b00000000000000000011100100001010;
assign LUT_1[40259] = 32'b11111111111111111100110110000110;
assign LUT_1[40260] = 32'b00000000000000001111101111010000;
assign LUT_1[40261] = 32'b00000000000000001001000001001100;
assign LUT_1[40262] = 32'b00000000000000001011011101100001;
assign LUT_1[40263] = 32'b00000000000000000100101111011101;
assign LUT_1[40264] = 32'b00000000000000000111000011101110;
assign LUT_1[40265] = 32'b00000000000000000000010101101010;
assign LUT_1[40266] = 32'b00000000000000000010110001111111;
assign LUT_1[40267] = 32'b11111111111111111100000011111011;
assign LUT_1[40268] = 32'b00000000000000001110111101000101;
assign LUT_1[40269] = 32'b00000000000000001000001111000001;
assign LUT_1[40270] = 32'b00000000000000001010101011010110;
assign LUT_1[40271] = 32'b00000000000000000011111101010010;
assign LUT_1[40272] = 32'b00000000000000001001110001011011;
assign LUT_1[40273] = 32'b00000000000000000011000011010111;
assign LUT_1[40274] = 32'b00000000000000000101011111101100;
assign LUT_1[40275] = 32'b11111111111111111110110001101000;
assign LUT_1[40276] = 32'b00000000000000010001101010110010;
assign LUT_1[40277] = 32'b00000000000000001010111100101110;
assign LUT_1[40278] = 32'b00000000000000001101011001000011;
assign LUT_1[40279] = 32'b00000000000000000110101010111111;
assign LUT_1[40280] = 32'b00000000000000001000111111010000;
assign LUT_1[40281] = 32'b00000000000000000010010001001100;
assign LUT_1[40282] = 32'b00000000000000000100101101100001;
assign LUT_1[40283] = 32'b11111111111111111101111111011101;
assign LUT_1[40284] = 32'b00000000000000010000111000100111;
assign LUT_1[40285] = 32'b00000000000000001010001010100011;
assign LUT_1[40286] = 32'b00000000000000001100100110111000;
assign LUT_1[40287] = 32'b00000000000000000101111000110100;
assign LUT_1[40288] = 32'b00000000000000001000110000111000;
assign LUT_1[40289] = 32'b00000000000000000010000010110100;
assign LUT_1[40290] = 32'b00000000000000000100011111001001;
assign LUT_1[40291] = 32'b11111111111111111101110001000101;
assign LUT_1[40292] = 32'b00000000000000010000101010001111;
assign LUT_1[40293] = 32'b00000000000000001001111100001011;
assign LUT_1[40294] = 32'b00000000000000001100011000100000;
assign LUT_1[40295] = 32'b00000000000000000101101010011100;
assign LUT_1[40296] = 32'b00000000000000000111111110101101;
assign LUT_1[40297] = 32'b00000000000000000001010000101001;
assign LUT_1[40298] = 32'b00000000000000000011101100111110;
assign LUT_1[40299] = 32'b11111111111111111100111110111010;
assign LUT_1[40300] = 32'b00000000000000001111111000000100;
assign LUT_1[40301] = 32'b00000000000000001001001010000000;
assign LUT_1[40302] = 32'b00000000000000001011100110010101;
assign LUT_1[40303] = 32'b00000000000000000100111000010001;
assign LUT_1[40304] = 32'b00000000000000001010101100011010;
assign LUT_1[40305] = 32'b00000000000000000011111110010110;
assign LUT_1[40306] = 32'b00000000000000000110011010101011;
assign LUT_1[40307] = 32'b11111111111111111111101100100111;
assign LUT_1[40308] = 32'b00000000000000010010100101110001;
assign LUT_1[40309] = 32'b00000000000000001011110111101101;
assign LUT_1[40310] = 32'b00000000000000001110010100000010;
assign LUT_1[40311] = 32'b00000000000000000111100101111110;
assign LUT_1[40312] = 32'b00000000000000001001111010001111;
assign LUT_1[40313] = 32'b00000000000000000011001100001011;
assign LUT_1[40314] = 32'b00000000000000000101101000100000;
assign LUT_1[40315] = 32'b11111111111111111110111010011100;
assign LUT_1[40316] = 32'b00000000000000010001110011100110;
assign LUT_1[40317] = 32'b00000000000000001011000101100010;
assign LUT_1[40318] = 32'b00000000000000001101100001110111;
assign LUT_1[40319] = 32'b00000000000000000110110011110011;
assign LUT_1[40320] = 32'b00000000000000001000111000010100;
assign LUT_1[40321] = 32'b00000000000000000010001010010000;
assign LUT_1[40322] = 32'b00000000000000000100100110100101;
assign LUT_1[40323] = 32'b11111111111111111101111000100001;
assign LUT_1[40324] = 32'b00000000000000010000110001101011;
assign LUT_1[40325] = 32'b00000000000000001010000011100111;
assign LUT_1[40326] = 32'b00000000000000001100011111111100;
assign LUT_1[40327] = 32'b00000000000000000101110001111000;
assign LUT_1[40328] = 32'b00000000000000001000000110001001;
assign LUT_1[40329] = 32'b00000000000000000001011000000101;
assign LUT_1[40330] = 32'b00000000000000000011110100011010;
assign LUT_1[40331] = 32'b11111111111111111101000110010110;
assign LUT_1[40332] = 32'b00000000000000001111111111100000;
assign LUT_1[40333] = 32'b00000000000000001001010001011100;
assign LUT_1[40334] = 32'b00000000000000001011101101110001;
assign LUT_1[40335] = 32'b00000000000000000100111111101101;
assign LUT_1[40336] = 32'b00000000000000001010110011110110;
assign LUT_1[40337] = 32'b00000000000000000100000101110010;
assign LUT_1[40338] = 32'b00000000000000000110100010000111;
assign LUT_1[40339] = 32'b11111111111111111111110100000011;
assign LUT_1[40340] = 32'b00000000000000010010101101001101;
assign LUT_1[40341] = 32'b00000000000000001011111111001001;
assign LUT_1[40342] = 32'b00000000000000001110011011011110;
assign LUT_1[40343] = 32'b00000000000000000111101101011010;
assign LUT_1[40344] = 32'b00000000000000001010000001101011;
assign LUT_1[40345] = 32'b00000000000000000011010011100111;
assign LUT_1[40346] = 32'b00000000000000000101101111111100;
assign LUT_1[40347] = 32'b11111111111111111111000001111000;
assign LUT_1[40348] = 32'b00000000000000010001111011000010;
assign LUT_1[40349] = 32'b00000000000000001011001100111110;
assign LUT_1[40350] = 32'b00000000000000001101101001010011;
assign LUT_1[40351] = 32'b00000000000000000110111011001111;
assign LUT_1[40352] = 32'b00000000000000001001110011010011;
assign LUT_1[40353] = 32'b00000000000000000011000101001111;
assign LUT_1[40354] = 32'b00000000000000000101100001100100;
assign LUT_1[40355] = 32'b11111111111111111110110011100000;
assign LUT_1[40356] = 32'b00000000000000010001101100101010;
assign LUT_1[40357] = 32'b00000000000000001010111110100110;
assign LUT_1[40358] = 32'b00000000000000001101011010111011;
assign LUT_1[40359] = 32'b00000000000000000110101100110111;
assign LUT_1[40360] = 32'b00000000000000001001000001001000;
assign LUT_1[40361] = 32'b00000000000000000010010011000100;
assign LUT_1[40362] = 32'b00000000000000000100101111011001;
assign LUT_1[40363] = 32'b11111111111111111110000001010101;
assign LUT_1[40364] = 32'b00000000000000010000111010011111;
assign LUT_1[40365] = 32'b00000000000000001010001100011011;
assign LUT_1[40366] = 32'b00000000000000001100101000110000;
assign LUT_1[40367] = 32'b00000000000000000101111010101100;
assign LUT_1[40368] = 32'b00000000000000001011101110110101;
assign LUT_1[40369] = 32'b00000000000000000101000000110001;
assign LUT_1[40370] = 32'b00000000000000000111011101000110;
assign LUT_1[40371] = 32'b00000000000000000000101111000010;
assign LUT_1[40372] = 32'b00000000000000010011101000001100;
assign LUT_1[40373] = 32'b00000000000000001100111010001000;
assign LUT_1[40374] = 32'b00000000000000001111010110011101;
assign LUT_1[40375] = 32'b00000000000000001000101000011001;
assign LUT_1[40376] = 32'b00000000000000001010111100101010;
assign LUT_1[40377] = 32'b00000000000000000100001110100110;
assign LUT_1[40378] = 32'b00000000000000000110101010111011;
assign LUT_1[40379] = 32'b11111111111111111111111100110111;
assign LUT_1[40380] = 32'b00000000000000010010110110000001;
assign LUT_1[40381] = 32'b00000000000000001100000111111101;
assign LUT_1[40382] = 32'b00000000000000001110100100010010;
assign LUT_1[40383] = 32'b00000000000000000111110110001110;
assign LUT_1[40384] = 32'b00000000000000001010110101111100;
assign LUT_1[40385] = 32'b00000000000000000100000111111000;
assign LUT_1[40386] = 32'b00000000000000000110100100001101;
assign LUT_1[40387] = 32'b11111111111111111111110110001001;
assign LUT_1[40388] = 32'b00000000000000010010101111010011;
assign LUT_1[40389] = 32'b00000000000000001100000001001111;
assign LUT_1[40390] = 32'b00000000000000001110011101100100;
assign LUT_1[40391] = 32'b00000000000000000111101111100000;
assign LUT_1[40392] = 32'b00000000000000001010000011110001;
assign LUT_1[40393] = 32'b00000000000000000011010101101101;
assign LUT_1[40394] = 32'b00000000000000000101110010000010;
assign LUT_1[40395] = 32'b11111111111111111111000011111110;
assign LUT_1[40396] = 32'b00000000000000010001111101001000;
assign LUT_1[40397] = 32'b00000000000000001011001111000100;
assign LUT_1[40398] = 32'b00000000000000001101101011011001;
assign LUT_1[40399] = 32'b00000000000000000110111101010101;
assign LUT_1[40400] = 32'b00000000000000001100110001011110;
assign LUT_1[40401] = 32'b00000000000000000110000011011010;
assign LUT_1[40402] = 32'b00000000000000001000011111101111;
assign LUT_1[40403] = 32'b00000000000000000001110001101011;
assign LUT_1[40404] = 32'b00000000000000010100101010110101;
assign LUT_1[40405] = 32'b00000000000000001101111100110001;
assign LUT_1[40406] = 32'b00000000000000010000011001000110;
assign LUT_1[40407] = 32'b00000000000000001001101011000010;
assign LUT_1[40408] = 32'b00000000000000001011111111010011;
assign LUT_1[40409] = 32'b00000000000000000101010001001111;
assign LUT_1[40410] = 32'b00000000000000000111101101100100;
assign LUT_1[40411] = 32'b00000000000000000000111111100000;
assign LUT_1[40412] = 32'b00000000000000010011111000101010;
assign LUT_1[40413] = 32'b00000000000000001101001010100110;
assign LUT_1[40414] = 32'b00000000000000001111100110111011;
assign LUT_1[40415] = 32'b00000000000000001000111000110111;
assign LUT_1[40416] = 32'b00000000000000001011110000111011;
assign LUT_1[40417] = 32'b00000000000000000101000010110111;
assign LUT_1[40418] = 32'b00000000000000000111011111001100;
assign LUT_1[40419] = 32'b00000000000000000000110001001000;
assign LUT_1[40420] = 32'b00000000000000010011101010010010;
assign LUT_1[40421] = 32'b00000000000000001100111100001110;
assign LUT_1[40422] = 32'b00000000000000001111011000100011;
assign LUT_1[40423] = 32'b00000000000000001000101010011111;
assign LUT_1[40424] = 32'b00000000000000001010111110110000;
assign LUT_1[40425] = 32'b00000000000000000100010000101100;
assign LUT_1[40426] = 32'b00000000000000000110101101000001;
assign LUT_1[40427] = 32'b11111111111111111111111110111101;
assign LUT_1[40428] = 32'b00000000000000010010111000000111;
assign LUT_1[40429] = 32'b00000000000000001100001010000011;
assign LUT_1[40430] = 32'b00000000000000001110100110011000;
assign LUT_1[40431] = 32'b00000000000000000111111000010100;
assign LUT_1[40432] = 32'b00000000000000001101101100011101;
assign LUT_1[40433] = 32'b00000000000000000110111110011001;
assign LUT_1[40434] = 32'b00000000000000001001011010101110;
assign LUT_1[40435] = 32'b00000000000000000010101100101010;
assign LUT_1[40436] = 32'b00000000000000010101100101110100;
assign LUT_1[40437] = 32'b00000000000000001110110111110000;
assign LUT_1[40438] = 32'b00000000000000010001010100000101;
assign LUT_1[40439] = 32'b00000000000000001010100110000001;
assign LUT_1[40440] = 32'b00000000000000001100111010010010;
assign LUT_1[40441] = 32'b00000000000000000110001100001110;
assign LUT_1[40442] = 32'b00000000000000001000101000100011;
assign LUT_1[40443] = 32'b00000000000000000001111010011111;
assign LUT_1[40444] = 32'b00000000000000010100110011101001;
assign LUT_1[40445] = 32'b00000000000000001110000101100101;
assign LUT_1[40446] = 32'b00000000000000010000100001111010;
assign LUT_1[40447] = 32'b00000000000000001001110011110110;
assign LUT_1[40448] = 32'b00000000000000000001110010100010;
assign LUT_1[40449] = 32'b11111111111111111011000100011110;
assign LUT_1[40450] = 32'b11111111111111111101100000110011;
assign LUT_1[40451] = 32'b11111111111111110110110010101111;
assign LUT_1[40452] = 32'b00000000000000001001101011111001;
assign LUT_1[40453] = 32'b00000000000000000010111101110101;
assign LUT_1[40454] = 32'b00000000000000000101011010001010;
assign LUT_1[40455] = 32'b11111111111111111110101100000110;
assign LUT_1[40456] = 32'b00000000000000000001000000010111;
assign LUT_1[40457] = 32'b11111111111111111010010010010011;
assign LUT_1[40458] = 32'b11111111111111111100101110101000;
assign LUT_1[40459] = 32'b11111111111111110110000000100100;
assign LUT_1[40460] = 32'b00000000000000001000111001101110;
assign LUT_1[40461] = 32'b00000000000000000010001011101010;
assign LUT_1[40462] = 32'b00000000000000000100100111111111;
assign LUT_1[40463] = 32'b11111111111111111101111001111011;
assign LUT_1[40464] = 32'b00000000000000000011101110000100;
assign LUT_1[40465] = 32'b11111111111111111101000000000000;
assign LUT_1[40466] = 32'b11111111111111111111011100010101;
assign LUT_1[40467] = 32'b11111111111111111000101110010001;
assign LUT_1[40468] = 32'b00000000000000001011100111011011;
assign LUT_1[40469] = 32'b00000000000000000100111001010111;
assign LUT_1[40470] = 32'b00000000000000000111010101101100;
assign LUT_1[40471] = 32'b00000000000000000000100111101000;
assign LUT_1[40472] = 32'b00000000000000000010111011111001;
assign LUT_1[40473] = 32'b11111111111111111100001101110101;
assign LUT_1[40474] = 32'b11111111111111111110101010001010;
assign LUT_1[40475] = 32'b11111111111111110111111100000110;
assign LUT_1[40476] = 32'b00000000000000001010110101010000;
assign LUT_1[40477] = 32'b00000000000000000100000111001100;
assign LUT_1[40478] = 32'b00000000000000000110100011100001;
assign LUT_1[40479] = 32'b11111111111111111111110101011101;
assign LUT_1[40480] = 32'b00000000000000000010101101100001;
assign LUT_1[40481] = 32'b11111111111111111011111111011101;
assign LUT_1[40482] = 32'b11111111111111111110011011110010;
assign LUT_1[40483] = 32'b11111111111111110111101101101110;
assign LUT_1[40484] = 32'b00000000000000001010100110111000;
assign LUT_1[40485] = 32'b00000000000000000011111000110100;
assign LUT_1[40486] = 32'b00000000000000000110010101001001;
assign LUT_1[40487] = 32'b11111111111111111111100111000101;
assign LUT_1[40488] = 32'b00000000000000000001111011010110;
assign LUT_1[40489] = 32'b11111111111111111011001101010010;
assign LUT_1[40490] = 32'b11111111111111111101101001100111;
assign LUT_1[40491] = 32'b11111111111111110110111011100011;
assign LUT_1[40492] = 32'b00000000000000001001110100101101;
assign LUT_1[40493] = 32'b00000000000000000011000110101001;
assign LUT_1[40494] = 32'b00000000000000000101100010111110;
assign LUT_1[40495] = 32'b11111111111111111110110100111010;
assign LUT_1[40496] = 32'b00000000000000000100101001000011;
assign LUT_1[40497] = 32'b11111111111111111101111010111111;
assign LUT_1[40498] = 32'b00000000000000000000010111010100;
assign LUT_1[40499] = 32'b11111111111111111001101001010000;
assign LUT_1[40500] = 32'b00000000000000001100100010011010;
assign LUT_1[40501] = 32'b00000000000000000101110100010110;
assign LUT_1[40502] = 32'b00000000000000001000010000101011;
assign LUT_1[40503] = 32'b00000000000000000001100010100111;
assign LUT_1[40504] = 32'b00000000000000000011110110111000;
assign LUT_1[40505] = 32'b11111111111111111101001000110100;
assign LUT_1[40506] = 32'b11111111111111111111100101001001;
assign LUT_1[40507] = 32'b11111111111111111000110111000101;
assign LUT_1[40508] = 32'b00000000000000001011110000001111;
assign LUT_1[40509] = 32'b00000000000000000101000010001011;
assign LUT_1[40510] = 32'b00000000000000000111011110100000;
assign LUT_1[40511] = 32'b00000000000000000000110000011100;
assign LUT_1[40512] = 32'b00000000000000000011110000001010;
assign LUT_1[40513] = 32'b11111111111111111101000010000110;
assign LUT_1[40514] = 32'b11111111111111111111011110011011;
assign LUT_1[40515] = 32'b11111111111111111000110000010111;
assign LUT_1[40516] = 32'b00000000000000001011101001100001;
assign LUT_1[40517] = 32'b00000000000000000100111011011101;
assign LUT_1[40518] = 32'b00000000000000000111010111110010;
assign LUT_1[40519] = 32'b00000000000000000000101001101110;
assign LUT_1[40520] = 32'b00000000000000000010111101111111;
assign LUT_1[40521] = 32'b11111111111111111100001111111011;
assign LUT_1[40522] = 32'b11111111111111111110101100010000;
assign LUT_1[40523] = 32'b11111111111111110111111110001100;
assign LUT_1[40524] = 32'b00000000000000001010110111010110;
assign LUT_1[40525] = 32'b00000000000000000100001001010010;
assign LUT_1[40526] = 32'b00000000000000000110100101100111;
assign LUT_1[40527] = 32'b11111111111111111111110111100011;
assign LUT_1[40528] = 32'b00000000000000000101101011101100;
assign LUT_1[40529] = 32'b11111111111111111110111101101000;
assign LUT_1[40530] = 32'b00000000000000000001011001111101;
assign LUT_1[40531] = 32'b11111111111111111010101011111001;
assign LUT_1[40532] = 32'b00000000000000001101100101000011;
assign LUT_1[40533] = 32'b00000000000000000110110110111111;
assign LUT_1[40534] = 32'b00000000000000001001010011010100;
assign LUT_1[40535] = 32'b00000000000000000010100101010000;
assign LUT_1[40536] = 32'b00000000000000000100111001100001;
assign LUT_1[40537] = 32'b11111111111111111110001011011101;
assign LUT_1[40538] = 32'b00000000000000000000100111110010;
assign LUT_1[40539] = 32'b11111111111111111001111001101110;
assign LUT_1[40540] = 32'b00000000000000001100110010111000;
assign LUT_1[40541] = 32'b00000000000000000110000100110100;
assign LUT_1[40542] = 32'b00000000000000001000100001001001;
assign LUT_1[40543] = 32'b00000000000000000001110011000101;
assign LUT_1[40544] = 32'b00000000000000000100101011001001;
assign LUT_1[40545] = 32'b11111111111111111101111101000101;
assign LUT_1[40546] = 32'b00000000000000000000011001011010;
assign LUT_1[40547] = 32'b11111111111111111001101011010110;
assign LUT_1[40548] = 32'b00000000000000001100100100100000;
assign LUT_1[40549] = 32'b00000000000000000101110110011100;
assign LUT_1[40550] = 32'b00000000000000001000010010110001;
assign LUT_1[40551] = 32'b00000000000000000001100100101101;
assign LUT_1[40552] = 32'b00000000000000000011111000111110;
assign LUT_1[40553] = 32'b11111111111111111101001010111010;
assign LUT_1[40554] = 32'b11111111111111111111100111001111;
assign LUT_1[40555] = 32'b11111111111111111000111001001011;
assign LUT_1[40556] = 32'b00000000000000001011110010010101;
assign LUT_1[40557] = 32'b00000000000000000101000100010001;
assign LUT_1[40558] = 32'b00000000000000000111100000100110;
assign LUT_1[40559] = 32'b00000000000000000000110010100010;
assign LUT_1[40560] = 32'b00000000000000000110100110101011;
assign LUT_1[40561] = 32'b11111111111111111111111000100111;
assign LUT_1[40562] = 32'b00000000000000000010010100111100;
assign LUT_1[40563] = 32'b11111111111111111011100110111000;
assign LUT_1[40564] = 32'b00000000000000001110100000000010;
assign LUT_1[40565] = 32'b00000000000000000111110001111110;
assign LUT_1[40566] = 32'b00000000000000001010001110010011;
assign LUT_1[40567] = 32'b00000000000000000011100000001111;
assign LUT_1[40568] = 32'b00000000000000000101110100100000;
assign LUT_1[40569] = 32'b11111111111111111111000110011100;
assign LUT_1[40570] = 32'b00000000000000000001100010110001;
assign LUT_1[40571] = 32'b11111111111111111010110100101101;
assign LUT_1[40572] = 32'b00000000000000001101101101110111;
assign LUT_1[40573] = 32'b00000000000000000110111111110011;
assign LUT_1[40574] = 32'b00000000000000001001011100001000;
assign LUT_1[40575] = 32'b00000000000000000010101110000100;
assign LUT_1[40576] = 32'b00000000000000000100110010100101;
assign LUT_1[40577] = 32'b11111111111111111110000100100001;
assign LUT_1[40578] = 32'b00000000000000000000100000110110;
assign LUT_1[40579] = 32'b11111111111111111001110010110010;
assign LUT_1[40580] = 32'b00000000000000001100101011111100;
assign LUT_1[40581] = 32'b00000000000000000101111101111000;
assign LUT_1[40582] = 32'b00000000000000001000011010001101;
assign LUT_1[40583] = 32'b00000000000000000001101100001001;
assign LUT_1[40584] = 32'b00000000000000000100000000011010;
assign LUT_1[40585] = 32'b11111111111111111101010010010110;
assign LUT_1[40586] = 32'b11111111111111111111101110101011;
assign LUT_1[40587] = 32'b11111111111111111001000000100111;
assign LUT_1[40588] = 32'b00000000000000001011111001110001;
assign LUT_1[40589] = 32'b00000000000000000101001011101101;
assign LUT_1[40590] = 32'b00000000000000000111101000000010;
assign LUT_1[40591] = 32'b00000000000000000000111001111110;
assign LUT_1[40592] = 32'b00000000000000000110101110000111;
assign LUT_1[40593] = 32'b00000000000000000000000000000011;
assign LUT_1[40594] = 32'b00000000000000000010011100011000;
assign LUT_1[40595] = 32'b11111111111111111011101110010100;
assign LUT_1[40596] = 32'b00000000000000001110100111011110;
assign LUT_1[40597] = 32'b00000000000000000111111001011010;
assign LUT_1[40598] = 32'b00000000000000001010010101101111;
assign LUT_1[40599] = 32'b00000000000000000011100111101011;
assign LUT_1[40600] = 32'b00000000000000000101111011111100;
assign LUT_1[40601] = 32'b11111111111111111111001101111000;
assign LUT_1[40602] = 32'b00000000000000000001101010001101;
assign LUT_1[40603] = 32'b11111111111111111010111100001001;
assign LUT_1[40604] = 32'b00000000000000001101110101010011;
assign LUT_1[40605] = 32'b00000000000000000111000111001111;
assign LUT_1[40606] = 32'b00000000000000001001100011100100;
assign LUT_1[40607] = 32'b00000000000000000010110101100000;
assign LUT_1[40608] = 32'b00000000000000000101101101100100;
assign LUT_1[40609] = 32'b11111111111111111110111111100000;
assign LUT_1[40610] = 32'b00000000000000000001011011110101;
assign LUT_1[40611] = 32'b11111111111111111010101101110001;
assign LUT_1[40612] = 32'b00000000000000001101100110111011;
assign LUT_1[40613] = 32'b00000000000000000110111000110111;
assign LUT_1[40614] = 32'b00000000000000001001010101001100;
assign LUT_1[40615] = 32'b00000000000000000010100111001000;
assign LUT_1[40616] = 32'b00000000000000000100111011011001;
assign LUT_1[40617] = 32'b11111111111111111110001101010101;
assign LUT_1[40618] = 32'b00000000000000000000101001101010;
assign LUT_1[40619] = 32'b11111111111111111001111011100110;
assign LUT_1[40620] = 32'b00000000000000001100110100110000;
assign LUT_1[40621] = 32'b00000000000000000110000110101100;
assign LUT_1[40622] = 32'b00000000000000001000100011000001;
assign LUT_1[40623] = 32'b00000000000000000001110100111101;
assign LUT_1[40624] = 32'b00000000000000000111101001000110;
assign LUT_1[40625] = 32'b00000000000000000000111011000010;
assign LUT_1[40626] = 32'b00000000000000000011010111010111;
assign LUT_1[40627] = 32'b11111111111111111100101001010011;
assign LUT_1[40628] = 32'b00000000000000001111100010011101;
assign LUT_1[40629] = 32'b00000000000000001000110100011001;
assign LUT_1[40630] = 32'b00000000000000001011010000101110;
assign LUT_1[40631] = 32'b00000000000000000100100010101010;
assign LUT_1[40632] = 32'b00000000000000000110110110111011;
assign LUT_1[40633] = 32'b00000000000000000000001000110111;
assign LUT_1[40634] = 32'b00000000000000000010100101001100;
assign LUT_1[40635] = 32'b11111111111111111011110111001000;
assign LUT_1[40636] = 32'b00000000000000001110110000010010;
assign LUT_1[40637] = 32'b00000000000000001000000010001110;
assign LUT_1[40638] = 32'b00000000000000001010011110100011;
assign LUT_1[40639] = 32'b00000000000000000011110000011111;
assign LUT_1[40640] = 32'b00000000000000000110110000001101;
assign LUT_1[40641] = 32'b00000000000000000000000010001001;
assign LUT_1[40642] = 32'b00000000000000000010011110011110;
assign LUT_1[40643] = 32'b11111111111111111011110000011010;
assign LUT_1[40644] = 32'b00000000000000001110101001100100;
assign LUT_1[40645] = 32'b00000000000000000111111011100000;
assign LUT_1[40646] = 32'b00000000000000001010010111110101;
assign LUT_1[40647] = 32'b00000000000000000011101001110001;
assign LUT_1[40648] = 32'b00000000000000000101111110000010;
assign LUT_1[40649] = 32'b11111111111111111111001111111110;
assign LUT_1[40650] = 32'b00000000000000000001101100010011;
assign LUT_1[40651] = 32'b11111111111111111010111110001111;
assign LUT_1[40652] = 32'b00000000000000001101110111011001;
assign LUT_1[40653] = 32'b00000000000000000111001001010101;
assign LUT_1[40654] = 32'b00000000000000001001100101101010;
assign LUT_1[40655] = 32'b00000000000000000010110111100110;
assign LUT_1[40656] = 32'b00000000000000001000101011101111;
assign LUT_1[40657] = 32'b00000000000000000001111101101011;
assign LUT_1[40658] = 32'b00000000000000000100011010000000;
assign LUT_1[40659] = 32'b11111111111111111101101011111100;
assign LUT_1[40660] = 32'b00000000000000010000100101000110;
assign LUT_1[40661] = 32'b00000000000000001001110111000010;
assign LUT_1[40662] = 32'b00000000000000001100010011010111;
assign LUT_1[40663] = 32'b00000000000000000101100101010011;
assign LUT_1[40664] = 32'b00000000000000000111111001100100;
assign LUT_1[40665] = 32'b00000000000000000001001011100000;
assign LUT_1[40666] = 32'b00000000000000000011100111110101;
assign LUT_1[40667] = 32'b11111111111111111100111001110001;
assign LUT_1[40668] = 32'b00000000000000001111110010111011;
assign LUT_1[40669] = 32'b00000000000000001001000100110111;
assign LUT_1[40670] = 32'b00000000000000001011100001001100;
assign LUT_1[40671] = 32'b00000000000000000100110011001000;
assign LUT_1[40672] = 32'b00000000000000000111101011001100;
assign LUT_1[40673] = 32'b00000000000000000000111101001000;
assign LUT_1[40674] = 32'b00000000000000000011011001011101;
assign LUT_1[40675] = 32'b11111111111111111100101011011001;
assign LUT_1[40676] = 32'b00000000000000001111100100100011;
assign LUT_1[40677] = 32'b00000000000000001000110110011111;
assign LUT_1[40678] = 32'b00000000000000001011010010110100;
assign LUT_1[40679] = 32'b00000000000000000100100100110000;
assign LUT_1[40680] = 32'b00000000000000000110111001000001;
assign LUT_1[40681] = 32'b00000000000000000000001010111101;
assign LUT_1[40682] = 32'b00000000000000000010100111010010;
assign LUT_1[40683] = 32'b11111111111111111011111001001110;
assign LUT_1[40684] = 32'b00000000000000001110110010011000;
assign LUT_1[40685] = 32'b00000000000000001000000100010100;
assign LUT_1[40686] = 32'b00000000000000001010100000101001;
assign LUT_1[40687] = 32'b00000000000000000011110010100101;
assign LUT_1[40688] = 32'b00000000000000001001100110101110;
assign LUT_1[40689] = 32'b00000000000000000010111000101010;
assign LUT_1[40690] = 32'b00000000000000000101010100111111;
assign LUT_1[40691] = 32'b11111111111111111110100110111011;
assign LUT_1[40692] = 32'b00000000000000010001100000000101;
assign LUT_1[40693] = 32'b00000000000000001010110010000001;
assign LUT_1[40694] = 32'b00000000000000001101001110010110;
assign LUT_1[40695] = 32'b00000000000000000110100000010010;
assign LUT_1[40696] = 32'b00000000000000001000110100100011;
assign LUT_1[40697] = 32'b00000000000000000010000110011111;
assign LUT_1[40698] = 32'b00000000000000000100100010110100;
assign LUT_1[40699] = 32'b11111111111111111101110100110000;
assign LUT_1[40700] = 32'b00000000000000010000101101111010;
assign LUT_1[40701] = 32'b00000000000000001001111111110110;
assign LUT_1[40702] = 32'b00000000000000001100011100001011;
assign LUT_1[40703] = 32'b00000000000000000101101110000111;
assign LUT_1[40704] = 32'b11111111111111111111100110101110;
assign LUT_1[40705] = 32'b11111111111111111000111000101010;
assign LUT_1[40706] = 32'b11111111111111111011010100111111;
assign LUT_1[40707] = 32'b11111111111111110100100110111011;
assign LUT_1[40708] = 32'b00000000000000000111100000000101;
assign LUT_1[40709] = 32'b00000000000000000000110010000001;
assign LUT_1[40710] = 32'b00000000000000000011001110010110;
assign LUT_1[40711] = 32'b11111111111111111100100000010010;
assign LUT_1[40712] = 32'b11111111111111111110110100100011;
assign LUT_1[40713] = 32'b11111111111111111000000110011111;
assign LUT_1[40714] = 32'b11111111111111111010100010110100;
assign LUT_1[40715] = 32'b11111111111111110011110100110000;
assign LUT_1[40716] = 32'b00000000000000000110101101111010;
assign LUT_1[40717] = 32'b11111111111111111111111111110110;
assign LUT_1[40718] = 32'b00000000000000000010011100001011;
assign LUT_1[40719] = 32'b11111111111111111011101110000111;
assign LUT_1[40720] = 32'b00000000000000000001100010010000;
assign LUT_1[40721] = 32'b11111111111111111010110100001100;
assign LUT_1[40722] = 32'b11111111111111111101010000100001;
assign LUT_1[40723] = 32'b11111111111111110110100010011101;
assign LUT_1[40724] = 32'b00000000000000001001011011100111;
assign LUT_1[40725] = 32'b00000000000000000010101101100011;
assign LUT_1[40726] = 32'b00000000000000000101001001111000;
assign LUT_1[40727] = 32'b11111111111111111110011011110100;
assign LUT_1[40728] = 32'b00000000000000000000110000000101;
assign LUT_1[40729] = 32'b11111111111111111010000010000001;
assign LUT_1[40730] = 32'b11111111111111111100011110010110;
assign LUT_1[40731] = 32'b11111111111111110101110000010010;
assign LUT_1[40732] = 32'b00000000000000001000101001011100;
assign LUT_1[40733] = 32'b00000000000000000001111011011000;
assign LUT_1[40734] = 32'b00000000000000000100010111101101;
assign LUT_1[40735] = 32'b11111111111111111101101001101001;
assign LUT_1[40736] = 32'b00000000000000000000100001101101;
assign LUT_1[40737] = 32'b11111111111111111001110011101001;
assign LUT_1[40738] = 32'b11111111111111111100001111111110;
assign LUT_1[40739] = 32'b11111111111111110101100001111010;
assign LUT_1[40740] = 32'b00000000000000001000011011000100;
assign LUT_1[40741] = 32'b00000000000000000001101101000000;
assign LUT_1[40742] = 32'b00000000000000000100001001010101;
assign LUT_1[40743] = 32'b11111111111111111101011011010001;
assign LUT_1[40744] = 32'b11111111111111111111101111100010;
assign LUT_1[40745] = 32'b11111111111111111001000001011110;
assign LUT_1[40746] = 32'b11111111111111111011011101110011;
assign LUT_1[40747] = 32'b11111111111111110100101111101111;
assign LUT_1[40748] = 32'b00000000000000000111101000111001;
assign LUT_1[40749] = 32'b00000000000000000000111010110101;
assign LUT_1[40750] = 32'b00000000000000000011010111001010;
assign LUT_1[40751] = 32'b11111111111111111100101001000110;
assign LUT_1[40752] = 32'b00000000000000000010011101001111;
assign LUT_1[40753] = 32'b11111111111111111011101111001011;
assign LUT_1[40754] = 32'b11111111111111111110001011100000;
assign LUT_1[40755] = 32'b11111111111111110111011101011100;
assign LUT_1[40756] = 32'b00000000000000001010010110100110;
assign LUT_1[40757] = 32'b00000000000000000011101000100010;
assign LUT_1[40758] = 32'b00000000000000000110000100110111;
assign LUT_1[40759] = 32'b11111111111111111111010110110011;
assign LUT_1[40760] = 32'b00000000000000000001101011000100;
assign LUT_1[40761] = 32'b11111111111111111010111101000000;
assign LUT_1[40762] = 32'b11111111111111111101011001010101;
assign LUT_1[40763] = 32'b11111111111111110110101011010001;
assign LUT_1[40764] = 32'b00000000000000001001100100011011;
assign LUT_1[40765] = 32'b00000000000000000010110110010111;
assign LUT_1[40766] = 32'b00000000000000000101010010101100;
assign LUT_1[40767] = 32'b11111111111111111110100100101000;
assign LUT_1[40768] = 32'b00000000000000000001100100010110;
assign LUT_1[40769] = 32'b11111111111111111010110110010010;
assign LUT_1[40770] = 32'b11111111111111111101010010100111;
assign LUT_1[40771] = 32'b11111111111111110110100100100011;
assign LUT_1[40772] = 32'b00000000000000001001011101101101;
assign LUT_1[40773] = 32'b00000000000000000010101111101001;
assign LUT_1[40774] = 32'b00000000000000000101001011111110;
assign LUT_1[40775] = 32'b11111111111111111110011101111010;
assign LUT_1[40776] = 32'b00000000000000000000110010001011;
assign LUT_1[40777] = 32'b11111111111111111010000100000111;
assign LUT_1[40778] = 32'b11111111111111111100100000011100;
assign LUT_1[40779] = 32'b11111111111111110101110010011000;
assign LUT_1[40780] = 32'b00000000000000001000101011100010;
assign LUT_1[40781] = 32'b00000000000000000001111101011110;
assign LUT_1[40782] = 32'b00000000000000000100011001110011;
assign LUT_1[40783] = 32'b11111111111111111101101011101111;
assign LUT_1[40784] = 32'b00000000000000000011011111111000;
assign LUT_1[40785] = 32'b11111111111111111100110001110100;
assign LUT_1[40786] = 32'b11111111111111111111001110001001;
assign LUT_1[40787] = 32'b11111111111111111000100000000101;
assign LUT_1[40788] = 32'b00000000000000001011011001001111;
assign LUT_1[40789] = 32'b00000000000000000100101011001011;
assign LUT_1[40790] = 32'b00000000000000000111000111100000;
assign LUT_1[40791] = 32'b00000000000000000000011001011100;
assign LUT_1[40792] = 32'b00000000000000000010101101101101;
assign LUT_1[40793] = 32'b11111111111111111011111111101001;
assign LUT_1[40794] = 32'b11111111111111111110011011111110;
assign LUT_1[40795] = 32'b11111111111111110111101101111010;
assign LUT_1[40796] = 32'b00000000000000001010100111000100;
assign LUT_1[40797] = 32'b00000000000000000011111001000000;
assign LUT_1[40798] = 32'b00000000000000000110010101010101;
assign LUT_1[40799] = 32'b11111111111111111111100111010001;
assign LUT_1[40800] = 32'b00000000000000000010011111010101;
assign LUT_1[40801] = 32'b11111111111111111011110001010001;
assign LUT_1[40802] = 32'b11111111111111111110001101100110;
assign LUT_1[40803] = 32'b11111111111111110111011111100010;
assign LUT_1[40804] = 32'b00000000000000001010011000101100;
assign LUT_1[40805] = 32'b00000000000000000011101010101000;
assign LUT_1[40806] = 32'b00000000000000000110000110111101;
assign LUT_1[40807] = 32'b11111111111111111111011000111001;
assign LUT_1[40808] = 32'b00000000000000000001101101001010;
assign LUT_1[40809] = 32'b11111111111111111010111111000110;
assign LUT_1[40810] = 32'b11111111111111111101011011011011;
assign LUT_1[40811] = 32'b11111111111111110110101101010111;
assign LUT_1[40812] = 32'b00000000000000001001100110100001;
assign LUT_1[40813] = 32'b00000000000000000010111000011101;
assign LUT_1[40814] = 32'b00000000000000000101010100110010;
assign LUT_1[40815] = 32'b11111111111111111110100110101110;
assign LUT_1[40816] = 32'b00000000000000000100011010110111;
assign LUT_1[40817] = 32'b11111111111111111101101100110011;
assign LUT_1[40818] = 32'b00000000000000000000001001001000;
assign LUT_1[40819] = 32'b11111111111111111001011011000100;
assign LUT_1[40820] = 32'b00000000000000001100010100001110;
assign LUT_1[40821] = 32'b00000000000000000101100110001010;
assign LUT_1[40822] = 32'b00000000000000001000000010011111;
assign LUT_1[40823] = 32'b00000000000000000001010100011011;
assign LUT_1[40824] = 32'b00000000000000000011101000101100;
assign LUT_1[40825] = 32'b11111111111111111100111010101000;
assign LUT_1[40826] = 32'b11111111111111111111010110111101;
assign LUT_1[40827] = 32'b11111111111111111000101000111001;
assign LUT_1[40828] = 32'b00000000000000001011100010000011;
assign LUT_1[40829] = 32'b00000000000000000100110011111111;
assign LUT_1[40830] = 32'b00000000000000000111010000010100;
assign LUT_1[40831] = 32'b00000000000000000000100010010000;
assign LUT_1[40832] = 32'b00000000000000000010100110110001;
assign LUT_1[40833] = 32'b11111111111111111011111000101101;
assign LUT_1[40834] = 32'b11111111111111111110010101000010;
assign LUT_1[40835] = 32'b11111111111111110111100110111110;
assign LUT_1[40836] = 32'b00000000000000001010100000001000;
assign LUT_1[40837] = 32'b00000000000000000011110010000100;
assign LUT_1[40838] = 32'b00000000000000000110001110011001;
assign LUT_1[40839] = 32'b11111111111111111111100000010101;
assign LUT_1[40840] = 32'b00000000000000000001110100100110;
assign LUT_1[40841] = 32'b11111111111111111011000110100010;
assign LUT_1[40842] = 32'b11111111111111111101100010110111;
assign LUT_1[40843] = 32'b11111111111111110110110100110011;
assign LUT_1[40844] = 32'b00000000000000001001101101111101;
assign LUT_1[40845] = 32'b00000000000000000010111111111001;
assign LUT_1[40846] = 32'b00000000000000000101011100001110;
assign LUT_1[40847] = 32'b11111111111111111110101110001010;
assign LUT_1[40848] = 32'b00000000000000000100100010010011;
assign LUT_1[40849] = 32'b11111111111111111101110100001111;
assign LUT_1[40850] = 32'b00000000000000000000010000100100;
assign LUT_1[40851] = 32'b11111111111111111001100010100000;
assign LUT_1[40852] = 32'b00000000000000001100011011101010;
assign LUT_1[40853] = 32'b00000000000000000101101101100110;
assign LUT_1[40854] = 32'b00000000000000001000001001111011;
assign LUT_1[40855] = 32'b00000000000000000001011011110111;
assign LUT_1[40856] = 32'b00000000000000000011110000001000;
assign LUT_1[40857] = 32'b11111111111111111101000010000100;
assign LUT_1[40858] = 32'b11111111111111111111011110011001;
assign LUT_1[40859] = 32'b11111111111111111000110000010101;
assign LUT_1[40860] = 32'b00000000000000001011101001011111;
assign LUT_1[40861] = 32'b00000000000000000100111011011011;
assign LUT_1[40862] = 32'b00000000000000000111010111110000;
assign LUT_1[40863] = 32'b00000000000000000000101001101100;
assign LUT_1[40864] = 32'b00000000000000000011100001110000;
assign LUT_1[40865] = 32'b11111111111111111100110011101100;
assign LUT_1[40866] = 32'b11111111111111111111010000000001;
assign LUT_1[40867] = 32'b11111111111111111000100001111101;
assign LUT_1[40868] = 32'b00000000000000001011011011000111;
assign LUT_1[40869] = 32'b00000000000000000100101101000011;
assign LUT_1[40870] = 32'b00000000000000000111001001011000;
assign LUT_1[40871] = 32'b00000000000000000000011011010100;
assign LUT_1[40872] = 32'b00000000000000000010101111100101;
assign LUT_1[40873] = 32'b11111111111111111100000001100001;
assign LUT_1[40874] = 32'b11111111111111111110011101110110;
assign LUT_1[40875] = 32'b11111111111111110111101111110010;
assign LUT_1[40876] = 32'b00000000000000001010101000111100;
assign LUT_1[40877] = 32'b00000000000000000011111010111000;
assign LUT_1[40878] = 32'b00000000000000000110010111001101;
assign LUT_1[40879] = 32'b11111111111111111111101001001001;
assign LUT_1[40880] = 32'b00000000000000000101011101010010;
assign LUT_1[40881] = 32'b11111111111111111110101111001110;
assign LUT_1[40882] = 32'b00000000000000000001001011100011;
assign LUT_1[40883] = 32'b11111111111111111010011101011111;
assign LUT_1[40884] = 32'b00000000000000001101010110101001;
assign LUT_1[40885] = 32'b00000000000000000110101000100101;
assign LUT_1[40886] = 32'b00000000000000001001000100111010;
assign LUT_1[40887] = 32'b00000000000000000010010110110110;
assign LUT_1[40888] = 32'b00000000000000000100101011000111;
assign LUT_1[40889] = 32'b11111111111111111101111101000011;
assign LUT_1[40890] = 32'b00000000000000000000011001011000;
assign LUT_1[40891] = 32'b11111111111111111001101011010100;
assign LUT_1[40892] = 32'b00000000000000001100100100011110;
assign LUT_1[40893] = 32'b00000000000000000101110110011010;
assign LUT_1[40894] = 32'b00000000000000001000010010101111;
assign LUT_1[40895] = 32'b00000000000000000001100100101011;
assign LUT_1[40896] = 32'b00000000000000000100100100011001;
assign LUT_1[40897] = 32'b11111111111111111101110110010101;
assign LUT_1[40898] = 32'b00000000000000000000010010101010;
assign LUT_1[40899] = 32'b11111111111111111001100100100110;
assign LUT_1[40900] = 32'b00000000000000001100011101110000;
assign LUT_1[40901] = 32'b00000000000000000101101111101100;
assign LUT_1[40902] = 32'b00000000000000001000001100000001;
assign LUT_1[40903] = 32'b00000000000000000001011101111101;
assign LUT_1[40904] = 32'b00000000000000000011110010001110;
assign LUT_1[40905] = 32'b11111111111111111101000100001010;
assign LUT_1[40906] = 32'b11111111111111111111100000011111;
assign LUT_1[40907] = 32'b11111111111111111000110010011011;
assign LUT_1[40908] = 32'b00000000000000001011101011100101;
assign LUT_1[40909] = 32'b00000000000000000100111101100001;
assign LUT_1[40910] = 32'b00000000000000000111011001110110;
assign LUT_1[40911] = 32'b00000000000000000000101011110010;
assign LUT_1[40912] = 32'b00000000000000000110011111111011;
assign LUT_1[40913] = 32'b11111111111111111111110001110111;
assign LUT_1[40914] = 32'b00000000000000000010001110001100;
assign LUT_1[40915] = 32'b11111111111111111011100000001000;
assign LUT_1[40916] = 32'b00000000000000001110011001010010;
assign LUT_1[40917] = 32'b00000000000000000111101011001110;
assign LUT_1[40918] = 32'b00000000000000001010000111100011;
assign LUT_1[40919] = 32'b00000000000000000011011001011111;
assign LUT_1[40920] = 32'b00000000000000000101101101110000;
assign LUT_1[40921] = 32'b11111111111111111110111111101100;
assign LUT_1[40922] = 32'b00000000000000000001011100000001;
assign LUT_1[40923] = 32'b11111111111111111010101101111101;
assign LUT_1[40924] = 32'b00000000000000001101100111000111;
assign LUT_1[40925] = 32'b00000000000000000110111001000011;
assign LUT_1[40926] = 32'b00000000000000001001010101011000;
assign LUT_1[40927] = 32'b00000000000000000010100111010100;
assign LUT_1[40928] = 32'b00000000000000000101011111011000;
assign LUT_1[40929] = 32'b11111111111111111110110001010100;
assign LUT_1[40930] = 32'b00000000000000000001001101101001;
assign LUT_1[40931] = 32'b11111111111111111010011111100101;
assign LUT_1[40932] = 32'b00000000000000001101011000101111;
assign LUT_1[40933] = 32'b00000000000000000110101010101011;
assign LUT_1[40934] = 32'b00000000000000001001000111000000;
assign LUT_1[40935] = 32'b00000000000000000010011000111100;
assign LUT_1[40936] = 32'b00000000000000000100101101001101;
assign LUT_1[40937] = 32'b11111111111111111101111111001001;
assign LUT_1[40938] = 32'b00000000000000000000011011011110;
assign LUT_1[40939] = 32'b11111111111111111001101101011010;
assign LUT_1[40940] = 32'b00000000000000001100100110100100;
assign LUT_1[40941] = 32'b00000000000000000101111000100000;
assign LUT_1[40942] = 32'b00000000000000001000010100110101;
assign LUT_1[40943] = 32'b00000000000000000001100110110001;
assign LUT_1[40944] = 32'b00000000000000000111011010111010;
assign LUT_1[40945] = 32'b00000000000000000000101100110110;
assign LUT_1[40946] = 32'b00000000000000000011001001001011;
assign LUT_1[40947] = 32'b11111111111111111100011011000111;
assign LUT_1[40948] = 32'b00000000000000001111010100010001;
assign LUT_1[40949] = 32'b00000000000000001000100110001101;
assign LUT_1[40950] = 32'b00000000000000001011000010100010;
assign LUT_1[40951] = 32'b00000000000000000100010100011110;
assign LUT_1[40952] = 32'b00000000000000000110101000101111;
assign LUT_1[40953] = 32'b11111111111111111111111010101011;
assign LUT_1[40954] = 32'b00000000000000000010010111000000;
assign LUT_1[40955] = 32'b11111111111111111011101000111100;
assign LUT_1[40956] = 32'b00000000000000001110100010000110;
assign LUT_1[40957] = 32'b00000000000000000111110100000010;
assign LUT_1[40958] = 32'b00000000000000001010010000010111;
assign LUT_1[40959] = 32'b00000000000000000011100010010011;
assign LUT_1[40960] = 32'b00000000000000000011111110110111;
assign LUT_1[40961] = 32'b11111111111111111101010000110011;
assign LUT_1[40962] = 32'b11111111111111111111101101001000;
assign LUT_1[40963] = 32'b11111111111111111000111111000100;
assign LUT_1[40964] = 32'b00000000000000001011111000001110;
assign LUT_1[40965] = 32'b00000000000000000101001010001010;
assign LUT_1[40966] = 32'b00000000000000000111100110011111;
assign LUT_1[40967] = 32'b00000000000000000000111000011011;
assign LUT_1[40968] = 32'b00000000000000000011001100101100;
assign LUT_1[40969] = 32'b11111111111111111100011110101000;
assign LUT_1[40970] = 32'b11111111111111111110111010111101;
assign LUT_1[40971] = 32'b11111111111111111000001100111001;
assign LUT_1[40972] = 32'b00000000000000001011000110000011;
assign LUT_1[40973] = 32'b00000000000000000100010111111111;
assign LUT_1[40974] = 32'b00000000000000000110110100010100;
assign LUT_1[40975] = 32'b00000000000000000000000110010000;
assign LUT_1[40976] = 32'b00000000000000000101111010011001;
assign LUT_1[40977] = 32'b11111111111111111111001100010101;
assign LUT_1[40978] = 32'b00000000000000000001101000101010;
assign LUT_1[40979] = 32'b11111111111111111010111010100110;
assign LUT_1[40980] = 32'b00000000000000001101110011110000;
assign LUT_1[40981] = 32'b00000000000000000111000101101100;
assign LUT_1[40982] = 32'b00000000000000001001100010000001;
assign LUT_1[40983] = 32'b00000000000000000010110011111101;
assign LUT_1[40984] = 32'b00000000000000000101001000001110;
assign LUT_1[40985] = 32'b11111111111111111110011010001010;
assign LUT_1[40986] = 32'b00000000000000000000110110011111;
assign LUT_1[40987] = 32'b11111111111111111010001000011011;
assign LUT_1[40988] = 32'b00000000000000001101000001100101;
assign LUT_1[40989] = 32'b00000000000000000110010011100001;
assign LUT_1[40990] = 32'b00000000000000001000101111110110;
assign LUT_1[40991] = 32'b00000000000000000010000001110010;
assign LUT_1[40992] = 32'b00000000000000000100111001110110;
assign LUT_1[40993] = 32'b11111111111111111110001011110010;
assign LUT_1[40994] = 32'b00000000000000000000101000000111;
assign LUT_1[40995] = 32'b11111111111111111001111010000011;
assign LUT_1[40996] = 32'b00000000000000001100110011001101;
assign LUT_1[40997] = 32'b00000000000000000110000101001001;
assign LUT_1[40998] = 32'b00000000000000001000100001011110;
assign LUT_1[40999] = 32'b00000000000000000001110011011010;
assign LUT_1[41000] = 32'b00000000000000000100000111101011;
assign LUT_1[41001] = 32'b11111111111111111101011001100111;
assign LUT_1[41002] = 32'b11111111111111111111110101111100;
assign LUT_1[41003] = 32'b11111111111111111001000111111000;
assign LUT_1[41004] = 32'b00000000000000001100000001000010;
assign LUT_1[41005] = 32'b00000000000000000101010010111110;
assign LUT_1[41006] = 32'b00000000000000000111101111010011;
assign LUT_1[41007] = 32'b00000000000000000001000001001111;
assign LUT_1[41008] = 32'b00000000000000000110110101011000;
assign LUT_1[41009] = 32'b00000000000000000000000111010100;
assign LUT_1[41010] = 32'b00000000000000000010100011101001;
assign LUT_1[41011] = 32'b11111111111111111011110101100101;
assign LUT_1[41012] = 32'b00000000000000001110101110101111;
assign LUT_1[41013] = 32'b00000000000000001000000000101011;
assign LUT_1[41014] = 32'b00000000000000001010011101000000;
assign LUT_1[41015] = 32'b00000000000000000011101110111100;
assign LUT_1[41016] = 32'b00000000000000000110000011001101;
assign LUT_1[41017] = 32'b11111111111111111111010101001001;
assign LUT_1[41018] = 32'b00000000000000000001110001011110;
assign LUT_1[41019] = 32'b11111111111111111011000011011010;
assign LUT_1[41020] = 32'b00000000000000001101111100100100;
assign LUT_1[41021] = 32'b00000000000000000111001110100000;
assign LUT_1[41022] = 32'b00000000000000001001101010110101;
assign LUT_1[41023] = 32'b00000000000000000010111100110001;
assign LUT_1[41024] = 32'b00000000000000000101111100011111;
assign LUT_1[41025] = 32'b11111111111111111111001110011011;
assign LUT_1[41026] = 32'b00000000000000000001101010110000;
assign LUT_1[41027] = 32'b11111111111111111010111100101100;
assign LUT_1[41028] = 32'b00000000000000001101110101110110;
assign LUT_1[41029] = 32'b00000000000000000111000111110010;
assign LUT_1[41030] = 32'b00000000000000001001100100000111;
assign LUT_1[41031] = 32'b00000000000000000010110110000011;
assign LUT_1[41032] = 32'b00000000000000000101001010010100;
assign LUT_1[41033] = 32'b11111111111111111110011100010000;
assign LUT_1[41034] = 32'b00000000000000000000111000100101;
assign LUT_1[41035] = 32'b11111111111111111010001010100001;
assign LUT_1[41036] = 32'b00000000000000001101000011101011;
assign LUT_1[41037] = 32'b00000000000000000110010101100111;
assign LUT_1[41038] = 32'b00000000000000001000110001111100;
assign LUT_1[41039] = 32'b00000000000000000010000011111000;
assign LUT_1[41040] = 32'b00000000000000000111111000000001;
assign LUT_1[41041] = 32'b00000000000000000001001001111101;
assign LUT_1[41042] = 32'b00000000000000000011100110010010;
assign LUT_1[41043] = 32'b11111111111111111100111000001110;
assign LUT_1[41044] = 32'b00000000000000001111110001011000;
assign LUT_1[41045] = 32'b00000000000000001001000011010100;
assign LUT_1[41046] = 32'b00000000000000001011011111101001;
assign LUT_1[41047] = 32'b00000000000000000100110001100101;
assign LUT_1[41048] = 32'b00000000000000000111000101110110;
assign LUT_1[41049] = 32'b00000000000000000000010111110010;
assign LUT_1[41050] = 32'b00000000000000000010110100000111;
assign LUT_1[41051] = 32'b11111111111111111100000110000011;
assign LUT_1[41052] = 32'b00000000000000001110111111001101;
assign LUT_1[41053] = 32'b00000000000000001000010001001001;
assign LUT_1[41054] = 32'b00000000000000001010101101011110;
assign LUT_1[41055] = 32'b00000000000000000011111111011010;
assign LUT_1[41056] = 32'b00000000000000000110110111011110;
assign LUT_1[41057] = 32'b00000000000000000000001001011010;
assign LUT_1[41058] = 32'b00000000000000000010100101101111;
assign LUT_1[41059] = 32'b11111111111111111011110111101011;
assign LUT_1[41060] = 32'b00000000000000001110110000110101;
assign LUT_1[41061] = 32'b00000000000000001000000010110001;
assign LUT_1[41062] = 32'b00000000000000001010011111000110;
assign LUT_1[41063] = 32'b00000000000000000011110001000010;
assign LUT_1[41064] = 32'b00000000000000000110000101010011;
assign LUT_1[41065] = 32'b11111111111111111111010111001111;
assign LUT_1[41066] = 32'b00000000000000000001110011100100;
assign LUT_1[41067] = 32'b11111111111111111011000101100000;
assign LUT_1[41068] = 32'b00000000000000001101111110101010;
assign LUT_1[41069] = 32'b00000000000000000111010000100110;
assign LUT_1[41070] = 32'b00000000000000001001101100111011;
assign LUT_1[41071] = 32'b00000000000000000010111110110111;
assign LUT_1[41072] = 32'b00000000000000001000110011000000;
assign LUT_1[41073] = 32'b00000000000000000010000100111100;
assign LUT_1[41074] = 32'b00000000000000000100100001010001;
assign LUT_1[41075] = 32'b11111111111111111101110011001101;
assign LUT_1[41076] = 32'b00000000000000010000101100010111;
assign LUT_1[41077] = 32'b00000000000000001001111110010011;
assign LUT_1[41078] = 32'b00000000000000001100011010101000;
assign LUT_1[41079] = 32'b00000000000000000101101100100100;
assign LUT_1[41080] = 32'b00000000000000001000000000110101;
assign LUT_1[41081] = 32'b00000000000000000001010010110001;
assign LUT_1[41082] = 32'b00000000000000000011101111000110;
assign LUT_1[41083] = 32'b11111111111111111101000001000010;
assign LUT_1[41084] = 32'b00000000000000001111111010001100;
assign LUT_1[41085] = 32'b00000000000000001001001100001000;
assign LUT_1[41086] = 32'b00000000000000001011101000011101;
assign LUT_1[41087] = 32'b00000000000000000100111010011001;
assign LUT_1[41088] = 32'b00000000000000000110111110111010;
assign LUT_1[41089] = 32'b00000000000000000000010000110110;
assign LUT_1[41090] = 32'b00000000000000000010101101001011;
assign LUT_1[41091] = 32'b11111111111111111011111111000111;
assign LUT_1[41092] = 32'b00000000000000001110111000010001;
assign LUT_1[41093] = 32'b00000000000000001000001010001101;
assign LUT_1[41094] = 32'b00000000000000001010100110100010;
assign LUT_1[41095] = 32'b00000000000000000011111000011110;
assign LUT_1[41096] = 32'b00000000000000000110001100101111;
assign LUT_1[41097] = 32'b11111111111111111111011110101011;
assign LUT_1[41098] = 32'b00000000000000000001111011000000;
assign LUT_1[41099] = 32'b11111111111111111011001100111100;
assign LUT_1[41100] = 32'b00000000000000001110000110000110;
assign LUT_1[41101] = 32'b00000000000000000111011000000010;
assign LUT_1[41102] = 32'b00000000000000001001110100010111;
assign LUT_1[41103] = 32'b00000000000000000011000110010011;
assign LUT_1[41104] = 32'b00000000000000001000111010011100;
assign LUT_1[41105] = 32'b00000000000000000010001100011000;
assign LUT_1[41106] = 32'b00000000000000000100101000101101;
assign LUT_1[41107] = 32'b11111111111111111101111010101001;
assign LUT_1[41108] = 32'b00000000000000010000110011110011;
assign LUT_1[41109] = 32'b00000000000000001010000101101111;
assign LUT_1[41110] = 32'b00000000000000001100100010000100;
assign LUT_1[41111] = 32'b00000000000000000101110100000000;
assign LUT_1[41112] = 32'b00000000000000001000001000010001;
assign LUT_1[41113] = 32'b00000000000000000001011010001101;
assign LUT_1[41114] = 32'b00000000000000000011110110100010;
assign LUT_1[41115] = 32'b11111111111111111101001000011110;
assign LUT_1[41116] = 32'b00000000000000010000000001101000;
assign LUT_1[41117] = 32'b00000000000000001001010011100100;
assign LUT_1[41118] = 32'b00000000000000001011101111111001;
assign LUT_1[41119] = 32'b00000000000000000101000001110101;
assign LUT_1[41120] = 32'b00000000000000000111111001111001;
assign LUT_1[41121] = 32'b00000000000000000001001011110101;
assign LUT_1[41122] = 32'b00000000000000000011101000001010;
assign LUT_1[41123] = 32'b11111111111111111100111010000110;
assign LUT_1[41124] = 32'b00000000000000001111110011010000;
assign LUT_1[41125] = 32'b00000000000000001001000101001100;
assign LUT_1[41126] = 32'b00000000000000001011100001100001;
assign LUT_1[41127] = 32'b00000000000000000100110011011101;
assign LUT_1[41128] = 32'b00000000000000000111000111101110;
assign LUT_1[41129] = 32'b00000000000000000000011001101010;
assign LUT_1[41130] = 32'b00000000000000000010110101111111;
assign LUT_1[41131] = 32'b11111111111111111100000111111011;
assign LUT_1[41132] = 32'b00000000000000001111000001000101;
assign LUT_1[41133] = 32'b00000000000000001000010011000001;
assign LUT_1[41134] = 32'b00000000000000001010101111010110;
assign LUT_1[41135] = 32'b00000000000000000100000001010010;
assign LUT_1[41136] = 32'b00000000000000001001110101011011;
assign LUT_1[41137] = 32'b00000000000000000011000111010111;
assign LUT_1[41138] = 32'b00000000000000000101100011101100;
assign LUT_1[41139] = 32'b11111111111111111110110101101000;
assign LUT_1[41140] = 32'b00000000000000010001101110110010;
assign LUT_1[41141] = 32'b00000000000000001011000000101110;
assign LUT_1[41142] = 32'b00000000000000001101011101000011;
assign LUT_1[41143] = 32'b00000000000000000110101110111111;
assign LUT_1[41144] = 32'b00000000000000001001000011010000;
assign LUT_1[41145] = 32'b00000000000000000010010101001100;
assign LUT_1[41146] = 32'b00000000000000000100110001100001;
assign LUT_1[41147] = 32'b11111111111111111110000011011101;
assign LUT_1[41148] = 32'b00000000000000010000111100100111;
assign LUT_1[41149] = 32'b00000000000000001010001110100011;
assign LUT_1[41150] = 32'b00000000000000001100101010111000;
assign LUT_1[41151] = 32'b00000000000000000101111100110100;
assign LUT_1[41152] = 32'b00000000000000001000111100100010;
assign LUT_1[41153] = 32'b00000000000000000010001110011110;
assign LUT_1[41154] = 32'b00000000000000000100101010110011;
assign LUT_1[41155] = 32'b11111111111111111101111100101111;
assign LUT_1[41156] = 32'b00000000000000010000110101111001;
assign LUT_1[41157] = 32'b00000000000000001010000111110101;
assign LUT_1[41158] = 32'b00000000000000001100100100001010;
assign LUT_1[41159] = 32'b00000000000000000101110110000110;
assign LUT_1[41160] = 32'b00000000000000001000001010010111;
assign LUT_1[41161] = 32'b00000000000000000001011100010011;
assign LUT_1[41162] = 32'b00000000000000000011111000101000;
assign LUT_1[41163] = 32'b11111111111111111101001010100100;
assign LUT_1[41164] = 32'b00000000000000010000000011101110;
assign LUT_1[41165] = 32'b00000000000000001001010101101010;
assign LUT_1[41166] = 32'b00000000000000001011110001111111;
assign LUT_1[41167] = 32'b00000000000000000101000011111011;
assign LUT_1[41168] = 32'b00000000000000001010111000000100;
assign LUT_1[41169] = 32'b00000000000000000100001010000000;
assign LUT_1[41170] = 32'b00000000000000000110100110010101;
assign LUT_1[41171] = 32'b11111111111111111111111000010001;
assign LUT_1[41172] = 32'b00000000000000010010110001011011;
assign LUT_1[41173] = 32'b00000000000000001100000011010111;
assign LUT_1[41174] = 32'b00000000000000001110011111101100;
assign LUT_1[41175] = 32'b00000000000000000111110001101000;
assign LUT_1[41176] = 32'b00000000000000001010000101111001;
assign LUT_1[41177] = 32'b00000000000000000011010111110101;
assign LUT_1[41178] = 32'b00000000000000000101110100001010;
assign LUT_1[41179] = 32'b11111111111111111111000110000110;
assign LUT_1[41180] = 32'b00000000000000010001111111010000;
assign LUT_1[41181] = 32'b00000000000000001011010001001100;
assign LUT_1[41182] = 32'b00000000000000001101101101100001;
assign LUT_1[41183] = 32'b00000000000000000110111111011101;
assign LUT_1[41184] = 32'b00000000000000001001110111100001;
assign LUT_1[41185] = 32'b00000000000000000011001001011101;
assign LUT_1[41186] = 32'b00000000000000000101100101110010;
assign LUT_1[41187] = 32'b11111111111111111110110111101110;
assign LUT_1[41188] = 32'b00000000000000010001110000111000;
assign LUT_1[41189] = 32'b00000000000000001011000010110100;
assign LUT_1[41190] = 32'b00000000000000001101011111001001;
assign LUT_1[41191] = 32'b00000000000000000110110001000101;
assign LUT_1[41192] = 32'b00000000000000001001000101010110;
assign LUT_1[41193] = 32'b00000000000000000010010111010010;
assign LUT_1[41194] = 32'b00000000000000000100110011100111;
assign LUT_1[41195] = 32'b11111111111111111110000101100011;
assign LUT_1[41196] = 32'b00000000000000010000111110101101;
assign LUT_1[41197] = 32'b00000000000000001010010000101001;
assign LUT_1[41198] = 32'b00000000000000001100101100111110;
assign LUT_1[41199] = 32'b00000000000000000101111110111010;
assign LUT_1[41200] = 32'b00000000000000001011110011000011;
assign LUT_1[41201] = 32'b00000000000000000101000100111111;
assign LUT_1[41202] = 32'b00000000000000000111100001010100;
assign LUT_1[41203] = 32'b00000000000000000000110011010000;
assign LUT_1[41204] = 32'b00000000000000010011101100011010;
assign LUT_1[41205] = 32'b00000000000000001100111110010110;
assign LUT_1[41206] = 32'b00000000000000001111011010101011;
assign LUT_1[41207] = 32'b00000000000000001000101100100111;
assign LUT_1[41208] = 32'b00000000000000001011000000111000;
assign LUT_1[41209] = 32'b00000000000000000100010010110100;
assign LUT_1[41210] = 32'b00000000000000000110101111001001;
assign LUT_1[41211] = 32'b00000000000000000000000001000101;
assign LUT_1[41212] = 32'b00000000000000010010111010001111;
assign LUT_1[41213] = 32'b00000000000000001100001100001011;
assign LUT_1[41214] = 32'b00000000000000001110101000100000;
assign LUT_1[41215] = 32'b00000000000000000111111010011100;
assign LUT_1[41216] = 32'b00000000000000000001110011000011;
assign LUT_1[41217] = 32'b11111111111111111011000100111111;
assign LUT_1[41218] = 32'b11111111111111111101100001010100;
assign LUT_1[41219] = 32'b11111111111111110110110011010000;
assign LUT_1[41220] = 32'b00000000000000001001101100011010;
assign LUT_1[41221] = 32'b00000000000000000010111110010110;
assign LUT_1[41222] = 32'b00000000000000000101011010101011;
assign LUT_1[41223] = 32'b11111111111111111110101100100111;
assign LUT_1[41224] = 32'b00000000000000000001000000111000;
assign LUT_1[41225] = 32'b11111111111111111010010010110100;
assign LUT_1[41226] = 32'b11111111111111111100101111001001;
assign LUT_1[41227] = 32'b11111111111111110110000001000101;
assign LUT_1[41228] = 32'b00000000000000001000111010001111;
assign LUT_1[41229] = 32'b00000000000000000010001100001011;
assign LUT_1[41230] = 32'b00000000000000000100101000100000;
assign LUT_1[41231] = 32'b11111111111111111101111010011100;
assign LUT_1[41232] = 32'b00000000000000000011101110100101;
assign LUT_1[41233] = 32'b11111111111111111101000000100001;
assign LUT_1[41234] = 32'b11111111111111111111011100110110;
assign LUT_1[41235] = 32'b11111111111111111000101110110010;
assign LUT_1[41236] = 32'b00000000000000001011100111111100;
assign LUT_1[41237] = 32'b00000000000000000100111001111000;
assign LUT_1[41238] = 32'b00000000000000000111010110001101;
assign LUT_1[41239] = 32'b00000000000000000000101000001001;
assign LUT_1[41240] = 32'b00000000000000000010111100011010;
assign LUT_1[41241] = 32'b11111111111111111100001110010110;
assign LUT_1[41242] = 32'b11111111111111111110101010101011;
assign LUT_1[41243] = 32'b11111111111111110111111100100111;
assign LUT_1[41244] = 32'b00000000000000001010110101110001;
assign LUT_1[41245] = 32'b00000000000000000100000111101101;
assign LUT_1[41246] = 32'b00000000000000000110100100000010;
assign LUT_1[41247] = 32'b11111111111111111111110101111110;
assign LUT_1[41248] = 32'b00000000000000000010101110000010;
assign LUT_1[41249] = 32'b11111111111111111011111111111110;
assign LUT_1[41250] = 32'b11111111111111111110011100010011;
assign LUT_1[41251] = 32'b11111111111111110111101110001111;
assign LUT_1[41252] = 32'b00000000000000001010100111011001;
assign LUT_1[41253] = 32'b00000000000000000011111001010101;
assign LUT_1[41254] = 32'b00000000000000000110010101101010;
assign LUT_1[41255] = 32'b11111111111111111111100111100110;
assign LUT_1[41256] = 32'b00000000000000000001111011110111;
assign LUT_1[41257] = 32'b11111111111111111011001101110011;
assign LUT_1[41258] = 32'b11111111111111111101101010001000;
assign LUT_1[41259] = 32'b11111111111111110110111100000100;
assign LUT_1[41260] = 32'b00000000000000001001110101001110;
assign LUT_1[41261] = 32'b00000000000000000011000111001010;
assign LUT_1[41262] = 32'b00000000000000000101100011011111;
assign LUT_1[41263] = 32'b11111111111111111110110101011011;
assign LUT_1[41264] = 32'b00000000000000000100101001100100;
assign LUT_1[41265] = 32'b11111111111111111101111011100000;
assign LUT_1[41266] = 32'b00000000000000000000010111110101;
assign LUT_1[41267] = 32'b11111111111111111001101001110001;
assign LUT_1[41268] = 32'b00000000000000001100100010111011;
assign LUT_1[41269] = 32'b00000000000000000101110100110111;
assign LUT_1[41270] = 32'b00000000000000001000010001001100;
assign LUT_1[41271] = 32'b00000000000000000001100011001000;
assign LUT_1[41272] = 32'b00000000000000000011110111011001;
assign LUT_1[41273] = 32'b11111111111111111101001001010101;
assign LUT_1[41274] = 32'b11111111111111111111100101101010;
assign LUT_1[41275] = 32'b11111111111111111000110111100110;
assign LUT_1[41276] = 32'b00000000000000001011110000110000;
assign LUT_1[41277] = 32'b00000000000000000101000010101100;
assign LUT_1[41278] = 32'b00000000000000000111011111000001;
assign LUT_1[41279] = 32'b00000000000000000000110000111101;
assign LUT_1[41280] = 32'b00000000000000000011110000101011;
assign LUT_1[41281] = 32'b11111111111111111101000010100111;
assign LUT_1[41282] = 32'b11111111111111111111011110111100;
assign LUT_1[41283] = 32'b11111111111111111000110000111000;
assign LUT_1[41284] = 32'b00000000000000001011101010000010;
assign LUT_1[41285] = 32'b00000000000000000100111011111110;
assign LUT_1[41286] = 32'b00000000000000000111011000010011;
assign LUT_1[41287] = 32'b00000000000000000000101010001111;
assign LUT_1[41288] = 32'b00000000000000000010111110100000;
assign LUT_1[41289] = 32'b11111111111111111100010000011100;
assign LUT_1[41290] = 32'b11111111111111111110101100110001;
assign LUT_1[41291] = 32'b11111111111111110111111110101101;
assign LUT_1[41292] = 32'b00000000000000001010110111110111;
assign LUT_1[41293] = 32'b00000000000000000100001001110011;
assign LUT_1[41294] = 32'b00000000000000000110100110001000;
assign LUT_1[41295] = 32'b11111111111111111111111000000100;
assign LUT_1[41296] = 32'b00000000000000000101101100001101;
assign LUT_1[41297] = 32'b11111111111111111110111110001001;
assign LUT_1[41298] = 32'b00000000000000000001011010011110;
assign LUT_1[41299] = 32'b11111111111111111010101100011010;
assign LUT_1[41300] = 32'b00000000000000001101100101100100;
assign LUT_1[41301] = 32'b00000000000000000110110111100000;
assign LUT_1[41302] = 32'b00000000000000001001010011110101;
assign LUT_1[41303] = 32'b00000000000000000010100101110001;
assign LUT_1[41304] = 32'b00000000000000000100111010000010;
assign LUT_1[41305] = 32'b11111111111111111110001011111110;
assign LUT_1[41306] = 32'b00000000000000000000101000010011;
assign LUT_1[41307] = 32'b11111111111111111001111010001111;
assign LUT_1[41308] = 32'b00000000000000001100110011011001;
assign LUT_1[41309] = 32'b00000000000000000110000101010101;
assign LUT_1[41310] = 32'b00000000000000001000100001101010;
assign LUT_1[41311] = 32'b00000000000000000001110011100110;
assign LUT_1[41312] = 32'b00000000000000000100101011101010;
assign LUT_1[41313] = 32'b11111111111111111101111101100110;
assign LUT_1[41314] = 32'b00000000000000000000011001111011;
assign LUT_1[41315] = 32'b11111111111111111001101011110111;
assign LUT_1[41316] = 32'b00000000000000001100100101000001;
assign LUT_1[41317] = 32'b00000000000000000101110110111101;
assign LUT_1[41318] = 32'b00000000000000001000010011010010;
assign LUT_1[41319] = 32'b00000000000000000001100101001110;
assign LUT_1[41320] = 32'b00000000000000000011111001011111;
assign LUT_1[41321] = 32'b11111111111111111101001011011011;
assign LUT_1[41322] = 32'b11111111111111111111100111110000;
assign LUT_1[41323] = 32'b11111111111111111000111001101100;
assign LUT_1[41324] = 32'b00000000000000001011110010110110;
assign LUT_1[41325] = 32'b00000000000000000101000100110010;
assign LUT_1[41326] = 32'b00000000000000000111100001000111;
assign LUT_1[41327] = 32'b00000000000000000000110011000011;
assign LUT_1[41328] = 32'b00000000000000000110100111001100;
assign LUT_1[41329] = 32'b11111111111111111111111001001000;
assign LUT_1[41330] = 32'b00000000000000000010010101011101;
assign LUT_1[41331] = 32'b11111111111111111011100111011001;
assign LUT_1[41332] = 32'b00000000000000001110100000100011;
assign LUT_1[41333] = 32'b00000000000000000111110010011111;
assign LUT_1[41334] = 32'b00000000000000001010001110110100;
assign LUT_1[41335] = 32'b00000000000000000011100000110000;
assign LUT_1[41336] = 32'b00000000000000000101110101000001;
assign LUT_1[41337] = 32'b11111111111111111111000110111101;
assign LUT_1[41338] = 32'b00000000000000000001100011010010;
assign LUT_1[41339] = 32'b11111111111111111010110101001110;
assign LUT_1[41340] = 32'b00000000000000001101101110011000;
assign LUT_1[41341] = 32'b00000000000000000111000000010100;
assign LUT_1[41342] = 32'b00000000000000001001011100101001;
assign LUT_1[41343] = 32'b00000000000000000010101110100101;
assign LUT_1[41344] = 32'b00000000000000000100110011000110;
assign LUT_1[41345] = 32'b11111111111111111110000101000010;
assign LUT_1[41346] = 32'b00000000000000000000100001010111;
assign LUT_1[41347] = 32'b11111111111111111001110011010011;
assign LUT_1[41348] = 32'b00000000000000001100101100011101;
assign LUT_1[41349] = 32'b00000000000000000101111110011001;
assign LUT_1[41350] = 32'b00000000000000001000011010101110;
assign LUT_1[41351] = 32'b00000000000000000001101100101010;
assign LUT_1[41352] = 32'b00000000000000000100000000111011;
assign LUT_1[41353] = 32'b11111111111111111101010010110111;
assign LUT_1[41354] = 32'b11111111111111111111101111001100;
assign LUT_1[41355] = 32'b11111111111111111001000001001000;
assign LUT_1[41356] = 32'b00000000000000001011111010010010;
assign LUT_1[41357] = 32'b00000000000000000101001100001110;
assign LUT_1[41358] = 32'b00000000000000000111101000100011;
assign LUT_1[41359] = 32'b00000000000000000000111010011111;
assign LUT_1[41360] = 32'b00000000000000000110101110101000;
assign LUT_1[41361] = 32'b00000000000000000000000000100100;
assign LUT_1[41362] = 32'b00000000000000000010011100111001;
assign LUT_1[41363] = 32'b11111111111111111011101110110101;
assign LUT_1[41364] = 32'b00000000000000001110100111111111;
assign LUT_1[41365] = 32'b00000000000000000111111001111011;
assign LUT_1[41366] = 32'b00000000000000001010010110010000;
assign LUT_1[41367] = 32'b00000000000000000011101000001100;
assign LUT_1[41368] = 32'b00000000000000000101111100011101;
assign LUT_1[41369] = 32'b11111111111111111111001110011001;
assign LUT_1[41370] = 32'b00000000000000000001101010101110;
assign LUT_1[41371] = 32'b11111111111111111010111100101010;
assign LUT_1[41372] = 32'b00000000000000001101110101110100;
assign LUT_1[41373] = 32'b00000000000000000111000111110000;
assign LUT_1[41374] = 32'b00000000000000001001100100000101;
assign LUT_1[41375] = 32'b00000000000000000010110110000001;
assign LUT_1[41376] = 32'b00000000000000000101101110000101;
assign LUT_1[41377] = 32'b11111111111111111111000000000001;
assign LUT_1[41378] = 32'b00000000000000000001011100010110;
assign LUT_1[41379] = 32'b11111111111111111010101110010010;
assign LUT_1[41380] = 32'b00000000000000001101100111011100;
assign LUT_1[41381] = 32'b00000000000000000110111001011000;
assign LUT_1[41382] = 32'b00000000000000001001010101101101;
assign LUT_1[41383] = 32'b00000000000000000010100111101001;
assign LUT_1[41384] = 32'b00000000000000000100111011111010;
assign LUT_1[41385] = 32'b11111111111111111110001101110110;
assign LUT_1[41386] = 32'b00000000000000000000101010001011;
assign LUT_1[41387] = 32'b11111111111111111001111100000111;
assign LUT_1[41388] = 32'b00000000000000001100110101010001;
assign LUT_1[41389] = 32'b00000000000000000110000111001101;
assign LUT_1[41390] = 32'b00000000000000001000100011100010;
assign LUT_1[41391] = 32'b00000000000000000001110101011110;
assign LUT_1[41392] = 32'b00000000000000000111101001100111;
assign LUT_1[41393] = 32'b00000000000000000000111011100011;
assign LUT_1[41394] = 32'b00000000000000000011010111111000;
assign LUT_1[41395] = 32'b11111111111111111100101001110100;
assign LUT_1[41396] = 32'b00000000000000001111100010111110;
assign LUT_1[41397] = 32'b00000000000000001000110100111010;
assign LUT_1[41398] = 32'b00000000000000001011010001001111;
assign LUT_1[41399] = 32'b00000000000000000100100011001011;
assign LUT_1[41400] = 32'b00000000000000000110110111011100;
assign LUT_1[41401] = 32'b00000000000000000000001001011000;
assign LUT_1[41402] = 32'b00000000000000000010100101101101;
assign LUT_1[41403] = 32'b11111111111111111011110111101001;
assign LUT_1[41404] = 32'b00000000000000001110110000110011;
assign LUT_1[41405] = 32'b00000000000000001000000010101111;
assign LUT_1[41406] = 32'b00000000000000001010011111000100;
assign LUT_1[41407] = 32'b00000000000000000011110001000000;
assign LUT_1[41408] = 32'b00000000000000000110110000101110;
assign LUT_1[41409] = 32'b00000000000000000000000010101010;
assign LUT_1[41410] = 32'b00000000000000000010011110111111;
assign LUT_1[41411] = 32'b11111111111111111011110000111011;
assign LUT_1[41412] = 32'b00000000000000001110101010000101;
assign LUT_1[41413] = 32'b00000000000000000111111100000001;
assign LUT_1[41414] = 32'b00000000000000001010011000010110;
assign LUT_1[41415] = 32'b00000000000000000011101010010010;
assign LUT_1[41416] = 32'b00000000000000000101111110100011;
assign LUT_1[41417] = 32'b11111111111111111111010000011111;
assign LUT_1[41418] = 32'b00000000000000000001101100110100;
assign LUT_1[41419] = 32'b11111111111111111010111110110000;
assign LUT_1[41420] = 32'b00000000000000001101110111111010;
assign LUT_1[41421] = 32'b00000000000000000111001001110110;
assign LUT_1[41422] = 32'b00000000000000001001100110001011;
assign LUT_1[41423] = 32'b00000000000000000010111000000111;
assign LUT_1[41424] = 32'b00000000000000001000101100010000;
assign LUT_1[41425] = 32'b00000000000000000001111110001100;
assign LUT_1[41426] = 32'b00000000000000000100011010100001;
assign LUT_1[41427] = 32'b11111111111111111101101100011101;
assign LUT_1[41428] = 32'b00000000000000010000100101100111;
assign LUT_1[41429] = 32'b00000000000000001001110111100011;
assign LUT_1[41430] = 32'b00000000000000001100010011111000;
assign LUT_1[41431] = 32'b00000000000000000101100101110100;
assign LUT_1[41432] = 32'b00000000000000000111111010000101;
assign LUT_1[41433] = 32'b00000000000000000001001100000001;
assign LUT_1[41434] = 32'b00000000000000000011101000010110;
assign LUT_1[41435] = 32'b11111111111111111100111010010010;
assign LUT_1[41436] = 32'b00000000000000001111110011011100;
assign LUT_1[41437] = 32'b00000000000000001001000101011000;
assign LUT_1[41438] = 32'b00000000000000001011100001101101;
assign LUT_1[41439] = 32'b00000000000000000100110011101001;
assign LUT_1[41440] = 32'b00000000000000000111101011101101;
assign LUT_1[41441] = 32'b00000000000000000000111101101001;
assign LUT_1[41442] = 32'b00000000000000000011011001111110;
assign LUT_1[41443] = 32'b11111111111111111100101011111010;
assign LUT_1[41444] = 32'b00000000000000001111100101000100;
assign LUT_1[41445] = 32'b00000000000000001000110111000000;
assign LUT_1[41446] = 32'b00000000000000001011010011010101;
assign LUT_1[41447] = 32'b00000000000000000100100101010001;
assign LUT_1[41448] = 32'b00000000000000000110111001100010;
assign LUT_1[41449] = 32'b00000000000000000000001011011110;
assign LUT_1[41450] = 32'b00000000000000000010100111110011;
assign LUT_1[41451] = 32'b11111111111111111011111001101111;
assign LUT_1[41452] = 32'b00000000000000001110110010111001;
assign LUT_1[41453] = 32'b00000000000000001000000100110101;
assign LUT_1[41454] = 32'b00000000000000001010100001001010;
assign LUT_1[41455] = 32'b00000000000000000011110011000110;
assign LUT_1[41456] = 32'b00000000000000001001100111001111;
assign LUT_1[41457] = 32'b00000000000000000010111001001011;
assign LUT_1[41458] = 32'b00000000000000000101010101100000;
assign LUT_1[41459] = 32'b11111111111111111110100111011100;
assign LUT_1[41460] = 32'b00000000000000010001100000100110;
assign LUT_1[41461] = 32'b00000000000000001010110010100010;
assign LUT_1[41462] = 32'b00000000000000001101001110110111;
assign LUT_1[41463] = 32'b00000000000000000110100000110011;
assign LUT_1[41464] = 32'b00000000000000001000110101000100;
assign LUT_1[41465] = 32'b00000000000000000010000111000000;
assign LUT_1[41466] = 32'b00000000000000000100100011010101;
assign LUT_1[41467] = 32'b11111111111111111101110101010001;
assign LUT_1[41468] = 32'b00000000000000010000101110011011;
assign LUT_1[41469] = 32'b00000000000000001010000000010111;
assign LUT_1[41470] = 32'b00000000000000001100011100101100;
assign LUT_1[41471] = 32'b00000000000000000101101110101000;
assign LUT_1[41472] = 32'b11111111111111111101101101010100;
assign LUT_1[41473] = 32'b11111111111111110110111111010000;
assign LUT_1[41474] = 32'b11111111111111111001011011100101;
assign LUT_1[41475] = 32'b11111111111111110010101101100001;
assign LUT_1[41476] = 32'b00000000000000000101100110101011;
assign LUT_1[41477] = 32'b11111111111111111110111000100111;
assign LUT_1[41478] = 32'b00000000000000000001010100111100;
assign LUT_1[41479] = 32'b11111111111111111010100110111000;
assign LUT_1[41480] = 32'b11111111111111111100111011001001;
assign LUT_1[41481] = 32'b11111111111111110110001101000101;
assign LUT_1[41482] = 32'b11111111111111111000101001011010;
assign LUT_1[41483] = 32'b11111111111111110001111011010110;
assign LUT_1[41484] = 32'b00000000000000000100110100100000;
assign LUT_1[41485] = 32'b11111111111111111110000110011100;
assign LUT_1[41486] = 32'b00000000000000000000100010110001;
assign LUT_1[41487] = 32'b11111111111111111001110100101101;
assign LUT_1[41488] = 32'b11111111111111111111101000110110;
assign LUT_1[41489] = 32'b11111111111111111000111010110010;
assign LUT_1[41490] = 32'b11111111111111111011010111000111;
assign LUT_1[41491] = 32'b11111111111111110100101001000011;
assign LUT_1[41492] = 32'b00000000000000000111100010001101;
assign LUT_1[41493] = 32'b00000000000000000000110100001001;
assign LUT_1[41494] = 32'b00000000000000000011010000011110;
assign LUT_1[41495] = 32'b11111111111111111100100010011010;
assign LUT_1[41496] = 32'b11111111111111111110110110101011;
assign LUT_1[41497] = 32'b11111111111111111000001000100111;
assign LUT_1[41498] = 32'b11111111111111111010100100111100;
assign LUT_1[41499] = 32'b11111111111111110011110110111000;
assign LUT_1[41500] = 32'b00000000000000000110110000000010;
assign LUT_1[41501] = 32'b00000000000000000000000001111110;
assign LUT_1[41502] = 32'b00000000000000000010011110010011;
assign LUT_1[41503] = 32'b11111111111111111011110000001111;
assign LUT_1[41504] = 32'b11111111111111111110101000010011;
assign LUT_1[41505] = 32'b11111111111111110111111010001111;
assign LUT_1[41506] = 32'b11111111111111111010010110100100;
assign LUT_1[41507] = 32'b11111111111111110011101000100000;
assign LUT_1[41508] = 32'b00000000000000000110100001101010;
assign LUT_1[41509] = 32'b11111111111111111111110011100110;
assign LUT_1[41510] = 32'b00000000000000000010001111111011;
assign LUT_1[41511] = 32'b11111111111111111011100001110111;
assign LUT_1[41512] = 32'b11111111111111111101110110001000;
assign LUT_1[41513] = 32'b11111111111111110111001000000100;
assign LUT_1[41514] = 32'b11111111111111111001100100011001;
assign LUT_1[41515] = 32'b11111111111111110010110110010101;
assign LUT_1[41516] = 32'b00000000000000000101101111011111;
assign LUT_1[41517] = 32'b11111111111111111111000001011011;
assign LUT_1[41518] = 32'b00000000000000000001011101110000;
assign LUT_1[41519] = 32'b11111111111111111010101111101100;
assign LUT_1[41520] = 32'b00000000000000000000100011110101;
assign LUT_1[41521] = 32'b11111111111111111001110101110001;
assign LUT_1[41522] = 32'b11111111111111111100010010000110;
assign LUT_1[41523] = 32'b11111111111111110101100100000010;
assign LUT_1[41524] = 32'b00000000000000001000011101001100;
assign LUT_1[41525] = 32'b00000000000000000001101111001000;
assign LUT_1[41526] = 32'b00000000000000000100001011011101;
assign LUT_1[41527] = 32'b11111111111111111101011101011001;
assign LUT_1[41528] = 32'b11111111111111111111110001101010;
assign LUT_1[41529] = 32'b11111111111111111001000011100110;
assign LUT_1[41530] = 32'b11111111111111111011011111111011;
assign LUT_1[41531] = 32'b11111111111111110100110001110111;
assign LUT_1[41532] = 32'b00000000000000000111101011000001;
assign LUT_1[41533] = 32'b00000000000000000000111100111101;
assign LUT_1[41534] = 32'b00000000000000000011011001010010;
assign LUT_1[41535] = 32'b11111111111111111100101011001110;
assign LUT_1[41536] = 32'b11111111111111111111101010111100;
assign LUT_1[41537] = 32'b11111111111111111000111100111000;
assign LUT_1[41538] = 32'b11111111111111111011011001001101;
assign LUT_1[41539] = 32'b11111111111111110100101011001001;
assign LUT_1[41540] = 32'b00000000000000000111100100010011;
assign LUT_1[41541] = 32'b00000000000000000000110110001111;
assign LUT_1[41542] = 32'b00000000000000000011010010100100;
assign LUT_1[41543] = 32'b11111111111111111100100100100000;
assign LUT_1[41544] = 32'b11111111111111111110111000110001;
assign LUT_1[41545] = 32'b11111111111111111000001010101101;
assign LUT_1[41546] = 32'b11111111111111111010100111000010;
assign LUT_1[41547] = 32'b11111111111111110011111000111110;
assign LUT_1[41548] = 32'b00000000000000000110110010001000;
assign LUT_1[41549] = 32'b00000000000000000000000100000100;
assign LUT_1[41550] = 32'b00000000000000000010100000011001;
assign LUT_1[41551] = 32'b11111111111111111011110010010101;
assign LUT_1[41552] = 32'b00000000000000000001100110011110;
assign LUT_1[41553] = 32'b11111111111111111010111000011010;
assign LUT_1[41554] = 32'b11111111111111111101010100101111;
assign LUT_1[41555] = 32'b11111111111111110110100110101011;
assign LUT_1[41556] = 32'b00000000000000001001011111110101;
assign LUT_1[41557] = 32'b00000000000000000010110001110001;
assign LUT_1[41558] = 32'b00000000000000000101001110000110;
assign LUT_1[41559] = 32'b11111111111111111110100000000010;
assign LUT_1[41560] = 32'b00000000000000000000110100010011;
assign LUT_1[41561] = 32'b11111111111111111010000110001111;
assign LUT_1[41562] = 32'b11111111111111111100100010100100;
assign LUT_1[41563] = 32'b11111111111111110101110100100000;
assign LUT_1[41564] = 32'b00000000000000001000101101101010;
assign LUT_1[41565] = 32'b00000000000000000001111111100110;
assign LUT_1[41566] = 32'b00000000000000000100011011111011;
assign LUT_1[41567] = 32'b11111111111111111101101101110111;
assign LUT_1[41568] = 32'b00000000000000000000100101111011;
assign LUT_1[41569] = 32'b11111111111111111001110111110111;
assign LUT_1[41570] = 32'b11111111111111111100010100001100;
assign LUT_1[41571] = 32'b11111111111111110101100110001000;
assign LUT_1[41572] = 32'b00000000000000001000011111010010;
assign LUT_1[41573] = 32'b00000000000000000001110001001110;
assign LUT_1[41574] = 32'b00000000000000000100001101100011;
assign LUT_1[41575] = 32'b11111111111111111101011111011111;
assign LUT_1[41576] = 32'b11111111111111111111110011110000;
assign LUT_1[41577] = 32'b11111111111111111001000101101100;
assign LUT_1[41578] = 32'b11111111111111111011100010000001;
assign LUT_1[41579] = 32'b11111111111111110100110011111101;
assign LUT_1[41580] = 32'b00000000000000000111101101000111;
assign LUT_1[41581] = 32'b00000000000000000000111111000011;
assign LUT_1[41582] = 32'b00000000000000000011011011011000;
assign LUT_1[41583] = 32'b11111111111111111100101101010100;
assign LUT_1[41584] = 32'b00000000000000000010100001011101;
assign LUT_1[41585] = 32'b11111111111111111011110011011001;
assign LUT_1[41586] = 32'b11111111111111111110001111101110;
assign LUT_1[41587] = 32'b11111111111111110111100001101010;
assign LUT_1[41588] = 32'b00000000000000001010011010110100;
assign LUT_1[41589] = 32'b00000000000000000011101100110000;
assign LUT_1[41590] = 32'b00000000000000000110001001000101;
assign LUT_1[41591] = 32'b11111111111111111111011011000001;
assign LUT_1[41592] = 32'b00000000000000000001101111010010;
assign LUT_1[41593] = 32'b11111111111111111011000001001110;
assign LUT_1[41594] = 32'b11111111111111111101011101100011;
assign LUT_1[41595] = 32'b11111111111111110110101111011111;
assign LUT_1[41596] = 32'b00000000000000001001101000101001;
assign LUT_1[41597] = 32'b00000000000000000010111010100101;
assign LUT_1[41598] = 32'b00000000000000000101010110111010;
assign LUT_1[41599] = 32'b11111111111111111110101000110110;
assign LUT_1[41600] = 32'b00000000000000000000101101010111;
assign LUT_1[41601] = 32'b11111111111111111001111111010011;
assign LUT_1[41602] = 32'b11111111111111111100011011101000;
assign LUT_1[41603] = 32'b11111111111111110101101101100100;
assign LUT_1[41604] = 32'b00000000000000001000100110101110;
assign LUT_1[41605] = 32'b00000000000000000001111000101010;
assign LUT_1[41606] = 32'b00000000000000000100010100111111;
assign LUT_1[41607] = 32'b11111111111111111101100110111011;
assign LUT_1[41608] = 32'b11111111111111111111111011001100;
assign LUT_1[41609] = 32'b11111111111111111001001101001000;
assign LUT_1[41610] = 32'b11111111111111111011101001011101;
assign LUT_1[41611] = 32'b11111111111111110100111011011001;
assign LUT_1[41612] = 32'b00000000000000000111110100100011;
assign LUT_1[41613] = 32'b00000000000000000001000110011111;
assign LUT_1[41614] = 32'b00000000000000000011100010110100;
assign LUT_1[41615] = 32'b11111111111111111100110100110000;
assign LUT_1[41616] = 32'b00000000000000000010101000111001;
assign LUT_1[41617] = 32'b11111111111111111011111010110101;
assign LUT_1[41618] = 32'b11111111111111111110010111001010;
assign LUT_1[41619] = 32'b11111111111111110111101001000110;
assign LUT_1[41620] = 32'b00000000000000001010100010010000;
assign LUT_1[41621] = 32'b00000000000000000011110100001100;
assign LUT_1[41622] = 32'b00000000000000000110010000100001;
assign LUT_1[41623] = 32'b11111111111111111111100010011101;
assign LUT_1[41624] = 32'b00000000000000000001110110101110;
assign LUT_1[41625] = 32'b11111111111111111011001000101010;
assign LUT_1[41626] = 32'b11111111111111111101100100111111;
assign LUT_1[41627] = 32'b11111111111111110110110110111011;
assign LUT_1[41628] = 32'b00000000000000001001110000000101;
assign LUT_1[41629] = 32'b00000000000000000011000010000001;
assign LUT_1[41630] = 32'b00000000000000000101011110010110;
assign LUT_1[41631] = 32'b11111111111111111110110000010010;
assign LUT_1[41632] = 32'b00000000000000000001101000010110;
assign LUT_1[41633] = 32'b11111111111111111010111010010010;
assign LUT_1[41634] = 32'b11111111111111111101010110100111;
assign LUT_1[41635] = 32'b11111111111111110110101000100011;
assign LUT_1[41636] = 32'b00000000000000001001100001101101;
assign LUT_1[41637] = 32'b00000000000000000010110011101001;
assign LUT_1[41638] = 32'b00000000000000000101001111111110;
assign LUT_1[41639] = 32'b11111111111111111110100001111010;
assign LUT_1[41640] = 32'b00000000000000000000110110001011;
assign LUT_1[41641] = 32'b11111111111111111010001000000111;
assign LUT_1[41642] = 32'b11111111111111111100100100011100;
assign LUT_1[41643] = 32'b11111111111111110101110110011000;
assign LUT_1[41644] = 32'b00000000000000001000101111100010;
assign LUT_1[41645] = 32'b00000000000000000010000001011110;
assign LUT_1[41646] = 32'b00000000000000000100011101110011;
assign LUT_1[41647] = 32'b11111111111111111101101111101111;
assign LUT_1[41648] = 32'b00000000000000000011100011111000;
assign LUT_1[41649] = 32'b11111111111111111100110101110100;
assign LUT_1[41650] = 32'b11111111111111111111010010001001;
assign LUT_1[41651] = 32'b11111111111111111000100100000101;
assign LUT_1[41652] = 32'b00000000000000001011011101001111;
assign LUT_1[41653] = 32'b00000000000000000100101111001011;
assign LUT_1[41654] = 32'b00000000000000000111001011100000;
assign LUT_1[41655] = 32'b00000000000000000000011101011100;
assign LUT_1[41656] = 32'b00000000000000000010110001101101;
assign LUT_1[41657] = 32'b11111111111111111100000011101001;
assign LUT_1[41658] = 32'b11111111111111111110011111111110;
assign LUT_1[41659] = 32'b11111111111111110111110001111010;
assign LUT_1[41660] = 32'b00000000000000001010101011000100;
assign LUT_1[41661] = 32'b00000000000000000011111101000000;
assign LUT_1[41662] = 32'b00000000000000000110011001010101;
assign LUT_1[41663] = 32'b11111111111111111111101011010001;
assign LUT_1[41664] = 32'b00000000000000000010101010111111;
assign LUT_1[41665] = 32'b11111111111111111011111100111011;
assign LUT_1[41666] = 32'b11111111111111111110011001010000;
assign LUT_1[41667] = 32'b11111111111111110111101011001100;
assign LUT_1[41668] = 32'b00000000000000001010100100010110;
assign LUT_1[41669] = 32'b00000000000000000011110110010010;
assign LUT_1[41670] = 32'b00000000000000000110010010100111;
assign LUT_1[41671] = 32'b11111111111111111111100100100011;
assign LUT_1[41672] = 32'b00000000000000000001111000110100;
assign LUT_1[41673] = 32'b11111111111111111011001010110000;
assign LUT_1[41674] = 32'b11111111111111111101100111000101;
assign LUT_1[41675] = 32'b11111111111111110110111001000001;
assign LUT_1[41676] = 32'b00000000000000001001110010001011;
assign LUT_1[41677] = 32'b00000000000000000011000100000111;
assign LUT_1[41678] = 32'b00000000000000000101100000011100;
assign LUT_1[41679] = 32'b11111111111111111110110010011000;
assign LUT_1[41680] = 32'b00000000000000000100100110100001;
assign LUT_1[41681] = 32'b11111111111111111101111000011101;
assign LUT_1[41682] = 32'b00000000000000000000010100110010;
assign LUT_1[41683] = 32'b11111111111111111001100110101110;
assign LUT_1[41684] = 32'b00000000000000001100011111111000;
assign LUT_1[41685] = 32'b00000000000000000101110001110100;
assign LUT_1[41686] = 32'b00000000000000001000001110001001;
assign LUT_1[41687] = 32'b00000000000000000001100000000101;
assign LUT_1[41688] = 32'b00000000000000000011110100010110;
assign LUT_1[41689] = 32'b11111111111111111101000110010010;
assign LUT_1[41690] = 32'b11111111111111111111100010100111;
assign LUT_1[41691] = 32'b11111111111111111000110100100011;
assign LUT_1[41692] = 32'b00000000000000001011101101101101;
assign LUT_1[41693] = 32'b00000000000000000100111111101001;
assign LUT_1[41694] = 32'b00000000000000000111011011111110;
assign LUT_1[41695] = 32'b00000000000000000000101101111010;
assign LUT_1[41696] = 32'b00000000000000000011100101111110;
assign LUT_1[41697] = 32'b11111111111111111100110111111010;
assign LUT_1[41698] = 32'b11111111111111111111010100001111;
assign LUT_1[41699] = 32'b11111111111111111000100110001011;
assign LUT_1[41700] = 32'b00000000000000001011011111010101;
assign LUT_1[41701] = 32'b00000000000000000100110001010001;
assign LUT_1[41702] = 32'b00000000000000000111001101100110;
assign LUT_1[41703] = 32'b00000000000000000000011111100010;
assign LUT_1[41704] = 32'b00000000000000000010110011110011;
assign LUT_1[41705] = 32'b11111111111111111100000101101111;
assign LUT_1[41706] = 32'b11111111111111111110100010000100;
assign LUT_1[41707] = 32'b11111111111111110111110100000000;
assign LUT_1[41708] = 32'b00000000000000001010101101001010;
assign LUT_1[41709] = 32'b00000000000000000011111111000110;
assign LUT_1[41710] = 32'b00000000000000000110011011011011;
assign LUT_1[41711] = 32'b11111111111111111111101101010111;
assign LUT_1[41712] = 32'b00000000000000000101100001100000;
assign LUT_1[41713] = 32'b11111111111111111110110011011100;
assign LUT_1[41714] = 32'b00000000000000000001001111110001;
assign LUT_1[41715] = 32'b11111111111111111010100001101101;
assign LUT_1[41716] = 32'b00000000000000001101011010110111;
assign LUT_1[41717] = 32'b00000000000000000110101100110011;
assign LUT_1[41718] = 32'b00000000000000001001001001001000;
assign LUT_1[41719] = 32'b00000000000000000010011011000100;
assign LUT_1[41720] = 32'b00000000000000000100101111010101;
assign LUT_1[41721] = 32'b11111111111111111110000001010001;
assign LUT_1[41722] = 32'b00000000000000000000011101100110;
assign LUT_1[41723] = 32'b11111111111111111001101111100010;
assign LUT_1[41724] = 32'b00000000000000001100101000101100;
assign LUT_1[41725] = 32'b00000000000000000101111010101000;
assign LUT_1[41726] = 32'b00000000000000001000010110111101;
assign LUT_1[41727] = 32'b00000000000000000001101000111001;
assign LUT_1[41728] = 32'b11111111111111111011100001100000;
assign LUT_1[41729] = 32'b11111111111111110100110011011100;
assign LUT_1[41730] = 32'b11111111111111110111001111110001;
assign LUT_1[41731] = 32'b11111111111111110000100001101101;
assign LUT_1[41732] = 32'b00000000000000000011011010110111;
assign LUT_1[41733] = 32'b11111111111111111100101100110011;
assign LUT_1[41734] = 32'b11111111111111111111001001001000;
assign LUT_1[41735] = 32'b11111111111111111000011011000100;
assign LUT_1[41736] = 32'b11111111111111111010101111010101;
assign LUT_1[41737] = 32'b11111111111111110100000001010001;
assign LUT_1[41738] = 32'b11111111111111110110011101100110;
assign LUT_1[41739] = 32'b11111111111111101111101111100010;
assign LUT_1[41740] = 32'b00000000000000000010101000101100;
assign LUT_1[41741] = 32'b11111111111111111011111010101000;
assign LUT_1[41742] = 32'b11111111111111111110010110111101;
assign LUT_1[41743] = 32'b11111111111111110111101000111001;
assign LUT_1[41744] = 32'b11111111111111111101011101000010;
assign LUT_1[41745] = 32'b11111111111111110110101110111110;
assign LUT_1[41746] = 32'b11111111111111111001001011010011;
assign LUT_1[41747] = 32'b11111111111111110010011101001111;
assign LUT_1[41748] = 32'b00000000000000000101010110011001;
assign LUT_1[41749] = 32'b11111111111111111110101000010101;
assign LUT_1[41750] = 32'b00000000000000000001000100101010;
assign LUT_1[41751] = 32'b11111111111111111010010110100110;
assign LUT_1[41752] = 32'b11111111111111111100101010110111;
assign LUT_1[41753] = 32'b11111111111111110101111100110011;
assign LUT_1[41754] = 32'b11111111111111111000011001001000;
assign LUT_1[41755] = 32'b11111111111111110001101011000100;
assign LUT_1[41756] = 32'b00000000000000000100100100001110;
assign LUT_1[41757] = 32'b11111111111111111101110110001010;
assign LUT_1[41758] = 32'b00000000000000000000010010011111;
assign LUT_1[41759] = 32'b11111111111111111001100100011011;
assign LUT_1[41760] = 32'b11111111111111111100011100011111;
assign LUT_1[41761] = 32'b11111111111111110101101110011011;
assign LUT_1[41762] = 32'b11111111111111111000001010110000;
assign LUT_1[41763] = 32'b11111111111111110001011100101100;
assign LUT_1[41764] = 32'b00000000000000000100010101110110;
assign LUT_1[41765] = 32'b11111111111111111101100111110010;
assign LUT_1[41766] = 32'b00000000000000000000000100000111;
assign LUT_1[41767] = 32'b11111111111111111001010110000011;
assign LUT_1[41768] = 32'b11111111111111111011101010010100;
assign LUT_1[41769] = 32'b11111111111111110100111100010000;
assign LUT_1[41770] = 32'b11111111111111110111011000100101;
assign LUT_1[41771] = 32'b11111111111111110000101010100001;
assign LUT_1[41772] = 32'b00000000000000000011100011101011;
assign LUT_1[41773] = 32'b11111111111111111100110101100111;
assign LUT_1[41774] = 32'b11111111111111111111010001111100;
assign LUT_1[41775] = 32'b11111111111111111000100011111000;
assign LUT_1[41776] = 32'b11111111111111111110011000000001;
assign LUT_1[41777] = 32'b11111111111111110111101001111101;
assign LUT_1[41778] = 32'b11111111111111111010000110010010;
assign LUT_1[41779] = 32'b11111111111111110011011000001110;
assign LUT_1[41780] = 32'b00000000000000000110010001011000;
assign LUT_1[41781] = 32'b11111111111111111111100011010100;
assign LUT_1[41782] = 32'b00000000000000000001111111101001;
assign LUT_1[41783] = 32'b11111111111111111011010001100101;
assign LUT_1[41784] = 32'b11111111111111111101100101110110;
assign LUT_1[41785] = 32'b11111111111111110110110111110010;
assign LUT_1[41786] = 32'b11111111111111111001010100000111;
assign LUT_1[41787] = 32'b11111111111111110010100110000011;
assign LUT_1[41788] = 32'b00000000000000000101011111001101;
assign LUT_1[41789] = 32'b11111111111111111110110001001001;
assign LUT_1[41790] = 32'b00000000000000000001001101011110;
assign LUT_1[41791] = 32'b11111111111111111010011111011010;
assign LUT_1[41792] = 32'b11111111111111111101011111001000;
assign LUT_1[41793] = 32'b11111111111111110110110001000100;
assign LUT_1[41794] = 32'b11111111111111111001001101011001;
assign LUT_1[41795] = 32'b11111111111111110010011111010101;
assign LUT_1[41796] = 32'b00000000000000000101011000011111;
assign LUT_1[41797] = 32'b11111111111111111110101010011011;
assign LUT_1[41798] = 32'b00000000000000000001000110110000;
assign LUT_1[41799] = 32'b11111111111111111010011000101100;
assign LUT_1[41800] = 32'b11111111111111111100101100111101;
assign LUT_1[41801] = 32'b11111111111111110101111110111001;
assign LUT_1[41802] = 32'b11111111111111111000011011001110;
assign LUT_1[41803] = 32'b11111111111111110001101101001010;
assign LUT_1[41804] = 32'b00000000000000000100100110010100;
assign LUT_1[41805] = 32'b11111111111111111101111000010000;
assign LUT_1[41806] = 32'b00000000000000000000010100100101;
assign LUT_1[41807] = 32'b11111111111111111001100110100001;
assign LUT_1[41808] = 32'b11111111111111111111011010101010;
assign LUT_1[41809] = 32'b11111111111111111000101100100110;
assign LUT_1[41810] = 32'b11111111111111111011001000111011;
assign LUT_1[41811] = 32'b11111111111111110100011010110111;
assign LUT_1[41812] = 32'b00000000000000000111010100000001;
assign LUT_1[41813] = 32'b00000000000000000000100101111101;
assign LUT_1[41814] = 32'b00000000000000000011000010010010;
assign LUT_1[41815] = 32'b11111111111111111100010100001110;
assign LUT_1[41816] = 32'b11111111111111111110101000011111;
assign LUT_1[41817] = 32'b11111111111111110111111010011011;
assign LUT_1[41818] = 32'b11111111111111111010010110110000;
assign LUT_1[41819] = 32'b11111111111111110011101000101100;
assign LUT_1[41820] = 32'b00000000000000000110100001110110;
assign LUT_1[41821] = 32'b11111111111111111111110011110010;
assign LUT_1[41822] = 32'b00000000000000000010010000000111;
assign LUT_1[41823] = 32'b11111111111111111011100010000011;
assign LUT_1[41824] = 32'b11111111111111111110011010000111;
assign LUT_1[41825] = 32'b11111111111111110111101100000011;
assign LUT_1[41826] = 32'b11111111111111111010001000011000;
assign LUT_1[41827] = 32'b11111111111111110011011010010100;
assign LUT_1[41828] = 32'b00000000000000000110010011011110;
assign LUT_1[41829] = 32'b11111111111111111111100101011010;
assign LUT_1[41830] = 32'b00000000000000000010000001101111;
assign LUT_1[41831] = 32'b11111111111111111011010011101011;
assign LUT_1[41832] = 32'b11111111111111111101100111111100;
assign LUT_1[41833] = 32'b11111111111111110110111001111000;
assign LUT_1[41834] = 32'b11111111111111111001010110001101;
assign LUT_1[41835] = 32'b11111111111111110010101000001001;
assign LUT_1[41836] = 32'b00000000000000000101100001010011;
assign LUT_1[41837] = 32'b11111111111111111110110011001111;
assign LUT_1[41838] = 32'b00000000000000000001001111100100;
assign LUT_1[41839] = 32'b11111111111111111010100001100000;
assign LUT_1[41840] = 32'b00000000000000000000010101101001;
assign LUT_1[41841] = 32'b11111111111111111001100111100101;
assign LUT_1[41842] = 32'b11111111111111111100000011111010;
assign LUT_1[41843] = 32'b11111111111111110101010101110110;
assign LUT_1[41844] = 32'b00000000000000001000001111000000;
assign LUT_1[41845] = 32'b00000000000000000001100000111100;
assign LUT_1[41846] = 32'b00000000000000000011111101010001;
assign LUT_1[41847] = 32'b11111111111111111101001111001101;
assign LUT_1[41848] = 32'b11111111111111111111100011011110;
assign LUT_1[41849] = 32'b11111111111111111000110101011010;
assign LUT_1[41850] = 32'b11111111111111111011010001101111;
assign LUT_1[41851] = 32'b11111111111111110100100011101011;
assign LUT_1[41852] = 32'b00000000000000000111011100110101;
assign LUT_1[41853] = 32'b00000000000000000000101110110001;
assign LUT_1[41854] = 32'b00000000000000000011001011000110;
assign LUT_1[41855] = 32'b11111111111111111100011101000010;
assign LUT_1[41856] = 32'b11111111111111111110100001100011;
assign LUT_1[41857] = 32'b11111111111111110111110011011111;
assign LUT_1[41858] = 32'b11111111111111111010001111110100;
assign LUT_1[41859] = 32'b11111111111111110011100001110000;
assign LUT_1[41860] = 32'b00000000000000000110011010111010;
assign LUT_1[41861] = 32'b11111111111111111111101100110110;
assign LUT_1[41862] = 32'b00000000000000000010001001001011;
assign LUT_1[41863] = 32'b11111111111111111011011011000111;
assign LUT_1[41864] = 32'b11111111111111111101101111011000;
assign LUT_1[41865] = 32'b11111111111111110111000001010100;
assign LUT_1[41866] = 32'b11111111111111111001011101101001;
assign LUT_1[41867] = 32'b11111111111111110010101111100101;
assign LUT_1[41868] = 32'b00000000000000000101101000101111;
assign LUT_1[41869] = 32'b11111111111111111110111010101011;
assign LUT_1[41870] = 32'b00000000000000000001010111000000;
assign LUT_1[41871] = 32'b11111111111111111010101000111100;
assign LUT_1[41872] = 32'b00000000000000000000011101000101;
assign LUT_1[41873] = 32'b11111111111111111001101111000001;
assign LUT_1[41874] = 32'b11111111111111111100001011010110;
assign LUT_1[41875] = 32'b11111111111111110101011101010010;
assign LUT_1[41876] = 32'b00000000000000001000010110011100;
assign LUT_1[41877] = 32'b00000000000000000001101000011000;
assign LUT_1[41878] = 32'b00000000000000000100000100101101;
assign LUT_1[41879] = 32'b11111111111111111101010110101001;
assign LUT_1[41880] = 32'b11111111111111111111101010111010;
assign LUT_1[41881] = 32'b11111111111111111000111100110110;
assign LUT_1[41882] = 32'b11111111111111111011011001001011;
assign LUT_1[41883] = 32'b11111111111111110100101011000111;
assign LUT_1[41884] = 32'b00000000000000000111100100010001;
assign LUT_1[41885] = 32'b00000000000000000000110110001101;
assign LUT_1[41886] = 32'b00000000000000000011010010100010;
assign LUT_1[41887] = 32'b11111111111111111100100100011110;
assign LUT_1[41888] = 32'b11111111111111111111011100100010;
assign LUT_1[41889] = 32'b11111111111111111000101110011110;
assign LUT_1[41890] = 32'b11111111111111111011001010110011;
assign LUT_1[41891] = 32'b11111111111111110100011100101111;
assign LUT_1[41892] = 32'b00000000000000000111010101111001;
assign LUT_1[41893] = 32'b00000000000000000000100111110101;
assign LUT_1[41894] = 32'b00000000000000000011000100001010;
assign LUT_1[41895] = 32'b11111111111111111100010110000110;
assign LUT_1[41896] = 32'b11111111111111111110101010010111;
assign LUT_1[41897] = 32'b11111111111111110111111100010011;
assign LUT_1[41898] = 32'b11111111111111111010011000101000;
assign LUT_1[41899] = 32'b11111111111111110011101010100100;
assign LUT_1[41900] = 32'b00000000000000000110100011101110;
assign LUT_1[41901] = 32'b11111111111111111111110101101010;
assign LUT_1[41902] = 32'b00000000000000000010010001111111;
assign LUT_1[41903] = 32'b11111111111111111011100011111011;
assign LUT_1[41904] = 32'b00000000000000000001011000000100;
assign LUT_1[41905] = 32'b11111111111111111010101010000000;
assign LUT_1[41906] = 32'b11111111111111111101000110010101;
assign LUT_1[41907] = 32'b11111111111111110110011000010001;
assign LUT_1[41908] = 32'b00000000000000001001010001011011;
assign LUT_1[41909] = 32'b00000000000000000010100011010111;
assign LUT_1[41910] = 32'b00000000000000000100111111101100;
assign LUT_1[41911] = 32'b11111111111111111110010001101000;
assign LUT_1[41912] = 32'b00000000000000000000100101111001;
assign LUT_1[41913] = 32'b11111111111111111001110111110101;
assign LUT_1[41914] = 32'b11111111111111111100010100001010;
assign LUT_1[41915] = 32'b11111111111111110101100110000110;
assign LUT_1[41916] = 32'b00000000000000001000011111010000;
assign LUT_1[41917] = 32'b00000000000000000001110001001100;
assign LUT_1[41918] = 32'b00000000000000000100001101100001;
assign LUT_1[41919] = 32'b11111111111111111101011111011101;
assign LUT_1[41920] = 32'b00000000000000000000011111001011;
assign LUT_1[41921] = 32'b11111111111111111001110001000111;
assign LUT_1[41922] = 32'b11111111111111111100001101011100;
assign LUT_1[41923] = 32'b11111111111111110101011111011000;
assign LUT_1[41924] = 32'b00000000000000001000011000100010;
assign LUT_1[41925] = 32'b00000000000000000001101010011110;
assign LUT_1[41926] = 32'b00000000000000000100000110110011;
assign LUT_1[41927] = 32'b11111111111111111101011000101111;
assign LUT_1[41928] = 32'b11111111111111111111101101000000;
assign LUT_1[41929] = 32'b11111111111111111000111110111100;
assign LUT_1[41930] = 32'b11111111111111111011011011010001;
assign LUT_1[41931] = 32'b11111111111111110100101101001101;
assign LUT_1[41932] = 32'b00000000000000000111100110010111;
assign LUT_1[41933] = 32'b00000000000000000000111000010011;
assign LUT_1[41934] = 32'b00000000000000000011010100101000;
assign LUT_1[41935] = 32'b11111111111111111100100110100100;
assign LUT_1[41936] = 32'b00000000000000000010011010101101;
assign LUT_1[41937] = 32'b11111111111111111011101100101001;
assign LUT_1[41938] = 32'b11111111111111111110001000111110;
assign LUT_1[41939] = 32'b11111111111111110111011010111010;
assign LUT_1[41940] = 32'b00000000000000001010010100000100;
assign LUT_1[41941] = 32'b00000000000000000011100110000000;
assign LUT_1[41942] = 32'b00000000000000000110000010010101;
assign LUT_1[41943] = 32'b11111111111111111111010100010001;
assign LUT_1[41944] = 32'b00000000000000000001101000100010;
assign LUT_1[41945] = 32'b11111111111111111010111010011110;
assign LUT_1[41946] = 32'b11111111111111111101010110110011;
assign LUT_1[41947] = 32'b11111111111111110110101000101111;
assign LUT_1[41948] = 32'b00000000000000001001100001111001;
assign LUT_1[41949] = 32'b00000000000000000010110011110101;
assign LUT_1[41950] = 32'b00000000000000000101010000001010;
assign LUT_1[41951] = 32'b11111111111111111110100010000110;
assign LUT_1[41952] = 32'b00000000000000000001011010001010;
assign LUT_1[41953] = 32'b11111111111111111010101100000110;
assign LUT_1[41954] = 32'b11111111111111111101001000011011;
assign LUT_1[41955] = 32'b11111111111111110110011010010111;
assign LUT_1[41956] = 32'b00000000000000001001010011100001;
assign LUT_1[41957] = 32'b00000000000000000010100101011101;
assign LUT_1[41958] = 32'b00000000000000000101000001110010;
assign LUT_1[41959] = 32'b11111111111111111110010011101110;
assign LUT_1[41960] = 32'b00000000000000000000100111111111;
assign LUT_1[41961] = 32'b11111111111111111001111001111011;
assign LUT_1[41962] = 32'b11111111111111111100010110010000;
assign LUT_1[41963] = 32'b11111111111111110101101000001100;
assign LUT_1[41964] = 32'b00000000000000001000100001010110;
assign LUT_1[41965] = 32'b00000000000000000001110011010010;
assign LUT_1[41966] = 32'b00000000000000000100001111100111;
assign LUT_1[41967] = 32'b11111111111111111101100001100011;
assign LUT_1[41968] = 32'b00000000000000000011010101101100;
assign LUT_1[41969] = 32'b11111111111111111100100111101000;
assign LUT_1[41970] = 32'b11111111111111111111000011111101;
assign LUT_1[41971] = 32'b11111111111111111000010101111001;
assign LUT_1[41972] = 32'b00000000000000001011001111000011;
assign LUT_1[41973] = 32'b00000000000000000100100000111111;
assign LUT_1[41974] = 32'b00000000000000000110111101010100;
assign LUT_1[41975] = 32'b00000000000000000000001111010000;
assign LUT_1[41976] = 32'b00000000000000000010100011100001;
assign LUT_1[41977] = 32'b11111111111111111011110101011101;
assign LUT_1[41978] = 32'b11111111111111111110010001110010;
assign LUT_1[41979] = 32'b11111111111111110111100011101110;
assign LUT_1[41980] = 32'b00000000000000001010011100111000;
assign LUT_1[41981] = 32'b00000000000000000011101110110100;
assign LUT_1[41982] = 32'b00000000000000000110001011001001;
assign LUT_1[41983] = 32'b11111111111111111111011101000101;
assign LUT_1[41984] = 32'b00000000000000001010010101100111;
assign LUT_1[41985] = 32'b00000000000000000011100111100011;
assign LUT_1[41986] = 32'b00000000000000000110000011111000;
assign LUT_1[41987] = 32'b11111111111111111111010101110100;
assign LUT_1[41988] = 32'b00000000000000010010001110111110;
assign LUT_1[41989] = 32'b00000000000000001011100000111010;
assign LUT_1[41990] = 32'b00000000000000001101111101001111;
assign LUT_1[41991] = 32'b00000000000000000111001111001011;
assign LUT_1[41992] = 32'b00000000000000001001100011011100;
assign LUT_1[41993] = 32'b00000000000000000010110101011000;
assign LUT_1[41994] = 32'b00000000000000000101010001101101;
assign LUT_1[41995] = 32'b11111111111111111110100011101001;
assign LUT_1[41996] = 32'b00000000000000010001011100110011;
assign LUT_1[41997] = 32'b00000000000000001010101110101111;
assign LUT_1[41998] = 32'b00000000000000001101001011000100;
assign LUT_1[41999] = 32'b00000000000000000110011101000000;
assign LUT_1[42000] = 32'b00000000000000001100010001001001;
assign LUT_1[42001] = 32'b00000000000000000101100011000101;
assign LUT_1[42002] = 32'b00000000000000000111111111011010;
assign LUT_1[42003] = 32'b00000000000000000001010001010110;
assign LUT_1[42004] = 32'b00000000000000010100001010100000;
assign LUT_1[42005] = 32'b00000000000000001101011100011100;
assign LUT_1[42006] = 32'b00000000000000001111111000110001;
assign LUT_1[42007] = 32'b00000000000000001001001010101101;
assign LUT_1[42008] = 32'b00000000000000001011011110111110;
assign LUT_1[42009] = 32'b00000000000000000100110000111010;
assign LUT_1[42010] = 32'b00000000000000000111001101001111;
assign LUT_1[42011] = 32'b00000000000000000000011111001011;
assign LUT_1[42012] = 32'b00000000000000010011011000010101;
assign LUT_1[42013] = 32'b00000000000000001100101010010001;
assign LUT_1[42014] = 32'b00000000000000001111000110100110;
assign LUT_1[42015] = 32'b00000000000000001000011000100010;
assign LUT_1[42016] = 32'b00000000000000001011010000100110;
assign LUT_1[42017] = 32'b00000000000000000100100010100010;
assign LUT_1[42018] = 32'b00000000000000000110111110110111;
assign LUT_1[42019] = 32'b00000000000000000000010000110011;
assign LUT_1[42020] = 32'b00000000000000010011001001111101;
assign LUT_1[42021] = 32'b00000000000000001100011011111001;
assign LUT_1[42022] = 32'b00000000000000001110111000001110;
assign LUT_1[42023] = 32'b00000000000000001000001010001010;
assign LUT_1[42024] = 32'b00000000000000001010011110011011;
assign LUT_1[42025] = 32'b00000000000000000011110000010111;
assign LUT_1[42026] = 32'b00000000000000000110001100101100;
assign LUT_1[42027] = 32'b11111111111111111111011110101000;
assign LUT_1[42028] = 32'b00000000000000010010010111110010;
assign LUT_1[42029] = 32'b00000000000000001011101001101110;
assign LUT_1[42030] = 32'b00000000000000001110000110000011;
assign LUT_1[42031] = 32'b00000000000000000111010111111111;
assign LUT_1[42032] = 32'b00000000000000001101001100001000;
assign LUT_1[42033] = 32'b00000000000000000110011110000100;
assign LUT_1[42034] = 32'b00000000000000001000111010011001;
assign LUT_1[42035] = 32'b00000000000000000010001100010101;
assign LUT_1[42036] = 32'b00000000000000010101000101011111;
assign LUT_1[42037] = 32'b00000000000000001110010111011011;
assign LUT_1[42038] = 32'b00000000000000010000110011110000;
assign LUT_1[42039] = 32'b00000000000000001010000101101100;
assign LUT_1[42040] = 32'b00000000000000001100011001111101;
assign LUT_1[42041] = 32'b00000000000000000101101011111001;
assign LUT_1[42042] = 32'b00000000000000001000001000001110;
assign LUT_1[42043] = 32'b00000000000000000001011010001010;
assign LUT_1[42044] = 32'b00000000000000010100010011010100;
assign LUT_1[42045] = 32'b00000000000000001101100101010000;
assign LUT_1[42046] = 32'b00000000000000010000000001100101;
assign LUT_1[42047] = 32'b00000000000000001001010011100001;
assign LUT_1[42048] = 32'b00000000000000001100010011001111;
assign LUT_1[42049] = 32'b00000000000000000101100101001011;
assign LUT_1[42050] = 32'b00000000000000001000000001100000;
assign LUT_1[42051] = 32'b00000000000000000001010011011100;
assign LUT_1[42052] = 32'b00000000000000010100001100100110;
assign LUT_1[42053] = 32'b00000000000000001101011110100010;
assign LUT_1[42054] = 32'b00000000000000001111111010110111;
assign LUT_1[42055] = 32'b00000000000000001001001100110011;
assign LUT_1[42056] = 32'b00000000000000001011100001000100;
assign LUT_1[42057] = 32'b00000000000000000100110011000000;
assign LUT_1[42058] = 32'b00000000000000000111001111010101;
assign LUT_1[42059] = 32'b00000000000000000000100001010001;
assign LUT_1[42060] = 32'b00000000000000010011011010011011;
assign LUT_1[42061] = 32'b00000000000000001100101100010111;
assign LUT_1[42062] = 32'b00000000000000001111001000101100;
assign LUT_1[42063] = 32'b00000000000000001000011010101000;
assign LUT_1[42064] = 32'b00000000000000001110001110110001;
assign LUT_1[42065] = 32'b00000000000000000111100000101101;
assign LUT_1[42066] = 32'b00000000000000001001111101000010;
assign LUT_1[42067] = 32'b00000000000000000011001110111110;
assign LUT_1[42068] = 32'b00000000000000010110001000001000;
assign LUT_1[42069] = 32'b00000000000000001111011010000100;
assign LUT_1[42070] = 32'b00000000000000010001110110011001;
assign LUT_1[42071] = 32'b00000000000000001011001000010101;
assign LUT_1[42072] = 32'b00000000000000001101011100100110;
assign LUT_1[42073] = 32'b00000000000000000110101110100010;
assign LUT_1[42074] = 32'b00000000000000001001001010110111;
assign LUT_1[42075] = 32'b00000000000000000010011100110011;
assign LUT_1[42076] = 32'b00000000000000010101010101111101;
assign LUT_1[42077] = 32'b00000000000000001110100111111001;
assign LUT_1[42078] = 32'b00000000000000010001000100001110;
assign LUT_1[42079] = 32'b00000000000000001010010110001010;
assign LUT_1[42080] = 32'b00000000000000001101001110001110;
assign LUT_1[42081] = 32'b00000000000000000110100000001010;
assign LUT_1[42082] = 32'b00000000000000001000111100011111;
assign LUT_1[42083] = 32'b00000000000000000010001110011011;
assign LUT_1[42084] = 32'b00000000000000010101000111100101;
assign LUT_1[42085] = 32'b00000000000000001110011001100001;
assign LUT_1[42086] = 32'b00000000000000010000110101110110;
assign LUT_1[42087] = 32'b00000000000000001010000111110010;
assign LUT_1[42088] = 32'b00000000000000001100011100000011;
assign LUT_1[42089] = 32'b00000000000000000101101101111111;
assign LUT_1[42090] = 32'b00000000000000001000001010010100;
assign LUT_1[42091] = 32'b00000000000000000001011100010000;
assign LUT_1[42092] = 32'b00000000000000010100010101011010;
assign LUT_1[42093] = 32'b00000000000000001101100111010110;
assign LUT_1[42094] = 32'b00000000000000010000000011101011;
assign LUT_1[42095] = 32'b00000000000000001001010101100111;
assign LUT_1[42096] = 32'b00000000000000001111001001110000;
assign LUT_1[42097] = 32'b00000000000000001000011011101100;
assign LUT_1[42098] = 32'b00000000000000001010111000000001;
assign LUT_1[42099] = 32'b00000000000000000100001001111101;
assign LUT_1[42100] = 32'b00000000000000010111000011000111;
assign LUT_1[42101] = 32'b00000000000000010000010101000011;
assign LUT_1[42102] = 32'b00000000000000010010110001011000;
assign LUT_1[42103] = 32'b00000000000000001100000011010100;
assign LUT_1[42104] = 32'b00000000000000001110010111100101;
assign LUT_1[42105] = 32'b00000000000000000111101001100001;
assign LUT_1[42106] = 32'b00000000000000001010000101110110;
assign LUT_1[42107] = 32'b00000000000000000011010111110010;
assign LUT_1[42108] = 32'b00000000000000010110010000111100;
assign LUT_1[42109] = 32'b00000000000000001111100010111000;
assign LUT_1[42110] = 32'b00000000000000010001111111001101;
assign LUT_1[42111] = 32'b00000000000000001011010001001001;
assign LUT_1[42112] = 32'b00000000000000001101010101101010;
assign LUT_1[42113] = 32'b00000000000000000110100111100110;
assign LUT_1[42114] = 32'b00000000000000001001000011111011;
assign LUT_1[42115] = 32'b00000000000000000010010101110111;
assign LUT_1[42116] = 32'b00000000000000010101001111000001;
assign LUT_1[42117] = 32'b00000000000000001110100000111101;
assign LUT_1[42118] = 32'b00000000000000010000111101010010;
assign LUT_1[42119] = 32'b00000000000000001010001111001110;
assign LUT_1[42120] = 32'b00000000000000001100100011011111;
assign LUT_1[42121] = 32'b00000000000000000101110101011011;
assign LUT_1[42122] = 32'b00000000000000001000010001110000;
assign LUT_1[42123] = 32'b00000000000000000001100011101100;
assign LUT_1[42124] = 32'b00000000000000010100011100110110;
assign LUT_1[42125] = 32'b00000000000000001101101110110010;
assign LUT_1[42126] = 32'b00000000000000010000001011000111;
assign LUT_1[42127] = 32'b00000000000000001001011101000011;
assign LUT_1[42128] = 32'b00000000000000001111010001001100;
assign LUT_1[42129] = 32'b00000000000000001000100011001000;
assign LUT_1[42130] = 32'b00000000000000001010111111011101;
assign LUT_1[42131] = 32'b00000000000000000100010001011001;
assign LUT_1[42132] = 32'b00000000000000010111001010100011;
assign LUT_1[42133] = 32'b00000000000000010000011100011111;
assign LUT_1[42134] = 32'b00000000000000010010111000110100;
assign LUT_1[42135] = 32'b00000000000000001100001010110000;
assign LUT_1[42136] = 32'b00000000000000001110011111000001;
assign LUT_1[42137] = 32'b00000000000000000111110000111101;
assign LUT_1[42138] = 32'b00000000000000001010001101010010;
assign LUT_1[42139] = 32'b00000000000000000011011111001110;
assign LUT_1[42140] = 32'b00000000000000010110011000011000;
assign LUT_1[42141] = 32'b00000000000000001111101010010100;
assign LUT_1[42142] = 32'b00000000000000010010000110101001;
assign LUT_1[42143] = 32'b00000000000000001011011000100101;
assign LUT_1[42144] = 32'b00000000000000001110010000101001;
assign LUT_1[42145] = 32'b00000000000000000111100010100101;
assign LUT_1[42146] = 32'b00000000000000001001111110111010;
assign LUT_1[42147] = 32'b00000000000000000011010000110110;
assign LUT_1[42148] = 32'b00000000000000010110001010000000;
assign LUT_1[42149] = 32'b00000000000000001111011011111100;
assign LUT_1[42150] = 32'b00000000000000010001111000010001;
assign LUT_1[42151] = 32'b00000000000000001011001010001101;
assign LUT_1[42152] = 32'b00000000000000001101011110011110;
assign LUT_1[42153] = 32'b00000000000000000110110000011010;
assign LUT_1[42154] = 32'b00000000000000001001001100101111;
assign LUT_1[42155] = 32'b00000000000000000010011110101011;
assign LUT_1[42156] = 32'b00000000000000010101010111110101;
assign LUT_1[42157] = 32'b00000000000000001110101001110001;
assign LUT_1[42158] = 32'b00000000000000010001000110000110;
assign LUT_1[42159] = 32'b00000000000000001010011000000010;
assign LUT_1[42160] = 32'b00000000000000010000001100001011;
assign LUT_1[42161] = 32'b00000000000000001001011110000111;
assign LUT_1[42162] = 32'b00000000000000001011111010011100;
assign LUT_1[42163] = 32'b00000000000000000101001100011000;
assign LUT_1[42164] = 32'b00000000000000011000000101100010;
assign LUT_1[42165] = 32'b00000000000000010001010111011110;
assign LUT_1[42166] = 32'b00000000000000010011110011110011;
assign LUT_1[42167] = 32'b00000000000000001101000101101111;
assign LUT_1[42168] = 32'b00000000000000001111011010000000;
assign LUT_1[42169] = 32'b00000000000000001000101011111100;
assign LUT_1[42170] = 32'b00000000000000001011001000010001;
assign LUT_1[42171] = 32'b00000000000000000100011010001101;
assign LUT_1[42172] = 32'b00000000000000010111010011010111;
assign LUT_1[42173] = 32'b00000000000000010000100101010011;
assign LUT_1[42174] = 32'b00000000000000010011000001101000;
assign LUT_1[42175] = 32'b00000000000000001100010011100100;
assign LUT_1[42176] = 32'b00000000000000001111010011010010;
assign LUT_1[42177] = 32'b00000000000000001000100101001110;
assign LUT_1[42178] = 32'b00000000000000001011000001100011;
assign LUT_1[42179] = 32'b00000000000000000100010011011111;
assign LUT_1[42180] = 32'b00000000000000010111001100101001;
assign LUT_1[42181] = 32'b00000000000000010000011110100101;
assign LUT_1[42182] = 32'b00000000000000010010111010111010;
assign LUT_1[42183] = 32'b00000000000000001100001100110110;
assign LUT_1[42184] = 32'b00000000000000001110100001000111;
assign LUT_1[42185] = 32'b00000000000000000111110011000011;
assign LUT_1[42186] = 32'b00000000000000001010001111011000;
assign LUT_1[42187] = 32'b00000000000000000011100001010100;
assign LUT_1[42188] = 32'b00000000000000010110011010011110;
assign LUT_1[42189] = 32'b00000000000000001111101100011010;
assign LUT_1[42190] = 32'b00000000000000010010001000101111;
assign LUT_1[42191] = 32'b00000000000000001011011010101011;
assign LUT_1[42192] = 32'b00000000000000010001001110110100;
assign LUT_1[42193] = 32'b00000000000000001010100000110000;
assign LUT_1[42194] = 32'b00000000000000001100111101000101;
assign LUT_1[42195] = 32'b00000000000000000110001111000001;
assign LUT_1[42196] = 32'b00000000000000011001001000001011;
assign LUT_1[42197] = 32'b00000000000000010010011010000111;
assign LUT_1[42198] = 32'b00000000000000010100110110011100;
assign LUT_1[42199] = 32'b00000000000000001110001000011000;
assign LUT_1[42200] = 32'b00000000000000010000011100101001;
assign LUT_1[42201] = 32'b00000000000000001001101110100101;
assign LUT_1[42202] = 32'b00000000000000001100001010111010;
assign LUT_1[42203] = 32'b00000000000000000101011100110110;
assign LUT_1[42204] = 32'b00000000000000011000010110000000;
assign LUT_1[42205] = 32'b00000000000000010001100111111100;
assign LUT_1[42206] = 32'b00000000000000010100000100010001;
assign LUT_1[42207] = 32'b00000000000000001101010110001101;
assign LUT_1[42208] = 32'b00000000000000010000001110010001;
assign LUT_1[42209] = 32'b00000000000000001001100000001101;
assign LUT_1[42210] = 32'b00000000000000001011111100100010;
assign LUT_1[42211] = 32'b00000000000000000101001110011110;
assign LUT_1[42212] = 32'b00000000000000011000000111101000;
assign LUT_1[42213] = 32'b00000000000000010001011001100100;
assign LUT_1[42214] = 32'b00000000000000010011110101111001;
assign LUT_1[42215] = 32'b00000000000000001101000111110101;
assign LUT_1[42216] = 32'b00000000000000001111011100000110;
assign LUT_1[42217] = 32'b00000000000000001000101110000010;
assign LUT_1[42218] = 32'b00000000000000001011001010010111;
assign LUT_1[42219] = 32'b00000000000000000100011100010011;
assign LUT_1[42220] = 32'b00000000000000010111010101011101;
assign LUT_1[42221] = 32'b00000000000000010000100111011001;
assign LUT_1[42222] = 32'b00000000000000010011000011101110;
assign LUT_1[42223] = 32'b00000000000000001100010101101010;
assign LUT_1[42224] = 32'b00000000000000010010001001110011;
assign LUT_1[42225] = 32'b00000000000000001011011011101111;
assign LUT_1[42226] = 32'b00000000000000001101111000000100;
assign LUT_1[42227] = 32'b00000000000000000111001010000000;
assign LUT_1[42228] = 32'b00000000000000011010000011001010;
assign LUT_1[42229] = 32'b00000000000000010011010101000110;
assign LUT_1[42230] = 32'b00000000000000010101110001011011;
assign LUT_1[42231] = 32'b00000000000000001111000011010111;
assign LUT_1[42232] = 32'b00000000000000010001010111101000;
assign LUT_1[42233] = 32'b00000000000000001010101001100100;
assign LUT_1[42234] = 32'b00000000000000001101000101111001;
assign LUT_1[42235] = 32'b00000000000000000110010111110101;
assign LUT_1[42236] = 32'b00000000000000011001010000111111;
assign LUT_1[42237] = 32'b00000000000000010010100010111011;
assign LUT_1[42238] = 32'b00000000000000010100111111010000;
assign LUT_1[42239] = 32'b00000000000000001110010001001100;
assign LUT_1[42240] = 32'b00000000000000001000001001110011;
assign LUT_1[42241] = 32'b00000000000000000001011011101111;
assign LUT_1[42242] = 32'b00000000000000000011111000000100;
assign LUT_1[42243] = 32'b11111111111111111101001010000000;
assign LUT_1[42244] = 32'b00000000000000010000000011001010;
assign LUT_1[42245] = 32'b00000000000000001001010101000110;
assign LUT_1[42246] = 32'b00000000000000001011110001011011;
assign LUT_1[42247] = 32'b00000000000000000101000011010111;
assign LUT_1[42248] = 32'b00000000000000000111010111101000;
assign LUT_1[42249] = 32'b00000000000000000000101001100100;
assign LUT_1[42250] = 32'b00000000000000000011000101111001;
assign LUT_1[42251] = 32'b11111111111111111100010111110101;
assign LUT_1[42252] = 32'b00000000000000001111010000111111;
assign LUT_1[42253] = 32'b00000000000000001000100010111011;
assign LUT_1[42254] = 32'b00000000000000001010111111010000;
assign LUT_1[42255] = 32'b00000000000000000100010001001100;
assign LUT_1[42256] = 32'b00000000000000001010000101010101;
assign LUT_1[42257] = 32'b00000000000000000011010111010001;
assign LUT_1[42258] = 32'b00000000000000000101110011100110;
assign LUT_1[42259] = 32'b11111111111111111111000101100010;
assign LUT_1[42260] = 32'b00000000000000010001111110101100;
assign LUT_1[42261] = 32'b00000000000000001011010000101000;
assign LUT_1[42262] = 32'b00000000000000001101101100111101;
assign LUT_1[42263] = 32'b00000000000000000110111110111001;
assign LUT_1[42264] = 32'b00000000000000001001010011001010;
assign LUT_1[42265] = 32'b00000000000000000010100101000110;
assign LUT_1[42266] = 32'b00000000000000000101000001011011;
assign LUT_1[42267] = 32'b11111111111111111110010011010111;
assign LUT_1[42268] = 32'b00000000000000010001001100100001;
assign LUT_1[42269] = 32'b00000000000000001010011110011101;
assign LUT_1[42270] = 32'b00000000000000001100111010110010;
assign LUT_1[42271] = 32'b00000000000000000110001100101110;
assign LUT_1[42272] = 32'b00000000000000001001000100110010;
assign LUT_1[42273] = 32'b00000000000000000010010110101110;
assign LUT_1[42274] = 32'b00000000000000000100110011000011;
assign LUT_1[42275] = 32'b11111111111111111110000100111111;
assign LUT_1[42276] = 32'b00000000000000010000111110001001;
assign LUT_1[42277] = 32'b00000000000000001010010000000101;
assign LUT_1[42278] = 32'b00000000000000001100101100011010;
assign LUT_1[42279] = 32'b00000000000000000101111110010110;
assign LUT_1[42280] = 32'b00000000000000001000010010100111;
assign LUT_1[42281] = 32'b00000000000000000001100100100011;
assign LUT_1[42282] = 32'b00000000000000000100000000111000;
assign LUT_1[42283] = 32'b11111111111111111101010010110100;
assign LUT_1[42284] = 32'b00000000000000010000001011111110;
assign LUT_1[42285] = 32'b00000000000000001001011101111010;
assign LUT_1[42286] = 32'b00000000000000001011111010001111;
assign LUT_1[42287] = 32'b00000000000000000101001100001011;
assign LUT_1[42288] = 32'b00000000000000001011000000010100;
assign LUT_1[42289] = 32'b00000000000000000100010010010000;
assign LUT_1[42290] = 32'b00000000000000000110101110100101;
assign LUT_1[42291] = 32'b00000000000000000000000000100001;
assign LUT_1[42292] = 32'b00000000000000010010111001101011;
assign LUT_1[42293] = 32'b00000000000000001100001011100111;
assign LUT_1[42294] = 32'b00000000000000001110100111111100;
assign LUT_1[42295] = 32'b00000000000000000111111001111000;
assign LUT_1[42296] = 32'b00000000000000001010001110001001;
assign LUT_1[42297] = 32'b00000000000000000011100000000101;
assign LUT_1[42298] = 32'b00000000000000000101111100011010;
assign LUT_1[42299] = 32'b11111111111111111111001110010110;
assign LUT_1[42300] = 32'b00000000000000010010000111100000;
assign LUT_1[42301] = 32'b00000000000000001011011001011100;
assign LUT_1[42302] = 32'b00000000000000001101110101110001;
assign LUT_1[42303] = 32'b00000000000000000111000111101101;
assign LUT_1[42304] = 32'b00000000000000001010000111011011;
assign LUT_1[42305] = 32'b00000000000000000011011001010111;
assign LUT_1[42306] = 32'b00000000000000000101110101101100;
assign LUT_1[42307] = 32'b11111111111111111111000111101000;
assign LUT_1[42308] = 32'b00000000000000010010000000110010;
assign LUT_1[42309] = 32'b00000000000000001011010010101110;
assign LUT_1[42310] = 32'b00000000000000001101101111000011;
assign LUT_1[42311] = 32'b00000000000000000111000000111111;
assign LUT_1[42312] = 32'b00000000000000001001010101010000;
assign LUT_1[42313] = 32'b00000000000000000010100111001100;
assign LUT_1[42314] = 32'b00000000000000000101000011100001;
assign LUT_1[42315] = 32'b11111111111111111110010101011101;
assign LUT_1[42316] = 32'b00000000000000010001001110100111;
assign LUT_1[42317] = 32'b00000000000000001010100000100011;
assign LUT_1[42318] = 32'b00000000000000001100111100111000;
assign LUT_1[42319] = 32'b00000000000000000110001110110100;
assign LUT_1[42320] = 32'b00000000000000001100000010111101;
assign LUT_1[42321] = 32'b00000000000000000101010100111001;
assign LUT_1[42322] = 32'b00000000000000000111110001001110;
assign LUT_1[42323] = 32'b00000000000000000001000011001010;
assign LUT_1[42324] = 32'b00000000000000010011111100010100;
assign LUT_1[42325] = 32'b00000000000000001101001110010000;
assign LUT_1[42326] = 32'b00000000000000001111101010100101;
assign LUT_1[42327] = 32'b00000000000000001000111100100001;
assign LUT_1[42328] = 32'b00000000000000001011010000110010;
assign LUT_1[42329] = 32'b00000000000000000100100010101110;
assign LUT_1[42330] = 32'b00000000000000000110111111000011;
assign LUT_1[42331] = 32'b00000000000000000000010000111111;
assign LUT_1[42332] = 32'b00000000000000010011001010001001;
assign LUT_1[42333] = 32'b00000000000000001100011100000101;
assign LUT_1[42334] = 32'b00000000000000001110111000011010;
assign LUT_1[42335] = 32'b00000000000000001000001010010110;
assign LUT_1[42336] = 32'b00000000000000001011000010011010;
assign LUT_1[42337] = 32'b00000000000000000100010100010110;
assign LUT_1[42338] = 32'b00000000000000000110110000101011;
assign LUT_1[42339] = 32'b00000000000000000000000010100111;
assign LUT_1[42340] = 32'b00000000000000010010111011110001;
assign LUT_1[42341] = 32'b00000000000000001100001101101101;
assign LUT_1[42342] = 32'b00000000000000001110101010000010;
assign LUT_1[42343] = 32'b00000000000000000111111011111110;
assign LUT_1[42344] = 32'b00000000000000001010010000001111;
assign LUT_1[42345] = 32'b00000000000000000011100010001011;
assign LUT_1[42346] = 32'b00000000000000000101111110100000;
assign LUT_1[42347] = 32'b11111111111111111111010000011100;
assign LUT_1[42348] = 32'b00000000000000010010001001100110;
assign LUT_1[42349] = 32'b00000000000000001011011011100010;
assign LUT_1[42350] = 32'b00000000000000001101110111110111;
assign LUT_1[42351] = 32'b00000000000000000111001001110011;
assign LUT_1[42352] = 32'b00000000000000001100111101111100;
assign LUT_1[42353] = 32'b00000000000000000110001111111000;
assign LUT_1[42354] = 32'b00000000000000001000101100001101;
assign LUT_1[42355] = 32'b00000000000000000001111110001001;
assign LUT_1[42356] = 32'b00000000000000010100110111010011;
assign LUT_1[42357] = 32'b00000000000000001110001001001111;
assign LUT_1[42358] = 32'b00000000000000010000100101100100;
assign LUT_1[42359] = 32'b00000000000000001001110111100000;
assign LUT_1[42360] = 32'b00000000000000001100001011110001;
assign LUT_1[42361] = 32'b00000000000000000101011101101101;
assign LUT_1[42362] = 32'b00000000000000000111111010000010;
assign LUT_1[42363] = 32'b00000000000000000001001011111110;
assign LUT_1[42364] = 32'b00000000000000010100000101001000;
assign LUT_1[42365] = 32'b00000000000000001101010111000100;
assign LUT_1[42366] = 32'b00000000000000001111110011011001;
assign LUT_1[42367] = 32'b00000000000000001001000101010101;
assign LUT_1[42368] = 32'b00000000000000001011001001110110;
assign LUT_1[42369] = 32'b00000000000000000100011011110010;
assign LUT_1[42370] = 32'b00000000000000000110111000000111;
assign LUT_1[42371] = 32'b00000000000000000000001010000011;
assign LUT_1[42372] = 32'b00000000000000010011000011001101;
assign LUT_1[42373] = 32'b00000000000000001100010101001001;
assign LUT_1[42374] = 32'b00000000000000001110110001011110;
assign LUT_1[42375] = 32'b00000000000000001000000011011010;
assign LUT_1[42376] = 32'b00000000000000001010010111101011;
assign LUT_1[42377] = 32'b00000000000000000011101001100111;
assign LUT_1[42378] = 32'b00000000000000000110000101111100;
assign LUT_1[42379] = 32'b11111111111111111111010111111000;
assign LUT_1[42380] = 32'b00000000000000010010010001000010;
assign LUT_1[42381] = 32'b00000000000000001011100010111110;
assign LUT_1[42382] = 32'b00000000000000001101111111010011;
assign LUT_1[42383] = 32'b00000000000000000111010001001111;
assign LUT_1[42384] = 32'b00000000000000001101000101011000;
assign LUT_1[42385] = 32'b00000000000000000110010111010100;
assign LUT_1[42386] = 32'b00000000000000001000110011101001;
assign LUT_1[42387] = 32'b00000000000000000010000101100101;
assign LUT_1[42388] = 32'b00000000000000010100111110101111;
assign LUT_1[42389] = 32'b00000000000000001110010000101011;
assign LUT_1[42390] = 32'b00000000000000010000101101000000;
assign LUT_1[42391] = 32'b00000000000000001001111110111100;
assign LUT_1[42392] = 32'b00000000000000001100010011001101;
assign LUT_1[42393] = 32'b00000000000000000101100101001001;
assign LUT_1[42394] = 32'b00000000000000001000000001011110;
assign LUT_1[42395] = 32'b00000000000000000001010011011010;
assign LUT_1[42396] = 32'b00000000000000010100001100100100;
assign LUT_1[42397] = 32'b00000000000000001101011110100000;
assign LUT_1[42398] = 32'b00000000000000001111111010110101;
assign LUT_1[42399] = 32'b00000000000000001001001100110001;
assign LUT_1[42400] = 32'b00000000000000001100000100110101;
assign LUT_1[42401] = 32'b00000000000000000101010110110001;
assign LUT_1[42402] = 32'b00000000000000000111110011000110;
assign LUT_1[42403] = 32'b00000000000000000001000101000010;
assign LUT_1[42404] = 32'b00000000000000010011111110001100;
assign LUT_1[42405] = 32'b00000000000000001101010000001000;
assign LUT_1[42406] = 32'b00000000000000001111101100011101;
assign LUT_1[42407] = 32'b00000000000000001000111110011001;
assign LUT_1[42408] = 32'b00000000000000001011010010101010;
assign LUT_1[42409] = 32'b00000000000000000100100100100110;
assign LUT_1[42410] = 32'b00000000000000000111000000111011;
assign LUT_1[42411] = 32'b00000000000000000000010010110111;
assign LUT_1[42412] = 32'b00000000000000010011001100000001;
assign LUT_1[42413] = 32'b00000000000000001100011101111101;
assign LUT_1[42414] = 32'b00000000000000001110111010010010;
assign LUT_1[42415] = 32'b00000000000000001000001100001110;
assign LUT_1[42416] = 32'b00000000000000001110000000010111;
assign LUT_1[42417] = 32'b00000000000000000111010010010011;
assign LUT_1[42418] = 32'b00000000000000001001101110101000;
assign LUT_1[42419] = 32'b00000000000000000011000000100100;
assign LUT_1[42420] = 32'b00000000000000010101111001101110;
assign LUT_1[42421] = 32'b00000000000000001111001011101010;
assign LUT_1[42422] = 32'b00000000000000010001100111111111;
assign LUT_1[42423] = 32'b00000000000000001010111001111011;
assign LUT_1[42424] = 32'b00000000000000001101001110001100;
assign LUT_1[42425] = 32'b00000000000000000110100000001000;
assign LUT_1[42426] = 32'b00000000000000001000111100011101;
assign LUT_1[42427] = 32'b00000000000000000010001110011001;
assign LUT_1[42428] = 32'b00000000000000010101000111100011;
assign LUT_1[42429] = 32'b00000000000000001110011001011111;
assign LUT_1[42430] = 32'b00000000000000010000110101110100;
assign LUT_1[42431] = 32'b00000000000000001010000111110000;
assign LUT_1[42432] = 32'b00000000000000001101000111011110;
assign LUT_1[42433] = 32'b00000000000000000110011001011010;
assign LUT_1[42434] = 32'b00000000000000001000110101101111;
assign LUT_1[42435] = 32'b00000000000000000010000111101011;
assign LUT_1[42436] = 32'b00000000000000010101000000110101;
assign LUT_1[42437] = 32'b00000000000000001110010010110001;
assign LUT_1[42438] = 32'b00000000000000010000101111000110;
assign LUT_1[42439] = 32'b00000000000000001010000001000010;
assign LUT_1[42440] = 32'b00000000000000001100010101010011;
assign LUT_1[42441] = 32'b00000000000000000101100111001111;
assign LUT_1[42442] = 32'b00000000000000001000000011100100;
assign LUT_1[42443] = 32'b00000000000000000001010101100000;
assign LUT_1[42444] = 32'b00000000000000010100001110101010;
assign LUT_1[42445] = 32'b00000000000000001101100000100110;
assign LUT_1[42446] = 32'b00000000000000001111111100111011;
assign LUT_1[42447] = 32'b00000000000000001001001110110111;
assign LUT_1[42448] = 32'b00000000000000001111000011000000;
assign LUT_1[42449] = 32'b00000000000000001000010100111100;
assign LUT_1[42450] = 32'b00000000000000001010110001010001;
assign LUT_1[42451] = 32'b00000000000000000100000011001101;
assign LUT_1[42452] = 32'b00000000000000010110111100010111;
assign LUT_1[42453] = 32'b00000000000000010000001110010011;
assign LUT_1[42454] = 32'b00000000000000010010101010101000;
assign LUT_1[42455] = 32'b00000000000000001011111100100100;
assign LUT_1[42456] = 32'b00000000000000001110010000110101;
assign LUT_1[42457] = 32'b00000000000000000111100010110001;
assign LUT_1[42458] = 32'b00000000000000001001111111000110;
assign LUT_1[42459] = 32'b00000000000000000011010001000010;
assign LUT_1[42460] = 32'b00000000000000010110001010001100;
assign LUT_1[42461] = 32'b00000000000000001111011100001000;
assign LUT_1[42462] = 32'b00000000000000010001111000011101;
assign LUT_1[42463] = 32'b00000000000000001011001010011001;
assign LUT_1[42464] = 32'b00000000000000001110000010011101;
assign LUT_1[42465] = 32'b00000000000000000111010100011001;
assign LUT_1[42466] = 32'b00000000000000001001110000101110;
assign LUT_1[42467] = 32'b00000000000000000011000010101010;
assign LUT_1[42468] = 32'b00000000000000010101111011110100;
assign LUT_1[42469] = 32'b00000000000000001111001101110000;
assign LUT_1[42470] = 32'b00000000000000010001101010000101;
assign LUT_1[42471] = 32'b00000000000000001010111100000001;
assign LUT_1[42472] = 32'b00000000000000001101010000010010;
assign LUT_1[42473] = 32'b00000000000000000110100010001110;
assign LUT_1[42474] = 32'b00000000000000001000111110100011;
assign LUT_1[42475] = 32'b00000000000000000010010000011111;
assign LUT_1[42476] = 32'b00000000000000010101001001101001;
assign LUT_1[42477] = 32'b00000000000000001110011011100101;
assign LUT_1[42478] = 32'b00000000000000010000110111111010;
assign LUT_1[42479] = 32'b00000000000000001010001001110110;
assign LUT_1[42480] = 32'b00000000000000001111111101111111;
assign LUT_1[42481] = 32'b00000000000000001001001111111011;
assign LUT_1[42482] = 32'b00000000000000001011101100010000;
assign LUT_1[42483] = 32'b00000000000000000100111110001100;
assign LUT_1[42484] = 32'b00000000000000010111110111010110;
assign LUT_1[42485] = 32'b00000000000000010001001001010010;
assign LUT_1[42486] = 32'b00000000000000010011100101100111;
assign LUT_1[42487] = 32'b00000000000000001100110111100011;
assign LUT_1[42488] = 32'b00000000000000001111001011110100;
assign LUT_1[42489] = 32'b00000000000000001000011101110000;
assign LUT_1[42490] = 32'b00000000000000001010111010000101;
assign LUT_1[42491] = 32'b00000000000000000100001100000001;
assign LUT_1[42492] = 32'b00000000000000010111000101001011;
assign LUT_1[42493] = 32'b00000000000000010000010111000111;
assign LUT_1[42494] = 32'b00000000000000010010110011011100;
assign LUT_1[42495] = 32'b00000000000000001100000101011000;
assign LUT_1[42496] = 32'b00000000000000000100000100000100;
assign LUT_1[42497] = 32'b11111111111111111101010110000000;
assign LUT_1[42498] = 32'b11111111111111111111110010010101;
assign LUT_1[42499] = 32'b11111111111111111001000100010001;
assign LUT_1[42500] = 32'b00000000000000001011111101011011;
assign LUT_1[42501] = 32'b00000000000000000101001111010111;
assign LUT_1[42502] = 32'b00000000000000000111101011101100;
assign LUT_1[42503] = 32'b00000000000000000000111101101000;
assign LUT_1[42504] = 32'b00000000000000000011010001111001;
assign LUT_1[42505] = 32'b11111111111111111100100011110101;
assign LUT_1[42506] = 32'b11111111111111111111000000001010;
assign LUT_1[42507] = 32'b11111111111111111000010010000110;
assign LUT_1[42508] = 32'b00000000000000001011001011010000;
assign LUT_1[42509] = 32'b00000000000000000100011101001100;
assign LUT_1[42510] = 32'b00000000000000000110111001100001;
assign LUT_1[42511] = 32'b00000000000000000000001011011101;
assign LUT_1[42512] = 32'b00000000000000000101111111100110;
assign LUT_1[42513] = 32'b11111111111111111111010001100010;
assign LUT_1[42514] = 32'b00000000000000000001101101110111;
assign LUT_1[42515] = 32'b11111111111111111010111111110011;
assign LUT_1[42516] = 32'b00000000000000001101111000111101;
assign LUT_1[42517] = 32'b00000000000000000111001010111001;
assign LUT_1[42518] = 32'b00000000000000001001100111001110;
assign LUT_1[42519] = 32'b00000000000000000010111001001010;
assign LUT_1[42520] = 32'b00000000000000000101001101011011;
assign LUT_1[42521] = 32'b11111111111111111110011111010111;
assign LUT_1[42522] = 32'b00000000000000000000111011101100;
assign LUT_1[42523] = 32'b11111111111111111010001101101000;
assign LUT_1[42524] = 32'b00000000000000001101000110110010;
assign LUT_1[42525] = 32'b00000000000000000110011000101110;
assign LUT_1[42526] = 32'b00000000000000001000110101000011;
assign LUT_1[42527] = 32'b00000000000000000010000110111111;
assign LUT_1[42528] = 32'b00000000000000000100111111000011;
assign LUT_1[42529] = 32'b11111111111111111110010000111111;
assign LUT_1[42530] = 32'b00000000000000000000101101010100;
assign LUT_1[42531] = 32'b11111111111111111001111111010000;
assign LUT_1[42532] = 32'b00000000000000001100111000011010;
assign LUT_1[42533] = 32'b00000000000000000110001010010110;
assign LUT_1[42534] = 32'b00000000000000001000100110101011;
assign LUT_1[42535] = 32'b00000000000000000001111000100111;
assign LUT_1[42536] = 32'b00000000000000000100001100111000;
assign LUT_1[42537] = 32'b11111111111111111101011110110100;
assign LUT_1[42538] = 32'b11111111111111111111111011001001;
assign LUT_1[42539] = 32'b11111111111111111001001101000101;
assign LUT_1[42540] = 32'b00000000000000001100000110001111;
assign LUT_1[42541] = 32'b00000000000000000101011000001011;
assign LUT_1[42542] = 32'b00000000000000000111110100100000;
assign LUT_1[42543] = 32'b00000000000000000001000110011100;
assign LUT_1[42544] = 32'b00000000000000000110111010100101;
assign LUT_1[42545] = 32'b00000000000000000000001100100001;
assign LUT_1[42546] = 32'b00000000000000000010101000110110;
assign LUT_1[42547] = 32'b11111111111111111011111010110010;
assign LUT_1[42548] = 32'b00000000000000001110110011111100;
assign LUT_1[42549] = 32'b00000000000000001000000101111000;
assign LUT_1[42550] = 32'b00000000000000001010100010001101;
assign LUT_1[42551] = 32'b00000000000000000011110100001001;
assign LUT_1[42552] = 32'b00000000000000000110001000011010;
assign LUT_1[42553] = 32'b11111111111111111111011010010110;
assign LUT_1[42554] = 32'b00000000000000000001110110101011;
assign LUT_1[42555] = 32'b11111111111111111011001000100111;
assign LUT_1[42556] = 32'b00000000000000001110000001110001;
assign LUT_1[42557] = 32'b00000000000000000111010011101101;
assign LUT_1[42558] = 32'b00000000000000001001110000000010;
assign LUT_1[42559] = 32'b00000000000000000011000001111110;
assign LUT_1[42560] = 32'b00000000000000000110000001101100;
assign LUT_1[42561] = 32'b11111111111111111111010011101000;
assign LUT_1[42562] = 32'b00000000000000000001101111111101;
assign LUT_1[42563] = 32'b11111111111111111011000001111001;
assign LUT_1[42564] = 32'b00000000000000001101111011000011;
assign LUT_1[42565] = 32'b00000000000000000111001100111111;
assign LUT_1[42566] = 32'b00000000000000001001101001010100;
assign LUT_1[42567] = 32'b00000000000000000010111011010000;
assign LUT_1[42568] = 32'b00000000000000000101001111100001;
assign LUT_1[42569] = 32'b11111111111111111110100001011101;
assign LUT_1[42570] = 32'b00000000000000000000111101110010;
assign LUT_1[42571] = 32'b11111111111111111010001111101110;
assign LUT_1[42572] = 32'b00000000000000001101001000111000;
assign LUT_1[42573] = 32'b00000000000000000110011010110100;
assign LUT_1[42574] = 32'b00000000000000001000110111001001;
assign LUT_1[42575] = 32'b00000000000000000010001001000101;
assign LUT_1[42576] = 32'b00000000000000000111111101001110;
assign LUT_1[42577] = 32'b00000000000000000001001111001010;
assign LUT_1[42578] = 32'b00000000000000000011101011011111;
assign LUT_1[42579] = 32'b11111111111111111100111101011011;
assign LUT_1[42580] = 32'b00000000000000001111110110100101;
assign LUT_1[42581] = 32'b00000000000000001001001000100001;
assign LUT_1[42582] = 32'b00000000000000001011100100110110;
assign LUT_1[42583] = 32'b00000000000000000100110110110010;
assign LUT_1[42584] = 32'b00000000000000000111001011000011;
assign LUT_1[42585] = 32'b00000000000000000000011100111111;
assign LUT_1[42586] = 32'b00000000000000000010111001010100;
assign LUT_1[42587] = 32'b11111111111111111100001011010000;
assign LUT_1[42588] = 32'b00000000000000001111000100011010;
assign LUT_1[42589] = 32'b00000000000000001000010110010110;
assign LUT_1[42590] = 32'b00000000000000001010110010101011;
assign LUT_1[42591] = 32'b00000000000000000100000100100111;
assign LUT_1[42592] = 32'b00000000000000000110111100101011;
assign LUT_1[42593] = 32'b00000000000000000000001110100111;
assign LUT_1[42594] = 32'b00000000000000000010101010111100;
assign LUT_1[42595] = 32'b11111111111111111011111100111000;
assign LUT_1[42596] = 32'b00000000000000001110110110000010;
assign LUT_1[42597] = 32'b00000000000000001000000111111110;
assign LUT_1[42598] = 32'b00000000000000001010100100010011;
assign LUT_1[42599] = 32'b00000000000000000011110110001111;
assign LUT_1[42600] = 32'b00000000000000000110001010100000;
assign LUT_1[42601] = 32'b11111111111111111111011100011100;
assign LUT_1[42602] = 32'b00000000000000000001111000110001;
assign LUT_1[42603] = 32'b11111111111111111011001010101101;
assign LUT_1[42604] = 32'b00000000000000001110000011110111;
assign LUT_1[42605] = 32'b00000000000000000111010101110011;
assign LUT_1[42606] = 32'b00000000000000001001110010001000;
assign LUT_1[42607] = 32'b00000000000000000011000100000100;
assign LUT_1[42608] = 32'b00000000000000001000111000001101;
assign LUT_1[42609] = 32'b00000000000000000010001010001001;
assign LUT_1[42610] = 32'b00000000000000000100100110011110;
assign LUT_1[42611] = 32'b11111111111111111101111000011010;
assign LUT_1[42612] = 32'b00000000000000010000110001100100;
assign LUT_1[42613] = 32'b00000000000000001010000011100000;
assign LUT_1[42614] = 32'b00000000000000001100011111110101;
assign LUT_1[42615] = 32'b00000000000000000101110001110001;
assign LUT_1[42616] = 32'b00000000000000001000000110000010;
assign LUT_1[42617] = 32'b00000000000000000001010111111110;
assign LUT_1[42618] = 32'b00000000000000000011110100010011;
assign LUT_1[42619] = 32'b11111111111111111101000110001111;
assign LUT_1[42620] = 32'b00000000000000001111111111011001;
assign LUT_1[42621] = 32'b00000000000000001001010001010101;
assign LUT_1[42622] = 32'b00000000000000001011101101101010;
assign LUT_1[42623] = 32'b00000000000000000100111111100110;
assign LUT_1[42624] = 32'b00000000000000000111000100000111;
assign LUT_1[42625] = 32'b00000000000000000000010110000011;
assign LUT_1[42626] = 32'b00000000000000000010110010011000;
assign LUT_1[42627] = 32'b11111111111111111100000100010100;
assign LUT_1[42628] = 32'b00000000000000001110111101011110;
assign LUT_1[42629] = 32'b00000000000000001000001111011010;
assign LUT_1[42630] = 32'b00000000000000001010101011101111;
assign LUT_1[42631] = 32'b00000000000000000011111101101011;
assign LUT_1[42632] = 32'b00000000000000000110010001111100;
assign LUT_1[42633] = 32'b11111111111111111111100011111000;
assign LUT_1[42634] = 32'b00000000000000000010000000001101;
assign LUT_1[42635] = 32'b11111111111111111011010010001001;
assign LUT_1[42636] = 32'b00000000000000001110001011010011;
assign LUT_1[42637] = 32'b00000000000000000111011101001111;
assign LUT_1[42638] = 32'b00000000000000001001111001100100;
assign LUT_1[42639] = 32'b00000000000000000011001011100000;
assign LUT_1[42640] = 32'b00000000000000001000111111101001;
assign LUT_1[42641] = 32'b00000000000000000010010001100101;
assign LUT_1[42642] = 32'b00000000000000000100101101111010;
assign LUT_1[42643] = 32'b11111111111111111101111111110110;
assign LUT_1[42644] = 32'b00000000000000010000111001000000;
assign LUT_1[42645] = 32'b00000000000000001010001010111100;
assign LUT_1[42646] = 32'b00000000000000001100100111010001;
assign LUT_1[42647] = 32'b00000000000000000101111001001101;
assign LUT_1[42648] = 32'b00000000000000001000001101011110;
assign LUT_1[42649] = 32'b00000000000000000001011111011010;
assign LUT_1[42650] = 32'b00000000000000000011111011101111;
assign LUT_1[42651] = 32'b11111111111111111101001101101011;
assign LUT_1[42652] = 32'b00000000000000010000000110110101;
assign LUT_1[42653] = 32'b00000000000000001001011000110001;
assign LUT_1[42654] = 32'b00000000000000001011110101000110;
assign LUT_1[42655] = 32'b00000000000000000101000111000010;
assign LUT_1[42656] = 32'b00000000000000000111111111000110;
assign LUT_1[42657] = 32'b00000000000000000001010001000010;
assign LUT_1[42658] = 32'b00000000000000000011101101010111;
assign LUT_1[42659] = 32'b11111111111111111100111111010011;
assign LUT_1[42660] = 32'b00000000000000001111111000011101;
assign LUT_1[42661] = 32'b00000000000000001001001010011001;
assign LUT_1[42662] = 32'b00000000000000001011100110101110;
assign LUT_1[42663] = 32'b00000000000000000100111000101010;
assign LUT_1[42664] = 32'b00000000000000000111001100111011;
assign LUT_1[42665] = 32'b00000000000000000000011110110111;
assign LUT_1[42666] = 32'b00000000000000000010111011001100;
assign LUT_1[42667] = 32'b11111111111111111100001101001000;
assign LUT_1[42668] = 32'b00000000000000001111000110010010;
assign LUT_1[42669] = 32'b00000000000000001000011000001110;
assign LUT_1[42670] = 32'b00000000000000001010110100100011;
assign LUT_1[42671] = 32'b00000000000000000100000110011111;
assign LUT_1[42672] = 32'b00000000000000001001111010101000;
assign LUT_1[42673] = 32'b00000000000000000011001100100100;
assign LUT_1[42674] = 32'b00000000000000000101101000111001;
assign LUT_1[42675] = 32'b11111111111111111110111010110101;
assign LUT_1[42676] = 32'b00000000000000010001110011111111;
assign LUT_1[42677] = 32'b00000000000000001011000101111011;
assign LUT_1[42678] = 32'b00000000000000001101100010010000;
assign LUT_1[42679] = 32'b00000000000000000110110100001100;
assign LUT_1[42680] = 32'b00000000000000001001001000011101;
assign LUT_1[42681] = 32'b00000000000000000010011010011001;
assign LUT_1[42682] = 32'b00000000000000000100110110101110;
assign LUT_1[42683] = 32'b11111111111111111110001000101010;
assign LUT_1[42684] = 32'b00000000000000010001000001110100;
assign LUT_1[42685] = 32'b00000000000000001010010011110000;
assign LUT_1[42686] = 32'b00000000000000001100110000000101;
assign LUT_1[42687] = 32'b00000000000000000110000010000001;
assign LUT_1[42688] = 32'b00000000000000001001000001101111;
assign LUT_1[42689] = 32'b00000000000000000010010011101011;
assign LUT_1[42690] = 32'b00000000000000000100110000000000;
assign LUT_1[42691] = 32'b11111111111111111110000001111100;
assign LUT_1[42692] = 32'b00000000000000010000111011000110;
assign LUT_1[42693] = 32'b00000000000000001010001101000010;
assign LUT_1[42694] = 32'b00000000000000001100101001010111;
assign LUT_1[42695] = 32'b00000000000000000101111011010011;
assign LUT_1[42696] = 32'b00000000000000001000001111100100;
assign LUT_1[42697] = 32'b00000000000000000001100001100000;
assign LUT_1[42698] = 32'b00000000000000000011111101110101;
assign LUT_1[42699] = 32'b11111111111111111101001111110001;
assign LUT_1[42700] = 32'b00000000000000010000001000111011;
assign LUT_1[42701] = 32'b00000000000000001001011010110111;
assign LUT_1[42702] = 32'b00000000000000001011110111001100;
assign LUT_1[42703] = 32'b00000000000000000101001001001000;
assign LUT_1[42704] = 32'b00000000000000001010111101010001;
assign LUT_1[42705] = 32'b00000000000000000100001111001101;
assign LUT_1[42706] = 32'b00000000000000000110101011100010;
assign LUT_1[42707] = 32'b11111111111111111111111101011110;
assign LUT_1[42708] = 32'b00000000000000010010110110101000;
assign LUT_1[42709] = 32'b00000000000000001100001000100100;
assign LUT_1[42710] = 32'b00000000000000001110100100111001;
assign LUT_1[42711] = 32'b00000000000000000111110110110101;
assign LUT_1[42712] = 32'b00000000000000001010001011000110;
assign LUT_1[42713] = 32'b00000000000000000011011101000010;
assign LUT_1[42714] = 32'b00000000000000000101111001010111;
assign LUT_1[42715] = 32'b11111111111111111111001011010011;
assign LUT_1[42716] = 32'b00000000000000010010000100011101;
assign LUT_1[42717] = 32'b00000000000000001011010110011001;
assign LUT_1[42718] = 32'b00000000000000001101110010101110;
assign LUT_1[42719] = 32'b00000000000000000111000100101010;
assign LUT_1[42720] = 32'b00000000000000001001111100101110;
assign LUT_1[42721] = 32'b00000000000000000011001110101010;
assign LUT_1[42722] = 32'b00000000000000000101101010111111;
assign LUT_1[42723] = 32'b11111111111111111110111100111011;
assign LUT_1[42724] = 32'b00000000000000010001110110000101;
assign LUT_1[42725] = 32'b00000000000000001011001000000001;
assign LUT_1[42726] = 32'b00000000000000001101100100010110;
assign LUT_1[42727] = 32'b00000000000000000110110110010010;
assign LUT_1[42728] = 32'b00000000000000001001001010100011;
assign LUT_1[42729] = 32'b00000000000000000010011100011111;
assign LUT_1[42730] = 32'b00000000000000000100111000110100;
assign LUT_1[42731] = 32'b11111111111111111110001010110000;
assign LUT_1[42732] = 32'b00000000000000010001000011111010;
assign LUT_1[42733] = 32'b00000000000000001010010101110110;
assign LUT_1[42734] = 32'b00000000000000001100110010001011;
assign LUT_1[42735] = 32'b00000000000000000110000100000111;
assign LUT_1[42736] = 32'b00000000000000001011111000010000;
assign LUT_1[42737] = 32'b00000000000000000101001010001100;
assign LUT_1[42738] = 32'b00000000000000000111100110100001;
assign LUT_1[42739] = 32'b00000000000000000000111000011101;
assign LUT_1[42740] = 32'b00000000000000010011110001100111;
assign LUT_1[42741] = 32'b00000000000000001101000011100011;
assign LUT_1[42742] = 32'b00000000000000001111011111111000;
assign LUT_1[42743] = 32'b00000000000000001000110001110100;
assign LUT_1[42744] = 32'b00000000000000001011000110000101;
assign LUT_1[42745] = 32'b00000000000000000100011000000001;
assign LUT_1[42746] = 32'b00000000000000000110110100010110;
assign LUT_1[42747] = 32'b00000000000000000000000110010010;
assign LUT_1[42748] = 32'b00000000000000010010111111011100;
assign LUT_1[42749] = 32'b00000000000000001100010001011000;
assign LUT_1[42750] = 32'b00000000000000001110101101101101;
assign LUT_1[42751] = 32'b00000000000000000111111111101001;
assign LUT_1[42752] = 32'b00000000000000000001111000010000;
assign LUT_1[42753] = 32'b11111111111111111011001010001100;
assign LUT_1[42754] = 32'b11111111111111111101100110100001;
assign LUT_1[42755] = 32'b11111111111111110110111000011101;
assign LUT_1[42756] = 32'b00000000000000001001110001100111;
assign LUT_1[42757] = 32'b00000000000000000011000011100011;
assign LUT_1[42758] = 32'b00000000000000000101011111111000;
assign LUT_1[42759] = 32'b11111111111111111110110001110100;
assign LUT_1[42760] = 32'b00000000000000000001000110000101;
assign LUT_1[42761] = 32'b11111111111111111010011000000001;
assign LUT_1[42762] = 32'b11111111111111111100110100010110;
assign LUT_1[42763] = 32'b11111111111111110110000110010010;
assign LUT_1[42764] = 32'b00000000000000001000111111011100;
assign LUT_1[42765] = 32'b00000000000000000010010001011000;
assign LUT_1[42766] = 32'b00000000000000000100101101101101;
assign LUT_1[42767] = 32'b11111111111111111101111111101001;
assign LUT_1[42768] = 32'b00000000000000000011110011110010;
assign LUT_1[42769] = 32'b11111111111111111101000101101110;
assign LUT_1[42770] = 32'b11111111111111111111100010000011;
assign LUT_1[42771] = 32'b11111111111111111000110011111111;
assign LUT_1[42772] = 32'b00000000000000001011101101001001;
assign LUT_1[42773] = 32'b00000000000000000100111111000101;
assign LUT_1[42774] = 32'b00000000000000000111011011011010;
assign LUT_1[42775] = 32'b00000000000000000000101101010110;
assign LUT_1[42776] = 32'b00000000000000000011000001100111;
assign LUT_1[42777] = 32'b11111111111111111100010011100011;
assign LUT_1[42778] = 32'b11111111111111111110101111111000;
assign LUT_1[42779] = 32'b11111111111111111000000001110100;
assign LUT_1[42780] = 32'b00000000000000001010111010111110;
assign LUT_1[42781] = 32'b00000000000000000100001100111010;
assign LUT_1[42782] = 32'b00000000000000000110101001001111;
assign LUT_1[42783] = 32'b11111111111111111111111011001011;
assign LUT_1[42784] = 32'b00000000000000000010110011001111;
assign LUT_1[42785] = 32'b11111111111111111100000101001011;
assign LUT_1[42786] = 32'b11111111111111111110100001100000;
assign LUT_1[42787] = 32'b11111111111111110111110011011100;
assign LUT_1[42788] = 32'b00000000000000001010101100100110;
assign LUT_1[42789] = 32'b00000000000000000011111110100010;
assign LUT_1[42790] = 32'b00000000000000000110011010110111;
assign LUT_1[42791] = 32'b11111111111111111111101100110011;
assign LUT_1[42792] = 32'b00000000000000000010000001000100;
assign LUT_1[42793] = 32'b11111111111111111011010011000000;
assign LUT_1[42794] = 32'b11111111111111111101101111010101;
assign LUT_1[42795] = 32'b11111111111111110111000001010001;
assign LUT_1[42796] = 32'b00000000000000001001111010011011;
assign LUT_1[42797] = 32'b00000000000000000011001100010111;
assign LUT_1[42798] = 32'b00000000000000000101101000101100;
assign LUT_1[42799] = 32'b11111111111111111110111010101000;
assign LUT_1[42800] = 32'b00000000000000000100101110110001;
assign LUT_1[42801] = 32'b11111111111111111110000000101101;
assign LUT_1[42802] = 32'b00000000000000000000011101000010;
assign LUT_1[42803] = 32'b11111111111111111001101110111110;
assign LUT_1[42804] = 32'b00000000000000001100101000001000;
assign LUT_1[42805] = 32'b00000000000000000101111010000100;
assign LUT_1[42806] = 32'b00000000000000001000010110011001;
assign LUT_1[42807] = 32'b00000000000000000001101000010101;
assign LUT_1[42808] = 32'b00000000000000000011111100100110;
assign LUT_1[42809] = 32'b11111111111111111101001110100010;
assign LUT_1[42810] = 32'b11111111111111111111101010110111;
assign LUT_1[42811] = 32'b11111111111111111000111100110011;
assign LUT_1[42812] = 32'b00000000000000001011110101111101;
assign LUT_1[42813] = 32'b00000000000000000101000111111001;
assign LUT_1[42814] = 32'b00000000000000000111100100001110;
assign LUT_1[42815] = 32'b00000000000000000000110110001010;
assign LUT_1[42816] = 32'b00000000000000000011110101111000;
assign LUT_1[42817] = 32'b11111111111111111101000111110100;
assign LUT_1[42818] = 32'b11111111111111111111100100001001;
assign LUT_1[42819] = 32'b11111111111111111000110110000101;
assign LUT_1[42820] = 32'b00000000000000001011101111001111;
assign LUT_1[42821] = 32'b00000000000000000101000001001011;
assign LUT_1[42822] = 32'b00000000000000000111011101100000;
assign LUT_1[42823] = 32'b00000000000000000000101111011100;
assign LUT_1[42824] = 32'b00000000000000000011000011101101;
assign LUT_1[42825] = 32'b11111111111111111100010101101001;
assign LUT_1[42826] = 32'b11111111111111111110110001111110;
assign LUT_1[42827] = 32'b11111111111111111000000011111010;
assign LUT_1[42828] = 32'b00000000000000001010111101000100;
assign LUT_1[42829] = 32'b00000000000000000100001111000000;
assign LUT_1[42830] = 32'b00000000000000000110101011010101;
assign LUT_1[42831] = 32'b11111111111111111111111101010001;
assign LUT_1[42832] = 32'b00000000000000000101110001011010;
assign LUT_1[42833] = 32'b11111111111111111111000011010110;
assign LUT_1[42834] = 32'b00000000000000000001011111101011;
assign LUT_1[42835] = 32'b11111111111111111010110001100111;
assign LUT_1[42836] = 32'b00000000000000001101101010110001;
assign LUT_1[42837] = 32'b00000000000000000110111100101101;
assign LUT_1[42838] = 32'b00000000000000001001011001000010;
assign LUT_1[42839] = 32'b00000000000000000010101010111110;
assign LUT_1[42840] = 32'b00000000000000000100111111001111;
assign LUT_1[42841] = 32'b11111111111111111110010001001011;
assign LUT_1[42842] = 32'b00000000000000000000101101100000;
assign LUT_1[42843] = 32'b11111111111111111001111111011100;
assign LUT_1[42844] = 32'b00000000000000001100111000100110;
assign LUT_1[42845] = 32'b00000000000000000110001010100010;
assign LUT_1[42846] = 32'b00000000000000001000100110110111;
assign LUT_1[42847] = 32'b00000000000000000001111000110011;
assign LUT_1[42848] = 32'b00000000000000000100110000110111;
assign LUT_1[42849] = 32'b11111111111111111110000010110011;
assign LUT_1[42850] = 32'b00000000000000000000011111001000;
assign LUT_1[42851] = 32'b11111111111111111001110001000100;
assign LUT_1[42852] = 32'b00000000000000001100101010001110;
assign LUT_1[42853] = 32'b00000000000000000101111100001010;
assign LUT_1[42854] = 32'b00000000000000001000011000011111;
assign LUT_1[42855] = 32'b00000000000000000001101010011011;
assign LUT_1[42856] = 32'b00000000000000000011111110101100;
assign LUT_1[42857] = 32'b11111111111111111101010000101000;
assign LUT_1[42858] = 32'b11111111111111111111101100111101;
assign LUT_1[42859] = 32'b11111111111111111000111110111001;
assign LUT_1[42860] = 32'b00000000000000001011111000000011;
assign LUT_1[42861] = 32'b00000000000000000101001001111111;
assign LUT_1[42862] = 32'b00000000000000000111100110010100;
assign LUT_1[42863] = 32'b00000000000000000000111000010000;
assign LUT_1[42864] = 32'b00000000000000000110101100011001;
assign LUT_1[42865] = 32'b11111111111111111111111110010101;
assign LUT_1[42866] = 32'b00000000000000000010011010101010;
assign LUT_1[42867] = 32'b11111111111111111011101100100110;
assign LUT_1[42868] = 32'b00000000000000001110100101110000;
assign LUT_1[42869] = 32'b00000000000000000111110111101100;
assign LUT_1[42870] = 32'b00000000000000001010010100000001;
assign LUT_1[42871] = 32'b00000000000000000011100101111101;
assign LUT_1[42872] = 32'b00000000000000000101111010001110;
assign LUT_1[42873] = 32'b11111111111111111111001100001010;
assign LUT_1[42874] = 32'b00000000000000000001101000011111;
assign LUT_1[42875] = 32'b11111111111111111010111010011011;
assign LUT_1[42876] = 32'b00000000000000001101110011100101;
assign LUT_1[42877] = 32'b00000000000000000111000101100001;
assign LUT_1[42878] = 32'b00000000000000001001100001110110;
assign LUT_1[42879] = 32'b00000000000000000010110011110010;
assign LUT_1[42880] = 32'b00000000000000000100111000010011;
assign LUT_1[42881] = 32'b11111111111111111110001010001111;
assign LUT_1[42882] = 32'b00000000000000000000100110100100;
assign LUT_1[42883] = 32'b11111111111111111001111000100000;
assign LUT_1[42884] = 32'b00000000000000001100110001101010;
assign LUT_1[42885] = 32'b00000000000000000110000011100110;
assign LUT_1[42886] = 32'b00000000000000001000011111111011;
assign LUT_1[42887] = 32'b00000000000000000001110001110111;
assign LUT_1[42888] = 32'b00000000000000000100000110001000;
assign LUT_1[42889] = 32'b11111111111111111101011000000100;
assign LUT_1[42890] = 32'b11111111111111111111110100011001;
assign LUT_1[42891] = 32'b11111111111111111001000110010101;
assign LUT_1[42892] = 32'b00000000000000001011111111011111;
assign LUT_1[42893] = 32'b00000000000000000101010001011011;
assign LUT_1[42894] = 32'b00000000000000000111101101110000;
assign LUT_1[42895] = 32'b00000000000000000000111111101100;
assign LUT_1[42896] = 32'b00000000000000000110110011110101;
assign LUT_1[42897] = 32'b00000000000000000000000101110001;
assign LUT_1[42898] = 32'b00000000000000000010100010000110;
assign LUT_1[42899] = 32'b11111111111111111011110100000010;
assign LUT_1[42900] = 32'b00000000000000001110101101001100;
assign LUT_1[42901] = 32'b00000000000000000111111111001000;
assign LUT_1[42902] = 32'b00000000000000001010011011011101;
assign LUT_1[42903] = 32'b00000000000000000011101101011001;
assign LUT_1[42904] = 32'b00000000000000000110000001101010;
assign LUT_1[42905] = 32'b11111111111111111111010011100110;
assign LUT_1[42906] = 32'b00000000000000000001101111111011;
assign LUT_1[42907] = 32'b11111111111111111011000001110111;
assign LUT_1[42908] = 32'b00000000000000001101111011000001;
assign LUT_1[42909] = 32'b00000000000000000111001100111101;
assign LUT_1[42910] = 32'b00000000000000001001101001010010;
assign LUT_1[42911] = 32'b00000000000000000010111011001110;
assign LUT_1[42912] = 32'b00000000000000000101110011010010;
assign LUT_1[42913] = 32'b11111111111111111111000101001110;
assign LUT_1[42914] = 32'b00000000000000000001100001100011;
assign LUT_1[42915] = 32'b11111111111111111010110011011111;
assign LUT_1[42916] = 32'b00000000000000001101101100101001;
assign LUT_1[42917] = 32'b00000000000000000110111110100101;
assign LUT_1[42918] = 32'b00000000000000001001011010111010;
assign LUT_1[42919] = 32'b00000000000000000010101100110110;
assign LUT_1[42920] = 32'b00000000000000000101000001000111;
assign LUT_1[42921] = 32'b11111111111111111110010011000011;
assign LUT_1[42922] = 32'b00000000000000000000101111011000;
assign LUT_1[42923] = 32'b11111111111111111010000001010100;
assign LUT_1[42924] = 32'b00000000000000001100111010011110;
assign LUT_1[42925] = 32'b00000000000000000110001100011010;
assign LUT_1[42926] = 32'b00000000000000001000101000101111;
assign LUT_1[42927] = 32'b00000000000000000001111010101011;
assign LUT_1[42928] = 32'b00000000000000000111101110110100;
assign LUT_1[42929] = 32'b00000000000000000001000000110000;
assign LUT_1[42930] = 32'b00000000000000000011011101000101;
assign LUT_1[42931] = 32'b11111111111111111100101111000001;
assign LUT_1[42932] = 32'b00000000000000001111101000001011;
assign LUT_1[42933] = 32'b00000000000000001000111010000111;
assign LUT_1[42934] = 32'b00000000000000001011010110011100;
assign LUT_1[42935] = 32'b00000000000000000100101000011000;
assign LUT_1[42936] = 32'b00000000000000000110111100101001;
assign LUT_1[42937] = 32'b00000000000000000000001110100101;
assign LUT_1[42938] = 32'b00000000000000000010101010111010;
assign LUT_1[42939] = 32'b11111111111111111011111100110110;
assign LUT_1[42940] = 32'b00000000000000001110110110000000;
assign LUT_1[42941] = 32'b00000000000000001000000111111100;
assign LUT_1[42942] = 32'b00000000000000001010100100010001;
assign LUT_1[42943] = 32'b00000000000000000011110110001101;
assign LUT_1[42944] = 32'b00000000000000000110110101111011;
assign LUT_1[42945] = 32'b00000000000000000000000111110111;
assign LUT_1[42946] = 32'b00000000000000000010100100001100;
assign LUT_1[42947] = 32'b11111111111111111011110110001000;
assign LUT_1[42948] = 32'b00000000000000001110101111010010;
assign LUT_1[42949] = 32'b00000000000000001000000001001110;
assign LUT_1[42950] = 32'b00000000000000001010011101100011;
assign LUT_1[42951] = 32'b00000000000000000011101111011111;
assign LUT_1[42952] = 32'b00000000000000000110000011110000;
assign LUT_1[42953] = 32'b11111111111111111111010101101100;
assign LUT_1[42954] = 32'b00000000000000000001110010000001;
assign LUT_1[42955] = 32'b11111111111111111011000011111101;
assign LUT_1[42956] = 32'b00000000000000001101111101000111;
assign LUT_1[42957] = 32'b00000000000000000111001111000011;
assign LUT_1[42958] = 32'b00000000000000001001101011011000;
assign LUT_1[42959] = 32'b00000000000000000010111101010100;
assign LUT_1[42960] = 32'b00000000000000001000110001011101;
assign LUT_1[42961] = 32'b00000000000000000010000011011001;
assign LUT_1[42962] = 32'b00000000000000000100011111101110;
assign LUT_1[42963] = 32'b11111111111111111101110001101010;
assign LUT_1[42964] = 32'b00000000000000010000101010110100;
assign LUT_1[42965] = 32'b00000000000000001001111100110000;
assign LUT_1[42966] = 32'b00000000000000001100011001000101;
assign LUT_1[42967] = 32'b00000000000000000101101011000001;
assign LUT_1[42968] = 32'b00000000000000000111111111010010;
assign LUT_1[42969] = 32'b00000000000000000001010001001110;
assign LUT_1[42970] = 32'b00000000000000000011101101100011;
assign LUT_1[42971] = 32'b11111111111111111100111111011111;
assign LUT_1[42972] = 32'b00000000000000001111111000101001;
assign LUT_1[42973] = 32'b00000000000000001001001010100101;
assign LUT_1[42974] = 32'b00000000000000001011100110111010;
assign LUT_1[42975] = 32'b00000000000000000100111000110110;
assign LUT_1[42976] = 32'b00000000000000000111110000111010;
assign LUT_1[42977] = 32'b00000000000000000001000010110110;
assign LUT_1[42978] = 32'b00000000000000000011011111001011;
assign LUT_1[42979] = 32'b11111111111111111100110001000111;
assign LUT_1[42980] = 32'b00000000000000001111101010010001;
assign LUT_1[42981] = 32'b00000000000000001000111100001101;
assign LUT_1[42982] = 32'b00000000000000001011011000100010;
assign LUT_1[42983] = 32'b00000000000000000100101010011110;
assign LUT_1[42984] = 32'b00000000000000000110111110101111;
assign LUT_1[42985] = 32'b00000000000000000000010000101011;
assign LUT_1[42986] = 32'b00000000000000000010101101000000;
assign LUT_1[42987] = 32'b11111111111111111011111110111100;
assign LUT_1[42988] = 32'b00000000000000001110111000000110;
assign LUT_1[42989] = 32'b00000000000000001000001010000010;
assign LUT_1[42990] = 32'b00000000000000001010100110010111;
assign LUT_1[42991] = 32'b00000000000000000011111000010011;
assign LUT_1[42992] = 32'b00000000000000001001101100011100;
assign LUT_1[42993] = 32'b00000000000000000010111110011000;
assign LUT_1[42994] = 32'b00000000000000000101011010101101;
assign LUT_1[42995] = 32'b11111111111111111110101100101001;
assign LUT_1[42996] = 32'b00000000000000010001100101110011;
assign LUT_1[42997] = 32'b00000000000000001010110111101111;
assign LUT_1[42998] = 32'b00000000000000001101010100000100;
assign LUT_1[42999] = 32'b00000000000000000110100110000000;
assign LUT_1[43000] = 32'b00000000000000001000111010010001;
assign LUT_1[43001] = 32'b00000000000000000010001100001101;
assign LUT_1[43002] = 32'b00000000000000000100101000100010;
assign LUT_1[43003] = 32'b11111111111111111101111010011110;
assign LUT_1[43004] = 32'b00000000000000010000110011101000;
assign LUT_1[43005] = 32'b00000000000000001010000101100100;
assign LUT_1[43006] = 32'b00000000000000001100100001111001;
assign LUT_1[43007] = 32'b00000000000000000101110011110101;
assign LUT_1[43008] = 32'b00000000000000000101000000110010;
assign LUT_1[43009] = 32'b11111111111111111110010010101110;
assign LUT_1[43010] = 32'b00000000000000000000101111000011;
assign LUT_1[43011] = 32'b11111111111111111010000000111111;
assign LUT_1[43012] = 32'b00000000000000001100111010001001;
assign LUT_1[43013] = 32'b00000000000000000110001100000101;
assign LUT_1[43014] = 32'b00000000000000001000101000011010;
assign LUT_1[43015] = 32'b00000000000000000001111010010110;
assign LUT_1[43016] = 32'b00000000000000000100001110100111;
assign LUT_1[43017] = 32'b11111111111111111101100000100011;
assign LUT_1[43018] = 32'b11111111111111111111111100111000;
assign LUT_1[43019] = 32'b11111111111111111001001110110100;
assign LUT_1[43020] = 32'b00000000000000001100000111111110;
assign LUT_1[43021] = 32'b00000000000000000101011001111010;
assign LUT_1[43022] = 32'b00000000000000000111110110001111;
assign LUT_1[43023] = 32'b00000000000000000001001000001011;
assign LUT_1[43024] = 32'b00000000000000000110111100010100;
assign LUT_1[43025] = 32'b00000000000000000000001110010000;
assign LUT_1[43026] = 32'b00000000000000000010101010100101;
assign LUT_1[43027] = 32'b11111111111111111011111100100001;
assign LUT_1[43028] = 32'b00000000000000001110110101101011;
assign LUT_1[43029] = 32'b00000000000000001000000111100111;
assign LUT_1[43030] = 32'b00000000000000001010100011111100;
assign LUT_1[43031] = 32'b00000000000000000011110101111000;
assign LUT_1[43032] = 32'b00000000000000000110001010001001;
assign LUT_1[43033] = 32'b11111111111111111111011100000101;
assign LUT_1[43034] = 32'b00000000000000000001111000011010;
assign LUT_1[43035] = 32'b11111111111111111011001010010110;
assign LUT_1[43036] = 32'b00000000000000001110000011100000;
assign LUT_1[43037] = 32'b00000000000000000111010101011100;
assign LUT_1[43038] = 32'b00000000000000001001110001110001;
assign LUT_1[43039] = 32'b00000000000000000011000011101101;
assign LUT_1[43040] = 32'b00000000000000000101111011110001;
assign LUT_1[43041] = 32'b11111111111111111111001101101101;
assign LUT_1[43042] = 32'b00000000000000000001101010000010;
assign LUT_1[43043] = 32'b11111111111111111010111011111110;
assign LUT_1[43044] = 32'b00000000000000001101110101001000;
assign LUT_1[43045] = 32'b00000000000000000111000111000100;
assign LUT_1[43046] = 32'b00000000000000001001100011011001;
assign LUT_1[43047] = 32'b00000000000000000010110101010101;
assign LUT_1[43048] = 32'b00000000000000000101001001100110;
assign LUT_1[43049] = 32'b11111111111111111110011011100010;
assign LUT_1[43050] = 32'b00000000000000000000110111110111;
assign LUT_1[43051] = 32'b11111111111111111010001001110011;
assign LUT_1[43052] = 32'b00000000000000001101000010111101;
assign LUT_1[43053] = 32'b00000000000000000110010100111001;
assign LUT_1[43054] = 32'b00000000000000001000110001001110;
assign LUT_1[43055] = 32'b00000000000000000010000011001010;
assign LUT_1[43056] = 32'b00000000000000000111110111010011;
assign LUT_1[43057] = 32'b00000000000000000001001001001111;
assign LUT_1[43058] = 32'b00000000000000000011100101100100;
assign LUT_1[43059] = 32'b11111111111111111100110111100000;
assign LUT_1[43060] = 32'b00000000000000001111110000101010;
assign LUT_1[43061] = 32'b00000000000000001001000010100110;
assign LUT_1[43062] = 32'b00000000000000001011011110111011;
assign LUT_1[43063] = 32'b00000000000000000100110000110111;
assign LUT_1[43064] = 32'b00000000000000000111000101001000;
assign LUT_1[43065] = 32'b00000000000000000000010111000100;
assign LUT_1[43066] = 32'b00000000000000000010110011011001;
assign LUT_1[43067] = 32'b11111111111111111100000101010101;
assign LUT_1[43068] = 32'b00000000000000001110111110011111;
assign LUT_1[43069] = 32'b00000000000000001000010000011011;
assign LUT_1[43070] = 32'b00000000000000001010101100110000;
assign LUT_1[43071] = 32'b00000000000000000011111110101100;
assign LUT_1[43072] = 32'b00000000000000000110111110011010;
assign LUT_1[43073] = 32'b00000000000000000000010000010110;
assign LUT_1[43074] = 32'b00000000000000000010101100101011;
assign LUT_1[43075] = 32'b11111111111111111011111110100111;
assign LUT_1[43076] = 32'b00000000000000001110110111110001;
assign LUT_1[43077] = 32'b00000000000000001000001001101101;
assign LUT_1[43078] = 32'b00000000000000001010100110000010;
assign LUT_1[43079] = 32'b00000000000000000011110111111110;
assign LUT_1[43080] = 32'b00000000000000000110001100001111;
assign LUT_1[43081] = 32'b11111111111111111111011110001011;
assign LUT_1[43082] = 32'b00000000000000000001111010100000;
assign LUT_1[43083] = 32'b11111111111111111011001100011100;
assign LUT_1[43084] = 32'b00000000000000001110000101100110;
assign LUT_1[43085] = 32'b00000000000000000111010111100010;
assign LUT_1[43086] = 32'b00000000000000001001110011110111;
assign LUT_1[43087] = 32'b00000000000000000011000101110011;
assign LUT_1[43088] = 32'b00000000000000001000111001111100;
assign LUT_1[43089] = 32'b00000000000000000010001011111000;
assign LUT_1[43090] = 32'b00000000000000000100101000001101;
assign LUT_1[43091] = 32'b11111111111111111101111010001001;
assign LUT_1[43092] = 32'b00000000000000010000110011010011;
assign LUT_1[43093] = 32'b00000000000000001010000101001111;
assign LUT_1[43094] = 32'b00000000000000001100100001100100;
assign LUT_1[43095] = 32'b00000000000000000101110011100000;
assign LUT_1[43096] = 32'b00000000000000001000000111110001;
assign LUT_1[43097] = 32'b00000000000000000001011001101101;
assign LUT_1[43098] = 32'b00000000000000000011110110000010;
assign LUT_1[43099] = 32'b11111111111111111101000111111110;
assign LUT_1[43100] = 32'b00000000000000010000000001001000;
assign LUT_1[43101] = 32'b00000000000000001001010011000100;
assign LUT_1[43102] = 32'b00000000000000001011101111011001;
assign LUT_1[43103] = 32'b00000000000000000101000001010101;
assign LUT_1[43104] = 32'b00000000000000000111111001011001;
assign LUT_1[43105] = 32'b00000000000000000001001011010101;
assign LUT_1[43106] = 32'b00000000000000000011100111101010;
assign LUT_1[43107] = 32'b11111111111111111100111001100110;
assign LUT_1[43108] = 32'b00000000000000001111110010110000;
assign LUT_1[43109] = 32'b00000000000000001001000100101100;
assign LUT_1[43110] = 32'b00000000000000001011100001000001;
assign LUT_1[43111] = 32'b00000000000000000100110010111101;
assign LUT_1[43112] = 32'b00000000000000000111000111001110;
assign LUT_1[43113] = 32'b00000000000000000000011001001010;
assign LUT_1[43114] = 32'b00000000000000000010110101011111;
assign LUT_1[43115] = 32'b11111111111111111100000111011011;
assign LUT_1[43116] = 32'b00000000000000001111000000100101;
assign LUT_1[43117] = 32'b00000000000000001000010010100001;
assign LUT_1[43118] = 32'b00000000000000001010101110110110;
assign LUT_1[43119] = 32'b00000000000000000100000000110010;
assign LUT_1[43120] = 32'b00000000000000001001110100111011;
assign LUT_1[43121] = 32'b00000000000000000011000110110111;
assign LUT_1[43122] = 32'b00000000000000000101100011001100;
assign LUT_1[43123] = 32'b11111111111111111110110101001000;
assign LUT_1[43124] = 32'b00000000000000010001101110010010;
assign LUT_1[43125] = 32'b00000000000000001011000000001110;
assign LUT_1[43126] = 32'b00000000000000001101011100100011;
assign LUT_1[43127] = 32'b00000000000000000110101110011111;
assign LUT_1[43128] = 32'b00000000000000001001000010110000;
assign LUT_1[43129] = 32'b00000000000000000010010100101100;
assign LUT_1[43130] = 32'b00000000000000000100110001000001;
assign LUT_1[43131] = 32'b11111111111111111110000010111101;
assign LUT_1[43132] = 32'b00000000000000010000111100000111;
assign LUT_1[43133] = 32'b00000000000000001010001110000011;
assign LUT_1[43134] = 32'b00000000000000001100101010011000;
assign LUT_1[43135] = 32'b00000000000000000101111100010100;
assign LUT_1[43136] = 32'b00000000000000001000000000110101;
assign LUT_1[43137] = 32'b00000000000000000001010010110001;
assign LUT_1[43138] = 32'b00000000000000000011101111000110;
assign LUT_1[43139] = 32'b11111111111111111101000001000010;
assign LUT_1[43140] = 32'b00000000000000001111111010001100;
assign LUT_1[43141] = 32'b00000000000000001001001100001000;
assign LUT_1[43142] = 32'b00000000000000001011101000011101;
assign LUT_1[43143] = 32'b00000000000000000100111010011001;
assign LUT_1[43144] = 32'b00000000000000000111001110101010;
assign LUT_1[43145] = 32'b00000000000000000000100000100110;
assign LUT_1[43146] = 32'b00000000000000000010111100111011;
assign LUT_1[43147] = 32'b11111111111111111100001110110111;
assign LUT_1[43148] = 32'b00000000000000001111001000000001;
assign LUT_1[43149] = 32'b00000000000000001000011001111101;
assign LUT_1[43150] = 32'b00000000000000001010110110010010;
assign LUT_1[43151] = 32'b00000000000000000100001000001110;
assign LUT_1[43152] = 32'b00000000000000001001111100010111;
assign LUT_1[43153] = 32'b00000000000000000011001110010011;
assign LUT_1[43154] = 32'b00000000000000000101101010101000;
assign LUT_1[43155] = 32'b11111111111111111110111100100100;
assign LUT_1[43156] = 32'b00000000000000010001110101101110;
assign LUT_1[43157] = 32'b00000000000000001011000111101010;
assign LUT_1[43158] = 32'b00000000000000001101100011111111;
assign LUT_1[43159] = 32'b00000000000000000110110101111011;
assign LUT_1[43160] = 32'b00000000000000001001001010001100;
assign LUT_1[43161] = 32'b00000000000000000010011100001000;
assign LUT_1[43162] = 32'b00000000000000000100111000011101;
assign LUT_1[43163] = 32'b11111111111111111110001010011001;
assign LUT_1[43164] = 32'b00000000000000010001000011100011;
assign LUT_1[43165] = 32'b00000000000000001010010101011111;
assign LUT_1[43166] = 32'b00000000000000001100110001110100;
assign LUT_1[43167] = 32'b00000000000000000110000011110000;
assign LUT_1[43168] = 32'b00000000000000001000111011110100;
assign LUT_1[43169] = 32'b00000000000000000010001101110000;
assign LUT_1[43170] = 32'b00000000000000000100101010000101;
assign LUT_1[43171] = 32'b11111111111111111101111100000001;
assign LUT_1[43172] = 32'b00000000000000010000110101001011;
assign LUT_1[43173] = 32'b00000000000000001010000111000111;
assign LUT_1[43174] = 32'b00000000000000001100100011011100;
assign LUT_1[43175] = 32'b00000000000000000101110101011000;
assign LUT_1[43176] = 32'b00000000000000001000001001101001;
assign LUT_1[43177] = 32'b00000000000000000001011011100101;
assign LUT_1[43178] = 32'b00000000000000000011110111111010;
assign LUT_1[43179] = 32'b11111111111111111101001001110110;
assign LUT_1[43180] = 32'b00000000000000010000000011000000;
assign LUT_1[43181] = 32'b00000000000000001001010100111100;
assign LUT_1[43182] = 32'b00000000000000001011110001010001;
assign LUT_1[43183] = 32'b00000000000000000101000011001101;
assign LUT_1[43184] = 32'b00000000000000001010110111010110;
assign LUT_1[43185] = 32'b00000000000000000100001001010010;
assign LUT_1[43186] = 32'b00000000000000000110100101100111;
assign LUT_1[43187] = 32'b11111111111111111111110111100011;
assign LUT_1[43188] = 32'b00000000000000010010110000101101;
assign LUT_1[43189] = 32'b00000000000000001100000010101001;
assign LUT_1[43190] = 32'b00000000000000001110011110111110;
assign LUT_1[43191] = 32'b00000000000000000111110000111010;
assign LUT_1[43192] = 32'b00000000000000001010000101001011;
assign LUT_1[43193] = 32'b00000000000000000011010111000111;
assign LUT_1[43194] = 32'b00000000000000000101110011011100;
assign LUT_1[43195] = 32'b11111111111111111111000101011000;
assign LUT_1[43196] = 32'b00000000000000010001111110100010;
assign LUT_1[43197] = 32'b00000000000000001011010000011110;
assign LUT_1[43198] = 32'b00000000000000001101101100110011;
assign LUT_1[43199] = 32'b00000000000000000110111110101111;
assign LUT_1[43200] = 32'b00000000000000001001111110011101;
assign LUT_1[43201] = 32'b00000000000000000011010000011001;
assign LUT_1[43202] = 32'b00000000000000000101101100101110;
assign LUT_1[43203] = 32'b11111111111111111110111110101010;
assign LUT_1[43204] = 32'b00000000000000010001110111110100;
assign LUT_1[43205] = 32'b00000000000000001011001001110000;
assign LUT_1[43206] = 32'b00000000000000001101100110000101;
assign LUT_1[43207] = 32'b00000000000000000110111000000001;
assign LUT_1[43208] = 32'b00000000000000001001001100010010;
assign LUT_1[43209] = 32'b00000000000000000010011110001110;
assign LUT_1[43210] = 32'b00000000000000000100111010100011;
assign LUT_1[43211] = 32'b11111111111111111110001100011111;
assign LUT_1[43212] = 32'b00000000000000010001000101101001;
assign LUT_1[43213] = 32'b00000000000000001010010111100101;
assign LUT_1[43214] = 32'b00000000000000001100110011111010;
assign LUT_1[43215] = 32'b00000000000000000110000101110110;
assign LUT_1[43216] = 32'b00000000000000001011111001111111;
assign LUT_1[43217] = 32'b00000000000000000101001011111011;
assign LUT_1[43218] = 32'b00000000000000000111101000010000;
assign LUT_1[43219] = 32'b00000000000000000000111010001100;
assign LUT_1[43220] = 32'b00000000000000010011110011010110;
assign LUT_1[43221] = 32'b00000000000000001101000101010010;
assign LUT_1[43222] = 32'b00000000000000001111100001100111;
assign LUT_1[43223] = 32'b00000000000000001000110011100011;
assign LUT_1[43224] = 32'b00000000000000001011000111110100;
assign LUT_1[43225] = 32'b00000000000000000100011001110000;
assign LUT_1[43226] = 32'b00000000000000000110110110000101;
assign LUT_1[43227] = 32'b00000000000000000000001000000001;
assign LUT_1[43228] = 32'b00000000000000010011000001001011;
assign LUT_1[43229] = 32'b00000000000000001100010011000111;
assign LUT_1[43230] = 32'b00000000000000001110101111011100;
assign LUT_1[43231] = 32'b00000000000000001000000001011000;
assign LUT_1[43232] = 32'b00000000000000001010111001011100;
assign LUT_1[43233] = 32'b00000000000000000100001011011000;
assign LUT_1[43234] = 32'b00000000000000000110100111101101;
assign LUT_1[43235] = 32'b11111111111111111111111001101001;
assign LUT_1[43236] = 32'b00000000000000010010110010110011;
assign LUT_1[43237] = 32'b00000000000000001100000100101111;
assign LUT_1[43238] = 32'b00000000000000001110100001000100;
assign LUT_1[43239] = 32'b00000000000000000111110011000000;
assign LUT_1[43240] = 32'b00000000000000001010000111010001;
assign LUT_1[43241] = 32'b00000000000000000011011001001101;
assign LUT_1[43242] = 32'b00000000000000000101110101100010;
assign LUT_1[43243] = 32'b11111111111111111111000111011110;
assign LUT_1[43244] = 32'b00000000000000010010000000101000;
assign LUT_1[43245] = 32'b00000000000000001011010010100100;
assign LUT_1[43246] = 32'b00000000000000001101101110111001;
assign LUT_1[43247] = 32'b00000000000000000111000000110101;
assign LUT_1[43248] = 32'b00000000000000001100110100111110;
assign LUT_1[43249] = 32'b00000000000000000110000110111010;
assign LUT_1[43250] = 32'b00000000000000001000100011001111;
assign LUT_1[43251] = 32'b00000000000000000001110101001011;
assign LUT_1[43252] = 32'b00000000000000010100101110010101;
assign LUT_1[43253] = 32'b00000000000000001110000000010001;
assign LUT_1[43254] = 32'b00000000000000010000011100100110;
assign LUT_1[43255] = 32'b00000000000000001001101110100010;
assign LUT_1[43256] = 32'b00000000000000001100000010110011;
assign LUT_1[43257] = 32'b00000000000000000101010100101111;
assign LUT_1[43258] = 32'b00000000000000000111110001000100;
assign LUT_1[43259] = 32'b00000000000000000001000011000000;
assign LUT_1[43260] = 32'b00000000000000010011111100001010;
assign LUT_1[43261] = 32'b00000000000000001101001110000110;
assign LUT_1[43262] = 32'b00000000000000001111101010011011;
assign LUT_1[43263] = 32'b00000000000000001000111100010111;
assign LUT_1[43264] = 32'b00000000000000000010110100111110;
assign LUT_1[43265] = 32'b11111111111111111100000110111010;
assign LUT_1[43266] = 32'b11111111111111111110100011001111;
assign LUT_1[43267] = 32'b11111111111111110111110101001011;
assign LUT_1[43268] = 32'b00000000000000001010101110010101;
assign LUT_1[43269] = 32'b00000000000000000100000000010001;
assign LUT_1[43270] = 32'b00000000000000000110011100100110;
assign LUT_1[43271] = 32'b11111111111111111111101110100010;
assign LUT_1[43272] = 32'b00000000000000000010000010110011;
assign LUT_1[43273] = 32'b11111111111111111011010100101111;
assign LUT_1[43274] = 32'b11111111111111111101110001000100;
assign LUT_1[43275] = 32'b11111111111111110111000011000000;
assign LUT_1[43276] = 32'b00000000000000001001111100001010;
assign LUT_1[43277] = 32'b00000000000000000011001110000110;
assign LUT_1[43278] = 32'b00000000000000000101101010011011;
assign LUT_1[43279] = 32'b11111111111111111110111100010111;
assign LUT_1[43280] = 32'b00000000000000000100110000100000;
assign LUT_1[43281] = 32'b11111111111111111110000010011100;
assign LUT_1[43282] = 32'b00000000000000000000011110110001;
assign LUT_1[43283] = 32'b11111111111111111001110000101101;
assign LUT_1[43284] = 32'b00000000000000001100101001110111;
assign LUT_1[43285] = 32'b00000000000000000101111011110011;
assign LUT_1[43286] = 32'b00000000000000001000011000001000;
assign LUT_1[43287] = 32'b00000000000000000001101010000100;
assign LUT_1[43288] = 32'b00000000000000000011111110010101;
assign LUT_1[43289] = 32'b11111111111111111101010000010001;
assign LUT_1[43290] = 32'b11111111111111111111101100100110;
assign LUT_1[43291] = 32'b11111111111111111000111110100010;
assign LUT_1[43292] = 32'b00000000000000001011110111101100;
assign LUT_1[43293] = 32'b00000000000000000101001001101000;
assign LUT_1[43294] = 32'b00000000000000000111100101111101;
assign LUT_1[43295] = 32'b00000000000000000000110111111001;
assign LUT_1[43296] = 32'b00000000000000000011101111111101;
assign LUT_1[43297] = 32'b11111111111111111101000001111001;
assign LUT_1[43298] = 32'b11111111111111111111011110001110;
assign LUT_1[43299] = 32'b11111111111111111000110000001010;
assign LUT_1[43300] = 32'b00000000000000001011101001010100;
assign LUT_1[43301] = 32'b00000000000000000100111011010000;
assign LUT_1[43302] = 32'b00000000000000000111010111100101;
assign LUT_1[43303] = 32'b00000000000000000000101001100001;
assign LUT_1[43304] = 32'b00000000000000000010111101110010;
assign LUT_1[43305] = 32'b11111111111111111100001111101110;
assign LUT_1[43306] = 32'b11111111111111111110101100000011;
assign LUT_1[43307] = 32'b11111111111111110111111101111111;
assign LUT_1[43308] = 32'b00000000000000001010110111001001;
assign LUT_1[43309] = 32'b00000000000000000100001001000101;
assign LUT_1[43310] = 32'b00000000000000000110100101011010;
assign LUT_1[43311] = 32'b11111111111111111111110111010110;
assign LUT_1[43312] = 32'b00000000000000000101101011011111;
assign LUT_1[43313] = 32'b11111111111111111110111101011011;
assign LUT_1[43314] = 32'b00000000000000000001011001110000;
assign LUT_1[43315] = 32'b11111111111111111010101011101100;
assign LUT_1[43316] = 32'b00000000000000001101100100110110;
assign LUT_1[43317] = 32'b00000000000000000110110110110010;
assign LUT_1[43318] = 32'b00000000000000001001010011000111;
assign LUT_1[43319] = 32'b00000000000000000010100101000011;
assign LUT_1[43320] = 32'b00000000000000000100111001010100;
assign LUT_1[43321] = 32'b11111111111111111110001011010000;
assign LUT_1[43322] = 32'b00000000000000000000100111100101;
assign LUT_1[43323] = 32'b11111111111111111001111001100001;
assign LUT_1[43324] = 32'b00000000000000001100110010101011;
assign LUT_1[43325] = 32'b00000000000000000110000100100111;
assign LUT_1[43326] = 32'b00000000000000001000100000111100;
assign LUT_1[43327] = 32'b00000000000000000001110010111000;
assign LUT_1[43328] = 32'b00000000000000000100110010100110;
assign LUT_1[43329] = 32'b11111111111111111110000100100010;
assign LUT_1[43330] = 32'b00000000000000000000100000110111;
assign LUT_1[43331] = 32'b11111111111111111001110010110011;
assign LUT_1[43332] = 32'b00000000000000001100101011111101;
assign LUT_1[43333] = 32'b00000000000000000101111101111001;
assign LUT_1[43334] = 32'b00000000000000001000011010001110;
assign LUT_1[43335] = 32'b00000000000000000001101100001010;
assign LUT_1[43336] = 32'b00000000000000000100000000011011;
assign LUT_1[43337] = 32'b11111111111111111101010010010111;
assign LUT_1[43338] = 32'b11111111111111111111101110101100;
assign LUT_1[43339] = 32'b11111111111111111001000000101000;
assign LUT_1[43340] = 32'b00000000000000001011111001110010;
assign LUT_1[43341] = 32'b00000000000000000101001011101110;
assign LUT_1[43342] = 32'b00000000000000000111101000000011;
assign LUT_1[43343] = 32'b00000000000000000000111001111111;
assign LUT_1[43344] = 32'b00000000000000000110101110001000;
assign LUT_1[43345] = 32'b00000000000000000000000000000100;
assign LUT_1[43346] = 32'b00000000000000000010011100011001;
assign LUT_1[43347] = 32'b11111111111111111011101110010101;
assign LUT_1[43348] = 32'b00000000000000001110100111011111;
assign LUT_1[43349] = 32'b00000000000000000111111001011011;
assign LUT_1[43350] = 32'b00000000000000001010010101110000;
assign LUT_1[43351] = 32'b00000000000000000011100111101100;
assign LUT_1[43352] = 32'b00000000000000000101111011111101;
assign LUT_1[43353] = 32'b11111111111111111111001101111001;
assign LUT_1[43354] = 32'b00000000000000000001101010001110;
assign LUT_1[43355] = 32'b11111111111111111010111100001010;
assign LUT_1[43356] = 32'b00000000000000001101110101010100;
assign LUT_1[43357] = 32'b00000000000000000111000111010000;
assign LUT_1[43358] = 32'b00000000000000001001100011100101;
assign LUT_1[43359] = 32'b00000000000000000010110101100001;
assign LUT_1[43360] = 32'b00000000000000000101101101100101;
assign LUT_1[43361] = 32'b11111111111111111110111111100001;
assign LUT_1[43362] = 32'b00000000000000000001011011110110;
assign LUT_1[43363] = 32'b11111111111111111010101101110010;
assign LUT_1[43364] = 32'b00000000000000001101100110111100;
assign LUT_1[43365] = 32'b00000000000000000110111000111000;
assign LUT_1[43366] = 32'b00000000000000001001010101001101;
assign LUT_1[43367] = 32'b00000000000000000010100111001001;
assign LUT_1[43368] = 32'b00000000000000000100111011011010;
assign LUT_1[43369] = 32'b11111111111111111110001101010110;
assign LUT_1[43370] = 32'b00000000000000000000101001101011;
assign LUT_1[43371] = 32'b11111111111111111001111011100111;
assign LUT_1[43372] = 32'b00000000000000001100110100110001;
assign LUT_1[43373] = 32'b00000000000000000110000110101101;
assign LUT_1[43374] = 32'b00000000000000001000100011000010;
assign LUT_1[43375] = 32'b00000000000000000001110100111110;
assign LUT_1[43376] = 32'b00000000000000000111101001000111;
assign LUT_1[43377] = 32'b00000000000000000000111011000011;
assign LUT_1[43378] = 32'b00000000000000000011010111011000;
assign LUT_1[43379] = 32'b11111111111111111100101001010100;
assign LUT_1[43380] = 32'b00000000000000001111100010011110;
assign LUT_1[43381] = 32'b00000000000000001000110100011010;
assign LUT_1[43382] = 32'b00000000000000001011010000101111;
assign LUT_1[43383] = 32'b00000000000000000100100010101011;
assign LUT_1[43384] = 32'b00000000000000000110110110111100;
assign LUT_1[43385] = 32'b00000000000000000000001000111000;
assign LUT_1[43386] = 32'b00000000000000000010100101001101;
assign LUT_1[43387] = 32'b11111111111111111011110111001001;
assign LUT_1[43388] = 32'b00000000000000001110110000010011;
assign LUT_1[43389] = 32'b00000000000000001000000010001111;
assign LUT_1[43390] = 32'b00000000000000001010011110100100;
assign LUT_1[43391] = 32'b00000000000000000011110000100000;
assign LUT_1[43392] = 32'b00000000000000000101110101000001;
assign LUT_1[43393] = 32'b11111111111111111111000110111101;
assign LUT_1[43394] = 32'b00000000000000000001100011010010;
assign LUT_1[43395] = 32'b11111111111111111010110101001110;
assign LUT_1[43396] = 32'b00000000000000001101101110011000;
assign LUT_1[43397] = 32'b00000000000000000111000000010100;
assign LUT_1[43398] = 32'b00000000000000001001011100101001;
assign LUT_1[43399] = 32'b00000000000000000010101110100101;
assign LUT_1[43400] = 32'b00000000000000000101000010110110;
assign LUT_1[43401] = 32'b11111111111111111110010100110010;
assign LUT_1[43402] = 32'b00000000000000000000110001000111;
assign LUT_1[43403] = 32'b11111111111111111010000011000011;
assign LUT_1[43404] = 32'b00000000000000001100111100001101;
assign LUT_1[43405] = 32'b00000000000000000110001110001001;
assign LUT_1[43406] = 32'b00000000000000001000101010011110;
assign LUT_1[43407] = 32'b00000000000000000001111100011010;
assign LUT_1[43408] = 32'b00000000000000000111110000100011;
assign LUT_1[43409] = 32'b00000000000000000001000010011111;
assign LUT_1[43410] = 32'b00000000000000000011011110110100;
assign LUT_1[43411] = 32'b11111111111111111100110000110000;
assign LUT_1[43412] = 32'b00000000000000001111101001111010;
assign LUT_1[43413] = 32'b00000000000000001000111011110110;
assign LUT_1[43414] = 32'b00000000000000001011011000001011;
assign LUT_1[43415] = 32'b00000000000000000100101010000111;
assign LUT_1[43416] = 32'b00000000000000000110111110011000;
assign LUT_1[43417] = 32'b00000000000000000000010000010100;
assign LUT_1[43418] = 32'b00000000000000000010101100101001;
assign LUT_1[43419] = 32'b11111111111111111011111110100101;
assign LUT_1[43420] = 32'b00000000000000001110110111101111;
assign LUT_1[43421] = 32'b00000000000000001000001001101011;
assign LUT_1[43422] = 32'b00000000000000001010100110000000;
assign LUT_1[43423] = 32'b00000000000000000011110111111100;
assign LUT_1[43424] = 32'b00000000000000000110110000000000;
assign LUT_1[43425] = 32'b00000000000000000000000001111100;
assign LUT_1[43426] = 32'b00000000000000000010011110010001;
assign LUT_1[43427] = 32'b11111111111111111011110000001101;
assign LUT_1[43428] = 32'b00000000000000001110101001010111;
assign LUT_1[43429] = 32'b00000000000000000111111011010011;
assign LUT_1[43430] = 32'b00000000000000001010010111101000;
assign LUT_1[43431] = 32'b00000000000000000011101001100100;
assign LUT_1[43432] = 32'b00000000000000000101111101110101;
assign LUT_1[43433] = 32'b11111111111111111111001111110001;
assign LUT_1[43434] = 32'b00000000000000000001101100000110;
assign LUT_1[43435] = 32'b11111111111111111010111110000010;
assign LUT_1[43436] = 32'b00000000000000001101110111001100;
assign LUT_1[43437] = 32'b00000000000000000111001001001000;
assign LUT_1[43438] = 32'b00000000000000001001100101011101;
assign LUT_1[43439] = 32'b00000000000000000010110111011001;
assign LUT_1[43440] = 32'b00000000000000001000101011100010;
assign LUT_1[43441] = 32'b00000000000000000001111101011110;
assign LUT_1[43442] = 32'b00000000000000000100011001110011;
assign LUT_1[43443] = 32'b11111111111111111101101011101111;
assign LUT_1[43444] = 32'b00000000000000010000100100111001;
assign LUT_1[43445] = 32'b00000000000000001001110110110101;
assign LUT_1[43446] = 32'b00000000000000001100010011001010;
assign LUT_1[43447] = 32'b00000000000000000101100101000110;
assign LUT_1[43448] = 32'b00000000000000000111111001010111;
assign LUT_1[43449] = 32'b00000000000000000001001011010011;
assign LUT_1[43450] = 32'b00000000000000000011100111101000;
assign LUT_1[43451] = 32'b11111111111111111100111001100100;
assign LUT_1[43452] = 32'b00000000000000001111110010101110;
assign LUT_1[43453] = 32'b00000000000000001001000100101010;
assign LUT_1[43454] = 32'b00000000000000001011100000111111;
assign LUT_1[43455] = 32'b00000000000000000100110010111011;
assign LUT_1[43456] = 32'b00000000000000000111110010101001;
assign LUT_1[43457] = 32'b00000000000000000001000100100101;
assign LUT_1[43458] = 32'b00000000000000000011100000111010;
assign LUT_1[43459] = 32'b11111111111111111100110010110110;
assign LUT_1[43460] = 32'b00000000000000001111101100000000;
assign LUT_1[43461] = 32'b00000000000000001000111101111100;
assign LUT_1[43462] = 32'b00000000000000001011011010010001;
assign LUT_1[43463] = 32'b00000000000000000100101100001101;
assign LUT_1[43464] = 32'b00000000000000000111000000011110;
assign LUT_1[43465] = 32'b00000000000000000000010010011010;
assign LUT_1[43466] = 32'b00000000000000000010101110101111;
assign LUT_1[43467] = 32'b11111111111111111100000000101011;
assign LUT_1[43468] = 32'b00000000000000001110111001110101;
assign LUT_1[43469] = 32'b00000000000000001000001011110001;
assign LUT_1[43470] = 32'b00000000000000001010101000000110;
assign LUT_1[43471] = 32'b00000000000000000011111010000010;
assign LUT_1[43472] = 32'b00000000000000001001101110001011;
assign LUT_1[43473] = 32'b00000000000000000011000000000111;
assign LUT_1[43474] = 32'b00000000000000000101011100011100;
assign LUT_1[43475] = 32'b11111111111111111110101110011000;
assign LUT_1[43476] = 32'b00000000000000010001100111100010;
assign LUT_1[43477] = 32'b00000000000000001010111001011110;
assign LUT_1[43478] = 32'b00000000000000001101010101110011;
assign LUT_1[43479] = 32'b00000000000000000110100111101111;
assign LUT_1[43480] = 32'b00000000000000001000111100000000;
assign LUT_1[43481] = 32'b00000000000000000010001101111100;
assign LUT_1[43482] = 32'b00000000000000000100101010010001;
assign LUT_1[43483] = 32'b11111111111111111101111100001101;
assign LUT_1[43484] = 32'b00000000000000010000110101010111;
assign LUT_1[43485] = 32'b00000000000000001010000111010011;
assign LUT_1[43486] = 32'b00000000000000001100100011101000;
assign LUT_1[43487] = 32'b00000000000000000101110101100100;
assign LUT_1[43488] = 32'b00000000000000001000101101101000;
assign LUT_1[43489] = 32'b00000000000000000001111111100100;
assign LUT_1[43490] = 32'b00000000000000000100011011111001;
assign LUT_1[43491] = 32'b11111111111111111101101101110101;
assign LUT_1[43492] = 32'b00000000000000010000100110111111;
assign LUT_1[43493] = 32'b00000000000000001001111000111011;
assign LUT_1[43494] = 32'b00000000000000001100010101010000;
assign LUT_1[43495] = 32'b00000000000000000101100111001100;
assign LUT_1[43496] = 32'b00000000000000000111111011011101;
assign LUT_1[43497] = 32'b00000000000000000001001101011001;
assign LUT_1[43498] = 32'b00000000000000000011101001101110;
assign LUT_1[43499] = 32'b11111111111111111100111011101010;
assign LUT_1[43500] = 32'b00000000000000001111110100110100;
assign LUT_1[43501] = 32'b00000000000000001001000110110000;
assign LUT_1[43502] = 32'b00000000000000001011100011000101;
assign LUT_1[43503] = 32'b00000000000000000100110101000001;
assign LUT_1[43504] = 32'b00000000000000001010101001001010;
assign LUT_1[43505] = 32'b00000000000000000011111011000110;
assign LUT_1[43506] = 32'b00000000000000000110010111011011;
assign LUT_1[43507] = 32'b11111111111111111111101001010111;
assign LUT_1[43508] = 32'b00000000000000010010100010100001;
assign LUT_1[43509] = 32'b00000000000000001011110100011101;
assign LUT_1[43510] = 32'b00000000000000001110010000110010;
assign LUT_1[43511] = 32'b00000000000000000111100010101110;
assign LUT_1[43512] = 32'b00000000000000001001110110111111;
assign LUT_1[43513] = 32'b00000000000000000011001000111011;
assign LUT_1[43514] = 32'b00000000000000000101100101010000;
assign LUT_1[43515] = 32'b11111111111111111110110111001100;
assign LUT_1[43516] = 32'b00000000000000010001110000010110;
assign LUT_1[43517] = 32'b00000000000000001011000010010010;
assign LUT_1[43518] = 32'b00000000000000001101011110100111;
assign LUT_1[43519] = 32'b00000000000000000110110000100011;
assign LUT_1[43520] = 32'b11111111111111111110101111001111;
assign LUT_1[43521] = 32'b11111111111111111000000001001011;
assign LUT_1[43522] = 32'b11111111111111111010011101100000;
assign LUT_1[43523] = 32'b11111111111111110011101111011100;
assign LUT_1[43524] = 32'b00000000000000000110101000100110;
assign LUT_1[43525] = 32'b11111111111111111111111010100010;
assign LUT_1[43526] = 32'b00000000000000000010010110110111;
assign LUT_1[43527] = 32'b11111111111111111011101000110011;
assign LUT_1[43528] = 32'b11111111111111111101111101000100;
assign LUT_1[43529] = 32'b11111111111111110111001111000000;
assign LUT_1[43530] = 32'b11111111111111111001101011010101;
assign LUT_1[43531] = 32'b11111111111111110010111101010001;
assign LUT_1[43532] = 32'b00000000000000000101110110011011;
assign LUT_1[43533] = 32'b11111111111111111111001000010111;
assign LUT_1[43534] = 32'b00000000000000000001100100101100;
assign LUT_1[43535] = 32'b11111111111111111010110110101000;
assign LUT_1[43536] = 32'b00000000000000000000101010110001;
assign LUT_1[43537] = 32'b11111111111111111001111100101101;
assign LUT_1[43538] = 32'b11111111111111111100011001000010;
assign LUT_1[43539] = 32'b11111111111111110101101010111110;
assign LUT_1[43540] = 32'b00000000000000001000100100001000;
assign LUT_1[43541] = 32'b00000000000000000001110110000100;
assign LUT_1[43542] = 32'b00000000000000000100010010011001;
assign LUT_1[43543] = 32'b11111111111111111101100100010101;
assign LUT_1[43544] = 32'b11111111111111111111111000100110;
assign LUT_1[43545] = 32'b11111111111111111001001010100010;
assign LUT_1[43546] = 32'b11111111111111111011100110110111;
assign LUT_1[43547] = 32'b11111111111111110100111000110011;
assign LUT_1[43548] = 32'b00000000000000000111110001111101;
assign LUT_1[43549] = 32'b00000000000000000001000011111001;
assign LUT_1[43550] = 32'b00000000000000000011100000001110;
assign LUT_1[43551] = 32'b11111111111111111100110010001010;
assign LUT_1[43552] = 32'b11111111111111111111101010001110;
assign LUT_1[43553] = 32'b11111111111111111000111100001010;
assign LUT_1[43554] = 32'b11111111111111111011011000011111;
assign LUT_1[43555] = 32'b11111111111111110100101010011011;
assign LUT_1[43556] = 32'b00000000000000000111100011100101;
assign LUT_1[43557] = 32'b00000000000000000000110101100001;
assign LUT_1[43558] = 32'b00000000000000000011010001110110;
assign LUT_1[43559] = 32'b11111111111111111100100011110010;
assign LUT_1[43560] = 32'b11111111111111111110111000000011;
assign LUT_1[43561] = 32'b11111111111111111000001001111111;
assign LUT_1[43562] = 32'b11111111111111111010100110010100;
assign LUT_1[43563] = 32'b11111111111111110011111000010000;
assign LUT_1[43564] = 32'b00000000000000000110110001011010;
assign LUT_1[43565] = 32'b00000000000000000000000011010110;
assign LUT_1[43566] = 32'b00000000000000000010011111101011;
assign LUT_1[43567] = 32'b11111111111111111011110001100111;
assign LUT_1[43568] = 32'b00000000000000000001100101110000;
assign LUT_1[43569] = 32'b11111111111111111010110111101100;
assign LUT_1[43570] = 32'b11111111111111111101010100000001;
assign LUT_1[43571] = 32'b11111111111111110110100101111101;
assign LUT_1[43572] = 32'b00000000000000001001011111000111;
assign LUT_1[43573] = 32'b00000000000000000010110001000011;
assign LUT_1[43574] = 32'b00000000000000000101001101011000;
assign LUT_1[43575] = 32'b11111111111111111110011111010100;
assign LUT_1[43576] = 32'b00000000000000000000110011100101;
assign LUT_1[43577] = 32'b11111111111111111010000101100001;
assign LUT_1[43578] = 32'b11111111111111111100100001110110;
assign LUT_1[43579] = 32'b11111111111111110101110011110010;
assign LUT_1[43580] = 32'b00000000000000001000101100111100;
assign LUT_1[43581] = 32'b00000000000000000001111110111000;
assign LUT_1[43582] = 32'b00000000000000000100011011001101;
assign LUT_1[43583] = 32'b11111111111111111101101101001001;
assign LUT_1[43584] = 32'b00000000000000000000101100110111;
assign LUT_1[43585] = 32'b11111111111111111001111110110011;
assign LUT_1[43586] = 32'b11111111111111111100011011001000;
assign LUT_1[43587] = 32'b11111111111111110101101101000100;
assign LUT_1[43588] = 32'b00000000000000001000100110001110;
assign LUT_1[43589] = 32'b00000000000000000001111000001010;
assign LUT_1[43590] = 32'b00000000000000000100010100011111;
assign LUT_1[43591] = 32'b11111111111111111101100110011011;
assign LUT_1[43592] = 32'b11111111111111111111111010101100;
assign LUT_1[43593] = 32'b11111111111111111001001100101000;
assign LUT_1[43594] = 32'b11111111111111111011101000111101;
assign LUT_1[43595] = 32'b11111111111111110100111010111001;
assign LUT_1[43596] = 32'b00000000000000000111110100000011;
assign LUT_1[43597] = 32'b00000000000000000001000101111111;
assign LUT_1[43598] = 32'b00000000000000000011100010010100;
assign LUT_1[43599] = 32'b11111111111111111100110100010000;
assign LUT_1[43600] = 32'b00000000000000000010101000011001;
assign LUT_1[43601] = 32'b11111111111111111011111010010101;
assign LUT_1[43602] = 32'b11111111111111111110010110101010;
assign LUT_1[43603] = 32'b11111111111111110111101000100110;
assign LUT_1[43604] = 32'b00000000000000001010100001110000;
assign LUT_1[43605] = 32'b00000000000000000011110011101100;
assign LUT_1[43606] = 32'b00000000000000000110010000000001;
assign LUT_1[43607] = 32'b11111111111111111111100001111101;
assign LUT_1[43608] = 32'b00000000000000000001110110001110;
assign LUT_1[43609] = 32'b11111111111111111011001000001010;
assign LUT_1[43610] = 32'b11111111111111111101100100011111;
assign LUT_1[43611] = 32'b11111111111111110110110110011011;
assign LUT_1[43612] = 32'b00000000000000001001101111100101;
assign LUT_1[43613] = 32'b00000000000000000011000001100001;
assign LUT_1[43614] = 32'b00000000000000000101011101110110;
assign LUT_1[43615] = 32'b11111111111111111110101111110010;
assign LUT_1[43616] = 32'b00000000000000000001100111110110;
assign LUT_1[43617] = 32'b11111111111111111010111001110010;
assign LUT_1[43618] = 32'b11111111111111111101010110000111;
assign LUT_1[43619] = 32'b11111111111111110110101000000011;
assign LUT_1[43620] = 32'b00000000000000001001100001001101;
assign LUT_1[43621] = 32'b00000000000000000010110011001001;
assign LUT_1[43622] = 32'b00000000000000000101001111011110;
assign LUT_1[43623] = 32'b11111111111111111110100001011010;
assign LUT_1[43624] = 32'b00000000000000000000110101101011;
assign LUT_1[43625] = 32'b11111111111111111010000111100111;
assign LUT_1[43626] = 32'b11111111111111111100100011111100;
assign LUT_1[43627] = 32'b11111111111111110101110101111000;
assign LUT_1[43628] = 32'b00000000000000001000101111000010;
assign LUT_1[43629] = 32'b00000000000000000010000000111110;
assign LUT_1[43630] = 32'b00000000000000000100011101010011;
assign LUT_1[43631] = 32'b11111111111111111101101111001111;
assign LUT_1[43632] = 32'b00000000000000000011100011011000;
assign LUT_1[43633] = 32'b11111111111111111100110101010100;
assign LUT_1[43634] = 32'b11111111111111111111010001101001;
assign LUT_1[43635] = 32'b11111111111111111000100011100101;
assign LUT_1[43636] = 32'b00000000000000001011011100101111;
assign LUT_1[43637] = 32'b00000000000000000100101110101011;
assign LUT_1[43638] = 32'b00000000000000000111001011000000;
assign LUT_1[43639] = 32'b00000000000000000000011100111100;
assign LUT_1[43640] = 32'b00000000000000000010110001001101;
assign LUT_1[43641] = 32'b11111111111111111100000011001001;
assign LUT_1[43642] = 32'b11111111111111111110011111011110;
assign LUT_1[43643] = 32'b11111111111111110111110001011010;
assign LUT_1[43644] = 32'b00000000000000001010101010100100;
assign LUT_1[43645] = 32'b00000000000000000011111100100000;
assign LUT_1[43646] = 32'b00000000000000000110011000110101;
assign LUT_1[43647] = 32'b11111111111111111111101010110001;
assign LUT_1[43648] = 32'b00000000000000000001101111010010;
assign LUT_1[43649] = 32'b11111111111111111011000001001110;
assign LUT_1[43650] = 32'b11111111111111111101011101100011;
assign LUT_1[43651] = 32'b11111111111111110110101111011111;
assign LUT_1[43652] = 32'b00000000000000001001101000101001;
assign LUT_1[43653] = 32'b00000000000000000010111010100101;
assign LUT_1[43654] = 32'b00000000000000000101010110111010;
assign LUT_1[43655] = 32'b11111111111111111110101000110110;
assign LUT_1[43656] = 32'b00000000000000000000111101000111;
assign LUT_1[43657] = 32'b11111111111111111010001111000011;
assign LUT_1[43658] = 32'b11111111111111111100101011011000;
assign LUT_1[43659] = 32'b11111111111111110101111101010100;
assign LUT_1[43660] = 32'b00000000000000001000110110011110;
assign LUT_1[43661] = 32'b00000000000000000010001000011010;
assign LUT_1[43662] = 32'b00000000000000000100100100101111;
assign LUT_1[43663] = 32'b11111111111111111101110110101011;
assign LUT_1[43664] = 32'b00000000000000000011101010110100;
assign LUT_1[43665] = 32'b11111111111111111100111100110000;
assign LUT_1[43666] = 32'b11111111111111111111011001000101;
assign LUT_1[43667] = 32'b11111111111111111000101011000001;
assign LUT_1[43668] = 32'b00000000000000001011100100001011;
assign LUT_1[43669] = 32'b00000000000000000100110110000111;
assign LUT_1[43670] = 32'b00000000000000000111010010011100;
assign LUT_1[43671] = 32'b00000000000000000000100100011000;
assign LUT_1[43672] = 32'b00000000000000000010111000101001;
assign LUT_1[43673] = 32'b11111111111111111100001010100101;
assign LUT_1[43674] = 32'b11111111111111111110100110111010;
assign LUT_1[43675] = 32'b11111111111111110111111000110110;
assign LUT_1[43676] = 32'b00000000000000001010110010000000;
assign LUT_1[43677] = 32'b00000000000000000100000011111100;
assign LUT_1[43678] = 32'b00000000000000000110100000010001;
assign LUT_1[43679] = 32'b11111111111111111111110010001101;
assign LUT_1[43680] = 32'b00000000000000000010101010010001;
assign LUT_1[43681] = 32'b11111111111111111011111100001101;
assign LUT_1[43682] = 32'b11111111111111111110011000100010;
assign LUT_1[43683] = 32'b11111111111111110111101010011110;
assign LUT_1[43684] = 32'b00000000000000001010100011101000;
assign LUT_1[43685] = 32'b00000000000000000011110101100100;
assign LUT_1[43686] = 32'b00000000000000000110010001111001;
assign LUT_1[43687] = 32'b11111111111111111111100011110101;
assign LUT_1[43688] = 32'b00000000000000000001111000000110;
assign LUT_1[43689] = 32'b11111111111111111011001010000010;
assign LUT_1[43690] = 32'b11111111111111111101100110010111;
assign LUT_1[43691] = 32'b11111111111111110110111000010011;
assign LUT_1[43692] = 32'b00000000000000001001110001011101;
assign LUT_1[43693] = 32'b00000000000000000011000011011001;
assign LUT_1[43694] = 32'b00000000000000000101011111101110;
assign LUT_1[43695] = 32'b11111111111111111110110001101010;
assign LUT_1[43696] = 32'b00000000000000000100100101110011;
assign LUT_1[43697] = 32'b11111111111111111101110111101111;
assign LUT_1[43698] = 32'b00000000000000000000010100000100;
assign LUT_1[43699] = 32'b11111111111111111001100110000000;
assign LUT_1[43700] = 32'b00000000000000001100011111001010;
assign LUT_1[43701] = 32'b00000000000000000101110001000110;
assign LUT_1[43702] = 32'b00000000000000001000001101011011;
assign LUT_1[43703] = 32'b00000000000000000001011111010111;
assign LUT_1[43704] = 32'b00000000000000000011110011101000;
assign LUT_1[43705] = 32'b11111111111111111101000101100100;
assign LUT_1[43706] = 32'b11111111111111111111100001111001;
assign LUT_1[43707] = 32'b11111111111111111000110011110101;
assign LUT_1[43708] = 32'b00000000000000001011101100111111;
assign LUT_1[43709] = 32'b00000000000000000100111110111011;
assign LUT_1[43710] = 32'b00000000000000000111011011010000;
assign LUT_1[43711] = 32'b00000000000000000000101101001100;
assign LUT_1[43712] = 32'b00000000000000000011101100111010;
assign LUT_1[43713] = 32'b11111111111111111100111110110110;
assign LUT_1[43714] = 32'b11111111111111111111011011001011;
assign LUT_1[43715] = 32'b11111111111111111000101101000111;
assign LUT_1[43716] = 32'b00000000000000001011100110010001;
assign LUT_1[43717] = 32'b00000000000000000100111000001101;
assign LUT_1[43718] = 32'b00000000000000000111010100100010;
assign LUT_1[43719] = 32'b00000000000000000000100110011110;
assign LUT_1[43720] = 32'b00000000000000000010111010101111;
assign LUT_1[43721] = 32'b11111111111111111100001100101011;
assign LUT_1[43722] = 32'b11111111111111111110101001000000;
assign LUT_1[43723] = 32'b11111111111111110111111010111100;
assign LUT_1[43724] = 32'b00000000000000001010110100000110;
assign LUT_1[43725] = 32'b00000000000000000100000110000010;
assign LUT_1[43726] = 32'b00000000000000000110100010010111;
assign LUT_1[43727] = 32'b11111111111111111111110100010011;
assign LUT_1[43728] = 32'b00000000000000000101101000011100;
assign LUT_1[43729] = 32'b11111111111111111110111010011000;
assign LUT_1[43730] = 32'b00000000000000000001010110101101;
assign LUT_1[43731] = 32'b11111111111111111010101000101001;
assign LUT_1[43732] = 32'b00000000000000001101100001110011;
assign LUT_1[43733] = 32'b00000000000000000110110011101111;
assign LUT_1[43734] = 32'b00000000000000001001010000000100;
assign LUT_1[43735] = 32'b00000000000000000010100010000000;
assign LUT_1[43736] = 32'b00000000000000000100110110010001;
assign LUT_1[43737] = 32'b11111111111111111110001000001101;
assign LUT_1[43738] = 32'b00000000000000000000100100100010;
assign LUT_1[43739] = 32'b11111111111111111001110110011110;
assign LUT_1[43740] = 32'b00000000000000001100101111101000;
assign LUT_1[43741] = 32'b00000000000000000110000001100100;
assign LUT_1[43742] = 32'b00000000000000001000011101111001;
assign LUT_1[43743] = 32'b00000000000000000001101111110101;
assign LUT_1[43744] = 32'b00000000000000000100100111111001;
assign LUT_1[43745] = 32'b11111111111111111101111001110101;
assign LUT_1[43746] = 32'b00000000000000000000010110001010;
assign LUT_1[43747] = 32'b11111111111111111001101000000110;
assign LUT_1[43748] = 32'b00000000000000001100100001010000;
assign LUT_1[43749] = 32'b00000000000000000101110011001100;
assign LUT_1[43750] = 32'b00000000000000001000001111100001;
assign LUT_1[43751] = 32'b00000000000000000001100001011101;
assign LUT_1[43752] = 32'b00000000000000000011110101101110;
assign LUT_1[43753] = 32'b11111111111111111101000111101010;
assign LUT_1[43754] = 32'b11111111111111111111100011111111;
assign LUT_1[43755] = 32'b11111111111111111000110101111011;
assign LUT_1[43756] = 32'b00000000000000001011101111000101;
assign LUT_1[43757] = 32'b00000000000000000101000001000001;
assign LUT_1[43758] = 32'b00000000000000000111011101010110;
assign LUT_1[43759] = 32'b00000000000000000000101111010010;
assign LUT_1[43760] = 32'b00000000000000000110100011011011;
assign LUT_1[43761] = 32'b11111111111111111111110101010111;
assign LUT_1[43762] = 32'b00000000000000000010010001101100;
assign LUT_1[43763] = 32'b11111111111111111011100011101000;
assign LUT_1[43764] = 32'b00000000000000001110011100110010;
assign LUT_1[43765] = 32'b00000000000000000111101110101110;
assign LUT_1[43766] = 32'b00000000000000001010001011000011;
assign LUT_1[43767] = 32'b00000000000000000011011100111111;
assign LUT_1[43768] = 32'b00000000000000000101110001010000;
assign LUT_1[43769] = 32'b11111111111111111111000011001100;
assign LUT_1[43770] = 32'b00000000000000000001011111100001;
assign LUT_1[43771] = 32'b11111111111111111010110001011101;
assign LUT_1[43772] = 32'b00000000000000001101101010100111;
assign LUT_1[43773] = 32'b00000000000000000110111100100011;
assign LUT_1[43774] = 32'b00000000000000001001011000111000;
assign LUT_1[43775] = 32'b00000000000000000010101010110100;
assign LUT_1[43776] = 32'b11111111111111111100100011011011;
assign LUT_1[43777] = 32'b11111111111111110101110101010111;
assign LUT_1[43778] = 32'b11111111111111111000010001101100;
assign LUT_1[43779] = 32'b11111111111111110001100011101000;
assign LUT_1[43780] = 32'b00000000000000000100011100110010;
assign LUT_1[43781] = 32'b11111111111111111101101110101110;
assign LUT_1[43782] = 32'b00000000000000000000001011000011;
assign LUT_1[43783] = 32'b11111111111111111001011100111111;
assign LUT_1[43784] = 32'b11111111111111111011110001010000;
assign LUT_1[43785] = 32'b11111111111111110101000011001100;
assign LUT_1[43786] = 32'b11111111111111110111011111100001;
assign LUT_1[43787] = 32'b11111111111111110000110001011101;
assign LUT_1[43788] = 32'b00000000000000000011101010100111;
assign LUT_1[43789] = 32'b11111111111111111100111100100011;
assign LUT_1[43790] = 32'b11111111111111111111011000111000;
assign LUT_1[43791] = 32'b11111111111111111000101010110100;
assign LUT_1[43792] = 32'b11111111111111111110011110111101;
assign LUT_1[43793] = 32'b11111111111111110111110000111001;
assign LUT_1[43794] = 32'b11111111111111111010001101001110;
assign LUT_1[43795] = 32'b11111111111111110011011111001010;
assign LUT_1[43796] = 32'b00000000000000000110011000010100;
assign LUT_1[43797] = 32'b11111111111111111111101010010000;
assign LUT_1[43798] = 32'b00000000000000000010000110100101;
assign LUT_1[43799] = 32'b11111111111111111011011000100001;
assign LUT_1[43800] = 32'b11111111111111111101101100110010;
assign LUT_1[43801] = 32'b11111111111111110110111110101110;
assign LUT_1[43802] = 32'b11111111111111111001011011000011;
assign LUT_1[43803] = 32'b11111111111111110010101100111111;
assign LUT_1[43804] = 32'b00000000000000000101100110001001;
assign LUT_1[43805] = 32'b11111111111111111110111000000101;
assign LUT_1[43806] = 32'b00000000000000000001010100011010;
assign LUT_1[43807] = 32'b11111111111111111010100110010110;
assign LUT_1[43808] = 32'b11111111111111111101011110011010;
assign LUT_1[43809] = 32'b11111111111111110110110000010110;
assign LUT_1[43810] = 32'b11111111111111111001001100101011;
assign LUT_1[43811] = 32'b11111111111111110010011110100111;
assign LUT_1[43812] = 32'b00000000000000000101010111110001;
assign LUT_1[43813] = 32'b11111111111111111110101001101101;
assign LUT_1[43814] = 32'b00000000000000000001000110000010;
assign LUT_1[43815] = 32'b11111111111111111010010111111110;
assign LUT_1[43816] = 32'b11111111111111111100101100001111;
assign LUT_1[43817] = 32'b11111111111111110101111110001011;
assign LUT_1[43818] = 32'b11111111111111111000011010100000;
assign LUT_1[43819] = 32'b11111111111111110001101100011100;
assign LUT_1[43820] = 32'b00000000000000000100100101100110;
assign LUT_1[43821] = 32'b11111111111111111101110111100010;
assign LUT_1[43822] = 32'b00000000000000000000010011110111;
assign LUT_1[43823] = 32'b11111111111111111001100101110011;
assign LUT_1[43824] = 32'b11111111111111111111011001111100;
assign LUT_1[43825] = 32'b11111111111111111000101011111000;
assign LUT_1[43826] = 32'b11111111111111111011001000001101;
assign LUT_1[43827] = 32'b11111111111111110100011010001001;
assign LUT_1[43828] = 32'b00000000000000000111010011010011;
assign LUT_1[43829] = 32'b00000000000000000000100101001111;
assign LUT_1[43830] = 32'b00000000000000000011000001100100;
assign LUT_1[43831] = 32'b11111111111111111100010011100000;
assign LUT_1[43832] = 32'b11111111111111111110100111110001;
assign LUT_1[43833] = 32'b11111111111111110111111001101101;
assign LUT_1[43834] = 32'b11111111111111111010010110000010;
assign LUT_1[43835] = 32'b11111111111111110011100111111110;
assign LUT_1[43836] = 32'b00000000000000000110100001001000;
assign LUT_1[43837] = 32'b11111111111111111111110011000100;
assign LUT_1[43838] = 32'b00000000000000000010001111011001;
assign LUT_1[43839] = 32'b11111111111111111011100001010101;
assign LUT_1[43840] = 32'b11111111111111111110100001000011;
assign LUT_1[43841] = 32'b11111111111111110111110010111111;
assign LUT_1[43842] = 32'b11111111111111111010001111010100;
assign LUT_1[43843] = 32'b11111111111111110011100001010000;
assign LUT_1[43844] = 32'b00000000000000000110011010011010;
assign LUT_1[43845] = 32'b11111111111111111111101100010110;
assign LUT_1[43846] = 32'b00000000000000000010001000101011;
assign LUT_1[43847] = 32'b11111111111111111011011010100111;
assign LUT_1[43848] = 32'b11111111111111111101101110111000;
assign LUT_1[43849] = 32'b11111111111111110111000000110100;
assign LUT_1[43850] = 32'b11111111111111111001011101001001;
assign LUT_1[43851] = 32'b11111111111111110010101111000101;
assign LUT_1[43852] = 32'b00000000000000000101101000001111;
assign LUT_1[43853] = 32'b11111111111111111110111010001011;
assign LUT_1[43854] = 32'b00000000000000000001010110100000;
assign LUT_1[43855] = 32'b11111111111111111010101000011100;
assign LUT_1[43856] = 32'b00000000000000000000011100100101;
assign LUT_1[43857] = 32'b11111111111111111001101110100001;
assign LUT_1[43858] = 32'b11111111111111111100001010110110;
assign LUT_1[43859] = 32'b11111111111111110101011100110010;
assign LUT_1[43860] = 32'b00000000000000001000010101111100;
assign LUT_1[43861] = 32'b00000000000000000001100111111000;
assign LUT_1[43862] = 32'b00000000000000000100000100001101;
assign LUT_1[43863] = 32'b11111111111111111101010110001001;
assign LUT_1[43864] = 32'b11111111111111111111101010011010;
assign LUT_1[43865] = 32'b11111111111111111000111100010110;
assign LUT_1[43866] = 32'b11111111111111111011011000101011;
assign LUT_1[43867] = 32'b11111111111111110100101010100111;
assign LUT_1[43868] = 32'b00000000000000000111100011110001;
assign LUT_1[43869] = 32'b00000000000000000000110101101101;
assign LUT_1[43870] = 32'b00000000000000000011010010000010;
assign LUT_1[43871] = 32'b11111111111111111100100011111110;
assign LUT_1[43872] = 32'b11111111111111111111011100000010;
assign LUT_1[43873] = 32'b11111111111111111000101101111110;
assign LUT_1[43874] = 32'b11111111111111111011001010010011;
assign LUT_1[43875] = 32'b11111111111111110100011100001111;
assign LUT_1[43876] = 32'b00000000000000000111010101011001;
assign LUT_1[43877] = 32'b00000000000000000000100111010101;
assign LUT_1[43878] = 32'b00000000000000000011000011101010;
assign LUT_1[43879] = 32'b11111111111111111100010101100110;
assign LUT_1[43880] = 32'b11111111111111111110101001110111;
assign LUT_1[43881] = 32'b11111111111111110111111011110011;
assign LUT_1[43882] = 32'b11111111111111111010011000001000;
assign LUT_1[43883] = 32'b11111111111111110011101010000100;
assign LUT_1[43884] = 32'b00000000000000000110100011001110;
assign LUT_1[43885] = 32'b11111111111111111111110101001010;
assign LUT_1[43886] = 32'b00000000000000000010010001011111;
assign LUT_1[43887] = 32'b11111111111111111011100011011011;
assign LUT_1[43888] = 32'b00000000000000000001010111100100;
assign LUT_1[43889] = 32'b11111111111111111010101001100000;
assign LUT_1[43890] = 32'b11111111111111111101000101110101;
assign LUT_1[43891] = 32'b11111111111111110110010111110001;
assign LUT_1[43892] = 32'b00000000000000001001010000111011;
assign LUT_1[43893] = 32'b00000000000000000010100010110111;
assign LUT_1[43894] = 32'b00000000000000000100111111001100;
assign LUT_1[43895] = 32'b11111111111111111110010001001000;
assign LUT_1[43896] = 32'b00000000000000000000100101011001;
assign LUT_1[43897] = 32'b11111111111111111001110111010101;
assign LUT_1[43898] = 32'b11111111111111111100010011101010;
assign LUT_1[43899] = 32'b11111111111111110101100101100110;
assign LUT_1[43900] = 32'b00000000000000001000011110110000;
assign LUT_1[43901] = 32'b00000000000000000001110000101100;
assign LUT_1[43902] = 32'b00000000000000000100001101000001;
assign LUT_1[43903] = 32'b11111111111111111101011110111101;
assign LUT_1[43904] = 32'b11111111111111111111100011011110;
assign LUT_1[43905] = 32'b11111111111111111000110101011010;
assign LUT_1[43906] = 32'b11111111111111111011010001101111;
assign LUT_1[43907] = 32'b11111111111111110100100011101011;
assign LUT_1[43908] = 32'b00000000000000000111011100110101;
assign LUT_1[43909] = 32'b00000000000000000000101110110001;
assign LUT_1[43910] = 32'b00000000000000000011001011000110;
assign LUT_1[43911] = 32'b11111111111111111100011101000010;
assign LUT_1[43912] = 32'b11111111111111111110110001010011;
assign LUT_1[43913] = 32'b11111111111111111000000011001111;
assign LUT_1[43914] = 32'b11111111111111111010011111100100;
assign LUT_1[43915] = 32'b11111111111111110011110001100000;
assign LUT_1[43916] = 32'b00000000000000000110101010101010;
assign LUT_1[43917] = 32'b11111111111111111111111100100110;
assign LUT_1[43918] = 32'b00000000000000000010011000111011;
assign LUT_1[43919] = 32'b11111111111111111011101010110111;
assign LUT_1[43920] = 32'b00000000000000000001011111000000;
assign LUT_1[43921] = 32'b11111111111111111010110000111100;
assign LUT_1[43922] = 32'b11111111111111111101001101010001;
assign LUT_1[43923] = 32'b11111111111111110110011111001101;
assign LUT_1[43924] = 32'b00000000000000001001011000010111;
assign LUT_1[43925] = 32'b00000000000000000010101010010011;
assign LUT_1[43926] = 32'b00000000000000000101000110101000;
assign LUT_1[43927] = 32'b11111111111111111110011000100100;
assign LUT_1[43928] = 32'b00000000000000000000101100110101;
assign LUT_1[43929] = 32'b11111111111111111001111110110001;
assign LUT_1[43930] = 32'b11111111111111111100011011000110;
assign LUT_1[43931] = 32'b11111111111111110101101101000010;
assign LUT_1[43932] = 32'b00000000000000001000100110001100;
assign LUT_1[43933] = 32'b00000000000000000001111000001000;
assign LUT_1[43934] = 32'b00000000000000000100010100011101;
assign LUT_1[43935] = 32'b11111111111111111101100110011001;
assign LUT_1[43936] = 32'b00000000000000000000011110011101;
assign LUT_1[43937] = 32'b11111111111111111001110000011001;
assign LUT_1[43938] = 32'b11111111111111111100001100101110;
assign LUT_1[43939] = 32'b11111111111111110101011110101010;
assign LUT_1[43940] = 32'b00000000000000001000010111110100;
assign LUT_1[43941] = 32'b00000000000000000001101001110000;
assign LUT_1[43942] = 32'b00000000000000000100000110000101;
assign LUT_1[43943] = 32'b11111111111111111101011000000001;
assign LUT_1[43944] = 32'b11111111111111111111101100010010;
assign LUT_1[43945] = 32'b11111111111111111000111110001110;
assign LUT_1[43946] = 32'b11111111111111111011011010100011;
assign LUT_1[43947] = 32'b11111111111111110100101100011111;
assign LUT_1[43948] = 32'b00000000000000000111100101101001;
assign LUT_1[43949] = 32'b00000000000000000000110111100101;
assign LUT_1[43950] = 32'b00000000000000000011010011111010;
assign LUT_1[43951] = 32'b11111111111111111100100101110110;
assign LUT_1[43952] = 32'b00000000000000000010011001111111;
assign LUT_1[43953] = 32'b11111111111111111011101011111011;
assign LUT_1[43954] = 32'b11111111111111111110001000010000;
assign LUT_1[43955] = 32'b11111111111111110111011010001100;
assign LUT_1[43956] = 32'b00000000000000001010010011010110;
assign LUT_1[43957] = 32'b00000000000000000011100101010010;
assign LUT_1[43958] = 32'b00000000000000000110000001100111;
assign LUT_1[43959] = 32'b11111111111111111111010011100011;
assign LUT_1[43960] = 32'b00000000000000000001100111110100;
assign LUT_1[43961] = 32'b11111111111111111010111001110000;
assign LUT_1[43962] = 32'b11111111111111111101010110000101;
assign LUT_1[43963] = 32'b11111111111111110110101000000001;
assign LUT_1[43964] = 32'b00000000000000001001100001001011;
assign LUT_1[43965] = 32'b00000000000000000010110011000111;
assign LUT_1[43966] = 32'b00000000000000000101001111011100;
assign LUT_1[43967] = 32'b11111111111111111110100001011000;
assign LUT_1[43968] = 32'b00000000000000000001100001000110;
assign LUT_1[43969] = 32'b11111111111111111010110011000010;
assign LUT_1[43970] = 32'b11111111111111111101001111010111;
assign LUT_1[43971] = 32'b11111111111111110110100001010011;
assign LUT_1[43972] = 32'b00000000000000001001011010011101;
assign LUT_1[43973] = 32'b00000000000000000010101100011001;
assign LUT_1[43974] = 32'b00000000000000000101001000101110;
assign LUT_1[43975] = 32'b11111111111111111110011010101010;
assign LUT_1[43976] = 32'b00000000000000000000101110111011;
assign LUT_1[43977] = 32'b11111111111111111010000000110111;
assign LUT_1[43978] = 32'b11111111111111111100011101001100;
assign LUT_1[43979] = 32'b11111111111111110101101111001000;
assign LUT_1[43980] = 32'b00000000000000001000101000010010;
assign LUT_1[43981] = 32'b00000000000000000001111010001110;
assign LUT_1[43982] = 32'b00000000000000000100010110100011;
assign LUT_1[43983] = 32'b11111111111111111101101000011111;
assign LUT_1[43984] = 32'b00000000000000000011011100101000;
assign LUT_1[43985] = 32'b11111111111111111100101110100100;
assign LUT_1[43986] = 32'b11111111111111111111001010111001;
assign LUT_1[43987] = 32'b11111111111111111000011100110101;
assign LUT_1[43988] = 32'b00000000000000001011010101111111;
assign LUT_1[43989] = 32'b00000000000000000100100111111011;
assign LUT_1[43990] = 32'b00000000000000000111000100010000;
assign LUT_1[43991] = 32'b00000000000000000000010110001100;
assign LUT_1[43992] = 32'b00000000000000000010101010011101;
assign LUT_1[43993] = 32'b11111111111111111011111100011001;
assign LUT_1[43994] = 32'b11111111111111111110011000101110;
assign LUT_1[43995] = 32'b11111111111111110111101010101010;
assign LUT_1[43996] = 32'b00000000000000001010100011110100;
assign LUT_1[43997] = 32'b00000000000000000011110101110000;
assign LUT_1[43998] = 32'b00000000000000000110010010000101;
assign LUT_1[43999] = 32'b11111111111111111111100100000001;
assign LUT_1[44000] = 32'b00000000000000000010011100000101;
assign LUT_1[44001] = 32'b11111111111111111011101110000001;
assign LUT_1[44002] = 32'b11111111111111111110001010010110;
assign LUT_1[44003] = 32'b11111111111111110111011100010010;
assign LUT_1[44004] = 32'b00000000000000001010010101011100;
assign LUT_1[44005] = 32'b00000000000000000011100111011000;
assign LUT_1[44006] = 32'b00000000000000000110000011101101;
assign LUT_1[44007] = 32'b11111111111111111111010101101001;
assign LUT_1[44008] = 32'b00000000000000000001101001111010;
assign LUT_1[44009] = 32'b11111111111111111010111011110110;
assign LUT_1[44010] = 32'b11111111111111111101011000001011;
assign LUT_1[44011] = 32'b11111111111111110110101010000111;
assign LUT_1[44012] = 32'b00000000000000001001100011010001;
assign LUT_1[44013] = 32'b00000000000000000010110101001101;
assign LUT_1[44014] = 32'b00000000000000000101010001100010;
assign LUT_1[44015] = 32'b11111111111111111110100011011110;
assign LUT_1[44016] = 32'b00000000000000000100010111100111;
assign LUT_1[44017] = 32'b11111111111111111101101001100011;
assign LUT_1[44018] = 32'b00000000000000000000000101111000;
assign LUT_1[44019] = 32'b11111111111111111001010111110100;
assign LUT_1[44020] = 32'b00000000000000001100010000111110;
assign LUT_1[44021] = 32'b00000000000000000101100010111010;
assign LUT_1[44022] = 32'b00000000000000000111111111001111;
assign LUT_1[44023] = 32'b00000000000000000001010001001011;
assign LUT_1[44024] = 32'b00000000000000000011100101011100;
assign LUT_1[44025] = 32'b11111111111111111100110111011000;
assign LUT_1[44026] = 32'b11111111111111111111010011101101;
assign LUT_1[44027] = 32'b11111111111111111000100101101001;
assign LUT_1[44028] = 32'b00000000000000001011011110110011;
assign LUT_1[44029] = 32'b00000000000000000100110000101111;
assign LUT_1[44030] = 32'b00000000000000000111001101000100;
assign LUT_1[44031] = 32'b00000000000000000000011111000000;
assign LUT_1[44032] = 32'b00000000000000001011010111100010;
assign LUT_1[44033] = 32'b00000000000000000100101001011110;
assign LUT_1[44034] = 32'b00000000000000000111000101110011;
assign LUT_1[44035] = 32'b00000000000000000000010111101111;
assign LUT_1[44036] = 32'b00000000000000010011010000111001;
assign LUT_1[44037] = 32'b00000000000000001100100010110101;
assign LUT_1[44038] = 32'b00000000000000001110111111001010;
assign LUT_1[44039] = 32'b00000000000000001000010001000110;
assign LUT_1[44040] = 32'b00000000000000001010100101010111;
assign LUT_1[44041] = 32'b00000000000000000011110111010011;
assign LUT_1[44042] = 32'b00000000000000000110010011101000;
assign LUT_1[44043] = 32'b11111111111111111111100101100100;
assign LUT_1[44044] = 32'b00000000000000010010011110101110;
assign LUT_1[44045] = 32'b00000000000000001011110000101010;
assign LUT_1[44046] = 32'b00000000000000001110001100111111;
assign LUT_1[44047] = 32'b00000000000000000111011110111011;
assign LUT_1[44048] = 32'b00000000000000001101010011000100;
assign LUT_1[44049] = 32'b00000000000000000110100101000000;
assign LUT_1[44050] = 32'b00000000000000001001000001010101;
assign LUT_1[44051] = 32'b00000000000000000010010011010001;
assign LUT_1[44052] = 32'b00000000000000010101001100011011;
assign LUT_1[44053] = 32'b00000000000000001110011110010111;
assign LUT_1[44054] = 32'b00000000000000010000111010101100;
assign LUT_1[44055] = 32'b00000000000000001010001100101000;
assign LUT_1[44056] = 32'b00000000000000001100100000111001;
assign LUT_1[44057] = 32'b00000000000000000101110010110101;
assign LUT_1[44058] = 32'b00000000000000001000001111001010;
assign LUT_1[44059] = 32'b00000000000000000001100001000110;
assign LUT_1[44060] = 32'b00000000000000010100011010010000;
assign LUT_1[44061] = 32'b00000000000000001101101100001100;
assign LUT_1[44062] = 32'b00000000000000010000001000100001;
assign LUT_1[44063] = 32'b00000000000000001001011010011101;
assign LUT_1[44064] = 32'b00000000000000001100010010100001;
assign LUT_1[44065] = 32'b00000000000000000101100100011101;
assign LUT_1[44066] = 32'b00000000000000001000000000110010;
assign LUT_1[44067] = 32'b00000000000000000001010010101110;
assign LUT_1[44068] = 32'b00000000000000010100001011111000;
assign LUT_1[44069] = 32'b00000000000000001101011101110100;
assign LUT_1[44070] = 32'b00000000000000001111111010001001;
assign LUT_1[44071] = 32'b00000000000000001001001100000101;
assign LUT_1[44072] = 32'b00000000000000001011100000010110;
assign LUT_1[44073] = 32'b00000000000000000100110010010010;
assign LUT_1[44074] = 32'b00000000000000000111001110100111;
assign LUT_1[44075] = 32'b00000000000000000000100000100011;
assign LUT_1[44076] = 32'b00000000000000010011011001101101;
assign LUT_1[44077] = 32'b00000000000000001100101011101001;
assign LUT_1[44078] = 32'b00000000000000001111000111111110;
assign LUT_1[44079] = 32'b00000000000000001000011001111010;
assign LUT_1[44080] = 32'b00000000000000001110001110000011;
assign LUT_1[44081] = 32'b00000000000000000111011111111111;
assign LUT_1[44082] = 32'b00000000000000001001111100010100;
assign LUT_1[44083] = 32'b00000000000000000011001110010000;
assign LUT_1[44084] = 32'b00000000000000010110000111011010;
assign LUT_1[44085] = 32'b00000000000000001111011001010110;
assign LUT_1[44086] = 32'b00000000000000010001110101101011;
assign LUT_1[44087] = 32'b00000000000000001011000111100111;
assign LUT_1[44088] = 32'b00000000000000001101011011111000;
assign LUT_1[44089] = 32'b00000000000000000110101101110100;
assign LUT_1[44090] = 32'b00000000000000001001001010001001;
assign LUT_1[44091] = 32'b00000000000000000010011100000101;
assign LUT_1[44092] = 32'b00000000000000010101010101001111;
assign LUT_1[44093] = 32'b00000000000000001110100111001011;
assign LUT_1[44094] = 32'b00000000000000010001000011100000;
assign LUT_1[44095] = 32'b00000000000000001010010101011100;
assign LUT_1[44096] = 32'b00000000000000001101010101001010;
assign LUT_1[44097] = 32'b00000000000000000110100111000110;
assign LUT_1[44098] = 32'b00000000000000001001000011011011;
assign LUT_1[44099] = 32'b00000000000000000010010101010111;
assign LUT_1[44100] = 32'b00000000000000010101001110100001;
assign LUT_1[44101] = 32'b00000000000000001110100000011101;
assign LUT_1[44102] = 32'b00000000000000010000111100110010;
assign LUT_1[44103] = 32'b00000000000000001010001110101110;
assign LUT_1[44104] = 32'b00000000000000001100100010111111;
assign LUT_1[44105] = 32'b00000000000000000101110100111011;
assign LUT_1[44106] = 32'b00000000000000001000010001010000;
assign LUT_1[44107] = 32'b00000000000000000001100011001100;
assign LUT_1[44108] = 32'b00000000000000010100011100010110;
assign LUT_1[44109] = 32'b00000000000000001101101110010010;
assign LUT_1[44110] = 32'b00000000000000010000001010100111;
assign LUT_1[44111] = 32'b00000000000000001001011100100011;
assign LUT_1[44112] = 32'b00000000000000001111010000101100;
assign LUT_1[44113] = 32'b00000000000000001000100010101000;
assign LUT_1[44114] = 32'b00000000000000001010111110111101;
assign LUT_1[44115] = 32'b00000000000000000100010000111001;
assign LUT_1[44116] = 32'b00000000000000010111001010000011;
assign LUT_1[44117] = 32'b00000000000000010000011011111111;
assign LUT_1[44118] = 32'b00000000000000010010111000010100;
assign LUT_1[44119] = 32'b00000000000000001100001010010000;
assign LUT_1[44120] = 32'b00000000000000001110011110100001;
assign LUT_1[44121] = 32'b00000000000000000111110000011101;
assign LUT_1[44122] = 32'b00000000000000001010001100110010;
assign LUT_1[44123] = 32'b00000000000000000011011110101110;
assign LUT_1[44124] = 32'b00000000000000010110010111111000;
assign LUT_1[44125] = 32'b00000000000000001111101001110100;
assign LUT_1[44126] = 32'b00000000000000010010000110001001;
assign LUT_1[44127] = 32'b00000000000000001011011000000101;
assign LUT_1[44128] = 32'b00000000000000001110010000001001;
assign LUT_1[44129] = 32'b00000000000000000111100010000101;
assign LUT_1[44130] = 32'b00000000000000001001111110011010;
assign LUT_1[44131] = 32'b00000000000000000011010000010110;
assign LUT_1[44132] = 32'b00000000000000010110001001100000;
assign LUT_1[44133] = 32'b00000000000000001111011011011100;
assign LUT_1[44134] = 32'b00000000000000010001110111110001;
assign LUT_1[44135] = 32'b00000000000000001011001001101101;
assign LUT_1[44136] = 32'b00000000000000001101011101111110;
assign LUT_1[44137] = 32'b00000000000000000110101111111010;
assign LUT_1[44138] = 32'b00000000000000001001001100001111;
assign LUT_1[44139] = 32'b00000000000000000010011110001011;
assign LUT_1[44140] = 32'b00000000000000010101010111010101;
assign LUT_1[44141] = 32'b00000000000000001110101001010001;
assign LUT_1[44142] = 32'b00000000000000010001000101100110;
assign LUT_1[44143] = 32'b00000000000000001010010111100010;
assign LUT_1[44144] = 32'b00000000000000010000001011101011;
assign LUT_1[44145] = 32'b00000000000000001001011101100111;
assign LUT_1[44146] = 32'b00000000000000001011111001111100;
assign LUT_1[44147] = 32'b00000000000000000101001011111000;
assign LUT_1[44148] = 32'b00000000000000011000000101000010;
assign LUT_1[44149] = 32'b00000000000000010001010110111110;
assign LUT_1[44150] = 32'b00000000000000010011110011010011;
assign LUT_1[44151] = 32'b00000000000000001101000101001111;
assign LUT_1[44152] = 32'b00000000000000001111011001100000;
assign LUT_1[44153] = 32'b00000000000000001000101011011100;
assign LUT_1[44154] = 32'b00000000000000001011000111110001;
assign LUT_1[44155] = 32'b00000000000000000100011001101101;
assign LUT_1[44156] = 32'b00000000000000010111010010110111;
assign LUT_1[44157] = 32'b00000000000000010000100100110011;
assign LUT_1[44158] = 32'b00000000000000010011000001001000;
assign LUT_1[44159] = 32'b00000000000000001100010011000100;
assign LUT_1[44160] = 32'b00000000000000001110010111100101;
assign LUT_1[44161] = 32'b00000000000000000111101001100001;
assign LUT_1[44162] = 32'b00000000000000001010000101110110;
assign LUT_1[44163] = 32'b00000000000000000011010111110010;
assign LUT_1[44164] = 32'b00000000000000010110010000111100;
assign LUT_1[44165] = 32'b00000000000000001111100010111000;
assign LUT_1[44166] = 32'b00000000000000010001111111001101;
assign LUT_1[44167] = 32'b00000000000000001011010001001001;
assign LUT_1[44168] = 32'b00000000000000001101100101011010;
assign LUT_1[44169] = 32'b00000000000000000110110111010110;
assign LUT_1[44170] = 32'b00000000000000001001010011101011;
assign LUT_1[44171] = 32'b00000000000000000010100101100111;
assign LUT_1[44172] = 32'b00000000000000010101011110110001;
assign LUT_1[44173] = 32'b00000000000000001110110000101101;
assign LUT_1[44174] = 32'b00000000000000010001001101000010;
assign LUT_1[44175] = 32'b00000000000000001010011110111110;
assign LUT_1[44176] = 32'b00000000000000010000010011000111;
assign LUT_1[44177] = 32'b00000000000000001001100101000011;
assign LUT_1[44178] = 32'b00000000000000001100000001011000;
assign LUT_1[44179] = 32'b00000000000000000101010011010100;
assign LUT_1[44180] = 32'b00000000000000011000001100011110;
assign LUT_1[44181] = 32'b00000000000000010001011110011010;
assign LUT_1[44182] = 32'b00000000000000010011111010101111;
assign LUT_1[44183] = 32'b00000000000000001101001100101011;
assign LUT_1[44184] = 32'b00000000000000001111100000111100;
assign LUT_1[44185] = 32'b00000000000000001000110010111000;
assign LUT_1[44186] = 32'b00000000000000001011001111001101;
assign LUT_1[44187] = 32'b00000000000000000100100001001001;
assign LUT_1[44188] = 32'b00000000000000010111011010010011;
assign LUT_1[44189] = 32'b00000000000000010000101100001111;
assign LUT_1[44190] = 32'b00000000000000010011001000100100;
assign LUT_1[44191] = 32'b00000000000000001100011010100000;
assign LUT_1[44192] = 32'b00000000000000001111010010100100;
assign LUT_1[44193] = 32'b00000000000000001000100100100000;
assign LUT_1[44194] = 32'b00000000000000001011000000110101;
assign LUT_1[44195] = 32'b00000000000000000100010010110001;
assign LUT_1[44196] = 32'b00000000000000010111001011111011;
assign LUT_1[44197] = 32'b00000000000000010000011101110111;
assign LUT_1[44198] = 32'b00000000000000010010111010001100;
assign LUT_1[44199] = 32'b00000000000000001100001100001000;
assign LUT_1[44200] = 32'b00000000000000001110100000011001;
assign LUT_1[44201] = 32'b00000000000000000111110010010101;
assign LUT_1[44202] = 32'b00000000000000001010001110101010;
assign LUT_1[44203] = 32'b00000000000000000011100000100110;
assign LUT_1[44204] = 32'b00000000000000010110011001110000;
assign LUT_1[44205] = 32'b00000000000000001111101011101100;
assign LUT_1[44206] = 32'b00000000000000010010001000000001;
assign LUT_1[44207] = 32'b00000000000000001011011001111101;
assign LUT_1[44208] = 32'b00000000000000010001001110000110;
assign LUT_1[44209] = 32'b00000000000000001010100000000010;
assign LUT_1[44210] = 32'b00000000000000001100111100010111;
assign LUT_1[44211] = 32'b00000000000000000110001110010011;
assign LUT_1[44212] = 32'b00000000000000011001000111011101;
assign LUT_1[44213] = 32'b00000000000000010010011001011001;
assign LUT_1[44214] = 32'b00000000000000010100110101101110;
assign LUT_1[44215] = 32'b00000000000000001110000111101010;
assign LUT_1[44216] = 32'b00000000000000010000011011111011;
assign LUT_1[44217] = 32'b00000000000000001001101101110111;
assign LUT_1[44218] = 32'b00000000000000001100001010001100;
assign LUT_1[44219] = 32'b00000000000000000101011100001000;
assign LUT_1[44220] = 32'b00000000000000011000010101010010;
assign LUT_1[44221] = 32'b00000000000000010001100111001110;
assign LUT_1[44222] = 32'b00000000000000010100000011100011;
assign LUT_1[44223] = 32'b00000000000000001101010101011111;
assign LUT_1[44224] = 32'b00000000000000010000010101001101;
assign LUT_1[44225] = 32'b00000000000000001001100111001001;
assign LUT_1[44226] = 32'b00000000000000001100000011011110;
assign LUT_1[44227] = 32'b00000000000000000101010101011010;
assign LUT_1[44228] = 32'b00000000000000011000001110100100;
assign LUT_1[44229] = 32'b00000000000000010001100000100000;
assign LUT_1[44230] = 32'b00000000000000010011111100110101;
assign LUT_1[44231] = 32'b00000000000000001101001110110001;
assign LUT_1[44232] = 32'b00000000000000001111100011000010;
assign LUT_1[44233] = 32'b00000000000000001000110100111110;
assign LUT_1[44234] = 32'b00000000000000001011010001010011;
assign LUT_1[44235] = 32'b00000000000000000100100011001111;
assign LUT_1[44236] = 32'b00000000000000010111011100011001;
assign LUT_1[44237] = 32'b00000000000000010000101110010101;
assign LUT_1[44238] = 32'b00000000000000010011001010101010;
assign LUT_1[44239] = 32'b00000000000000001100011100100110;
assign LUT_1[44240] = 32'b00000000000000010010010000101111;
assign LUT_1[44241] = 32'b00000000000000001011100010101011;
assign LUT_1[44242] = 32'b00000000000000001101111111000000;
assign LUT_1[44243] = 32'b00000000000000000111010000111100;
assign LUT_1[44244] = 32'b00000000000000011010001010000110;
assign LUT_1[44245] = 32'b00000000000000010011011100000010;
assign LUT_1[44246] = 32'b00000000000000010101111000010111;
assign LUT_1[44247] = 32'b00000000000000001111001010010011;
assign LUT_1[44248] = 32'b00000000000000010001011110100100;
assign LUT_1[44249] = 32'b00000000000000001010110000100000;
assign LUT_1[44250] = 32'b00000000000000001101001100110101;
assign LUT_1[44251] = 32'b00000000000000000110011110110001;
assign LUT_1[44252] = 32'b00000000000000011001010111111011;
assign LUT_1[44253] = 32'b00000000000000010010101001110111;
assign LUT_1[44254] = 32'b00000000000000010101000110001100;
assign LUT_1[44255] = 32'b00000000000000001110011000001000;
assign LUT_1[44256] = 32'b00000000000000010001010000001100;
assign LUT_1[44257] = 32'b00000000000000001010100010001000;
assign LUT_1[44258] = 32'b00000000000000001100111110011101;
assign LUT_1[44259] = 32'b00000000000000000110010000011001;
assign LUT_1[44260] = 32'b00000000000000011001001001100011;
assign LUT_1[44261] = 32'b00000000000000010010011011011111;
assign LUT_1[44262] = 32'b00000000000000010100110111110100;
assign LUT_1[44263] = 32'b00000000000000001110001001110000;
assign LUT_1[44264] = 32'b00000000000000010000011110000001;
assign LUT_1[44265] = 32'b00000000000000001001101111111101;
assign LUT_1[44266] = 32'b00000000000000001100001100010010;
assign LUT_1[44267] = 32'b00000000000000000101011110001110;
assign LUT_1[44268] = 32'b00000000000000011000010111011000;
assign LUT_1[44269] = 32'b00000000000000010001101001010100;
assign LUT_1[44270] = 32'b00000000000000010100000101101001;
assign LUT_1[44271] = 32'b00000000000000001101010111100101;
assign LUT_1[44272] = 32'b00000000000000010011001011101110;
assign LUT_1[44273] = 32'b00000000000000001100011101101010;
assign LUT_1[44274] = 32'b00000000000000001110111001111111;
assign LUT_1[44275] = 32'b00000000000000001000001011111011;
assign LUT_1[44276] = 32'b00000000000000011011000101000101;
assign LUT_1[44277] = 32'b00000000000000010100010111000001;
assign LUT_1[44278] = 32'b00000000000000010110110011010110;
assign LUT_1[44279] = 32'b00000000000000010000000101010010;
assign LUT_1[44280] = 32'b00000000000000010010011001100011;
assign LUT_1[44281] = 32'b00000000000000001011101011011111;
assign LUT_1[44282] = 32'b00000000000000001110000111110100;
assign LUT_1[44283] = 32'b00000000000000000111011001110000;
assign LUT_1[44284] = 32'b00000000000000011010010010111010;
assign LUT_1[44285] = 32'b00000000000000010011100100110110;
assign LUT_1[44286] = 32'b00000000000000010110000001001011;
assign LUT_1[44287] = 32'b00000000000000001111010011000111;
assign LUT_1[44288] = 32'b00000000000000001001001011101110;
assign LUT_1[44289] = 32'b00000000000000000010011101101010;
assign LUT_1[44290] = 32'b00000000000000000100111001111111;
assign LUT_1[44291] = 32'b11111111111111111110001011111011;
assign LUT_1[44292] = 32'b00000000000000010001000101000101;
assign LUT_1[44293] = 32'b00000000000000001010010111000001;
assign LUT_1[44294] = 32'b00000000000000001100110011010110;
assign LUT_1[44295] = 32'b00000000000000000110000101010010;
assign LUT_1[44296] = 32'b00000000000000001000011001100011;
assign LUT_1[44297] = 32'b00000000000000000001101011011111;
assign LUT_1[44298] = 32'b00000000000000000100000111110100;
assign LUT_1[44299] = 32'b11111111111111111101011001110000;
assign LUT_1[44300] = 32'b00000000000000010000010010111010;
assign LUT_1[44301] = 32'b00000000000000001001100100110110;
assign LUT_1[44302] = 32'b00000000000000001100000001001011;
assign LUT_1[44303] = 32'b00000000000000000101010011000111;
assign LUT_1[44304] = 32'b00000000000000001011000111010000;
assign LUT_1[44305] = 32'b00000000000000000100011001001100;
assign LUT_1[44306] = 32'b00000000000000000110110101100001;
assign LUT_1[44307] = 32'b00000000000000000000000111011101;
assign LUT_1[44308] = 32'b00000000000000010011000000100111;
assign LUT_1[44309] = 32'b00000000000000001100010010100011;
assign LUT_1[44310] = 32'b00000000000000001110101110111000;
assign LUT_1[44311] = 32'b00000000000000001000000000110100;
assign LUT_1[44312] = 32'b00000000000000001010010101000101;
assign LUT_1[44313] = 32'b00000000000000000011100111000001;
assign LUT_1[44314] = 32'b00000000000000000110000011010110;
assign LUT_1[44315] = 32'b11111111111111111111010101010010;
assign LUT_1[44316] = 32'b00000000000000010010001110011100;
assign LUT_1[44317] = 32'b00000000000000001011100000011000;
assign LUT_1[44318] = 32'b00000000000000001101111100101101;
assign LUT_1[44319] = 32'b00000000000000000111001110101001;
assign LUT_1[44320] = 32'b00000000000000001010000110101101;
assign LUT_1[44321] = 32'b00000000000000000011011000101001;
assign LUT_1[44322] = 32'b00000000000000000101110100111110;
assign LUT_1[44323] = 32'b11111111111111111111000110111010;
assign LUT_1[44324] = 32'b00000000000000010010000000000100;
assign LUT_1[44325] = 32'b00000000000000001011010010000000;
assign LUT_1[44326] = 32'b00000000000000001101101110010101;
assign LUT_1[44327] = 32'b00000000000000000111000000010001;
assign LUT_1[44328] = 32'b00000000000000001001010100100010;
assign LUT_1[44329] = 32'b00000000000000000010100110011110;
assign LUT_1[44330] = 32'b00000000000000000101000010110011;
assign LUT_1[44331] = 32'b11111111111111111110010100101111;
assign LUT_1[44332] = 32'b00000000000000010001001101111001;
assign LUT_1[44333] = 32'b00000000000000001010011111110101;
assign LUT_1[44334] = 32'b00000000000000001100111100001010;
assign LUT_1[44335] = 32'b00000000000000000110001110000110;
assign LUT_1[44336] = 32'b00000000000000001100000010001111;
assign LUT_1[44337] = 32'b00000000000000000101010100001011;
assign LUT_1[44338] = 32'b00000000000000000111110000100000;
assign LUT_1[44339] = 32'b00000000000000000001000010011100;
assign LUT_1[44340] = 32'b00000000000000010011111011100110;
assign LUT_1[44341] = 32'b00000000000000001101001101100010;
assign LUT_1[44342] = 32'b00000000000000001111101001110111;
assign LUT_1[44343] = 32'b00000000000000001000111011110011;
assign LUT_1[44344] = 32'b00000000000000001011010000000100;
assign LUT_1[44345] = 32'b00000000000000000100100010000000;
assign LUT_1[44346] = 32'b00000000000000000110111110010101;
assign LUT_1[44347] = 32'b00000000000000000000010000010001;
assign LUT_1[44348] = 32'b00000000000000010011001001011011;
assign LUT_1[44349] = 32'b00000000000000001100011011010111;
assign LUT_1[44350] = 32'b00000000000000001110110111101100;
assign LUT_1[44351] = 32'b00000000000000001000001001101000;
assign LUT_1[44352] = 32'b00000000000000001011001001010110;
assign LUT_1[44353] = 32'b00000000000000000100011011010010;
assign LUT_1[44354] = 32'b00000000000000000110110111100111;
assign LUT_1[44355] = 32'b00000000000000000000001001100011;
assign LUT_1[44356] = 32'b00000000000000010011000010101101;
assign LUT_1[44357] = 32'b00000000000000001100010100101001;
assign LUT_1[44358] = 32'b00000000000000001110110000111110;
assign LUT_1[44359] = 32'b00000000000000001000000010111010;
assign LUT_1[44360] = 32'b00000000000000001010010111001011;
assign LUT_1[44361] = 32'b00000000000000000011101001000111;
assign LUT_1[44362] = 32'b00000000000000000110000101011100;
assign LUT_1[44363] = 32'b11111111111111111111010111011000;
assign LUT_1[44364] = 32'b00000000000000010010010000100010;
assign LUT_1[44365] = 32'b00000000000000001011100010011110;
assign LUT_1[44366] = 32'b00000000000000001101111110110011;
assign LUT_1[44367] = 32'b00000000000000000111010000101111;
assign LUT_1[44368] = 32'b00000000000000001101000100111000;
assign LUT_1[44369] = 32'b00000000000000000110010110110100;
assign LUT_1[44370] = 32'b00000000000000001000110011001001;
assign LUT_1[44371] = 32'b00000000000000000010000101000101;
assign LUT_1[44372] = 32'b00000000000000010100111110001111;
assign LUT_1[44373] = 32'b00000000000000001110010000001011;
assign LUT_1[44374] = 32'b00000000000000010000101100100000;
assign LUT_1[44375] = 32'b00000000000000001001111110011100;
assign LUT_1[44376] = 32'b00000000000000001100010010101101;
assign LUT_1[44377] = 32'b00000000000000000101100100101001;
assign LUT_1[44378] = 32'b00000000000000001000000000111110;
assign LUT_1[44379] = 32'b00000000000000000001010010111010;
assign LUT_1[44380] = 32'b00000000000000010100001100000100;
assign LUT_1[44381] = 32'b00000000000000001101011110000000;
assign LUT_1[44382] = 32'b00000000000000001111111010010101;
assign LUT_1[44383] = 32'b00000000000000001001001100010001;
assign LUT_1[44384] = 32'b00000000000000001100000100010101;
assign LUT_1[44385] = 32'b00000000000000000101010110010001;
assign LUT_1[44386] = 32'b00000000000000000111110010100110;
assign LUT_1[44387] = 32'b00000000000000000001000100100010;
assign LUT_1[44388] = 32'b00000000000000010011111101101100;
assign LUT_1[44389] = 32'b00000000000000001101001111101000;
assign LUT_1[44390] = 32'b00000000000000001111101011111101;
assign LUT_1[44391] = 32'b00000000000000001000111101111001;
assign LUT_1[44392] = 32'b00000000000000001011010010001010;
assign LUT_1[44393] = 32'b00000000000000000100100100000110;
assign LUT_1[44394] = 32'b00000000000000000111000000011011;
assign LUT_1[44395] = 32'b00000000000000000000010010010111;
assign LUT_1[44396] = 32'b00000000000000010011001011100001;
assign LUT_1[44397] = 32'b00000000000000001100011101011101;
assign LUT_1[44398] = 32'b00000000000000001110111001110010;
assign LUT_1[44399] = 32'b00000000000000001000001011101110;
assign LUT_1[44400] = 32'b00000000000000001101111111110111;
assign LUT_1[44401] = 32'b00000000000000000111010001110011;
assign LUT_1[44402] = 32'b00000000000000001001101110001000;
assign LUT_1[44403] = 32'b00000000000000000011000000000100;
assign LUT_1[44404] = 32'b00000000000000010101111001001110;
assign LUT_1[44405] = 32'b00000000000000001111001011001010;
assign LUT_1[44406] = 32'b00000000000000010001100111011111;
assign LUT_1[44407] = 32'b00000000000000001010111001011011;
assign LUT_1[44408] = 32'b00000000000000001101001101101100;
assign LUT_1[44409] = 32'b00000000000000000110011111101000;
assign LUT_1[44410] = 32'b00000000000000001000111011111101;
assign LUT_1[44411] = 32'b00000000000000000010001101111001;
assign LUT_1[44412] = 32'b00000000000000010101000111000011;
assign LUT_1[44413] = 32'b00000000000000001110011000111111;
assign LUT_1[44414] = 32'b00000000000000010000110101010100;
assign LUT_1[44415] = 32'b00000000000000001010000111010000;
assign LUT_1[44416] = 32'b00000000000000001100001011110001;
assign LUT_1[44417] = 32'b00000000000000000101011101101101;
assign LUT_1[44418] = 32'b00000000000000000111111010000010;
assign LUT_1[44419] = 32'b00000000000000000001001011111110;
assign LUT_1[44420] = 32'b00000000000000010100000101001000;
assign LUT_1[44421] = 32'b00000000000000001101010111000100;
assign LUT_1[44422] = 32'b00000000000000001111110011011001;
assign LUT_1[44423] = 32'b00000000000000001001000101010101;
assign LUT_1[44424] = 32'b00000000000000001011011001100110;
assign LUT_1[44425] = 32'b00000000000000000100101011100010;
assign LUT_1[44426] = 32'b00000000000000000111000111110111;
assign LUT_1[44427] = 32'b00000000000000000000011001110011;
assign LUT_1[44428] = 32'b00000000000000010011010010111101;
assign LUT_1[44429] = 32'b00000000000000001100100100111001;
assign LUT_1[44430] = 32'b00000000000000001111000001001110;
assign LUT_1[44431] = 32'b00000000000000001000010011001010;
assign LUT_1[44432] = 32'b00000000000000001110000111010011;
assign LUT_1[44433] = 32'b00000000000000000111011001001111;
assign LUT_1[44434] = 32'b00000000000000001001110101100100;
assign LUT_1[44435] = 32'b00000000000000000011000111100000;
assign LUT_1[44436] = 32'b00000000000000010110000000101010;
assign LUT_1[44437] = 32'b00000000000000001111010010100110;
assign LUT_1[44438] = 32'b00000000000000010001101110111011;
assign LUT_1[44439] = 32'b00000000000000001011000000110111;
assign LUT_1[44440] = 32'b00000000000000001101010101001000;
assign LUT_1[44441] = 32'b00000000000000000110100111000100;
assign LUT_1[44442] = 32'b00000000000000001001000011011001;
assign LUT_1[44443] = 32'b00000000000000000010010101010101;
assign LUT_1[44444] = 32'b00000000000000010101001110011111;
assign LUT_1[44445] = 32'b00000000000000001110100000011011;
assign LUT_1[44446] = 32'b00000000000000010000111100110000;
assign LUT_1[44447] = 32'b00000000000000001010001110101100;
assign LUT_1[44448] = 32'b00000000000000001101000110110000;
assign LUT_1[44449] = 32'b00000000000000000110011000101100;
assign LUT_1[44450] = 32'b00000000000000001000110101000001;
assign LUT_1[44451] = 32'b00000000000000000010000110111101;
assign LUT_1[44452] = 32'b00000000000000010101000000000111;
assign LUT_1[44453] = 32'b00000000000000001110010010000011;
assign LUT_1[44454] = 32'b00000000000000010000101110011000;
assign LUT_1[44455] = 32'b00000000000000001010000000010100;
assign LUT_1[44456] = 32'b00000000000000001100010100100101;
assign LUT_1[44457] = 32'b00000000000000000101100110100001;
assign LUT_1[44458] = 32'b00000000000000001000000010110110;
assign LUT_1[44459] = 32'b00000000000000000001010100110010;
assign LUT_1[44460] = 32'b00000000000000010100001101111100;
assign LUT_1[44461] = 32'b00000000000000001101011111111000;
assign LUT_1[44462] = 32'b00000000000000001111111100001101;
assign LUT_1[44463] = 32'b00000000000000001001001110001001;
assign LUT_1[44464] = 32'b00000000000000001111000010010010;
assign LUT_1[44465] = 32'b00000000000000001000010100001110;
assign LUT_1[44466] = 32'b00000000000000001010110000100011;
assign LUT_1[44467] = 32'b00000000000000000100000010011111;
assign LUT_1[44468] = 32'b00000000000000010110111011101001;
assign LUT_1[44469] = 32'b00000000000000010000001101100101;
assign LUT_1[44470] = 32'b00000000000000010010101001111010;
assign LUT_1[44471] = 32'b00000000000000001011111011110110;
assign LUT_1[44472] = 32'b00000000000000001110010000000111;
assign LUT_1[44473] = 32'b00000000000000000111100010000011;
assign LUT_1[44474] = 32'b00000000000000001001111110011000;
assign LUT_1[44475] = 32'b00000000000000000011010000010100;
assign LUT_1[44476] = 32'b00000000000000010110001001011110;
assign LUT_1[44477] = 32'b00000000000000001111011011011010;
assign LUT_1[44478] = 32'b00000000000000010001110111101111;
assign LUT_1[44479] = 32'b00000000000000001011001001101011;
assign LUT_1[44480] = 32'b00000000000000001110001001011001;
assign LUT_1[44481] = 32'b00000000000000000111011011010101;
assign LUT_1[44482] = 32'b00000000000000001001110111101010;
assign LUT_1[44483] = 32'b00000000000000000011001001100110;
assign LUT_1[44484] = 32'b00000000000000010110000010110000;
assign LUT_1[44485] = 32'b00000000000000001111010100101100;
assign LUT_1[44486] = 32'b00000000000000010001110001000001;
assign LUT_1[44487] = 32'b00000000000000001011000010111101;
assign LUT_1[44488] = 32'b00000000000000001101010111001110;
assign LUT_1[44489] = 32'b00000000000000000110101001001010;
assign LUT_1[44490] = 32'b00000000000000001001000101011111;
assign LUT_1[44491] = 32'b00000000000000000010010111011011;
assign LUT_1[44492] = 32'b00000000000000010101010000100101;
assign LUT_1[44493] = 32'b00000000000000001110100010100001;
assign LUT_1[44494] = 32'b00000000000000010000111110110110;
assign LUT_1[44495] = 32'b00000000000000001010010000110010;
assign LUT_1[44496] = 32'b00000000000000010000000100111011;
assign LUT_1[44497] = 32'b00000000000000001001010110110111;
assign LUT_1[44498] = 32'b00000000000000001011110011001100;
assign LUT_1[44499] = 32'b00000000000000000101000101001000;
assign LUT_1[44500] = 32'b00000000000000010111111110010010;
assign LUT_1[44501] = 32'b00000000000000010001010000001110;
assign LUT_1[44502] = 32'b00000000000000010011101100100011;
assign LUT_1[44503] = 32'b00000000000000001100111110011111;
assign LUT_1[44504] = 32'b00000000000000001111010010110000;
assign LUT_1[44505] = 32'b00000000000000001000100100101100;
assign LUT_1[44506] = 32'b00000000000000001011000001000001;
assign LUT_1[44507] = 32'b00000000000000000100010010111101;
assign LUT_1[44508] = 32'b00000000000000010111001100000111;
assign LUT_1[44509] = 32'b00000000000000010000011110000011;
assign LUT_1[44510] = 32'b00000000000000010010111010011000;
assign LUT_1[44511] = 32'b00000000000000001100001100010100;
assign LUT_1[44512] = 32'b00000000000000001111000100011000;
assign LUT_1[44513] = 32'b00000000000000001000010110010100;
assign LUT_1[44514] = 32'b00000000000000001010110010101001;
assign LUT_1[44515] = 32'b00000000000000000100000100100101;
assign LUT_1[44516] = 32'b00000000000000010110111101101111;
assign LUT_1[44517] = 32'b00000000000000010000001111101011;
assign LUT_1[44518] = 32'b00000000000000010010101100000000;
assign LUT_1[44519] = 32'b00000000000000001011111101111100;
assign LUT_1[44520] = 32'b00000000000000001110010010001101;
assign LUT_1[44521] = 32'b00000000000000000111100100001001;
assign LUT_1[44522] = 32'b00000000000000001010000000011110;
assign LUT_1[44523] = 32'b00000000000000000011010010011010;
assign LUT_1[44524] = 32'b00000000000000010110001011100100;
assign LUT_1[44525] = 32'b00000000000000001111011101100000;
assign LUT_1[44526] = 32'b00000000000000010001111001110101;
assign LUT_1[44527] = 32'b00000000000000001011001011110001;
assign LUT_1[44528] = 32'b00000000000000010000111111111010;
assign LUT_1[44529] = 32'b00000000000000001010010001110110;
assign LUT_1[44530] = 32'b00000000000000001100101110001011;
assign LUT_1[44531] = 32'b00000000000000000110000000000111;
assign LUT_1[44532] = 32'b00000000000000011000111001010001;
assign LUT_1[44533] = 32'b00000000000000010010001011001101;
assign LUT_1[44534] = 32'b00000000000000010100100111100010;
assign LUT_1[44535] = 32'b00000000000000001101111001011110;
assign LUT_1[44536] = 32'b00000000000000010000001101101111;
assign LUT_1[44537] = 32'b00000000000000001001011111101011;
assign LUT_1[44538] = 32'b00000000000000001011111100000000;
assign LUT_1[44539] = 32'b00000000000000000101001101111100;
assign LUT_1[44540] = 32'b00000000000000011000000111000110;
assign LUT_1[44541] = 32'b00000000000000010001011001000010;
assign LUT_1[44542] = 32'b00000000000000010011110101010111;
assign LUT_1[44543] = 32'b00000000000000001101000111010011;
assign LUT_1[44544] = 32'b00000000000000000101000101111111;
assign LUT_1[44545] = 32'b11111111111111111110010111111011;
assign LUT_1[44546] = 32'b00000000000000000000110100010000;
assign LUT_1[44547] = 32'b11111111111111111010000110001100;
assign LUT_1[44548] = 32'b00000000000000001100111111010110;
assign LUT_1[44549] = 32'b00000000000000000110010001010010;
assign LUT_1[44550] = 32'b00000000000000001000101101100111;
assign LUT_1[44551] = 32'b00000000000000000001111111100011;
assign LUT_1[44552] = 32'b00000000000000000100010011110100;
assign LUT_1[44553] = 32'b11111111111111111101100101110000;
assign LUT_1[44554] = 32'b00000000000000000000000010000101;
assign LUT_1[44555] = 32'b11111111111111111001010100000001;
assign LUT_1[44556] = 32'b00000000000000001100001101001011;
assign LUT_1[44557] = 32'b00000000000000000101011111000111;
assign LUT_1[44558] = 32'b00000000000000000111111011011100;
assign LUT_1[44559] = 32'b00000000000000000001001101011000;
assign LUT_1[44560] = 32'b00000000000000000111000001100001;
assign LUT_1[44561] = 32'b00000000000000000000010011011101;
assign LUT_1[44562] = 32'b00000000000000000010101111110010;
assign LUT_1[44563] = 32'b11111111111111111100000001101110;
assign LUT_1[44564] = 32'b00000000000000001110111010111000;
assign LUT_1[44565] = 32'b00000000000000001000001100110100;
assign LUT_1[44566] = 32'b00000000000000001010101001001001;
assign LUT_1[44567] = 32'b00000000000000000011111011000101;
assign LUT_1[44568] = 32'b00000000000000000110001111010110;
assign LUT_1[44569] = 32'b11111111111111111111100001010010;
assign LUT_1[44570] = 32'b00000000000000000001111101100111;
assign LUT_1[44571] = 32'b11111111111111111011001111100011;
assign LUT_1[44572] = 32'b00000000000000001110001000101101;
assign LUT_1[44573] = 32'b00000000000000000111011010101001;
assign LUT_1[44574] = 32'b00000000000000001001110110111110;
assign LUT_1[44575] = 32'b00000000000000000011001000111010;
assign LUT_1[44576] = 32'b00000000000000000110000000111110;
assign LUT_1[44577] = 32'b11111111111111111111010010111010;
assign LUT_1[44578] = 32'b00000000000000000001101111001111;
assign LUT_1[44579] = 32'b11111111111111111011000001001011;
assign LUT_1[44580] = 32'b00000000000000001101111010010101;
assign LUT_1[44581] = 32'b00000000000000000111001100010001;
assign LUT_1[44582] = 32'b00000000000000001001101000100110;
assign LUT_1[44583] = 32'b00000000000000000010111010100010;
assign LUT_1[44584] = 32'b00000000000000000101001110110011;
assign LUT_1[44585] = 32'b11111111111111111110100000101111;
assign LUT_1[44586] = 32'b00000000000000000000111101000100;
assign LUT_1[44587] = 32'b11111111111111111010001111000000;
assign LUT_1[44588] = 32'b00000000000000001101001000001010;
assign LUT_1[44589] = 32'b00000000000000000110011010000110;
assign LUT_1[44590] = 32'b00000000000000001000110110011011;
assign LUT_1[44591] = 32'b00000000000000000010001000010111;
assign LUT_1[44592] = 32'b00000000000000000111111100100000;
assign LUT_1[44593] = 32'b00000000000000000001001110011100;
assign LUT_1[44594] = 32'b00000000000000000011101010110001;
assign LUT_1[44595] = 32'b11111111111111111100111100101101;
assign LUT_1[44596] = 32'b00000000000000001111110101110111;
assign LUT_1[44597] = 32'b00000000000000001001000111110011;
assign LUT_1[44598] = 32'b00000000000000001011100100001000;
assign LUT_1[44599] = 32'b00000000000000000100110110000100;
assign LUT_1[44600] = 32'b00000000000000000111001010010101;
assign LUT_1[44601] = 32'b00000000000000000000011100010001;
assign LUT_1[44602] = 32'b00000000000000000010111000100110;
assign LUT_1[44603] = 32'b11111111111111111100001010100010;
assign LUT_1[44604] = 32'b00000000000000001111000011101100;
assign LUT_1[44605] = 32'b00000000000000001000010101101000;
assign LUT_1[44606] = 32'b00000000000000001010110001111101;
assign LUT_1[44607] = 32'b00000000000000000100000011111001;
assign LUT_1[44608] = 32'b00000000000000000111000011100111;
assign LUT_1[44609] = 32'b00000000000000000000010101100011;
assign LUT_1[44610] = 32'b00000000000000000010110001111000;
assign LUT_1[44611] = 32'b11111111111111111100000011110100;
assign LUT_1[44612] = 32'b00000000000000001110111100111110;
assign LUT_1[44613] = 32'b00000000000000001000001110111010;
assign LUT_1[44614] = 32'b00000000000000001010101011001111;
assign LUT_1[44615] = 32'b00000000000000000011111101001011;
assign LUT_1[44616] = 32'b00000000000000000110010001011100;
assign LUT_1[44617] = 32'b11111111111111111111100011011000;
assign LUT_1[44618] = 32'b00000000000000000001111111101101;
assign LUT_1[44619] = 32'b11111111111111111011010001101001;
assign LUT_1[44620] = 32'b00000000000000001110001010110011;
assign LUT_1[44621] = 32'b00000000000000000111011100101111;
assign LUT_1[44622] = 32'b00000000000000001001111001000100;
assign LUT_1[44623] = 32'b00000000000000000011001011000000;
assign LUT_1[44624] = 32'b00000000000000001000111111001001;
assign LUT_1[44625] = 32'b00000000000000000010010001000101;
assign LUT_1[44626] = 32'b00000000000000000100101101011010;
assign LUT_1[44627] = 32'b11111111111111111101111111010110;
assign LUT_1[44628] = 32'b00000000000000010000111000100000;
assign LUT_1[44629] = 32'b00000000000000001010001010011100;
assign LUT_1[44630] = 32'b00000000000000001100100110110001;
assign LUT_1[44631] = 32'b00000000000000000101111000101101;
assign LUT_1[44632] = 32'b00000000000000001000001100111110;
assign LUT_1[44633] = 32'b00000000000000000001011110111010;
assign LUT_1[44634] = 32'b00000000000000000011111011001111;
assign LUT_1[44635] = 32'b11111111111111111101001101001011;
assign LUT_1[44636] = 32'b00000000000000010000000110010101;
assign LUT_1[44637] = 32'b00000000000000001001011000010001;
assign LUT_1[44638] = 32'b00000000000000001011110100100110;
assign LUT_1[44639] = 32'b00000000000000000101000110100010;
assign LUT_1[44640] = 32'b00000000000000000111111110100110;
assign LUT_1[44641] = 32'b00000000000000000001010000100010;
assign LUT_1[44642] = 32'b00000000000000000011101100110111;
assign LUT_1[44643] = 32'b11111111111111111100111110110011;
assign LUT_1[44644] = 32'b00000000000000001111110111111101;
assign LUT_1[44645] = 32'b00000000000000001001001001111001;
assign LUT_1[44646] = 32'b00000000000000001011100110001110;
assign LUT_1[44647] = 32'b00000000000000000100111000001010;
assign LUT_1[44648] = 32'b00000000000000000111001100011011;
assign LUT_1[44649] = 32'b00000000000000000000011110010111;
assign LUT_1[44650] = 32'b00000000000000000010111010101100;
assign LUT_1[44651] = 32'b11111111111111111100001100101000;
assign LUT_1[44652] = 32'b00000000000000001111000101110010;
assign LUT_1[44653] = 32'b00000000000000001000010111101110;
assign LUT_1[44654] = 32'b00000000000000001010110100000011;
assign LUT_1[44655] = 32'b00000000000000000100000101111111;
assign LUT_1[44656] = 32'b00000000000000001001111010001000;
assign LUT_1[44657] = 32'b00000000000000000011001100000100;
assign LUT_1[44658] = 32'b00000000000000000101101000011001;
assign LUT_1[44659] = 32'b11111111111111111110111010010101;
assign LUT_1[44660] = 32'b00000000000000010001110011011111;
assign LUT_1[44661] = 32'b00000000000000001011000101011011;
assign LUT_1[44662] = 32'b00000000000000001101100001110000;
assign LUT_1[44663] = 32'b00000000000000000110110011101100;
assign LUT_1[44664] = 32'b00000000000000001001000111111101;
assign LUT_1[44665] = 32'b00000000000000000010011001111001;
assign LUT_1[44666] = 32'b00000000000000000100110110001110;
assign LUT_1[44667] = 32'b11111111111111111110001000001010;
assign LUT_1[44668] = 32'b00000000000000010001000001010100;
assign LUT_1[44669] = 32'b00000000000000001010010011010000;
assign LUT_1[44670] = 32'b00000000000000001100101111100101;
assign LUT_1[44671] = 32'b00000000000000000110000001100001;
assign LUT_1[44672] = 32'b00000000000000001000000110000010;
assign LUT_1[44673] = 32'b00000000000000000001010111111110;
assign LUT_1[44674] = 32'b00000000000000000011110100010011;
assign LUT_1[44675] = 32'b11111111111111111101000110001111;
assign LUT_1[44676] = 32'b00000000000000001111111111011001;
assign LUT_1[44677] = 32'b00000000000000001001010001010101;
assign LUT_1[44678] = 32'b00000000000000001011101101101010;
assign LUT_1[44679] = 32'b00000000000000000100111111100110;
assign LUT_1[44680] = 32'b00000000000000000111010011110111;
assign LUT_1[44681] = 32'b00000000000000000000100101110011;
assign LUT_1[44682] = 32'b00000000000000000011000010001000;
assign LUT_1[44683] = 32'b11111111111111111100010100000100;
assign LUT_1[44684] = 32'b00000000000000001111001101001110;
assign LUT_1[44685] = 32'b00000000000000001000011111001010;
assign LUT_1[44686] = 32'b00000000000000001010111011011111;
assign LUT_1[44687] = 32'b00000000000000000100001101011011;
assign LUT_1[44688] = 32'b00000000000000001010000001100100;
assign LUT_1[44689] = 32'b00000000000000000011010011100000;
assign LUT_1[44690] = 32'b00000000000000000101101111110101;
assign LUT_1[44691] = 32'b11111111111111111111000001110001;
assign LUT_1[44692] = 32'b00000000000000010001111010111011;
assign LUT_1[44693] = 32'b00000000000000001011001100110111;
assign LUT_1[44694] = 32'b00000000000000001101101001001100;
assign LUT_1[44695] = 32'b00000000000000000110111011001000;
assign LUT_1[44696] = 32'b00000000000000001001001111011001;
assign LUT_1[44697] = 32'b00000000000000000010100001010101;
assign LUT_1[44698] = 32'b00000000000000000100111101101010;
assign LUT_1[44699] = 32'b11111111111111111110001111100110;
assign LUT_1[44700] = 32'b00000000000000010001001000110000;
assign LUT_1[44701] = 32'b00000000000000001010011010101100;
assign LUT_1[44702] = 32'b00000000000000001100110111000001;
assign LUT_1[44703] = 32'b00000000000000000110001000111101;
assign LUT_1[44704] = 32'b00000000000000001001000001000001;
assign LUT_1[44705] = 32'b00000000000000000010010010111101;
assign LUT_1[44706] = 32'b00000000000000000100101111010010;
assign LUT_1[44707] = 32'b11111111111111111110000001001110;
assign LUT_1[44708] = 32'b00000000000000010000111010011000;
assign LUT_1[44709] = 32'b00000000000000001010001100010100;
assign LUT_1[44710] = 32'b00000000000000001100101000101001;
assign LUT_1[44711] = 32'b00000000000000000101111010100101;
assign LUT_1[44712] = 32'b00000000000000001000001110110110;
assign LUT_1[44713] = 32'b00000000000000000001100000110010;
assign LUT_1[44714] = 32'b00000000000000000011111101000111;
assign LUT_1[44715] = 32'b11111111111111111101001111000011;
assign LUT_1[44716] = 32'b00000000000000010000001000001101;
assign LUT_1[44717] = 32'b00000000000000001001011010001001;
assign LUT_1[44718] = 32'b00000000000000001011110110011110;
assign LUT_1[44719] = 32'b00000000000000000101001000011010;
assign LUT_1[44720] = 32'b00000000000000001010111100100011;
assign LUT_1[44721] = 32'b00000000000000000100001110011111;
assign LUT_1[44722] = 32'b00000000000000000110101010110100;
assign LUT_1[44723] = 32'b11111111111111111111111100110000;
assign LUT_1[44724] = 32'b00000000000000010010110101111010;
assign LUT_1[44725] = 32'b00000000000000001100000111110110;
assign LUT_1[44726] = 32'b00000000000000001110100100001011;
assign LUT_1[44727] = 32'b00000000000000000111110110000111;
assign LUT_1[44728] = 32'b00000000000000001010001010011000;
assign LUT_1[44729] = 32'b00000000000000000011011100010100;
assign LUT_1[44730] = 32'b00000000000000000101111000101001;
assign LUT_1[44731] = 32'b11111111111111111111001010100101;
assign LUT_1[44732] = 32'b00000000000000010010000011101111;
assign LUT_1[44733] = 32'b00000000000000001011010101101011;
assign LUT_1[44734] = 32'b00000000000000001101110010000000;
assign LUT_1[44735] = 32'b00000000000000000111000011111100;
assign LUT_1[44736] = 32'b00000000000000001010000011101010;
assign LUT_1[44737] = 32'b00000000000000000011010101100110;
assign LUT_1[44738] = 32'b00000000000000000101110001111011;
assign LUT_1[44739] = 32'b11111111111111111111000011110111;
assign LUT_1[44740] = 32'b00000000000000010001111101000001;
assign LUT_1[44741] = 32'b00000000000000001011001110111101;
assign LUT_1[44742] = 32'b00000000000000001101101011010010;
assign LUT_1[44743] = 32'b00000000000000000110111101001110;
assign LUT_1[44744] = 32'b00000000000000001001010001011111;
assign LUT_1[44745] = 32'b00000000000000000010100011011011;
assign LUT_1[44746] = 32'b00000000000000000100111111110000;
assign LUT_1[44747] = 32'b11111111111111111110010001101100;
assign LUT_1[44748] = 32'b00000000000000010001001010110110;
assign LUT_1[44749] = 32'b00000000000000001010011100110010;
assign LUT_1[44750] = 32'b00000000000000001100111001000111;
assign LUT_1[44751] = 32'b00000000000000000110001011000011;
assign LUT_1[44752] = 32'b00000000000000001011111111001100;
assign LUT_1[44753] = 32'b00000000000000000101010001001000;
assign LUT_1[44754] = 32'b00000000000000000111101101011101;
assign LUT_1[44755] = 32'b00000000000000000000111111011001;
assign LUT_1[44756] = 32'b00000000000000010011111000100011;
assign LUT_1[44757] = 32'b00000000000000001101001010011111;
assign LUT_1[44758] = 32'b00000000000000001111100110110100;
assign LUT_1[44759] = 32'b00000000000000001000111000110000;
assign LUT_1[44760] = 32'b00000000000000001011001101000001;
assign LUT_1[44761] = 32'b00000000000000000100011110111101;
assign LUT_1[44762] = 32'b00000000000000000110111011010010;
assign LUT_1[44763] = 32'b00000000000000000000001101001110;
assign LUT_1[44764] = 32'b00000000000000010011000110011000;
assign LUT_1[44765] = 32'b00000000000000001100011000010100;
assign LUT_1[44766] = 32'b00000000000000001110110100101001;
assign LUT_1[44767] = 32'b00000000000000001000000110100101;
assign LUT_1[44768] = 32'b00000000000000001010111110101001;
assign LUT_1[44769] = 32'b00000000000000000100010000100101;
assign LUT_1[44770] = 32'b00000000000000000110101100111010;
assign LUT_1[44771] = 32'b11111111111111111111111110110110;
assign LUT_1[44772] = 32'b00000000000000010010111000000000;
assign LUT_1[44773] = 32'b00000000000000001100001001111100;
assign LUT_1[44774] = 32'b00000000000000001110100110010001;
assign LUT_1[44775] = 32'b00000000000000000111111000001101;
assign LUT_1[44776] = 32'b00000000000000001010001100011110;
assign LUT_1[44777] = 32'b00000000000000000011011110011010;
assign LUT_1[44778] = 32'b00000000000000000101111010101111;
assign LUT_1[44779] = 32'b11111111111111111111001100101011;
assign LUT_1[44780] = 32'b00000000000000010010000101110101;
assign LUT_1[44781] = 32'b00000000000000001011010111110001;
assign LUT_1[44782] = 32'b00000000000000001101110100000110;
assign LUT_1[44783] = 32'b00000000000000000111000110000010;
assign LUT_1[44784] = 32'b00000000000000001100111010001011;
assign LUT_1[44785] = 32'b00000000000000000110001100000111;
assign LUT_1[44786] = 32'b00000000000000001000101000011100;
assign LUT_1[44787] = 32'b00000000000000000001111010011000;
assign LUT_1[44788] = 32'b00000000000000010100110011100010;
assign LUT_1[44789] = 32'b00000000000000001110000101011110;
assign LUT_1[44790] = 32'b00000000000000010000100001110011;
assign LUT_1[44791] = 32'b00000000000000001001110011101111;
assign LUT_1[44792] = 32'b00000000000000001100001000000000;
assign LUT_1[44793] = 32'b00000000000000000101011001111100;
assign LUT_1[44794] = 32'b00000000000000000111110110010001;
assign LUT_1[44795] = 32'b00000000000000000001001000001101;
assign LUT_1[44796] = 32'b00000000000000010100000001010111;
assign LUT_1[44797] = 32'b00000000000000001101010011010011;
assign LUT_1[44798] = 32'b00000000000000001111101111101000;
assign LUT_1[44799] = 32'b00000000000000001001000001100100;
assign LUT_1[44800] = 32'b00000000000000000010111010001011;
assign LUT_1[44801] = 32'b11111111111111111100001100000111;
assign LUT_1[44802] = 32'b11111111111111111110101000011100;
assign LUT_1[44803] = 32'b11111111111111110111111010011000;
assign LUT_1[44804] = 32'b00000000000000001010110011100010;
assign LUT_1[44805] = 32'b00000000000000000100000101011110;
assign LUT_1[44806] = 32'b00000000000000000110100001110011;
assign LUT_1[44807] = 32'b11111111111111111111110011101111;
assign LUT_1[44808] = 32'b00000000000000000010001000000000;
assign LUT_1[44809] = 32'b11111111111111111011011001111100;
assign LUT_1[44810] = 32'b11111111111111111101110110010001;
assign LUT_1[44811] = 32'b11111111111111110111001000001101;
assign LUT_1[44812] = 32'b00000000000000001010000001010111;
assign LUT_1[44813] = 32'b00000000000000000011010011010011;
assign LUT_1[44814] = 32'b00000000000000000101101111101000;
assign LUT_1[44815] = 32'b11111111111111111111000001100100;
assign LUT_1[44816] = 32'b00000000000000000100110101101101;
assign LUT_1[44817] = 32'b11111111111111111110000111101001;
assign LUT_1[44818] = 32'b00000000000000000000100011111110;
assign LUT_1[44819] = 32'b11111111111111111001110101111010;
assign LUT_1[44820] = 32'b00000000000000001100101111000100;
assign LUT_1[44821] = 32'b00000000000000000110000001000000;
assign LUT_1[44822] = 32'b00000000000000001000011101010101;
assign LUT_1[44823] = 32'b00000000000000000001101111010001;
assign LUT_1[44824] = 32'b00000000000000000100000011100010;
assign LUT_1[44825] = 32'b11111111111111111101010101011110;
assign LUT_1[44826] = 32'b11111111111111111111110001110011;
assign LUT_1[44827] = 32'b11111111111111111001000011101111;
assign LUT_1[44828] = 32'b00000000000000001011111100111001;
assign LUT_1[44829] = 32'b00000000000000000101001110110101;
assign LUT_1[44830] = 32'b00000000000000000111101011001010;
assign LUT_1[44831] = 32'b00000000000000000000111101000110;
assign LUT_1[44832] = 32'b00000000000000000011110101001010;
assign LUT_1[44833] = 32'b11111111111111111101000111000110;
assign LUT_1[44834] = 32'b11111111111111111111100011011011;
assign LUT_1[44835] = 32'b11111111111111111000110101010111;
assign LUT_1[44836] = 32'b00000000000000001011101110100001;
assign LUT_1[44837] = 32'b00000000000000000101000000011101;
assign LUT_1[44838] = 32'b00000000000000000111011100110010;
assign LUT_1[44839] = 32'b00000000000000000000101110101110;
assign LUT_1[44840] = 32'b00000000000000000011000010111111;
assign LUT_1[44841] = 32'b11111111111111111100010100111011;
assign LUT_1[44842] = 32'b11111111111111111110110001010000;
assign LUT_1[44843] = 32'b11111111111111111000000011001100;
assign LUT_1[44844] = 32'b00000000000000001010111100010110;
assign LUT_1[44845] = 32'b00000000000000000100001110010010;
assign LUT_1[44846] = 32'b00000000000000000110101010100111;
assign LUT_1[44847] = 32'b11111111111111111111111100100011;
assign LUT_1[44848] = 32'b00000000000000000101110000101100;
assign LUT_1[44849] = 32'b11111111111111111111000010101000;
assign LUT_1[44850] = 32'b00000000000000000001011110111101;
assign LUT_1[44851] = 32'b11111111111111111010110000111001;
assign LUT_1[44852] = 32'b00000000000000001101101010000011;
assign LUT_1[44853] = 32'b00000000000000000110111011111111;
assign LUT_1[44854] = 32'b00000000000000001001011000010100;
assign LUT_1[44855] = 32'b00000000000000000010101010010000;
assign LUT_1[44856] = 32'b00000000000000000100111110100001;
assign LUT_1[44857] = 32'b11111111111111111110010000011101;
assign LUT_1[44858] = 32'b00000000000000000000101100110010;
assign LUT_1[44859] = 32'b11111111111111111001111110101110;
assign LUT_1[44860] = 32'b00000000000000001100110111111000;
assign LUT_1[44861] = 32'b00000000000000000110001001110100;
assign LUT_1[44862] = 32'b00000000000000001000100110001001;
assign LUT_1[44863] = 32'b00000000000000000001111000000101;
assign LUT_1[44864] = 32'b00000000000000000100110111110011;
assign LUT_1[44865] = 32'b11111111111111111110001001101111;
assign LUT_1[44866] = 32'b00000000000000000000100110000100;
assign LUT_1[44867] = 32'b11111111111111111001111000000000;
assign LUT_1[44868] = 32'b00000000000000001100110001001010;
assign LUT_1[44869] = 32'b00000000000000000110000011000110;
assign LUT_1[44870] = 32'b00000000000000001000011111011011;
assign LUT_1[44871] = 32'b00000000000000000001110001010111;
assign LUT_1[44872] = 32'b00000000000000000100000101101000;
assign LUT_1[44873] = 32'b11111111111111111101010111100100;
assign LUT_1[44874] = 32'b11111111111111111111110011111001;
assign LUT_1[44875] = 32'b11111111111111111001000101110101;
assign LUT_1[44876] = 32'b00000000000000001011111110111111;
assign LUT_1[44877] = 32'b00000000000000000101010000111011;
assign LUT_1[44878] = 32'b00000000000000000111101101010000;
assign LUT_1[44879] = 32'b00000000000000000000111111001100;
assign LUT_1[44880] = 32'b00000000000000000110110011010101;
assign LUT_1[44881] = 32'b00000000000000000000000101010001;
assign LUT_1[44882] = 32'b00000000000000000010100001100110;
assign LUT_1[44883] = 32'b11111111111111111011110011100010;
assign LUT_1[44884] = 32'b00000000000000001110101100101100;
assign LUT_1[44885] = 32'b00000000000000000111111110101000;
assign LUT_1[44886] = 32'b00000000000000001010011010111101;
assign LUT_1[44887] = 32'b00000000000000000011101100111001;
assign LUT_1[44888] = 32'b00000000000000000110000001001010;
assign LUT_1[44889] = 32'b11111111111111111111010011000110;
assign LUT_1[44890] = 32'b00000000000000000001101111011011;
assign LUT_1[44891] = 32'b11111111111111111011000001010111;
assign LUT_1[44892] = 32'b00000000000000001101111010100001;
assign LUT_1[44893] = 32'b00000000000000000111001100011101;
assign LUT_1[44894] = 32'b00000000000000001001101000110010;
assign LUT_1[44895] = 32'b00000000000000000010111010101110;
assign LUT_1[44896] = 32'b00000000000000000101110010110010;
assign LUT_1[44897] = 32'b11111111111111111111000100101110;
assign LUT_1[44898] = 32'b00000000000000000001100001000011;
assign LUT_1[44899] = 32'b11111111111111111010110010111111;
assign LUT_1[44900] = 32'b00000000000000001101101100001001;
assign LUT_1[44901] = 32'b00000000000000000110111110000101;
assign LUT_1[44902] = 32'b00000000000000001001011010011010;
assign LUT_1[44903] = 32'b00000000000000000010101100010110;
assign LUT_1[44904] = 32'b00000000000000000101000000100111;
assign LUT_1[44905] = 32'b11111111111111111110010010100011;
assign LUT_1[44906] = 32'b00000000000000000000101110111000;
assign LUT_1[44907] = 32'b11111111111111111010000000110100;
assign LUT_1[44908] = 32'b00000000000000001100111001111110;
assign LUT_1[44909] = 32'b00000000000000000110001011111010;
assign LUT_1[44910] = 32'b00000000000000001000101000001111;
assign LUT_1[44911] = 32'b00000000000000000001111010001011;
assign LUT_1[44912] = 32'b00000000000000000111101110010100;
assign LUT_1[44913] = 32'b00000000000000000001000000010000;
assign LUT_1[44914] = 32'b00000000000000000011011100100101;
assign LUT_1[44915] = 32'b11111111111111111100101110100001;
assign LUT_1[44916] = 32'b00000000000000001111100111101011;
assign LUT_1[44917] = 32'b00000000000000001000111001100111;
assign LUT_1[44918] = 32'b00000000000000001011010101111100;
assign LUT_1[44919] = 32'b00000000000000000100100111111000;
assign LUT_1[44920] = 32'b00000000000000000110111100001001;
assign LUT_1[44921] = 32'b00000000000000000000001110000101;
assign LUT_1[44922] = 32'b00000000000000000010101010011010;
assign LUT_1[44923] = 32'b11111111111111111011111100010110;
assign LUT_1[44924] = 32'b00000000000000001110110101100000;
assign LUT_1[44925] = 32'b00000000000000001000000111011100;
assign LUT_1[44926] = 32'b00000000000000001010100011110001;
assign LUT_1[44927] = 32'b00000000000000000011110101101101;
assign LUT_1[44928] = 32'b00000000000000000101111010001110;
assign LUT_1[44929] = 32'b11111111111111111111001100001010;
assign LUT_1[44930] = 32'b00000000000000000001101000011111;
assign LUT_1[44931] = 32'b11111111111111111010111010011011;
assign LUT_1[44932] = 32'b00000000000000001101110011100101;
assign LUT_1[44933] = 32'b00000000000000000111000101100001;
assign LUT_1[44934] = 32'b00000000000000001001100001110110;
assign LUT_1[44935] = 32'b00000000000000000010110011110010;
assign LUT_1[44936] = 32'b00000000000000000101001000000011;
assign LUT_1[44937] = 32'b11111111111111111110011001111111;
assign LUT_1[44938] = 32'b00000000000000000000110110010100;
assign LUT_1[44939] = 32'b11111111111111111010001000010000;
assign LUT_1[44940] = 32'b00000000000000001101000001011010;
assign LUT_1[44941] = 32'b00000000000000000110010011010110;
assign LUT_1[44942] = 32'b00000000000000001000101111101011;
assign LUT_1[44943] = 32'b00000000000000000010000001100111;
assign LUT_1[44944] = 32'b00000000000000000111110101110000;
assign LUT_1[44945] = 32'b00000000000000000001000111101100;
assign LUT_1[44946] = 32'b00000000000000000011100100000001;
assign LUT_1[44947] = 32'b11111111111111111100110101111101;
assign LUT_1[44948] = 32'b00000000000000001111101111000111;
assign LUT_1[44949] = 32'b00000000000000001001000001000011;
assign LUT_1[44950] = 32'b00000000000000001011011101011000;
assign LUT_1[44951] = 32'b00000000000000000100101111010100;
assign LUT_1[44952] = 32'b00000000000000000111000011100101;
assign LUT_1[44953] = 32'b00000000000000000000010101100001;
assign LUT_1[44954] = 32'b00000000000000000010110001110110;
assign LUT_1[44955] = 32'b11111111111111111100000011110010;
assign LUT_1[44956] = 32'b00000000000000001110111100111100;
assign LUT_1[44957] = 32'b00000000000000001000001110111000;
assign LUT_1[44958] = 32'b00000000000000001010101011001101;
assign LUT_1[44959] = 32'b00000000000000000011111101001001;
assign LUT_1[44960] = 32'b00000000000000000110110101001101;
assign LUT_1[44961] = 32'b00000000000000000000000111001001;
assign LUT_1[44962] = 32'b00000000000000000010100011011110;
assign LUT_1[44963] = 32'b11111111111111111011110101011010;
assign LUT_1[44964] = 32'b00000000000000001110101110100100;
assign LUT_1[44965] = 32'b00000000000000001000000000100000;
assign LUT_1[44966] = 32'b00000000000000001010011100110101;
assign LUT_1[44967] = 32'b00000000000000000011101110110001;
assign LUT_1[44968] = 32'b00000000000000000110000011000010;
assign LUT_1[44969] = 32'b11111111111111111111010100111110;
assign LUT_1[44970] = 32'b00000000000000000001110001010011;
assign LUT_1[44971] = 32'b11111111111111111011000011001111;
assign LUT_1[44972] = 32'b00000000000000001101111100011001;
assign LUT_1[44973] = 32'b00000000000000000111001110010101;
assign LUT_1[44974] = 32'b00000000000000001001101010101010;
assign LUT_1[44975] = 32'b00000000000000000010111100100110;
assign LUT_1[44976] = 32'b00000000000000001000110000101111;
assign LUT_1[44977] = 32'b00000000000000000010000010101011;
assign LUT_1[44978] = 32'b00000000000000000100011111000000;
assign LUT_1[44979] = 32'b11111111111111111101110000111100;
assign LUT_1[44980] = 32'b00000000000000010000101010000110;
assign LUT_1[44981] = 32'b00000000000000001001111100000010;
assign LUT_1[44982] = 32'b00000000000000001100011000010111;
assign LUT_1[44983] = 32'b00000000000000000101101010010011;
assign LUT_1[44984] = 32'b00000000000000000111111110100100;
assign LUT_1[44985] = 32'b00000000000000000001010000100000;
assign LUT_1[44986] = 32'b00000000000000000011101100110101;
assign LUT_1[44987] = 32'b11111111111111111100111110110001;
assign LUT_1[44988] = 32'b00000000000000001111110111111011;
assign LUT_1[44989] = 32'b00000000000000001001001001110111;
assign LUT_1[44990] = 32'b00000000000000001011100110001100;
assign LUT_1[44991] = 32'b00000000000000000100111000001000;
assign LUT_1[44992] = 32'b00000000000000000111110111110110;
assign LUT_1[44993] = 32'b00000000000000000001001001110010;
assign LUT_1[44994] = 32'b00000000000000000011100110000111;
assign LUT_1[44995] = 32'b11111111111111111100111000000011;
assign LUT_1[44996] = 32'b00000000000000001111110001001101;
assign LUT_1[44997] = 32'b00000000000000001001000011001001;
assign LUT_1[44998] = 32'b00000000000000001011011111011110;
assign LUT_1[44999] = 32'b00000000000000000100110001011010;
assign LUT_1[45000] = 32'b00000000000000000111000101101011;
assign LUT_1[45001] = 32'b00000000000000000000010111100111;
assign LUT_1[45002] = 32'b00000000000000000010110011111100;
assign LUT_1[45003] = 32'b11111111111111111100000101111000;
assign LUT_1[45004] = 32'b00000000000000001110111111000010;
assign LUT_1[45005] = 32'b00000000000000001000010000111110;
assign LUT_1[45006] = 32'b00000000000000001010101101010011;
assign LUT_1[45007] = 32'b00000000000000000011111111001111;
assign LUT_1[45008] = 32'b00000000000000001001110011011000;
assign LUT_1[45009] = 32'b00000000000000000011000101010100;
assign LUT_1[45010] = 32'b00000000000000000101100001101001;
assign LUT_1[45011] = 32'b11111111111111111110110011100101;
assign LUT_1[45012] = 32'b00000000000000010001101100101111;
assign LUT_1[45013] = 32'b00000000000000001010111110101011;
assign LUT_1[45014] = 32'b00000000000000001101011011000000;
assign LUT_1[45015] = 32'b00000000000000000110101100111100;
assign LUT_1[45016] = 32'b00000000000000001001000001001101;
assign LUT_1[45017] = 32'b00000000000000000010010011001001;
assign LUT_1[45018] = 32'b00000000000000000100101111011110;
assign LUT_1[45019] = 32'b11111111111111111110000001011010;
assign LUT_1[45020] = 32'b00000000000000010000111010100100;
assign LUT_1[45021] = 32'b00000000000000001010001100100000;
assign LUT_1[45022] = 32'b00000000000000001100101000110101;
assign LUT_1[45023] = 32'b00000000000000000101111010110001;
assign LUT_1[45024] = 32'b00000000000000001000110010110101;
assign LUT_1[45025] = 32'b00000000000000000010000100110001;
assign LUT_1[45026] = 32'b00000000000000000100100001000110;
assign LUT_1[45027] = 32'b11111111111111111101110011000010;
assign LUT_1[45028] = 32'b00000000000000010000101100001100;
assign LUT_1[45029] = 32'b00000000000000001001111110001000;
assign LUT_1[45030] = 32'b00000000000000001100011010011101;
assign LUT_1[45031] = 32'b00000000000000000101101100011001;
assign LUT_1[45032] = 32'b00000000000000001000000000101010;
assign LUT_1[45033] = 32'b00000000000000000001010010100110;
assign LUT_1[45034] = 32'b00000000000000000011101110111011;
assign LUT_1[45035] = 32'b11111111111111111101000000110111;
assign LUT_1[45036] = 32'b00000000000000001111111010000001;
assign LUT_1[45037] = 32'b00000000000000001001001011111101;
assign LUT_1[45038] = 32'b00000000000000001011101000010010;
assign LUT_1[45039] = 32'b00000000000000000100111010001110;
assign LUT_1[45040] = 32'b00000000000000001010101110010111;
assign LUT_1[45041] = 32'b00000000000000000100000000010011;
assign LUT_1[45042] = 32'b00000000000000000110011100101000;
assign LUT_1[45043] = 32'b11111111111111111111101110100100;
assign LUT_1[45044] = 32'b00000000000000010010100111101110;
assign LUT_1[45045] = 32'b00000000000000001011111001101010;
assign LUT_1[45046] = 32'b00000000000000001110010101111111;
assign LUT_1[45047] = 32'b00000000000000000111100111111011;
assign LUT_1[45048] = 32'b00000000000000001001111100001100;
assign LUT_1[45049] = 32'b00000000000000000011001110001000;
assign LUT_1[45050] = 32'b00000000000000000101101010011101;
assign LUT_1[45051] = 32'b11111111111111111110111100011001;
assign LUT_1[45052] = 32'b00000000000000010001110101100011;
assign LUT_1[45053] = 32'b00000000000000001011000111011111;
assign LUT_1[45054] = 32'b00000000000000001101100011110100;
assign LUT_1[45055] = 32'b00000000000000000110110101110000;
assign LUT_1[45056] = 32'b00000000000000000011110011111101;
assign LUT_1[45057] = 32'b11111111111111111101000101111001;
assign LUT_1[45058] = 32'b11111111111111111111100010001110;
assign LUT_1[45059] = 32'b11111111111111111000110100001010;
assign LUT_1[45060] = 32'b00000000000000001011101101010100;
assign LUT_1[45061] = 32'b00000000000000000100111111010000;
assign LUT_1[45062] = 32'b00000000000000000111011011100101;
assign LUT_1[45063] = 32'b00000000000000000000101101100001;
assign LUT_1[45064] = 32'b00000000000000000011000001110010;
assign LUT_1[45065] = 32'b11111111111111111100010011101110;
assign LUT_1[45066] = 32'b11111111111111111110110000000011;
assign LUT_1[45067] = 32'b11111111111111111000000001111111;
assign LUT_1[45068] = 32'b00000000000000001010111011001001;
assign LUT_1[45069] = 32'b00000000000000000100001101000101;
assign LUT_1[45070] = 32'b00000000000000000110101001011010;
assign LUT_1[45071] = 32'b11111111111111111111111011010110;
assign LUT_1[45072] = 32'b00000000000000000101101111011111;
assign LUT_1[45073] = 32'b11111111111111111111000001011011;
assign LUT_1[45074] = 32'b00000000000000000001011101110000;
assign LUT_1[45075] = 32'b11111111111111111010101111101100;
assign LUT_1[45076] = 32'b00000000000000001101101000110110;
assign LUT_1[45077] = 32'b00000000000000000110111010110010;
assign LUT_1[45078] = 32'b00000000000000001001010111000111;
assign LUT_1[45079] = 32'b00000000000000000010101001000011;
assign LUT_1[45080] = 32'b00000000000000000100111101010100;
assign LUT_1[45081] = 32'b11111111111111111110001111010000;
assign LUT_1[45082] = 32'b00000000000000000000101011100101;
assign LUT_1[45083] = 32'b11111111111111111001111101100001;
assign LUT_1[45084] = 32'b00000000000000001100110110101011;
assign LUT_1[45085] = 32'b00000000000000000110001000100111;
assign LUT_1[45086] = 32'b00000000000000001000100100111100;
assign LUT_1[45087] = 32'b00000000000000000001110110111000;
assign LUT_1[45088] = 32'b00000000000000000100101110111100;
assign LUT_1[45089] = 32'b11111111111111111110000000111000;
assign LUT_1[45090] = 32'b00000000000000000000011101001101;
assign LUT_1[45091] = 32'b11111111111111111001101111001001;
assign LUT_1[45092] = 32'b00000000000000001100101000010011;
assign LUT_1[45093] = 32'b00000000000000000101111010001111;
assign LUT_1[45094] = 32'b00000000000000001000010110100100;
assign LUT_1[45095] = 32'b00000000000000000001101000100000;
assign LUT_1[45096] = 32'b00000000000000000011111100110001;
assign LUT_1[45097] = 32'b11111111111111111101001110101101;
assign LUT_1[45098] = 32'b11111111111111111111101011000010;
assign LUT_1[45099] = 32'b11111111111111111000111100111110;
assign LUT_1[45100] = 32'b00000000000000001011110110001000;
assign LUT_1[45101] = 32'b00000000000000000101001000000100;
assign LUT_1[45102] = 32'b00000000000000000111100100011001;
assign LUT_1[45103] = 32'b00000000000000000000110110010101;
assign LUT_1[45104] = 32'b00000000000000000110101010011110;
assign LUT_1[45105] = 32'b11111111111111111111111100011010;
assign LUT_1[45106] = 32'b00000000000000000010011000101111;
assign LUT_1[45107] = 32'b11111111111111111011101010101011;
assign LUT_1[45108] = 32'b00000000000000001110100011110101;
assign LUT_1[45109] = 32'b00000000000000000111110101110001;
assign LUT_1[45110] = 32'b00000000000000001010010010000110;
assign LUT_1[45111] = 32'b00000000000000000011100100000010;
assign LUT_1[45112] = 32'b00000000000000000101111000010011;
assign LUT_1[45113] = 32'b11111111111111111111001010001111;
assign LUT_1[45114] = 32'b00000000000000000001100110100100;
assign LUT_1[45115] = 32'b11111111111111111010111000100000;
assign LUT_1[45116] = 32'b00000000000000001101110001101010;
assign LUT_1[45117] = 32'b00000000000000000111000011100110;
assign LUT_1[45118] = 32'b00000000000000001001011111111011;
assign LUT_1[45119] = 32'b00000000000000000010110001110111;
assign LUT_1[45120] = 32'b00000000000000000101110001100101;
assign LUT_1[45121] = 32'b11111111111111111111000011100001;
assign LUT_1[45122] = 32'b00000000000000000001011111110110;
assign LUT_1[45123] = 32'b11111111111111111010110001110010;
assign LUT_1[45124] = 32'b00000000000000001101101010111100;
assign LUT_1[45125] = 32'b00000000000000000110111100111000;
assign LUT_1[45126] = 32'b00000000000000001001011001001101;
assign LUT_1[45127] = 32'b00000000000000000010101011001001;
assign LUT_1[45128] = 32'b00000000000000000100111111011010;
assign LUT_1[45129] = 32'b11111111111111111110010001010110;
assign LUT_1[45130] = 32'b00000000000000000000101101101011;
assign LUT_1[45131] = 32'b11111111111111111001111111100111;
assign LUT_1[45132] = 32'b00000000000000001100111000110001;
assign LUT_1[45133] = 32'b00000000000000000110001010101101;
assign LUT_1[45134] = 32'b00000000000000001000100111000010;
assign LUT_1[45135] = 32'b00000000000000000001111000111110;
assign LUT_1[45136] = 32'b00000000000000000111101101000111;
assign LUT_1[45137] = 32'b00000000000000000000111111000011;
assign LUT_1[45138] = 32'b00000000000000000011011011011000;
assign LUT_1[45139] = 32'b11111111111111111100101101010100;
assign LUT_1[45140] = 32'b00000000000000001111100110011110;
assign LUT_1[45141] = 32'b00000000000000001000111000011010;
assign LUT_1[45142] = 32'b00000000000000001011010100101111;
assign LUT_1[45143] = 32'b00000000000000000100100110101011;
assign LUT_1[45144] = 32'b00000000000000000110111010111100;
assign LUT_1[45145] = 32'b00000000000000000000001100111000;
assign LUT_1[45146] = 32'b00000000000000000010101001001101;
assign LUT_1[45147] = 32'b11111111111111111011111011001001;
assign LUT_1[45148] = 32'b00000000000000001110110100010011;
assign LUT_1[45149] = 32'b00000000000000001000000110001111;
assign LUT_1[45150] = 32'b00000000000000001010100010100100;
assign LUT_1[45151] = 32'b00000000000000000011110100100000;
assign LUT_1[45152] = 32'b00000000000000000110101100100100;
assign LUT_1[45153] = 32'b11111111111111111111111110100000;
assign LUT_1[45154] = 32'b00000000000000000010011010110101;
assign LUT_1[45155] = 32'b11111111111111111011101100110001;
assign LUT_1[45156] = 32'b00000000000000001110100101111011;
assign LUT_1[45157] = 32'b00000000000000000111110111110111;
assign LUT_1[45158] = 32'b00000000000000001010010100001100;
assign LUT_1[45159] = 32'b00000000000000000011100110001000;
assign LUT_1[45160] = 32'b00000000000000000101111010011001;
assign LUT_1[45161] = 32'b11111111111111111111001100010101;
assign LUT_1[45162] = 32'b00000000000000000001101000101010;
assign LUT_1[45163] = 32'b11111111111111111010111010100110;
assign LUT_1[45164] = 32'b00000000000000001101110011110000;
assign LUT_1[45165] = 32'b00000000000000000111000101101100;
assign LUT_1[45166] = 32'b00000000000000001001100010000001;
assign LUT_1[45167] = 32'b00000000000000000010110011111101;
assign LUT_1[45168] = 32'b00000000000000001000101000000110;
assign LUT_1[45169] = 32'b00000000000000000001111010000010;
assign LUT_1[45170] = 32'b00000000000000000100010110010111;
assign LUT_1[45171] = 32'b11111111111111111101101000010011;
assign LUT_1[45172] = 32'b00000000000000010000100001011101;
assign LUT_1[45173] = 32'b00000000000000001001110011011001;
assign LUT_1[45174] = 32'b00000000000000001100001111101110;
assign LUT_1[45175] = 32'b00000000000000000101100001101010;
assign LUT_1[45176] = 32'b00000000000000000111110101111011;
assign LUT_1[45177] = 32'b00000000000000000001000111110111;
assign LUT_1[45178] = 32'b00000000000000000011100100001100;
assign LUT_1[45179] = 32'b11111111111111111100110110001000;
assign LUT_1[45180] = 32'b00000000000000001111101111010010;
assign LUT_1[45181] = 32'b00000000000000001001000001001110;
assign LUT_1[45182] = 32'b00000000000000001011011101100011;
assign LUT_1[45183] = 32'b00000000000000000100101111011111;
assign LUT_1[45184] = 32'b00000000000000000110110100000000;
assign LUT_1[45185] = 32'b00000000000000000000000101111100;
assign LUT_1[45186] = 32'b00000000000000000010100010010001;
assign LUT_1[45187] = 32'b11111111111111111011110100001101;
assign LUT_1[45188] = 32'b00000000000000001110101101010111;
assign LUT_1[45189] = 32'b00000000000000000111111111010011;
assign LUT_1[45190] = 32'b00000000000000001010011011101000;
assign LUT_1[45191] = 32'b00000000000000000011101101100100;
assign LUT_1[45192] = 32'b00000000000000000110000001110101;
assign LUT_1[45193] = 32'b11111111111111111111010011110001;
assign LUT_1[45194] = 32'b00000000000000000001110000000110;
assign LUT_1[45195] = 32'b11111111111111111011000010000010;
assign LUT_1[45196] = 32'b00000000000000001101111011001100;
assign LUT_1[45197] = 32'b00000000000000000111001101001000;
assign LUT_1[45198] = 32'b00000000000000001001101001011101;
assign LUT_1[45199] = 32'b00000000000000000010111011011001;
assign LUT_1[45200] = 32'b00000000000000001000101111100010;
assign LUT_1[45201] = 32'b00000000000000000010000001011110;
assign LUT_1[45202] = 32'b00000000000000000100011101110011;
assign LUT_1[45203] = 32'b11111111111111111101101111101111;
assign LUT_1[45204] = 32'b00000000000000010000101000111001;
assign LUT_1[45205] = 32'b00000000000000001001111010110101;
assign LUT_1[45206] = 32'b00000000000000001100010111001010;
assign LUT_1[45207] = 32'b00000000000000000101101001000110;
assign LUT_1[45208] = 32'b00000000000000000111111101010111;
assign LUT_1[45209] = 32'b00000000000000000001001111010011;
assign LUT_1[45210] = 32'b00000000000000000011101011101000;
assign LUT_1[45211] = 32'b11111111111111111100111101100100;
assign LUT_1[45212] = 32'b00000000000000001111110110101110;
assign LUT_1[45213] = 32'b00000000000000001001001000101010;
assign LUT_1[45214] = 32'b00000000000000001011100100111111;
assign LUT_1[45215] = 32'b00000000000000000100110110111011;
assign LUT_1[45216] = 32'b00000000000000000111101110111111;
assign LUT_1[45217] = 32'b00000000000000000001000000111011;
assign LUT_1[45218] = 32'b00000000000000000011011101010000;
assign LUT_1[45219] = 32'b11111111111111111100101111001100;
assign LUT_1[45220] = 32'b00000000000000001111101000010110;
assign LUT_1[45221] = 32'b00000000000000001000111010010010;
assign LUT_1[45222] = 32'b00000000000000001011010110100111;
assign LUT_1[45223] = 32'b00000000000000000100101000100011;
assign LUT_1[45224] = 32'b00000000000000000110111100110100;
assign LUT_1[45225] = 32'b00000000000000000000001110110000;
assign LUT_1[45226] = 32'b00000000000000000010101011000101;
assign LUT_1[45227] = 32'b11111111111111111011111101000001;
assign LUT_1[45228] = 32'b00000000000000001110110110001011;
assign LUT_1[45229] = 32'b00000000000000001000001000000111;
assign LUT_1[45230] = 32'b00000000000000001010100100011100;
assign LUT_1[45231] = 32'b00000000000000000011110110011000;
assign LUT_1[45232] = 32'b00000000000000001001101010100001;
assign LUT_1[45233] = 32'b00000000000000000010111100011101;
assign LUT_1[45234] = 32'b00000000000000000101011000110010;
assign LUT_1[45235] = 32'b11111111111111111110101010101110;
assign LUT_1[45236] = 32'b00000000000000010001100011111000;
assign LUT_1[45237] = 32'b00000000000000001010110101110100;
assign LUT_1[45238] = 32'b00000000000000001101010010001001;
assign LUT_1[45239] = 32'b00000000000000000110100100000101;
assign LUT_1[45240] = 32'b00000000000000001000111000010110;
assign LUT_1[45241] = 32'b00000000000000000010001010010010;
assign LUT_1[45242] = 32'b00000000000000000100100110100111;
assign LUT_1[45243] = 32'b11111111111111111101111000100011;
assign LUT_1[45244] = 32'b00000000000000010000110001101101;
assign LUT_1[45245] = 32'b00000000000000001010000011101001;
assign LUT_1[45246] = 32'b00000000000000001100011111111110;
assign LUT_1[45247] = 32'b00000000000000000101110001111010;
assign LUT_1[45248] = 32'b00000000000000001000110001101000;
assign LUT_1[45249] = 32'b00000000000000000010000011100100;
assign LUT_1[45250] = 32'b00000000000000000100011111111001;
assign LUT_1[45251] = 32'b11111111111111111101110001110101;
assign LUT_1[45252] = 32'b00000000000000010000101010111111;
assign LUT_1[45253] = 32'b00000000000000001001111100111011;
assign LUT_1[45254] = 32'b00000000000000001100011001010000;
assign LUT_1[45255] = 32'b00000000000000000101101011001100;
assign LUT_1[45256] = 32'b00000000000000000111111111011101;
assign LUT_1[45257] = 32'b00000000000000000001010001011001;
assign LUT_1[45258] = 32'b00000000000000000011101101101110;
assign LUT_1[45259] = 32'b11111111111111111100111111101010;
assign LUT_1[45260] = 32'b00000000000000001111111000110100;
assign LUT_1[45261] = 32'b00000000000000001001001010110000;
assign LUT_1[45262] = 32'b00000000000000001011100111000101;
assign LUT_1[45263] = 32'b00000000000000000100111001000001;
assign LUT_1[45264] = 32'b00000000000000001010101101001010;
assign LUT_1[45265] = 32'b00000000000000000011111111000110;
assign LUT_1[45266] = 32'b00000000000000000110011011011011;
assign LUT_1[45267] = 32'b11111111111111111111101101010111;
assign LUT_1[45268] = 32'b00000000000000010010100110100001;
assign LUT_1[45269] = 32'b00000000000000001011111000011101;
assign LUT_1[45270] = 32'b00000000000000001110010100110010;
assign LUT_1[45271] = 32'b00000000000000000111100110101110;
assign LUT_1[45272] = 32'b00000000000000001001111010111111;
assign LUT_1[45273] = 32'b00000000000000000011001100111011;
assign LUT_1[45274] = 32'b00000000000000000101101001010000;
assign LUT_1[45275] = 32'b11111111111111111110111011001100;
assign LUT_1[45276] = 32'b00000000000000010001110100010110;
assign LUT_1[45277] = 32'b00000000000000001011000110010010;
assign LUT_1[45278] = 32'b00000000000000001101100010100111;
assign LUT_1[45279] = 32'b00000000000000000110110100100011;
assign LUT_1[45280] = 32'b00000000000000001001101100100111;
assign LUT_1[45281] = 32'b00000000000000000010111110100011;
assign LUT_1[45282] = 32'b00000000000000000101011010111000;
assign LUT_1[45283] = 32'b11111111111111111110101100110100;
assign LUT_1[45284] = 32'b00000000000000010001100101111110;
assign LUT_1[45285] = 32'b00000000000000001010110111111010;
assign LUT_1[45286] = 32'b00000000000000001101010100001111;
assign LUT_1[45287] = 32'b00000000000000000110100110001011;
assign LUT_1[45288] = 32'b00000000000000001000111010011100;
assign LUT_1[45289] = 32'b00000000000000000010001100011000;
assign LUT_1[45290] = 32'b00000000000000000100101000101101;
assign LUT_1[45291] = 32'b11111111111111111101111010101001;
assign LUT_1[45292] = 32'b00000000000000010000110011110011;
assign LUT_1[45293] = 32'b00000000000000001010000101101111;
assign LUT_1[45294] = 32'b00000000000000001100100010000100;
assign LUT_1[45295] = 32'b00000000000000000101110100000000;
assign LUT_1[45296] = 32'b00000000000000001011101000001001;
assign LUT_1[45297] = 32'b00000000000000000100111010000101;
assign LUT_1[45298] = 32'b00000000000000000111010110011010;
assign LUT_1[45299] = 32'b00000000000000000000101000010110;
assign LUT_1[45300] = 32'b00000000000000010011100001100000;
assign LUT_1[45301] = 32'b00000000000000001100110011011100;
assign LUT_1[45302] = 32'b00000000000000001111001111110001;
assign LUT_1[45303] = 32'b00000000000000001000100001101101;
assign LUT_1[45304] = 32'b00000000000000001010110101111110;
assign LUT_1[45305] = 32'b00000000000000000100000111111010;
assign LUT_1[45306] = 32'b00000000000000000110100100001111;
assign LUT_1[45307] = 32'b11111111111111111111110110001011;
assign LUT_1[45308] = 32'b00000000000000010010101111010101;
assign LUT_1[45309] = 32'b00000000000000001100000001010001;
assign LUT_1[45310] = 32'b00000000000000001110011101100110;
assign LUT_1[45311] = 32'b00000000000000000111101111100010;
assign LUT_1[45312] = 32'b00000000000000000001101000001001;
assign LUT_1[45313] = 32'b11111111111111111010111010000101;
assign LUT_1[45314] = 32'b11111111111111111101010110011010;
assign LUT_1[45315] = 32'b11111111111111110110101000010110;
assign LUT_1[45316] = 32'b00000000000000001001100001100000;
assign LUT_1[45317] = 32'b00000000000000000010110011011100;
assign LUT_1[45318] = 32'b00000000000000000101001111110001;
assign LUT_1[45319] = 32'b11111111111111111110100001101101;
assign LUT_1[45320] = 32'b00000000000000000000110101111110;
assign LUT_1[45321] = 32'b11111111111111111010000111111010;
assign LUT_1[45322] = 32'b11111111111111111100100100001111;
assign LUT_1[45323] = 32'b11111111111111110101110110001011;
assign LUT_1[45324] = 32'b00000000000000001000101111010101;
assign LUT_1[45325] = 32'b00000000000000000010000001010001;
assign LUT_1[45326] = 32'b00000000000000000100011101100110;
assign LUT_1[45327] = 32'b11111111111111111101101111100010;
assign LUT_1[45328] = 32'b00000000000000000011100011101011;
assign LUT_1[45329] = 32'b11111111111111111100110101100111;
assign LUT_1[45330] = 32'b11111111111111111111010001111100;
assign LUT_1[45331] = 32'b11111111111111111000100011111000;
assign LUT_1[45332] = 32'b00000000000000001011011101000010;
assign LUT_1[45333] = 32'b00000000000000000100101110111110;
assign LUT_1[45334] = 32'b00000000000000000111001011010011;
assign LUT_1[45335] = 32'b00000000000000000000011101001111;
assign LUT_1[45336] = 32'b00000000000000000010110001100000;
assign LUT_1[45337] = 32'b11111111111111111100000011011100;
assign LUT_1[45338] = 32'b11111111111111111110011111110001;
assign LUT_1[45339] = 32'b11111111111111110111110001101101;
assign LUT_1[45340] = 32'b00000000000000001010101010110111;
assign LUT_1[45341] = 32'b00000000000000000011111100110011;
assign LUT_1[45342] = 32'b00000000000000000110011001001000;
assign LUT_1[45343] = 32'b11111111111111111111101011000100;
assign LUT_1[45344] = 32'b00000000000000000010100011001000;
assign LUT_1[45345] = 32'b11111111111111111011110101000100;
assign LUT_1[45346] = 32'b11111111111111111110010001011001;
assign LUT_1[45347] = 32'b11111111111111110111100011010101;
assign LUT_1[45348] = 32'b00000000000000001010011100011111;
assign LUT_1[45349] = 32'b00000000000000000011101110011011;
assign LUT_1[45350] = 32'b00000000000000000110001010110000;
assign LUT_1[45351] = 32'b11111111111111111111011100101100;
assign LUT_1[45352] = 32'b00000000000000000001110000111101;
assign LUT_1[45353] = 32'b11111111111111111011000010111001;
assign LUT_1[45354] = 32'b11111111111111111101011111001110;
assign LUT_1[45355] = 32'b11111111111111110110110001001010;
assign LUT_1[45356] = 32'b00000000000000001001101010010100;
assign LUT_1[45357] = 32'b00000000000000000010111100010000;
assign LUT_1[45358] = 32'b00000000000000000101011000100101;
assign LUT_1[45359] = 32'b11111111111111111110101010100001;
assign LUT_1[45360] = 32'b00000000000000000100011110101010;
assign LUT_1[45361] = 32'b11111111111111111101110000100110;
assign LUT_1[45362] = 32'b00000000000000000000001100111011;
assign LUT_1[45363] = 32'b11111111111111111001011110110111;
assign LUT_1[45364] = 32'b00000000000000001100011000000001;
assign LUT_1[45365] = 32'b00000000000000000101101001111101;
assign LUT_1[45366] = 32'b00000000000000001000000110010010;
assign LUT_1[45367] = 32'b00000000000000000001011000001110;
assign LUT_1[45368] = 32'b00000000000000000011101100011111;
assign LUT_1[45369] = 32'b11111111111111111100111110011011;
assign LUT_1[45370] = 32'b11111111111111111111011010110000;
assign LUT_1[45371] = 32'b11111111111111111000101100101100;
assign LUT_1[45372] = 32'b00000000000000001011100101110110;
assign LUT_1[45373] = 32'b00000000000000000100110111110010;
assign LUT_1[45374] = 32'b00000000000000000111010100000111;
assign LUT_1[45375] = 32'b00000000000000000000100110000011;
assign LUT_1[45376] = 32'b00000000000000000011100101110001;
assign LUT_1[45377] = 32'b11111111111111111100110111101101;
assign LUT_1[45378] = 32'b11111111111111111111010100000010;
assign LUT_1[45379] = 32'b11111111111111111000100101111110;
assign LUT_1[45380] = 32'b00000000000000001011011111001000;
assign LUT_1[45381] = 32'b00000000000000000100110001000100;
assign LUT_1[45382] = 32'b00000000000000000111001101011001;
assign LUT_1[45383] = 32'b00000000000000000000011111010101;
assign LUT_1[45384] = 32'b00000000000000000010110011100110;
assign LUT_1[45385] = 32'b11111111111111111100000101100010;
assign LUT_1[45386] = 32'b11111111111111111110100001110111;
assign LUT_1[45387] = 32'b11111111111111110111110011110011;
assign LUT_1[45388] = 32'b00000000000000001010101100111101;
assign LUT_1[45389] = 32'b00000000000000000011111110111001;
assign LUT_1[45390] = 32'b00000000000000000110011011001110;
assign LUT_1[45391] = 32'b11111111111111111111101101001010;
assign LUT_1[45392] = 32'b00000000000000000101100001010011;
assign LUT_1[45393] = 32'b11111111111111111110110011001111;
assign LUT_1[45394] = 32'b00000000000000000001001111100100;
assign LUT_1[45395] = 32'b11111111111111111010100001100000;
assign LUT_1[45396] = 32'b00000000000000001101011010101010;
assign LUT_1[45397] = 32'b00000000000000000110101100100110;
assign LUT_1[45398] = 32'b00000000000000001001001000111011;
assign LUT_1[45399] = 32'b00000000000000000010011010110111;
assign LUT_1[45400] = 32'b00000000000000000100101111001000;
assign LUT_1[45401] = 32'b11111111111111111110000001000100;
assign LUT_1[45402] = 32'b00000000000000000000011101011001;
assign LUT_1[45403] = 32'b11111111111111111001101111010101;
assign LUT_1[45404] = 32'b00000000000000001100101000011111;
assign LUT_1[45405] = 32'b00000000000000000101111010011011;
assign LUT_1[45406] = 32'b00000000000000001000010110110000;
assign LUT_1[45407] = 32'b00000000000000000001101000101100;
assign LUT_1[45408] = 32'b00000000000000000100100000110000;
assign LUT_1[45409] = 32'b11111111111111111101110010101100;
assign LUT_1[45410] = 32'b00000000000000000000001111000001;
assign LUT_1[45411] = 32'b11111111111111111001100000111101;
assign LUT_1[45412] = 32'b00000000000000001100011010000111;
assign LUT_1[45413] = 32'b00000000000000000101101100000011;
assign LUT_1[45414] = 32'b00000000000000001000001000011000;
assign LUT_1[45415] = 32'b00000000000000000001011010010100;
assign LUT_1[45416] = 32'b00000000000000000011101110100101;
assign LUT_1[45417] = 32'b11111111111111111101000000100001;
assign LUT_1[45418] = 32'b11111111111111111111011100110110;
assign LUT_1[45419] = 32'b11111111111111111000101110110010;
assign LUT_1[45420] = 32'b00000000000000001011100111111100;
assign LUT_1[45421] = 32'b00000000000000000100111001111000;
assign LUT_1[45422] = 32'b00000000000000000111010110001101;
assign LUT_1[45423] = 32'b00000000000000000000101000001001;
assign LUT_1[45424] = 32'b00000000000000000110011100010010;
assign LUT_1[45425] = 32'b11111111111111111111101110001110;
assign LUT_1[45426] = 32'b00000000000000000010001010100011;
assign LUT_1[45427] = 32'b11111111111111111011011100011111;
assign LUT_1[45428] = 32'b00000000000000001110010101101001;
assign LUT_1[45429] = 32'b00000000000000000111100111100101;
assign LUT_1[45430] = 32'b00000000000000001010000011111010;
assign LUT_1[45431] = 32'b00000000000000000011010101110110;
assign LUT_1[45432] = 32'b00000000000000000101101010000111;
assign LUT_1[45433] = 32'b11111111111111111110111100000011;
assign LUT_1[45434] = 32'b00000000000000000001011000011000;
assign LUT_1[45435] = 32'b11111111111111111010101010010100;
assign LUT_1[45436] = 32'b00000000000000001101100011011110;
assign LUT_1[45437] = 32'b00000000000000000110110101011010;
assign LUT_1[45438] = 32'b00000000000000001001010001101111;
assign LUT_1[45439] = 32'b00000000000000000010100011101011;
assign LUT_1[45440] = 32'b00000000000000000100101000001100;
assign LUT_1[45441] = 32'b11111111111111111101111010001000;
assign LUT_1[45442] = 32'b00000000000000000000010110011101;
assign LUT_1[45443] = 32'b11111111111111111001101000011001;
assign LUT_1[45444] = 32'b00000000000000001100100001100011;
assign LUT_1[45445] = 32'b00000000000000000101110011011111;
assign LUT_1[45446] = 32'b00000000000000001000001111110100;
assign LUT_1[45447] = 32'b00000000000000000001100001110000;
assign LUT_1[45448] = 32'b00000000000000000011110110000001;
assign LUT_1[45449] = 32'b11111111111111111101000111111101;
assign LUT_1[45450] = 32'b11111111111111111111100100010010;
assign LUT_1[45451] = 32'b11111111111111111000110110001110;
assign LUT_1[45452] = 32'b00000000000000001011101111011000;
assign LUT_1[45453] = 32'b00000000000000000101000001010100;
assign LUT_1[45454] = 32'b00000000000000000111011101101001;
assign LUT_1[45455] = 32'b00000000000000000000101111100101;
assign LUT_1[45456] = 32'b00000000000000000110100011101110;
assign LUT_1[45457] = 32'b11111111111111111111110101101010;
assign LUT_1[45458] = 32'b00000000000000000010010001111111;
assign LUT_1[45459] = 32'b11111111111111111011100011111011;
assign LUT_1[45460] = 32'b00000000000000001110011101000101;
assign LUT_1[45461] = 32'b00000000000000000111101111000001;
assign LUT_1[45462] = 32'b00000000000000001010001011010110;
assign LUT_1[45463] = 32'b00000000000000000011011101010010;
assign LUT_1[45464] = 32'b00000000000000000101110001100011;
assign LUT_1[45465] = 32'b11111111111111111111000011011111;
assign LUT_1[45466] = 32'b00000000000000000001011111110100;
assign LUT_1[45467] = 32'b11111111111111111010110001110000;
assign LUT_1[45468] = 32'b00000000000000001101101010111010;
assign LUT_1[45469] = 32'b00000000000000000110111100110110;
assign LUT_1[45470] = 32'b00000000000000001001011001001011;
assign LUT_1[45471] = 32'b00000000000000000010101011000111;
assign LUT_1[45472] = 32'b00000000000000000101100011001011;
assign LUT_1[45473] = 32'b11111111111111111110110101000111;
assign LUT_1[45474] = 32'b00000000000000000001010001011100;
assign LUT_1[45475] = 32'b11111111111111111010100011011000;
assign LUT_1[45476] = 32'b00000000000000001101011100100010;
assign LUT_1[45477] = 32'b00000000000000000110101110011110;
assign LUT_1[45478] = 32'b00000000000000001001001010110011;
assign LUT_1[45479] = 32'b00000000000000000010011100101111;
assign LUT_1[45480] = 32'b00000000000000000100110001000000;
assign LUT_1[45481] = 32'b11111111111111111110000010111100;
assign LUT_1[45482] = 32'b00000000000000000000011111010001;
assign LUT_1[45483] = 32'b11111111111111111001110001001101;
assign LUT_1[45484] = 32'b00000000000000001100101010010111;
assign LUT_1[45485] = 32'b00000000000000000101111100010011;
assign LUT_1[45486] = 32'b00000000000000001000011000101000;
assign LUT_1[45487] = 32'b00000000000000000001101010100100;
assign LUT_1[45488] = 32'b00000000000000000111011110101101;
assign LUT_1[45489] = 32'b00000000000000000000110000101001;
assign LUT_1[45490] = 32'b00000000000000000011001100111110;
assign LUT_1[45491] = 32'b11111111111111111100011110111010;
assign LUT_1[45492] = 32'b00000000000000001111011000000100;
assign LUT_1[45493] = 32'b00000000000000001000101010000000;
assign LUT_1[45494] = 32'b00000000000000001011000110010101;
assign LUT_1[45495] = 32'b00000000000000000100011000010001;
assign LUT_1[45496] = 32'b00000000000000000110101100100010;
assign LUT_1[45497] = 32'b11111111111111111111111110011110;
assign LUT_1[45498] = 32'b00000000000000000010011010110011;
assign LUT_1[45499] = 32'b11111111111111111011101100101111;
assign LUT_1[45500] = 32'b00000000000000001110100101111001;
assign LUT_1[45501] = 32'b00000000000000000111110111110101;
assign LUT_1[45502] = 32'b00000000000000001010010100001010;
assign LUT_1[45503] = 32'b00000000000000000011100110000110;
assign LUT_1[45504] = 32'b00000000000000000110100101110100;
assign LUT_1[45505] = 32'b11111111111111111111110111110000;
assign LUT_1[45506] = 32'b00000000000000000010010100000101;
assign LUT_1[45507] = 32'b11111111111111111011100110000001;
assign LUT_1[45508] = 32'b00000000000000001110011111001011;
assign LUT_1[45509] = 32'b00000000000000000111110001000111;
assign LUT_1[45510] = 32'b00000000000000001010001101011100;
assign LUT_1[45511] = 32'b00000000000000000011011111011000;
assign LUT_1[45512] = 32'b00000000000000000101110011101001;
assign LUT_1[45513] = 32'b11111111111111111111000101100101;
assign LUT_1[45514] = 32'b00000000000000000001100001111010;
assign LUT_1[45515] = 32'b11111111111111111010110011110110;
assign LUT_1[45516] = 32'b00000000000000001101101101000000;
assign LUT_1[45517] = 32'b00000000000000000110111110111100;
assign LUT_1[45518] = 32'b00000000000000001001011011010001;
assign LUT_1[45519] = 32'b00000000000000000010101101001101;
assign LUT_1[45520] = 32'b00000000000000001000100001010110;
assign LUT_1[45521] = 32'b00000000000000000001110011010010;
assign LUT_1[45522] = 32'b00000000000000000100001111100111;
assign LUT_1[45523] = 32'b11111111111111111101100001100011;
assign LUT_1[45524] = 32'b00000000000000010000011010101101;
assign LUT_1[45525] = 32'b00000000000000001001101100101001;
assign LUT_1[45526] = 32'b00000000000000001100001000111110;
assign LUT_1[45527] = 32'b00000000000000000101011010111010;
assign LUT_1[45528] = 32'b00000000000000000111101111001011;
assign LUT_1[45529] = 32'b00000000000000000001000001000111;
assign LUT_1[45530] = 32'b00000000000000000011011101011100;
assign LUT_1[45531] = 32'b11111111111111111100101111011000;
assign LUT_1[45532] = 32'b00000000000000001111101000100010;
assign LUT_1[45533] = 32'b00000000000000001000111010011110;
assign LUT_1[45534] = 32'b00000000000000001011010110110011;
assign LUT_1[45535] = 32'b00000000000000000100101000101111;
assign LUT_1[45536] = 32'b00000000000000000111100000110011;
assign LUT_1[45537] = 32'b00000000000000000000110010101111;
assign LUT_1[45538] = 32'b00000000000000000011001111000100;
assign LUT_1[45539] = 32'b11111111111111111100100001000000;
assign LUT_1[45540] = 32'b00000000000000001111011010001010;
assign LUT_1[45541] = 32'b00000000000000001000101100000110;
assign LUT_1[45542] = 32'b00000000000000001011001000011011;
assign LUT_1[45543] = 32'b00000000000000000100011010010111;
assign LUT_1[45544] = 32'b00000000000000000110101110101000;
assign LUT_1[45545] = 32'b00000000000000000000000000100100;
assign LUT_1[45546] = 32'b00000000000000000010011100111001;
assign LUT_1[45547] = 32'b11111111111111111011101110110101;
assign LUT_1[45548] = 32'b00000000000000001110100111111111;
assign LUT_1[45549] = 32'b00000000000000000111111001111011;
assign LUT_1[45550] = 32'b00000000000000001010010110010000;
assign LUT_1[45551] = 32'b00000000000000000011101000001100;
assign LUT_1[45552] = 32'b00000000000000001001011100010101;
assign LUT_1[45553] = 32'b00000000000000000010101110010001;
assign LUT_1[45554] = 32'b00000000000000000101001010100110;
assign LUT_1[45555] = 32'b11111111111111111110011100100010;
assign LUT_1[45556] = 32'b00000000000000010001010101101100;
assign LUT_1[45557] = 32'b00000000000000001010100111101000;
assign LUT_1[45558] = 32'b00000000000000001101000011111101;
assign LUT_1[45559] = 32'b00000000000000000110010101111001;
assign LUT_1[45560] = 32'b00000000000000001000101010001010;
assign LUT_1[45561] = 32'b00000000000000000001111100000110;
assign LUT_1[45562] = 32'b00000000000000000100011000011011;
assign LUT_1[45563] = 32'b11111111111111111101101010010111;
assign LUT_1[45564] = 32'b00000000000000010000100011100001;
assign LUT_1[45565] = 32'b00000000000000001001110101011101;
assign LUT_1[45566] = 32'b00000000000000001100010001110010;
assign LUT_1[45567] = 32'b00000000000000000101100011101110;
assign LUT_1[45568] = 32'b11111111111111111101100010011010;
assign LUT_1[45569] = 32'b11111111111111110110110100010110;
assign LUT_1[45570] = 32'b11111111111111111001010000101011;
assign LUT_1[45571] = 32'b11111111111111110010100010100111;
assign LUT_1[45572] = 32'b00000000000000000101011011110001;
assign LUT_1[45573] = 32'b11111111111111111110101101101101;
assign LUT_1[45574] = 32'b00000000000000000001001010000010;
assign LUT_1[45575] = 32'b11111111111111111010011011111110;
assign LUT_1[45576] = 32'b11111111111111111100110000001111;
assign LUT_1[45577] = 32'b11111111111111110110000010001011;
assign LUT_1[45578] = 32'b11111111111111111000011110100000;
assign LUT_1[45579] = 32'b11111111111111110001110000011100;
assign LUT_1[45580] = 32'b00000000000000000100101001100110;
assign LUT_1[45581] = 32'b11111111111111111101111011100010;
assign LUT_1[45582] = 32'b00000000000000000000010111110111;
assign LUT_1[45583] = 32'b11111111111111111001101001110011;
assign LUT_1[45584] = 32'b11111111111111111111011101111100;
assign LUT_1[45585] = 32'b11111111111111111000101111111000;
assign LUT_1[45586] = 32'b11111111111111111011001100001101;
assign LUT_1[45587] = 32'b11111111111111110100011110001001;
assign LUT_1[45588] = 32'b00000000000000000111010111010011;
assign LUT_1[45589] = 32'b00000000000000000000101001001111;
assign LUT_1[45590] = 32'b00000000000000000011000101100100;
assign LUT_1[45591] = 32'b11111111111111111100010111100000;
assign LUT_1[45592] = 32'b11111111111111111110101011110001;
assign LUT_1[45593] = 32'b11111111111111110111111101101101;
assign LUT_1[45594] = 32'b11111111111111111010011010000010;
assign LUT_1[45595] = 32'b11111111111111110011101011111110;
assign LUT_1[45596] = 32'b00000000000000000110100101001000;
assign LUT_1[45597] = 32'b11111111111111111111110111000100;
assign LUT_1[45598] = 32'b00000000000000000010010011011001;
assign LUT_1[45599] = 32'b11111111111111111011100101010101;
assign LUT_1[45600] = 32'b11111111111111111110011101011001;
assign LUT_1[45601] = 32'b11111111111111110111101111010101;
assign LUT_1[45602] = 32'b11111111111111111010001011101010;
assign LUT_1[45603] = 32'b11111111111111110011011101100110;
assign LUT_1[45604] = 32'b00000000000000000110010110110000;
assign LUT_1[45605] = 32'b11111111111111111111101000101100;
assign LUT_1[45606] = 32'b00000000000000000010000101000001;
assign LUT_1[45607] = 32'b11111111111111111011010110111101;
assign LUT_1[45608] = 32'b11111111111111111101101011001110;
assign LUT_1[45609] = 32'b11111111111111110110111101001010;
assign LUT_1[45610] = 32'b11111111111111111001011001011111;
assign LUT_1[45611] = 32'b11111111111111110010101011011011;
assign LUT_1[45612] = 32'b00000000000000000101100100100101;
assign LUT_1[45613] = 32'b11111111111111111110110110100001;
assign LUT_1[45614] = 32'b00000000000000000001010010110110;
assign LUT_1[45615] = 32'b11111111111111111010100100110010;
assign LUT_1[45616] = 32'b00000000000000000000011000111011;
assign LUT_1[45617] = 32'b11111111111111111001101010110111;
assign LUT_1[45618] = 32'b11111111111111111100000111001100;
assign LUT_1[45619] = 32'b11111111111111110101011001001000;
assign LUT_1[45620] = 32'b00000000000000001000010010010010;
assign LUT_1[45621] = 32'b00000000000000000001100100001110;
assign LUT_1[45622] = 32'b00000000000000000100000000100011;
assign LUT_1[45623] = 32'b11111111111111111101010010011111;
assign LUT_1[45624] = 32'b11111111111111111111100110110000;
assign LUT_1[45625] = 32'b11111111111111111000111000101100;
assign LUT_1[45626] = 32'b11111111111111111011010101000001;
assign LUT_1[45627] = 32'b11111111111111110100100110111101;
assign LUT_1[45628] = 32'b00000000000000000111100000000111;
assign LUT_1[45629] = 32'b00000000000000000000110010000011;
assign LUT_1[45630] = 32'b00000000000000000011001110011000;
assign LUT_1[45631] = 32'b11111111111111111100100000010100;
assign LUT_1[45632] = 32'b11111111111111111111100000000010;
assign LUT_1[45633] = 32'b11111111111111111000110001111110;
assign LUT_1[45634] = 32'b11111111111111111011001110010011;
assign LUT_1[45635] = 32'b11111111111111110100100000001111;
assign LUT_1[45636] = 32'b00000000000000000111011001011001;
assign LUT_1[45637] = 32'b00000000000000000000101011010101;
assign LUT_1[45638] = 32'b00000000000000000011000111101010;
assign LUT_1[45639] = 32'b11111111111111111100011001100110;
assign LUT_1[45640] = 32'b11111111111111111110101101110111;
assign LUT_1[45641] = 32'b11111111111111110111111111110011;
assign LUT_1[45642] = 32'b11111111111111111010011100001000;
assign LUT_1[45643] = 32'b11111111111111110011101110000100;
assign LUT_1[45644] = 32'b00000000000000000110100111001110;
assign LUT_1[45645] = 32'b11111111111111111111111001001010;
assign LUT_1[45646] = 32'b00000000000000000010010101011111;
assign LUT_1[45647] = 32'b11111111111111111011100111011011;
assign LUT_1[45648] = 32'b00000000000000000001011011100100;
assign LUT_1[45649] = 32'b11111111111111111010101101100000;
assign LUT_1[45650] = 32'b11111111111111111101001001110101;
assign LUT_1[45651] = 32'b11111111111111110110011011110001;
assign LUT_1[45652] = 32'b00000000000000001001010100111011;
assign LUT_1[45653] = 32'b00000000000000000010100110110111;
assign LUT_1[45654] = 32'b00000000000000000101000011001100;
assign LUT_1[45655] = 32'b11111111111111111110010101001000;
assign LUT_1[45656] = 32'b00000000000000000000101001011001;
assign LUT_1[45657] = 32'b11111111111111111001111011010101;
assign LUT_1[45658] = 32'b11111111111111111100010111101010;
assign LUT_1[45659] = 32'b11111111111111110101101001100110;
assign LUT_1[45660] = 32'b00000000000000001000100010110000;
assign LUT_1[45661] = 32'b00000000000000000001110100101100;
assign LUT_1[45662] = 32'b00000000000000000100010001000001;
assign LUT_1[45663] = 32'b11111111111111111101100010111101;
assign LUT_1[45664] = 32'b00000000000000000000011011000001;
assign LUT_1[45665] = 32'b11111111111111111001101100111101;
assign LUT_1[45666] = 32'b11111111111111111100001001010010;
assign LUT_1[45667] = 32'b11111111111111110101011011001110;
assign LUT_1[45668] = 32'b00000000000000001000010100011000;
assign LUT_1[45669] = 32'b00000000000000000001100110010100;
assign LUT_1[45670] = 32'b00000000000000000100000010101001;
assign LUT_1[45671] = 32'b11111111111111111101010100100101;
assign LUT_1[45672] = 32'b11111111111111111111101000110110;
assign LUT_1[45673] = 32'b11111111111111111000111010110010;
assign LUT_1[45674] = 32'b11111111111111111011010111000111;
assign LUT_1[45675] = 32'b11111111111111110100101001000011;
assign LUT_1[45676] = 32'b00000000000000000111100010001101;
assign LUT_1[45677] = 32'b00000000000000000000110100001001;
assign LUT_1[45678] = 32'b00000000000000000011010000011110;
assign LUT_1[45679] = 32'b11111111111111111100100010011010;
assign LUT_1[45680] = 32'b00000000000000000010010110100011;
assign LUT_1[45681] = 32'b11111111111111111011101000011111;
assign LUT_1[45682] = 32'b11111111111111111110000100110100;
assign LUT_1[45683] = 32'b11111111111111110111010110110000;
assign LUT_1[45684] = 32'b00000000000000001010001111111010;
assign LUT_1[45685] = 32'b00000000000000000011100001110110;
assign LUT_1[45686] = 32'b00000000000000000101111110001011;
assign LUT_1[45687] = 32'b11111111111111111111010000000111;
assign LUT_1[45688] = 32'b00000000000000000001100100011000;
assign LUT_1[45689] = 32'b11111111111111111010110110010100;
assign LUT_1[45690] = 32'b11111111111111111101010010101001;
assign LUT_1[45691] = 32'b11111111111111110110100100100101;
assign LUT_1[45692] = 32'b00000000000000001001011101101111;
assign LUT_1[45693] = 32'b00000000000000000010101111101011;
assign LUT_1[45694] = 32'b00000000000000000101001100000000;
assign LUT_1[45695] = 32'b11111111111111111110011101111100;
assign LUT_1[45696] = 32'b00000000000000000000100010011101;
assign LUT_1[45697] = 32'b11111111111111111001110100011001;
assign LUT_1[45698] = 32'b11111111111111111100010000101110;
assign LUT_1[45699] = 32'b11111111111111110101100010101010;
assign LUT_1[45700] = 32'b00000000000000001000011011110100;
assign LUT_1[45701] = 32'b00000000000000000001101101110000;
assign LUT_1[45702] = 32'b00000000000000000100001010000101;
assign LUT_1[45703] = 32'b11111111111111111101011100000001;
assign LUT_1[45704] = 32'b11111111111111111111110000010010;
assign LUT_1[45705] = 32'b11111111111111111001000010001110;
assign LUT_1[45706] = 32'b11111111111111111011011110100011;
assign LUT_1[45707] = 32'b11111111111111110100110000011111;
assign LUT_1[45708] = 32'b00000000000000000111101001101001;
assign LUT_1[45709] = 32'b00000000000000000000111011100101;
assign LUT_1[45710] = 32'b00000000000000000011010111111010;
assign LUT_1[45711] = 32'b11111111111111111100101001110110;
assign LUT_1[45712] = 32'b00000000000000000010011101111111;
assign LUT_1[45713] = 32'b11111111111111111011101111111011;
assign LUT_1[45714] = 32'b11111111111111111110001100010000;
assign LUT_1[45715] = 32'b11111111111111110111011110001100;
assign LUT_1[45716] = 32'b00000000000000001010010111010110;
assign LUT_1[45717] = 32'b00000000000000000011101001010010;
assign LUT_1[45718] = 32'b00000000000000000110000101100111;
assign LUT_1[45719] = 32'b11111111111111111111010111100011;
assign LUT_1[45720] = 32'b00000000000000000001101011110100;
assign LUT_1[45721] = 32'b11111111111111111010111101110000;
assign LUT_1[45722] = 32'b11111111111111111101011010000101;
assign LUT_1[45723] = 32'b11111111111111110110101100000001;
assign LUT_1[45724] = 32'b00000000000000001001100101001011;
assign LUT_1[45725] = 32'b00000000000000000010110111000111;
assign LUT_1[45726] = 32'b00000000000000000101010011011100;
assign LUT_1[45727] = 32'b11111111111111111110100101011000;
assign LUT_1[45728] = 32'b00000000000000000001011101011100;
assign LUT_1[45729] = 32'b11111111111111111010101111011000;
assign LUT_1[45730] = 32'b11111111111111111101001011101101;
assign LUT_1[45731] = 32'b11111111111111110110011101101001;
assign LUT_1[45732] = 32'b00000000000000001001010110110011;
assign LUT_1[45733] = 32'b00000000000000000010101000101111;
assign LUT_1[45734] = 32'b00000000000000000101000101000100;
assign LUT_1[45735] = 32'b11111111111111111110010111000000;
assign LUT_1[45736] = 32'b00000000000000000000101011010001;
assign LUT_1[45737] = 32'b11111111111111111001111101001101;
assign LUT_1[45738] = 32'b11111111111111111100011001100010;
assign LUT_1[45739] = 32'b11111111111111110101101011011110;
assign LUT_1[45740] = 32'b00000000000000001000100100101000;
assign LUT_1[45741] = 32'b00000000000000000001110110100100;
assign LUT_1[45742] = 32'b00000000000000000100010010111001;
assign LUT_1[45743] = 32'b11111111111111111101100100110101;
assign LUT_1[45744] = 32'b00000000000000000011011000111110;
assign LUT_1[45745] = 32'b11111111111111111100101010111010;
assign LUT_1[45746] = 32'b11111111111111111111000111001111;
assign LUT_1[45747] = 32'b11111111111111111000011001001011;
assign LUT_1[45748] = 32'b00000000000000001011010010010101;
assign LUT_1[45749] = 32'b00000000000000000100100100010001;
assign LUT_1[45750] = 32'b00000000000000000111000000100110;
assign LUT_1[45751] = 32'b00000000000000000000010010100010;
assign LUT_1[45752] = 32'b00000000000000000010100110110011;
assign LUT_1[45753] = 32'b11111111111111111011111000101111;
assign LUT_1[45754] = 32'b11111111111111111110010101000100;
assign LUT_1[45755] = 32'b11111111111111110111100111000000;
assign LUT_1[45756] = 32'b00000000000000001010100000001010;
assign LUT_1[45757] = 32'b00000000000000000011110010000110;
assign LUT_1[45758] = 32'b00000000000000000110001110011011;
assign LUT_1[45759] = 32'b11111111111111111111100000010111;
assign LUT_1[45760] = 32'b00000000000000000010100000000101;
assign LUT_1[45761] = 32'b11111111111111111011110010000001;
assign LUT_1[45762] = 32'b11111111111111111110001110010110;
assign LUT_1[45763] = 32'b11111111111111110111100000010010;
assign LUT_1[45764] = 32'b00000000000000001010011001011100;
assign LUT_1[45765] = 32'b00000000000000000011101011011000;
assign LUT_1[45766] = 32'b00000000000000000110000111101101;
assign LUT_1[45767] = 32'b11111111111111111111011001101001;
assign LUT_1[45768] = 32'b00000000000000000001101101111010;
assign LUT_1[45769] = 32'b11111111111111111010111111110110;
assign LUT_1[45770] = 32'b11111111111111111101011100001011;
assign LUT_1[45771] = 32'b11111111111111110110101110000111;
assign LUT_1[45772] = 32'b00000000000000001001100111010001;
assign LUT_1[45773] = 32'b00000000000000000010111001001101;
assign LUT_1[45774] = 32'b00000000000000000101010101100010;
assign LUT_1[45775] = 32'b11111111111111111110100111011110;
assign LUT_1[45776] = 32'b00000000000000000100011011100111;
assign LUT_1[45777] = 32'b11111111111111111101101101100011;
assign LUT_1[45778] = 32'b00000000000000000000001001111000;
assign LUT_1[45779] = 32'b11111111111111111001011011110100;
assign LUT_1[45780] = 32'b00000000000000001100010100111110;
assign LUT_1[45781] = 32'b00000000000000000101100110111010;
assign LUT_1[45782] = 32'b00000000000000001000000011001111;
assign LUT_1[45783] = 32'b00000000000000000001010101001011;
assign LUT_1[45784] = 32'b00000000000000000011101001011100;
assign LUT_1[45785] = 32'b11111111111111111100111011011000;
assign LUT_1[45786] = 32'b11111111111111111111010111101101;
assign LUT_1[45787] = 32'b11111111111111111000101001101001;
assign LUT_1[45788] = 32'b00000000000000001011100010110011;
assign LUT_1[45789] = 32'b00000000000000000100110100101111;
assign LUT_1[45790] = 32'b00000000000000000111010001000100;
assign LUT_1[45791] = 32'b00000000000000000000100011000000;
assign LUT_1[45792] = 32'b00000000000000000011011011000100;
assign LUT_1[45793] = 32'b11111111111111111100101101000000;
assign LUT_1[45794] = 32'b11111111111111111111001001010101;
assign LUT_1[45795] = 32'b11111111111111111000011011010001;
assign LUT_1[45796] = 32'b00000000000000001011010100011011;
assign LUT_1[45797] = 32'b00000000000000000100100110010111;
assign LUT_1[45798] = 32'b00000000000000000111000010101100;
assign LUT_1[45799] = 32'b00000000000000000000010100101000;
assign LUT_1[45800] = 32'b00000000000000000010101000111001;
assign LUT_1[45801] = 32'b11111111111111111011111010110101;
assign LUT_1[45802] = 32'b11111111111111111110010111001010;
assign LUT_1[45803] = 32'b11111111111111110111101001000110;
assign LUT_1[45804] = 32'b00000000000000001010100010010000;
assign LUT_1[45805] = 32'b00000000000000000011110100001100;
assign LUT_1[45806] = 32'b00000000000000000110010000100001;
assign LUT_1[45807] = 32'b11111111111111111111100010011101;
assign LUT_1[45808] = 32'b00000000000000000101010110100110;
assign LUT_1[45809] = 32'b11111111111111111110101000100010;
assign LUT_1[45810] = 32'b00000000000000000001000100110111;
assign LUT_1[45811] = 32'b11111111111111111010010110110011;
assign LUT_1[45812] = 32'b00000000000000001101001111111101;
assign LUT_1[45813] = 32'b00000000000000000110100001111001;
assign LUT_1[45814] = 32'b00000000000000001000111110001110;
assign LUT_1[45815] = 32'b00000000000000000010010000001010;
assign LUT_1[45816] = 32'b00000000000000000100100100011011;
assign LUT_1[45817] = 32'b11111111111111111101110110010111;
assign LUT_1[45818] = 32'b00000000000000000000010010101100;
assign LUT_1[45819] = 32'b11111111111111111001100100101000;
assign LUT_1[45820] = 32'b00000000000000001100011101110010;
assign LUT_1[45821] = 32'b00000000000000000101101111101110;
assign LUT_1[45822] = 32'b00000000000000001000001100000011;
assign LUT_1[45823] = 32'b00000000000000000001011101111111;
assign LUT_1[45824] = 32'b11111111111111111011010110100110;
assign LUT_1[45825] = 32'b11111111111111110100101000100010;
assign LUT_1[45826] = 32'b11111111111111110111000100110111;
assign LUT_1[45827] = 32'b11111111111111110000010110110011;
assign LUT_1[45828] = 32'b00000000000000000011001111111101;
assign LUT_1[45829] = 32'b11111111111111111100100001111001;
assign LUT_1[45830] = 32'b11111111111111111110111110001110;
assign LUT_1[45831] = 32'b11111111111111111000010000001010;
assign LUT_1[45832] = 32'b11111111111111111010100100011011;
assign LUT_1[45833] = 32'b11111111111111110011110110010111;
assign LUT_1[45834] = 32'b11111111111111110110010010101100;
assign LUT_1[45835] = 32'b11111111111111101111100100101000;
assign LUT_1[45836] = 32'b00000000000000000010011101110010;
assign LUT_1[45837] = 32'b11111111111111111011101111101110;
assign LUT_1[45838] = 32'b11111111111111111110001100000011;
assign LUT_1[45839] = 32'b11111111111111110111011101111111;
assign LUT_1[45840] = 32'b11111111111111111101010010001000;
assign LUT_1[45841] = 32'b11111111111111110110100100000100;
assign LUT_1[45842] = 32'b11111111111111111001000000011001;
assign LUT_1[45843] = 32'b11111111111111110010010010010101;
assign LUT_1[45844] = 32'b00000000000000000101001011011111;
assign LUT_1[45845] = 32'b11111111111111111110011101011011;
assign LUT_1[45846] = 32'b00000000000000000000111001110000;
assign LUT_1[45847] = 32'b11111111111111111010001011101100;
assign LUT_1[45848] = 32'b11111111111111111100011111111101;
assign LUT_1[45849] = 32'b11111111111111110101110001111001;
assign LUT_1[45850] = 32'b11111111111111111000001110001110;
assign LUT_1[45851] = 32'b11111111111111110001100000001010;
assign LUT_1[45852] = 32'b00000000000000000100011001010100;
assign LUT_1[45853] = 32'b11111111111111111101101011010000;
assign LUT_1[45854] = 32'b00000000000000000000000111100101;
assign LUT_1[45855] = 32'b11111111111111111001011001100001;
assign LUT_1[45856] = 32'b11111111111111111100010001100101;
assign LUT_1[45857] = 32'b11111111111111110101100011100001;
assign LUT_1[45858] = 32'b11111111111111110111111111110110;
assign LUT_1[45859] = 32'b11111111111111110001010001110010;
assign LUT_1[45860] = 32'b00000000000000000100001010111100;
assign LUT_1[45861] = 32'b11111111111111111101011100111000;
assign LUT_1[45862] = 32'b11111111111111111111111001001101;
assign LUT_1[45863] = 32'b11111111111111111001001011001001;
assign LUT_1[45864] = 32'b11111111111111111011011111011010;
assign LUT_1[45865] = 32'b11111111111111110100110001010110;
assign LUT_1[45866] = 32'b11111111111111110111001101101011;
assign LUT_1[45867] = 32'b11111111111111110000011111100111;
assign LUT_1[45868] = 32'b00000000000000000011011000110001;
assign LUT_1[45869] = 32'b11111111111111111100101010101101;
assign LUT_1[45870] = 32'b11111111111111111111000111000010;
assign LUT_1[45871] = 32'b11111111111111111000011000111110;
assign LUT_1[45872] = 32'b11111111111111111110001101000111;
assign LUT_1[45873] = 32'b11111111111111110111011111000011;
assign LUT_1[45874] = 32'b11111111111111111001111011011000;
assign LUT_1[45875] = 32'b11111111111111110011001101010100;
assign LUT_1[45876] = 32'b00000000000000000110000110011110;
assign LUT_1[45877] = 32'b11111111111111111111011000011010;
assign LUT_1[45878] = 32'b00000000000000000001110100101111;
assign LUT_1[45879] = 32'b11111111111111111011000110101011;
assign LUT_1[45880] = 32'b11111111111111111101011010111100;
assign LUT_1[45881] = 32'b11111111111111110110101100111000;
assign LUT_1[45882] = 32'b11111111111111111001001001001101;
assign LUT_1[45883] = 32'b11111111111111110010011011001001;
assign LUT_1[45884] = 32'b00000000000000000101010100010011;
assign LUT_1[45885] = 32'b11111111111111111110100110001111;
assign LUT_1[45886] = 32'b00000000000000000001000010100100;
assign LUT_1[45887] = 32'b11111111111111111010010100100000;
assign LUT_1[45888] = 32'b11111111111111111101010100001110;
assign LUT_1[45889] = 32'b11111111111111110110100110001010;
assign LUT_1[45890] = 32'b11111111111111111001000010011111;
assign LUT_1[45891] = 32'b11111111111111110010010100011011;
assign LUT_1[45892] = 32'b00000000000000000101001101100101;
assign LUT_1[45893] = 32'b11111111111111111110011111100001;
assign LUT_1[45894] = 32'b00000000000000000000111011110110;
assign LUT_1[45895] = 32'b11111111111111111010001101110010;
assign LUT_1[45896] = 32'b11111111111111111100100010000011;
assign LUT_1[45897] = 32'b11111111111111110101110011111111;
assign LUT_1[45898] = 32'b11111111111111111000010000010100;
assign LUT_1[45899] = 32'b11111111111111110001100010010000;
assign LUT_1[45900] = 32'b00000000000000000100011011011010;
assign LUT_1[45901] = 32'b11111111111111111101101101010110;
assign LUT_1[45902] = 32'b00000000000000000000001001101011;
assign LUT_1[45903] = 32'b11111111111111111001011011100111;
assign LUT_1[45904] = 32'b11111111111111111111001111110000;
assign LUT_1[45905] = 32'b11111111111111111000100001101100;
assign LUT_1[45906] = 32'b11111111111111111010111110000001;
assign LUT_1[45907] = 32'b11111111111111110100001111111101;
assign LUT_1[45908] = 32'b00000000000000000111001001000111;
assign LUT_1[45909] = 32'b00000000000000000000011011000011;
assign LUT_1[45910] = 32'b00000000000000000010110111011000;
assign LUT_1[45911] = 32'b11111111111111111100001001010100;
assign LUT_1[45912] = 32'b11111111111111111110011101100101;
assign LUT_1[45913] = 32'b11111111111111110111101111100001;
assign LUT_1[45914] = 32'b11111111111111111010001011110110;
assign LUT_1[45915] = 32'b11111111111111110011011101110010;
assign LUT_1[45916] = 32'b00000000000000000110010110111100;
assign LUT_1[45917] = 32'b11111111111111111111101000111000;
assign LUT_1[45918] = 32'b00000000000000000010000101001101;
assign LUT_1[45919] = 32'b11111111111111111011010111001001;
assign LUT_1[45920] = 32'b11111111111111111110001111001101;
assign LUT_1[45921] = 32'b11111111111111110111100001001001;
assign LUT_1[45922] = 32'b11111111111111111001111101011110;
assign LUT_1[45923] = 32'b11111111111111110011001111011010;
assign LUT_1[45924] = 32'b00000000000000000110001000100100;
assign LUT_1[45925] = 32'b11111111111111111111011010100000;
assign LUT_1[45926] = 32'b00000000000000000001110110110101;
assign LUT_1[45927] = 32'b11111111111111111011001000110001;
assign LUT_1[45928] = 32'b11111111111111111101011101000010;
assign LUT_1[45929] = 32'b11111111111111110110101110111110;
assign LUT_1[45930] = 32'b11111111111111111001001011010011;
assign LUT_1[45931] = 32'b11111111111111110010011101001111;
assign LUT_1[45932] = 32'b00000000000000000101010110011001;
assign LUT_1[45933] = 32'b11111111111111111110101000010101;
assign LUT_1[45934] = 32'b00000000000000000001000100101010;
assign LUT_1[45935] = 32'b11111111111111111010010110100110;
assign LUT_1[45936] = 32'b00000000000000000000001010101111;
assign LUT_1[45937] = 32'b11111111111111111001011100101011;
assign LUT_1[45938] = 32'b11111111111111111011111001000000;
assign LUT_1[45939] = 32'b11111111111111110101001010111100;
assign LUT_1[45940] = 32'b00000000000000001000000100000110;
assign LUT_1[45941] = 32'b00000000000000000001010110000010;
assign LUT_1[45942] = 32'b00000000000000000011110010010111;
assign LUT_1[45943] = 32'b11111111111111111101000100010011;
assign LUT_1[45944] = 32'b11111111111111111111011000100100;
assign LUT_1[45945] = 32'b11111111111111111000101010100000;
assign LUT_1[45946] = 32'b11111111111111111011000110110101;
assign LUT_1[45947] = 32'b11111111111111110100011000110001;
assign LUT_1[45948] = 32'b00000000000000000111010001111011;
assign LUT_1[45949] = 32'b00000000000000000000100011110111;
assign LUT_1[45950] = 32'b00000000000000000011000000001100;
assign LUT_1[45951] = 32'b11111111111111111100010010001000;
assign LUT_1[45952] = 32'b11111111111111111110010110101001;
assign LUT_1[45953] = 32'b11111111111111110111101000100101;
assign LUT_1[45954] = 32'b11111111111111111010000100111010;
assign LUT_1[45955] = 32'b11111111111111110011010110110110;
assign LUT_1[45956] = 32'b00000000000000000110010000000000;
assign LUT_1[45957] = 32'b11111111111111111111100001111100;
assign LUT_1[45958] = 32'b00000000000000000001111110010001;
assign LUT_1[45959] = 32'b11111111111111111011010000001101;
assign LUT_1[45960] = 32'b11111111111111111101100100011110;
assign LUT_1[45961] = 32'b11111111111111110110110110011010;
assign LUT_1[45962] = 32'b11111111111111111001010010101111;
assign LUT_1[45963] = 32'b11111111111111110010100100101011;
assign LUT_1[45964] = 32'b00000000000000000101011101110101;
assign LUT_1[45965] = 32'b11111111111111111110101111110001;
assign LUT_1[45966] = 32'b00000000000000000001001100000110;
assign LUT_1[45967] = 32'b11111111111111111010011110000010;
assign LUT_1[45968] = 32'b00000000000000000000010010001011;
assign LUT_1[45969] = 32'b11111111111111111001100100000111;
assign LUT_1[45970] = 32'b11111111111111111100000000011100;
assign LUT_1[45971] = 32'b11111111111111110101010010011000;
assign LUT_1[45972] = 32'b00000000000000001000001011100010;
assign LUT_1[45973] = 32'b00000000000000000001011101011110;
assign LUT_1[45974] = 32'b00000000000000000011111001110011;
assign LUT_1[45975] = 32'b11111111111111111101001011101111;
assign LUT_1[45976] = 32'b11111111111111111111100000000000;
assign LUT_1[45977] = 32'b11111111111111111000110001111100;
assign LUT_1[45978] = 32'b11111111111111111011001110010001;
assign LUT_1[45979] = 32'b11111111111111110100100000001101;
assign LUT_1[45980] = 32'b00000000000000000111011001010111;
assign LUT_1[45981] = 32'b00000000000000000000101011010011;
assign LUT_1[45982] = 32'b00000000000000000011000111101000;
assign LUT_1[45983] = 32'b11111111111111111100011001100100;
assign LUT_1[45984] = 32'b11111111111111111111010001101000;
assign LUT_1[45985] = 32'b11111111111111111000100011100100;
assign LUT_1[45986] = 32'b11111111111111111010111111111001;
assign LUT_1[45987] = 32'b11111111111111110100010001110101;
assign LUT_1[45988] = 32'b00000000000000000111001010111111;
assign LUT_1[45989] = 32'b00000000000000000000011100111011;
assign LUT_1[45990] = 32'b00000000000000000010111001010000;
assign LUT_1[45991] = 32'b11111111111111111100001011001100;
assign LUT_1[45992] = 32'b11111111111111111110011111011101;
assign LUT_1[45993] = 32'b11111111111111110111110001011001;
assign LUT_1[45994] = 32'b11111111111111111010001101101110;
assign LUT_1[45995] = 32'b11111111111111110011011111101010;
assign LUT_1[45996] = 32'b00000000000000000110011000110100;
assign LUT_1[45997] = 32'b11111111111111111111101010110000;
assign LUT_1[45998] = 32'b00000000000000000010000111000101;
assign LUT_1[45999] = 32'b11111111111111111011011001000001;
assign LUT_1[46000] = 32'b00000000000000000001001101001010;
assign LUT_1[46001] = 32'b11111111111111111010011111000110;
assign LUT_1[46002] = 32'b11111111111111111100111011011011;
assign LUT_1[46003] = 32'b11111111111111110110001101010111;
assign LUT_1[46004] = 32'b00000000000000001001000110100001;
assign LUT_1[46005] = 32'b00000000000000000010011000011101;
assign LUT_1[46006] = 32'b00000000000000000100110100110010;
assign LUT_1[46007] = 32'b11111111111111111110000110101110;
assign LUT_1[46008] = 32'b00000000000000000000011010111111;
assign LUT_1[46009] = 32'b11111111111111111001101100111011;
assign LUT_1[46010] = 32'b11111111111111111100001001010000;
assign LUT_1[46011] = 32'b11111111111111110101011011001100;
assign LUT_1[46012] = 32'b00000000000000001000010100010110;
assign LUT_1[46013] = 32'b00000000000000000001100110010010;
assign LUT_1[46014] = 32'b00000000000000000100000010100111;
assign LUT_1[46015] = 32'b11111111111111111101010100100011;
assign LUT_1[46016] = 32'b00000000000000000000010100010001;
assign LUT_1[46017] = 32'b11111111111111111001100110001101;
assign LUT_1[46018] = 32'b11111111111111111100000010100010;
assign LUT_1[46019] = 32'b11111111111111110101010100011110;
assign LUT_1[46020] = 32'b00000000000000001000001101101000;
assign LUT_1[46021] = 32'b00000000000000000001011111100100;
assign LUT_1[46022] = 32'b00000000000000000011111011111001;
assign LUT_1[46023] = 32'b11111111111111111101001101110101;
assign LUT_1[46024] = 32'b11111111111111111111100010000110;
assign LUT_1[46025] = 32'b11111111111111111000110100000010;
assign LUT_1[46026] = 32'b11111111111111111011010000010111;
assign LUT_1[46027] = 32'b11111111111111110100100010010011;
assign LUT_1[46028] = 32'b00000000000000000111011011011101;
assign LUT_1[46029] = 32'b00000000000000000000101101011001;
assign LUT_1[46030] = 32'b00000000000000000011001001101110;
assign LUT_1[46031] = 32'b11111111111111111100011011101010;
assign LUT_1[46032] = 32'b00000000000000000010001111110011;
assign LUT_1[46033] = 32'b11111111111111111011100001101111;
assign LUT_1[46034] = 32'b11111111111111111101111110000100;
assign LUT_1[46035] = 32'b11111111111111110111010000000000;
assign LUT_1[46036] = 32'b00000000000000001010001001001010;
assign LUT_1[46037] = 32'b00000000000000000011011011000110;
assign LUT_1[46038] = 32'b00000000000000000101110111011011;
assign LUT_1[46039] = 32'b11111111111111111111001001010111;
assign LUT_1[46040] = 32'b00000000000000000001011101101000;
assign LUT_1[46041] = 32'b11111111111111111010101111100100;
assign LUT_1[46042] = 32'b11111111111111111101001011111001;
assign LUT_1[46043] = 32'b11111111111111110110011101110101;
assign LUT_1[46044] = 32'b00000000000000001001010110111111;
assign LUT_1[46045] = 32'b00000000000000000010101000111011;
assign LUT_1[46046] = 32'b00000000000000000101000101010000;
assign LUT_1[46047] = 32'b11111111111111111110010111001100;
assign LUT_1[46048] = 32'b00000000000000000001001111010000;
assign LUT_1[46049] = 32'b11111111111111111010100001001100;
assign LUT_1[46050] = 32'b11111111111111111100111101100001;
assign LUT_1[46051] = 32'b11111111111111110110001111011101;
assign LUT_1[46052] = 32'b00000000000000001001001000100111;
assign LUT_1[46053] = 32'b00000000000000000010011010100011;
assign LUT_1[46054] = 32'b00000000000000000100110110111000;
assign LUT_1[46055] = 32'b11111111111111111110001000110100;
assign LUT_1[46056] = 32'b00000000000000000000011101000101;
assign LUT_1[46057] = 32'b11111111111111111001101111000001;
assign LUT_1[46058] = 32'b11111111111111111100001011010110;
assign LUT_1[46059] = 32'b11111111111111110101011101010010;
assign LUT_1[46060] = 32'b00000000000000001000010110011100;
assign LUT_1[46061] = 32'b00000000000000000001101000011000;
assign LUT_1[46062] = 32'b00000000000000000100000100101101;
assign LUT_1[46063] = 32'b11111111111111111101010110101001;
assign LUT_1[46064] = 32'b00000000000000000011001010110010;
assign LUT_1[46065] = 32'b11111111111111111100011100101110;
assign LUT_1[46066] = 32'b11111111111111111110111001000011;
assign LUT_1[46067] = 32'b11111111111111111000001010111111;
assign LUT_1[46068] = 32'b00000000000000001011000100001001;
assign LUT_1[46069] = 32'b00000000000000000100010110000101;
assign LUT_1[46070] = 32'b00000000000000000110110010011010;
assign LUT_1[46071] = 32'b00000000000000000000000100010110;
assign LUT_1[46072] = 32'b00000000000000000010011000100111;
assign LUT_1[46073] = 32'b11111111111111111011101010100011;
assign LUT_1[46074] = 32'b11111111111111111110000110111000;
assign LUT_1[46075] = 32'b11111111111111110111011000110100;
assign LUT_1[46076] = 32'b00000000000000001010010001111110;
assign LUT_1[46077] = 32'b00000000000000000011100011111010;
assign LUT_1[46078] = 32'b00000000000000000110000000001111;
assign LUT_1[46079] = 32'b11111111111111111111010010001011;
assign LUT_1[46080] = 32'b00000000000000001010001010101101;
assign LUT_1[46081] = 32'b00000000000000000011011100101001;
assign LUT_1[46082] = 32'b00000000000000000101111000111110;
assign LUT_1[46083] = 32'b11111111111111111111001010111010;
assign LUT_1[46084] = 32'b00000000000000010010000100000100;
assign LUT_1[46085] = 32'b00000000000000001011010110000000;
assign LUT_1[46086] = 32'b00000000000000001101110010010101;
assign LUT_1[46087] = 32'b00000000000000000111000100010001;
assign LUT_1[46088] = 32'b00000000000000001001011000100010;
assign LUT_1[46089] = 32'b00000000000000000010101010011110;
assign LUT_1[46090] = 32'b00000000000000000101000110110011;
assign LUT_1[46091] = 32'b11111111111111111110011000101111;
assign LUT_1[46092] = 32'b00000000000000010001010001111001;
assign LUT_1[46093] = 32'b00000000000000001010100011110101;
assign LUT_1[46094] = 32'b00000000000000001101000000001010;
assign LUT_1[46095] = 32'b00000000000000000110010010000110;
assign LUT_1[46096] = 32'b00000000000000001100000110001111;
assign LUT_1[46097] = 32'b00000000000000000101011000001011;
assign LUT_1[46098] = 32'b00000000000000000111110100100000;
assign LUT_1[46099] = 32'b00000000000000000001000110011100;
assign LUT_1[46100] = 32'b00000000000000010011111111100110;
assign LUT_1[46101] = 32'b00000000000000001101010001100010;
assign LUT_1[46102] = 32'b00000000000000001111101101110111;
assign LUT_1[46103] = 32'b00000000000000001000111111110011;
assign LUT_1[46104] = 32'b00000000000000001011010100000100;
assign LUT_1[46105] = 32'b00000000000000000100100110000000;
assign LUT_1[46106] = 32'b00000000000000000111000010010101;
assign LUT_1[46107] = 32'b00000000000000000000010100010001;
assign LUT_1[46108] = 32'b00000000000000010011001101011011;
assign LUT_1[46109] = 32'b00000000000000001100011111010111;
assign LUT_1[46110] = 32'b00000000000000001110111011101100;
assign LUT_1[46111] = 32'b00000000000000001000001101101000;
assign LUT_1[46112] = 32'b00000000000000001011000101101100;
assign LUT_1[46113] = 32'b00000000000000000100010111101000;
assign LUT_1[46114] = 32'b00000000000000000110110011111101;
assign LUT_1[46115] = 32'b00000000000000000000000101111001;
assign LUT_1[46116] = 32'b00000000000000010010111111000011;
assign LUT_1[46117] = 32'b00000000000000001100010000111111;
assign LUT_1[46118] = 32'b00000000000000001110101101010100;
assign LUT_1[46119] = 32'b00000000000000000111111111010000;
assign LUT_1[46120] = 32'b00000000000000001010010011100001;
assign LUT_1[46121] = 32'b00000000000000000011100101011101;
assign LUT_1[46122] = 32'b00000000000000000110000001110010;
assign LUT_1[46123] = 32'b11111111111111111111010011101110;
assign LUT_1[46124] = 32'b00000000000000010010001100111000;
assign LUT_1[46125] = 32'b00000000000000001011011110110100;
assign LUT_1[46126] = 32'b00000000000000001101111011001001;
assign LUT_1[46127] = 32'b00000000000000000111001101000101;
assign LUT_1[46128] = 32'b00000000000000001101000001001110;
assign LUT_1[46129] = 32'b00000000000000000110010011001010;
assign LUT_1[46130] = 32'b00000000000000001000101111011111;
assign LUT_1[46131] = 32'b00000000000000000010000001011011;
assign LUT_1[46132] = 32'b00000000000000010100111010100101;
assign LUT_1[46133] = 32'b00000000000000001110001100100001;
assign LUT_1[46134] = 32'b00000000000000010000101000110110;
assign LUT_1[46135] = 32'b00000000000000001001111010110010;
assign LUT_1[46136] = 32'b00000000000000001100001111000011;
assign LUT_1[46137] = 32'b00000000000000000101100000111111;
assign LUT_1[46138] = 32'b00000000000000000111111101010100;
assign LUT_1[46139] = 32'b00000000000000000001001111010000;
assign LUT_1[46140] = 32'b00000000000000010100001000011010;
assign LUT_1[46141] = 32'b00000000000000001101011010010110;
assign LUT_1[46142] = 32'b00000000000000001111110110101011;
assign LUT_1[46143] = 32'b00000000000000001001001000100111;
assign LUT_1[46144] = 32'b00000000000000001100001000010101;
assign LUT_1[46145] = 32'b00000000000000000101011010010001;
assign LUT_1[46146] = 32'b00000000000000000111110110100110;
assign LUT_1[46147] = 32'b00000000000000000001001000100010;
assign LUT_1[46148] = 32'b00000000000000010100000001101100;
assign LUT_1[46149] = 32'b00000000000000001101010011101000;
assign LUT_1[46150] = 32'b00000000000000001111101111111101;
assign LUT_1[46151] = 32'b00000000000000001001000001111001;
assign LUT_1[46152] = 32'b00000000000000001011010110001010;
assign LUT_1[46153] = 32'b00000000000000000100101000000110;
assign LUT_1[46154] = 32'b00000000000000000111000100011011;
assign LUT_1[46155] = 32'b00000000000000000000010110010111;
assign LUT_1[46156] = 32'b00000000000000010011001111100001;
assign LUT_1[46157] = 32'b00000000000000001100100001011101;
assign LUT_1[46158] = 32'b00000000000000001110111101110010;
assign LUT_1[46159] = 32'b00000000000000001000001111101110;
assign LUT_1[46160] = 32'b00000000000000001110000011110111;
assign LUT_1[46161] = 32'b00000000000000000111010101110011;
assign LUT_1[46162] = 32'b00000000000000001001110010001000;
assign LUT_1[46163] = 32'b00000000000000000011000100000100;
assign LUT_1[46164] = 32'b00000000000000010101111101001110;
assign LUT_1[46165] = 32'b00000000000000001111001111001010;
assign LUT_1[46166] = 32'b00000000000000010001101011011111;
assign LUT_1[46167] = 32'b00000000000000001010111101011011;
assign LUT_1[46168] = 32'b00000000000000001101010001101100;
assign LUT_1[46169] = 32'b00000000000000000110100011101000;
assign LUT_1[46170] = 32'b00000000000000001000111111111101;
assign LUT_1[46171] = 32'b00000000000000000010010001111001;
assign LUT_1[46172] = 32'b00000000000000010101001011000011;
assign LUT_1[46173] = 32'b00000000000000001110011100111111;
assign LUT_1[46174] = 32'b00000000000000010000111001010100;
assign LUT_1[46175] = 32'b00000000000000001010001011010000;
assign LUT_1[46176] = 32'b00000000000000001101000011010100;
assign LUT_1[46177] = 32'b00000000000000000110010101010000;
assign LUT_1[46178] = 32'b00000000000000001000110001100101;
assign LUT_1[46179] = 32'b00000000000000000010000011100001;
assign LUT_1[46180] = 32'b00000000000000010100111100101011;
assign LUT_1[46181] = 32'b00000000000000001110001110100111;
assign LUT_1[46182] = 32'b00000000000000010000101010111100;
assign LUT_1[46183] = 32'b00000000000000001001111100111000;
assign LUT_1[46184] = 32'b00000000000000001100010001001001;
assign LUT_1[46185] = 32'b00000000000000000101100011000101;
assign LUT_1[46186] = 32'b00000000000000000111111111011010;
assign LUT_1[46187] = 32'b00000000000000000001010001010110;
assign LUT_1[46188] = 32'b00000000000000010100001010100000;
assign LUT_1[46189] = 32'b00000000000000001101011100011100;
assign LUT_1[46190] = 32'b00000000000000001111111000110001;
assign LUT_1[46191] = 32'b00000000000000001001001010101101;
assign LUT_1[46192] = 32'b00000000000000001110111110110110;
assign LUT_1[46193] = 32'b00000000000000001000010000110010;
assign LUT_1[46194] = 32'b00000000000000001010101101000111;
assign LUT_1[46195] = 32'b00000000000000000011111111000011;
assign LUT_1[46196] = 32'b00000000000000010110111000001101;
assign LUT_1[46197] = 32'b00000000000000010000001010001001;
assign LUT_1[46198] = 32'b00000000000000010010100110011110;
assign LUT_1[46199] = 32'b00000000000000001011111000011010;
assign LUT_1[46200] = 32'b00000000000000001110001100101011;
assign LUT_1[46201] = 32'b00000000000000000111011110100111;
assign LUT_1[46202] = 32'b00000000000000001001111010111100;
assign LUT_1[46203] = 32'b00000000000000000011001100111000;
assign LUT_1[46204] = 32'b00000000000000010110000110000010;
assign LUT_1[46205] = 32'b00000000000000001111010111111110;
assign LUT_1[46206] = 32'b00000000000000010001110100010011;
assign LUT_1[46207] = 32'b00000000000000001011000110001111;
assign LUT_1[46208] = 32'b00000000000000001101001010110000;
assign LUT_1[46209] = 32'b00000000000000000110011100101100;
assign LUT_1[46210] = 32'b00000000000000001000111001000001;
assign LUT_1[46211] = 32'b00000000000000000010001010111101;
assign LUT_1[46212] = 32'b00000000000000010101000100000111;
assign LUT_1[46213] = 32'b00000000000000001110010110000011;
assign LUT_1[46214] = 32'b00000000000000010000110010011000;
assign LUT_1[46215] = 32'b00000000000000001010000100010100;
assign LUT_1[46216] = 32'b00000000000000001100011000100101;
assign LUT_1[46217] = 32'b00000000000000000101101010100001;
assign LUT_1[46218] = 32'b00000000000000001000000110110110;
assign LUT_1[46219] = 32'b00000000000000000001011000110010;
assign LUT_1[46220] = 32'b00000000000000010100010001111100;
assign LUT_1[46221] = 32'b00000000000000001101100011111000;
assign LUT_1[46222] = 32'b00000000000000010000000000001101;
assign LUT_1[46223] = 32'b00000000000000001001010010001001;
assign LUT_1[46224] = 32'b00000000000000001111000110010010;
assign LUT_1[46225] = 32'b00000000000000001000011000001110;
assign LUT_1[46226] = 32'b00000000000000001010110100100011;
assign LUT_1[46227] = 32'b00000000000000000100000110011111;
assign LUT_1[46228] = 32'b00000000000000010110111111101001;
assign LUT_1[46229] = 32'b00000000000000010000010001100101;
assign LUT_1[46230] = 32'b00000000000000010010101101111010;
assign LUT_1[46231] = 32'b00000000000000001011111111110110;
assign LUT_1[46232] = 32'b00000000000000001110010100000111;
assign LUT_1[46233] = 32'b00000000000000000111100110000011;
assign LUT_1[46234] = 32'b00000000000000001010000010011000;
assign LUT_1[46235] = 32'b00000000000000000011010100010100;
assign LUT_1[46236] = 32'b00000000000000010110001101011110;
assign LUT_1[46237] = 32'b00000000000000001111011111011010;
assign LUT_1[46238] = 32'b00000000000000010001111011101111;
assign LUT_1[46239] = 32'b00000000000000001011001101101011;
assign LUT_1[46240] = 32'b00000000000000001110000101101111;
assign LUT_1[46241] = 32'b00000000000000000111010111101011;
assign LUT_1[46242] = 32'b00000000000000001001110100000000;
assign LUT_1[46243] = 32'b00000000000000000011000101111100;
assign LUT_1[46244] = 32'b00000000000000010101111111000110;
assign LUT_1[46245] = 32'b00000000000000001111010001000010;
assign LUT_1[46246] = 32'b00000000000000010001101101010111;
assign LUT_1[46247] = 32'b00000000000000001010111111010011;
assign LUT_1[46248] = 32'b00000000000000001101010011100100;
assign LUT_1[46249] = 32'b00000000000000000110100101100000;
assign LUT_1[46250] = 32'b00000000000000001001000001110101;
assign LUT_1[46251] = 32'b00000000000000000010010011110001;
assign LUT_1[46252] = 32'b00000000000000010101001100111011;
assign LUT_1[46253] = 32'b00000000000000001110011110110111;
assign LUT_1[46254] = 32'b00000000000000010000111011001100;
assign LUT_1[46255] = 32'b00000000000000001010001101001000;
assign LUT_1[46256] = 32'b00000000000000010000000001010001;
assign LUT_1[46257] = 32'b00000000000000001001010011001101;
assign LUT_1[46258] = 32'b00000000000000001011101111100010;
assign LUT_1[46259] = 32'b00000000000000000101000001011110;
assign LUT_1[46260] = 32'b00000000000000010111111010101000;
assign LUT_1[46261] = 32'b00000000000000010001001100100100;
assign LUT_1[46262] = 32'b00000000000000010011101000111001;
assign LUT_1[46263] = 32'b00000000000000001100111010110101;
assign LUT_1[46264] = 32'b00000000000000001111001111000110;
assign LUT_1[46265] = 32'b00000000000000001000100001000010;
assign LUT_1[46266] = 32'b00000000000000001010111101010111;
assign LUT_1[46267] = 32'b00000000000000000100001111010011;
assign LUT_1[46268] = 32'b00000000000000010111001000011101;
assign LUT_1[46269] = 32'b00000000000000010000011010011001;
assign LUT_1[46270] = 32'b00000000000000010010110110101110;
assign LUT_1[46271] = 32'b00000000000000001100001000101010;
assign LUT_1[46272] = 32'b00000000000000001111001000011000;
assign LUT_1[46273] = 32'b00000000000000001000011010010100;
assign LUT_1[46274] = 32'b00000000000000001010110110101001;
assign LUT_1[46275] = 32'b00000000000000000100001000100101;
assign LUT_1[46276] = 32'b00000000000000010111000001101111;
assign LUT_1[46277] = 32'b00000000000000010000010011101011;
assign LUT_1[46278] = 32'b00000000000000010010110000000000;
assign LUT_1[46279] = 32'b00000000000000001100000001111100;
assign LUT_1[46280] = 32'b00000000000000001110010110001101;
assign LUT_1[46281] = 32'b00000000000000000111101000001001;
assign LUT_1[46282] = 32'b00000000000000001010000100011110;
assign LUT_1[46283] = 32'b00000000000000000011010110011010;
assign LUT_1[46284] = 32'b00000000000000010110001111100100;
assign LUT_1[46285] = 32'b00000000000000001111100001100000;
assign LUT_1[46286] = 32'b00000000000000010001111101110101;
assign LUT_1[46287] = 32'b00000000000000001011001111110001;
assign LUT_1[46288] = 32'b00000000000000010001000011111010;
assign LUT_1[46289] = 32'b00000000000000001010010101110110;
assign LUT_1[46290] = 32'b00000000000000001100110010001011;
assign LUT_1[46291] = 32'b00000000000000000110000100000111;
assign LUT_1[46292] = 32'b00000000000000011000111101010001;
assign LUT_1[46293] = 32'b00000000000000010010001111001101;
assign LUT_1[46294] = 32'b00000000000000010100101011100010;
assign LUT_1[46295] = 32'b00000000000000001101111101011110;
assign LUT_1[46296] = 32'b00000000000000010000010001101111;
assign LUT_1[46297] = 32'b00000000000000001001100011101011;
assign LUT_1[46298] = 32'b00000000000000001100000000000000;
assign LUT_1[46299] = 32'b00000000000000000101010001111100;
assign LUT_1[46300] = 32'b00000000000000011000001011000110;
assign LUT_1[46301] = 32'b00000000000000010001011101000010;
assign LUT_1[46302] = 32'b00000000000000010011111001010111;
assign LUT_1[46303] = 32'b00000000000000001101001011010011;
assign LUT_1[46304] = 32'b00000000000000010000000011010111;
assign LUT_1[46305] = 32'b00000000000000001001010101010011;
assign LUT_1[46306] = 32'b00000000000000001011110001101000;
assign LUT_1[46307] = 32'b00000000000000000101000011100100;
assign LUT_1[46308] = 32'b00000000000000010111111100101110;
assign LUT_1[46309] = 32'b00000000000000010001001110101010;
assign LUT_1[46310] = 32'b00000000000000010011101010111111;
assign LUT_1[46311] = 32'b00000000000000001100111100111011;
assign LUT_1[46312] = 32'b00000000000000001111010001001100;
assign LUT_1[46313] = 32'b00000000000000001000100011001000;
assign LUT_1[46314] = 32'b00000000000000001010111111011101;
assign LUT_1[46315] = 32'b00000000000000000100010001011001;
assign LUT_1[46316] = 32'b00000000000000010111001010100011;
assign LUT_1[46317] = 32'b00000000000000010000011100011111;
assign LUT_1[46318] = 32'b00000000000000010010111000110100;
assign LUT_1[46319] = 32'b00000000000000001100001010110000;
assign LUT_1[46320] = 32'b00000000000000010001111110111001;
assign LUT_1[46321] = 32'b00000000000000001011010000110101;
assign LUT_1[46322] = 32'b00000000000000001101101101001010;
assign LUT_1[46323] = 32'b00000000000000000110111111000110;
assign LUT_1[46324] = 32'b00000000000000011001111000010000;
assign LUT_1[46325] = 32'b00000000000000010011001010001100;
assign LUT_1[46326] = 32'b00000000000000010101100110100001;
assign LUT_1[46327] = 32'b00000000000000001110111000011101;
assign LUT_1[46328] = 32'b00000000000000010001001100101110;
assign LUT_1[46329] = 32'b00000000000000001010011110101010;
assign LUT_1[46330] = 32'b00000000000000001100111010111111;
assign LUT_1[46331] = 32'b00000000000000000110001100111011;
assign LUT_1[46332] = 32'b00000000000000011001000110000101;
assign LUT_1[46333] = 32'b00000000000000010010011000000001;
assign LUT_1[46334] = 32'b00000000000000010100110100010110;
assign LUT_1[46335] = 32'b00000000000000001110000110010010;
assign LUT_1[46336] = 32'b00000000000000000111111110111001;
assign LUT_1[46337] = 32'b00000000000000000001010000110101;
assign LUT_1[46338] = 32'b00000000000000000011101101001010;
assign LUT_1[46339] = 32'b11111111111111111100111111000110;
assign LUT_1[46340] = 32'b00000000000000001111111000010000;
assign LUT_1[46341] = 32'b00000000000000001001001010001100;
assign LUT_1[46342] = 32'b00000000000000001011100110100001;
assign LUT_1[46343] = 32'b00000000000000000100111000011101;
assign LUT_1[46344] = 32'b00000000000000000111001100101110;
assign LUT_1[46345] = 32'b00000000000000000000011110101010;
assign LUT_1[46346] = 32'b00000000000000000010111010111111;
assign LUT_1[46347] = 32'b11111111111111111100001100111011;
assign LUT_1[46348] = 32'b00000000000000001111000110000101;
assign LUT_1[46349] = 32'b00000000000000001000011000000001;
assign LUT_1[46350] = 32'b00000000000000001010110100010110;
assign LUT_1[46351] = 32'b00000000000000000100000110010010;
assign LUT_1[46352] = 32'b00000000000000001001111010011011;
assign LUT_1[46353] = 32'b00000000000000000011001100010111;
assign LUT_1[46354] = 32'b00000000000000000101101000101100;
assign LUT_1[46355] = 32'b11111111111111111110111010101000;
assign LUT_1[46356] = 32'b00000000000000010001110011110010;
assign LUT_1[46357] = 32'b00000000000000001011000101101110;
assign LUT_1[46358] = 32'b00000000000000001101100010000011;
assign LUT_1[46359] = 32'b00000000000000000110110011111111;
assign LUT_1[46360] = 32'b00000000000000001001001000010000;
assign LUT_1[46361] = 32'b00000000000000000010011010001100;
assign LUT_1[46362] = 32'b00000000000000000100110110100001;
assign LUT_1[46363] = 32'b11111111111111111110001000011101;
assign LUT_1[46364] = 32'b00000000000000010001000001100111;
assign LUT_1[46365] = 32'b00000000000000001010010011100011;
assign LUT_1[46366] = 32'b00000000000000001100101111111000;
assign LUT_1[46367] = 32'b00000000000000000110000001110100;
assign LUT_1[46368] = 32'b00000000000000001000111001111000;
assign LUT_1[46369] = 32'b00000000000000000010001011110100;
assign LUT_1[46370] = 32'b00000000000000000100101000001001;
assign LUT_1[46371] = 32'b11111111111111111101111010000101;
assign LUT_1[46372] = 32'b00000000000000010000110011001111;
assign LUT_1[46373] = 32'b00000000000000001010000101001011;
assign LUT_1[46374] = 32'b00000000000000001100100001100000;
assign LUT_1[46375] = 32'b00000000000000000101110011011100;
assign LUT_1[46376] = 32'b00000000000000001000000111101101;
assign LUT_1[46377] = 32'b00000000000000000001011001101001;
assign LUT_1[46378] = 32'b00000000000000000011110101111110;
assign LUT_1[46379] = 32'b11111111111111111101000111111010;
assign LUT_1[46380] = 32'b00000000000000010000000001000100;
assign LUT_1[46381] = 32'b00000000000000001001010011000000;
assign LUT_1[46382] = 32'b00000000000000001011101111010101;
assign LUT_1[46383] = 32'b00000000000000000101000001010001;
assign LUT_1[46384] = 32'b00000000000000001010110101011010;
assign LUT_1[46385] = 32'b00000000000000000100000111010110;
assign LUT_1[46386] = 32'b00000000000000000110100011101011;
assign LUT_1[46387] = 32'b11111111111111111111110101100111;
assign LUT_1[46388] = 32'b00000000000000010010101110110001;
assign LUT_1[46389] = 32'b00000000000000001100000000101101;
assign LUT_1[46390] = 32'b00000000000000001110011101000010;
assign LUT_1[46391] = 32'b00000000000000000111101110111110;
assign LUT_1[46392] = 32'b00000000000000001010000011001111;
assign LUT_1[46393] = 32'b00000000000000000011010101001011;
assign LUT_1[46394] = 32'b00000000000000000101110001100000;
assign LUT_1[46395] = 32'b11111111111111111111000011011100;
assign LUT_1[46396] = 32'b00000000000000010001111100100110;
assign LUT_1[46397] = 32'b00000000000000001011001110100010;
assign LUT_1[46398] = 32'b00000000000000001101101010110111;
assign LUT_1[46399] = 32'b00000000000000000110111100110011;
assign LUT_1[46400] = 32'b00000000000000001001111100100001;
assign LUT_1[46401] = 32'b00000000000000000011001110011101;
assign LUT_1[46402] = 32'b00000000000000000101101010110010;
assign LUT_1[46403] = 32'b11111111111111111110111100101110;
assign LUT_1[46404] = 32'b00000000000000010001110101111000;
assign LUT_1[46405] = 32'b00000000000000001011000111110100;
assign LUT_1[46406] = 32'b00000000000000001101100100001001;
assign LUT_1[46407] = 32'b00000000000000000110110110000101;
assign LUT_1[46408] = 32'b00000000000000001001001010010110;
assign LUT_1[46409] = 32'b00000000000000000010011100010010;
assign LUT_1[46410] = 32'b00000000000000000100111000100111;
assign LUT_1[46411] = 32'b11111111111111111110001010100011;
assign LUT_1[46412] = 32'b00000000000000010001000011101101;
assign LUT_1[46413] = 32'b00000000000000001010010101101001;
assign LUT_1[46414] = 32'b00000000000000001100110001111110;
assign LUT_1[46415] = 32'b00000000000000000110000011111010;
assign LUT_1[46416] = 32'b00000000000000001011111000000011;
assign LUT_1[46417] = 32'b00000000000000000101001001111111;
assign LUT_1[46418] = 32'b00000000000000000111100110010100;
assign LUT_1[46419] = 32'b00000000000000000000111000010000;
assign LUT_1[46420] = 32'b00000000000000010011110001011010;
assign LUT_1[46421] = 32'b00000000000000001101000011010110;
assign LUT_1[46422] = 32'b00000000000000001111011111101011;
assign LUT_1[46423] = 32'b00000000000000001000110001100111;
assign LUT_1[46424] = 32'b00000000000000001011000101111000;
assign LUT_1[46425] = 32'b00000000000000000100010111110100;
assign LUT_1[46426] = 32'b00000000000000000110110100001001;
assign LUT_1[46427] = 32'b00000000000000000000000110000101;
assign LUT_1[46428] = 32'b00000000000000010010111111001111;
assign LUT_1[46429] = 32'b00000000000000001100010001001011;
assign LUT_1[46430] = 32'b00000000000000001110101101100000;
assign LUT_1[46431] = 32'b00000000000000000111111111011100;
assign LUT_1[46432] = 32'b00000000000000001010110111100000;
assign LUT_1[46433] = 32'b00000000000000000100001001011100;
assign LUT_1[46434] = 32'b00000000000000000110100101110001;
assign LUT_1[46435] = 32'b11111111111111111111110111101101;
assign LUT_1[46436] = 32'b00000000000000010010110000110111;
assign LUT_1[46437] = 32'b00000000000000001100000010110011;
assign LUT_1[46438] = 32'b00000000000000001110011111001000;
assign LUT_1[46439] = 32'b00000000000000000111110001000100;
assign LUT_1[46440] = 32'b00000000000000001010000101010101;
assign LUT_1[46441] = 32'b00000000000000000011010111010001;
assign LUT_1[46442] = 32'b00000000000000000101110011100110;
assign LUT_1[46443] = 32'b11111111111111111111000101100010;
assign LUT_1[46444] = 32'b00000000000000010001111110101100;
assign LUT_1[46445] = 32'b00000000000000001011010000101000;
assign LUT_1[46446] = 32'b00000000000000001101101100111101;
assign LUT_1[46447] = 32'b00000000000000000110111110111001;
assign LUT_1[46448] = 32'b00000000000000001100110011000010;
assign LUT_1[46449] = 32'b00000000000000000110000100111110;
assign LUT_1[46450] = 32'b00000000000000001000100001010011;
assign LUT_1[46451] = 32'b00000000000000000001110011001111;
assign LUT_1[46452] = 32'b00000000000000010100101100011001;
assign LUT_1[46453] = 32'b00000000000000001101111110010101;
assign LUT_1[46454] = 32'b00000000000000010000011010101010;
assign LUT_1[46455] = 32'b00000000000000001001101100100110;
assign LUT_1[46456] = 32'b00000000000000001100000000110111;
assign LUT_1[46457] = 32'b00000000000000000101010010110011;
assign LUT_1[46458] = 32'b00000000000000000111101111001000;
assign LUT_1[46459] = 32'b00000000000000000001000001000100;
assign LUT_1[46460] = 32'b00000000000000010011111010001110;
assign LUT_1[46461] = 32'b00000000000000001101001100001010;
assign LUT_1[46462] = 32'b00000000000000001111101000011111;
assign LUT_1[46463] = 32'b00000000000000001000111010011011;
assign LUT_1[46464] = 32'b00000000000000001010111110111100;
assign LUT_1[46465] = 32'b00000000000000000100010000111000;
assign LUT_1[46466] = 32'b00000000000000000110101101001101;
assign LUT_1[46467] = 32'b11111111111111111111111111001001;
assign LUT_1[46468] = 32'b00000000000000010010111000010011;
assign LUT_1[46469] = 32'b00000000000000001100001010001111;
assign LUT_1[46470] = 32'b00000000000000001110100110100100;
assign LUT_1[46471] = 32'b00000000000000000111111000100000;
assign LUT_1[46472] = 32'b00000000000000001010001100110001;
assign LUT_1[46473] = 32'b00000000000000000011011110101101;
assign LUT_1[46474] = 32'b00000000000000000101111011000010;
assign LUT_1[46475] = 32'b11111111111111111111001100111110;
assign LUT_1[46476] = 32'b00000000000000010010000110001000;
assign LUT_1[46477] = 32'b00000000000000001011011000000100;
assign LUT_1[46478] = 32'b00000000000000001101110100011001;
assign LUT_1[46479] = 32'b00000000000000000111000110010101;
assign LUT_1[46480] = 32'b00000000000000001100111010011110;
assign LUT_1[46481] = 32'b00000000000000000110001100011010;
assign LUT_1[46482] = 32'b00000000000000001000101000101111;
assign LUT_1[46483] = 32'b00000000000000000001111010101011;
assign LUT_1[46484] = 32'b00000000000000010100110011110101;
assign LUT_1[46485] = 32'b00000000000000001110000101110001;
assign LUT_1[46486] = 32'b00000000000000010000100010000110;
assign LUT_1[46487] = 32'b00000000000000001001110100000010;
assign LUT_1[46488] = 32'b00000000000000001100001000010011;
assign LUT_1[46489] = 32'b00000000000000000101011010001111;
assign LUT_1[46490] = 32'b00000000000000000111110110100100;
assign LUT_1[46491] = 32'b00000000000000000001001000100000;
assign LUT_1[46492] = 32'b00000000000000010100000001101010;
assign LUT_1[46493] = 32'b00000000000000001101010011100110;
assign LUT_1[46494] = 32'b00000000000000001111101111111011;
assign LUT_1[46495] = 32'b00000000000000001001000001110111;
assign LUT_1[46496] = 32'b00000000000000001011111001111011;
assign LUT_1[46497] = 32'b00000000000000000101001011110111;
assign LUT_1[46498] = 32'b00000000000000000111101000001100;
assign LUT_1[46499] = 32'b00000000000000000000111010001000;
assign LUT_1[46500] = 32'b00000000000000010011110011010010;
assign LUT_1[46501] = 32'b00000000000000001101000101001110;
assign LUT_1[46502] = 32'b00000000000000001111100001100011;
assign LUT_1[46503] = 32'b00000000000000001000110011011111;
assign LUT_1[46504] = 32'b00000000000000001011000111110000;
assign LUT_1[46505] = 32'b00000000000000000100011001101100;
assign LUT_1[46506] = 32'b00000000000000000110110110000001;
assign LUT_1[46507] = 32'b00000000000000000000000111111101;
assign LUT_1[46508] = 32'b00000000000000010011000001000111;
assign LUT_1[46509] = 32'b00000000000000001100010011000011;
assign LUT_1[46510] = 32'b00000000000000001110101111011000;
assign LUT_1[46511] = 32'b00000000000000001000000001010100;
assign LUT_1[46512] = 32'b00000000000000001101110101011101;
assign LUT_1[46513] = 32'b00000000000000000111000111011001;
assign LUT_1[46514] = 32'b00000000000000001001100011101110;
assign LUT_1[46515] = 32'b00000000000000000010110101101010;
assign LUT_1[46516] = 32'b00000000000000010101101110110100;
assign LUT_1[46517] = 32'b00000000000000001111000000110000;
assign LUT_1[46518] = 32'b00000000000000010001011101000101;
assign LUT_1[46519] = 32'b00000000000000001010101111000001;
assign LUT_1[46520] = 32'b00000000000000001101000011010010;
assign LUT_1[46521] = 32'b00000000000000000110010101001110;
assign LUT_1[46522] = 32'b00000000000000001000110001100011;
assign LUT_1[46523] = 32'b00000000000000000010000011011111;
assign LUT_1[46524] = 32'b00000000000000010100111100101001;
assign LUT_1[46525] = 32'b00000000000000001110001110100101;
assign LUT_1[46526] = 32'b00000000000000010000101010111010;
assign LUT_1[46527] = 32'b00000000000000001001111100110110;
assign LUT_1[46528] = 32'b00000000000000001100111100100100;
assign LUT_1[46529] = 32'b00000000000000000110001110100000;
assign LUT_1[46530] = 32'b00000000000000001000101010110101;
assign LUT_1[46531] = 32'b00000000000000000001111100110001;
assign LUT_1[46532] = 32'b00000000000000010100110101111011;
assign LUT_1[46533] = 32'b00000000000000001110000111110111;
assign LUT_1[46534] = 32'b00000000000000010000100100001100;
assign LUT_1[46535] = 32'b00000000000000001001110110001000;
assign LUT_1[46536] = 32'b00000000000000001100001010011001;
assign LUT_1[46537] = 32'b00000000000000000101011100010101;
assign LUT_1[46538] = 32'b00000000000000000111111000101010;
assign LUT_1[46539] = 32'b00000000000000000001001010100110;
assign LUT_1[46540] = 32'b00000000000000010100000011110000;
assign LUT_1[46541] = 32'b00000000000000001101010101101100;
assign LUT_1[46542] = 32'b00000000000000001111110010000001;
assign LUT_1[46543] = 32'b00000000000000001001000011111101;
assign LUT_1[46544] = 32'b00000000000000001110111000000110;
assign LUT_1[46545] = 32'b00000000000000001000001010000010;
assign LUT_1[46546] = 32'b00000000000000001010100110010111;
assign LUT_1[46547] = 32'b00000000000000000011111000010011;
assign LUT_1[46548] = 32'b00000000000000010110110001011101;
assign LUT_1[46549] = 32'b00000000000000010000000011011001;
assign LUT_1[46550] = 32'b00000000000000010010011111101110;
assign LUT_1[46551] = 32'b00000000000000001011110001101010;
assign LUT_1[46552] = 32'b00000000000000001110000101111011;
assign LUT_1[46553] = 32'b00000000000000000111010111110111;
assign LUT_1[46554] = 32'b00000000000000001001110100001100;
assign LUT_1[46555] = 32'b00000000000000000011000110001000;
assign LUT_1[46556] = 32'b00000000000000010101111111010010;
assign LUT_1[46557] = 32'b00000000000000001111010001001110;
assign LUT_1[46558] = 32'b00000000000000010001101101100011;
assign LUT_1[46559] = 32'b00000000000000001010111111011111;
assign LUT_1[46560] = 32'b00000000000000001101110111100011;
assign LUT_1[46561] = 32'b00000000000000000111001001011111;
assign LUT_1[46562] = 32'b00000000000000001001100101110100;
assign LUT_1[46563] = 32'b00000000000000000010110111110000;
assign LUT_1[46564] = 32'b00000000000000010101110000111010;
assign LUT_1[46565] = 32'b00000000000000001111000010110110;
assign LUT_1[46566] = 32'b00000000000000010001011111001011;
assign LUT_1[46567] = 32'b00000000000000001010110001000111;
assign LUT_1[46568] = 32'b00000000000000001101000101011000;
assign LUT_1[46569] = 32'b00000000000000000110010111010100;
assign LUT_1[46570] = 32'b00000000000000001000110011101001;
assign LUT_1[46571] = 32'b00000000000000000010000101100101;
assign LUT_1[46572] = 32'b00000000000000010100111110101111;
assign LUT_1[46573] = 32'b00000000000000001110010000101011;
assign LUT_1[46574] = 32'b00000000000000010000101101000000;
assign LUT_1[46575] = 32'b00000000000000001001111110111100;
assign LUT_1[46576] = 32'b00000000000000001111110011000101;
assign LUT_1[46577] = 32'b00000000000000001001000101000001;
assign LUT_1[46578] = 32'b00000000000000001011100001010110;
assign LUT_1[46579] = 32'b00000000000000000100110011010010;
assign LUT_1[46580] = 32'b00000000000000010111101100011100;
assign LUT_1[46581] = 32'b00000000000000010000111110011000;
assign LUT_1[46582] = 32'b00000000000000010011011010101101;
assign LUT_1[46583] = 32'b00000000000000001100101100101001;
assign LUT_1[46584] = 32'b00000000000000001111000000111010;
assign LUT_1[46585] = 32'b00000000000000001000010010110110;
assign LUT_1[46586] = 32'b00000000000000001010101111001011;
assign LUT_1[46587] = 32'b00000000000000000100000001000111;
assign LUT_1[46588] = 32'b00000000000000010110111010010001;
assign LUT_1[46589] = 32'b00000000000000010000001100001101;
assign LUT_1[46590] = 32'b00000000000000010010101000100010;
assign LUT_1[46591] = 32'b00000000000000001011111010011110;
assign LUT_1[46592] = 32'b00000000000000000011111001001010;
assign LUT_1[46593] = 32'b11111111111111111101001011000110;
assign LUT_1[46594] = 32'b11111111111111111111100111011011;
assign LUT_1[46595] = 32'b11111111111111111000111001010111;
assign LUT_1[46596] = 32'b00000000000000001011110010100001;
assign LUT_1[46597] = 32'b00000000000000000101000100011101;
assign LUT_1[46598] = 32'b00000000000000000111100000110010;
assign LUT_1[46599] = 32'b00000000000000000000110010101110;
assign LUT_1[46600] = 32'b00000000000000000011000110111111;
assign LUT_1[46601] = 32'b11111111111111111100011000111011;
assign LUT_1[46602] = 32'b11111111111111111110110101010000;
assign LUT_1[46603] = 32'b11111111111111111000000111001100;
assign LUT_1[46604] = 32'b00000000000000001011000000010110;
assign LUT_1[46605] = 32'b00000000000000000100010010010010;
assign LUT_1[46606] = 32'b00000000000000000110101110100111;
assign LUT_1[46607] = 32'b00000000000000000000000000100011;
assign LUT_1[46608] = 32'b00000000000000000101110100101100;
assign LUT_1[46609] = 32'b11111111111111111111000110101000;
assign LUT_1[46610] = 32'b00000000000000000001100010111101;
assign LUT_1[46611] = 32'b11111111111111111010110100111001;
assign LUT_1[46612] = 32'b00000000000000001101101110000011;
assign LUT_1[46613] = 32'b00000000000000000110111111111111;
assign LUT_1[46614] = 32'b00000000000000001001011100010100;
assign LUT_1[46615] = 32'b00000000000000000010101110010000;
assign LUT_1[46616] = 32'b00000000000000000101000010100001;
assign LUT_1[46617] = 32'b11111111111111111110010100011101;
assign LUT_1[46618] = 32'b00000000000000000000110000110010;
assign LUT_1[46619] = 32'b11111111111111111010000010101110;
assign LUT_1[46620] = 32'b00000000000000001100111011111000;
assign LUT_1[46621] = 32'b00000000000000000110001101110100;
assign LUT_1[46622] = 32'b00000000000000001000101010001001;
assign LUT_1[46623] = 32'b00000000000000000001111100000101;
assign LUT_1[46624] = 32'b00000000000000000100110100001001;
assign LUT_1[46625] = 32'b11111111111111111110000110000101;
assign LUT_1[46626] = 32'b00000000000000000000100010011010;
assign LUT_1[46627] = 32'b11111111111111111001110100010110;
assign LUT_1[46628] = 32'b00000000000000001100101101100000;
assign LUT_1[46629] = 32'b00000000000000000101111111011100;
assign LUT_1[46630] = 32'b00000000000000001000011011110001;
assign LUT_1[46631] = 32'b00000000000000000001101101101101;
assign LUT_1[46632] = 32'b00000000000000000100000001111110;
assign LUT_1[46633] = 32'b11111111111111111101010011111010;
assign LUT_1[46634] = 32'b11111111111111111111110000001111;
assign LUT_1[46635] = 32'b11111111111111111001000010001011;
assign LUT_1[46636] = 32'b00000000000000001011111011010101;
assign LUT_1[46637] = 32'b00000000000000000101001101010001;
assign LUT_1[46638] = 32'b00000000000000000111101001100110;
assign LUT_1[46639] = 32'b00000000000000000000111011100010;
assign LUT_1[46640] = 32'b00000000000000000110101111101011;
assign LUT_1[46641] = 32'b00000000000000000000000001100111;
assign LUT_1[46642] = 32'b00000000000000000010011101111100;
assign LUT_1[46643] = 32'b11111111111111111011101111111000;
assign LUT_1[46644] = 32'b00000000000000001110101001000010;
assign LUT_1[46645] = 32'b00000000000000000111111010111110;
assign LUT_1[46646] = 32'b00000000000000001010010111010011;
assign LUT_1[46647] = 32'b00000000000000000011101001001111;
assign LUT_1[46648] = 32'b00000000000000000101111101100000;
assign LUT_1[46649] = 32'b11111111111111111111001111011100;
assign LUT_1[46650] = 32'b00000000000000000001101011110001;
assign LUT_1[46651] = 32'b11111111111111111010111101101101;
assign LUT_1[46652] = 32'b00000000000000001101110110110111;
assign LUT_1[46653] = 32'b00000000000000000111001000110011;
assign LUT_1[46654] = 32'b00000000000000001001100101001000;
assign LUT_1[46655] = 32'b00000000000000000010110111000100;
assign LUT_1[46656] = 32'b00000000000000000101110110110010;
assign LUT_1[46657] = 32'b11111111111111111111001000101110;
assign LUT_1[46658] = 32'b00000000000000000001100101000011;
assign LUT_1[46659] = 32'b11111111111111111010110110111111;
assign LUT_1[46660] = 32'b00000000000000001101110000001001;
assign LUT_1[46661] = 32'b00000000000000000111000010000101;
assign LUT_1[46662] = 32'b00000000000000001001011110011010;
assign LUT_1[46663] = 32'b00000000000000000010110000010110;
assign LUT_1[46664] = 32'b00000000000000000101000100100111;
assign LUT_1[46665] = 32'b11111111111111111110010110100011;
assign LUT_1[46666] = 32'b00000000000000000000110010111000;
assign LUT_1[46667] = 32'b11111111111111111010000100110100;
assign LUT_1[46668] = 32'b00000000000000001100111101111110;
assign LUT_1[46669] = 32'b00000000000000000110001111111010;
assign LUT_1[46670] = 32'b00000000000000001000101100001111;
assign LUT_1[46671] = 32'b00000000000000000001111110001011;
assign LUT_1[46672] = 32'b00000000000000000111110010010100;
assign LUT_1[46673] = 32'b00000000000000000001000100010000;
assign LUT_1[46674] = 32'b00000000000000000011100000100101;
assign LUT_1[46675] = 32'b11111111111111111100110010100001;
assign LUT_1[46676] = 32'b00000000000000001111101011101011;
assign LUT_1[46677] = 32'b00000000000000001000111101100111;
assign LUT_1[46678] = 32'b00000000000000001011011001111100;
assign LUT_1[46679] = 32'b00000000000000000100101011111000;
assign LUT_1[46680] = 32'b00000000000000000111000000001001;
assign LUT_1[46681] = 32'b00000000000000000000010010000101;
assign LUT_1[46682] = 32'b00000000000000000010101110011010;
assign LUT_1[46683] = 32'b11111111111111111100000000010110;
assign LUT_1[46684] = 32'b00000000000000001110111001100000;
assign LUT_1[46685] = 32'b00000000000000001000001011011100;
assign LUT_1[46686] = 32'b00000000000000001010100111110001;
assign LUT_1[46687] = 32'b00000000000000000011111001101101;
assign LUT_1[46688] = 32'b00000000000000000110110001110001;
assign LUT_1[46689] = 32'b00000000000000000000000011101101;
assign LUT_1[46690] = 32'b00000000000000000010100000000010;
assign LUT_1[46691] = 32'b11111111111111111011110001111110;
assign LUT_1[46692] = 32'b00000000000000001110101011001000;
assign LUT_1[46693] = 32'b00000000000000000111111101000100;
assign LUT_1[46694] = 32'b00000000000000001010011001011001;
assign LUT_1[46695] = 32'b00000000000000000011101011010101;
assign LUT_1[46696] = 32'b00000000000000000101111111100110;
assign LUT_1[46697] = 32'b11111111111111111111010001100010;
assign LUT_1[46698] = 32'b00000000000000000001101101110111;
assign LUT_1[46699] = 32'b11111111111111111010111111110011;
assign LUT_1[46700] = 32'b00000000000000001101111000111101;
assign LUT_1[46701] = 32'b00000000000000000111001010111001;
assign LUT_1[46702] = 32'b00000000000000001001100111001110;
assign LUT_1[46703] = 32'b00000000000000000010111001001010;
assign LUT_1[46704] = 32'b00000000000000001000101101010011;
assign LUT_1[46705] = 32'b00000000000000000001111111001111;
assign LUT_1[46706] = 32'b00000000000000000100011011100100;
assign LUT_1[46707] = 32'b11111111111111111101101101100000;
assign LUT_1[46708] = 32'b00000000000000010000100110101010;
assign LUT_1[46709] = 32'b00000000000000001001111000100110;
assign LUT_1[46710] = 32'b00000000000000001100010100111011;
assign LUT_1[46711] = 32'b00000000000000000101100110110111;
assign LUT_1[46712] = 32'b00000000000000000111111011001000;
assign LUT_1[46713] = 32'b00000000000000000001001101000100;
assign LUT_1[46714] = 32'b00000000000000000011101001011001;
assign LUT_1[46715] = 32'b11111111111111111100111011010101;
assign LUT_1[46716] = 32'b00000000000000001111110100011111;
assign LUT_1[46717] = 32'b00000000000000001001000110011011;
assign LUT_1[46718] = 32'b00000000000000001011100010110000;
assign LUT_1[46719] = 32'b00000000000000000100110100101100;
assign LUT_1[46720] = 32'b00000000000000000110111001001101;
assign LUT_1[46721] = 32'b00000000000000000000001011001001;
assign LUT_1[46722] = 32'b00000000000000000010100111011110;
assign LUT_1[46723] = 32'b11111111111111111011111001011010;
assign LUT_1[46724] = 32'b00000000000000001110110010100100;
assign LUT_1[46725] = 32'b00000000000000001000000100100000;
assign LUT_1[46726] = 32'b00000000000000001010100000110101;
assign LUT_1[46727] = 32'b00000000000000000011110010110001;
assign LUT_1[46728] = 32'b00000000000000000110000111000010;
assign LUT_1[46729] = 32'b11111111111111111111011000111110;
assign LUT_1[46730] = 32'b00000000000000000001110101010011;
assign LUT_1[46731] = 32'b11111111111111111011000111001111;
assign LUT_1[46732] = 32'b00000000000000001110000000011001;
assign LUT_1[46733] = 32'b00000000000000000111010010010101;
assign LUT_1[46734] = 32'b00000000000000001001101110101010;
assign LUT_1[46735] = 32'b00000000000000000011000000100110;
assign LUT_1[46736] = 32'b00000000000000001000110100101111;
assign LUT_1[46737] = 32'b00000000000000000010000110101011;
assign LUT_1[46738] = 32'b00000000000000000100100011000000;
assign LUT_1[46739] = 32'b11111111111111111101110100111100;
assign LUT_1[46740] = 32'b00000000000000010000101110000110;
assign LUT_1[46741] = 32'b00000000000000001010000000000010;
assign LUT_1[46742] = 32'b00000000000000001100011100010111;
assign LUT_1[46743] = 32'b00000000000000000101101110010011;
assign LUT_1[46744] = 32'b00000000000000001000000010100100;
assign LUT_1[46745] = 32'b00000000000000000001010100100000;
assign LUT_1[46746] = 32'b00000000000000000011110000110101;
assign LUT_1[46747] = 32'b11111111111111111101000010110001;
assign LUT_1[46748] = 32'b00000000000000001111111011111011;
assign LUT_1[46749] = 32'b00000000000000001001001101110111;
assign LUT_1[46750] = 32'b00000000000000001011101010001100;
assign LUT_1[46751] = 32'b00000000000000000100111100001000;
assign LUT_1[46752] = 32'b00000000000000000111110100001100;
assign LUT_1[46753] = 32'b00000000000000000001000110001000;
assign LUT_1[46754] = 32'b00000000000000000011100010011101;
assign LUT_1[46755] = 32'b11111111111111111100110100011001;
assign LUT_1[46756] = 32'b00000000000000001111101101100011;
assign LUT_1[46757] = 32'b00000000000000001000111111011111;
assign LUT_1[46758] = 32'b00000000000000001011011011110100;
assign LUT_1[46759] = 32'b00000000000000000100101101110000;
assign LUT_1[46760] = 32'b00000000000000000111000010000001;
assign LUT_1[46761] = 32'b00000000000000000000010011111101;
assign LUT_1[46762] = 32'b00000000000000000010110000010010;
assign LUT_1[46763] = 32'b11111111111111111100000010001110;
assign LUT_1[46764] = 32'b00000000000000001110111011011000;
assign LUT_1[46765] = 32'b00000000000000001000001101010100;
assign LUT_1[46766] = 32'b00000000000000001010101001101001;
assign LUT_1[46767] = 32'b00000000000000000011111011100101;
assign LUT_1[46768] = 32'b00000000000000001001101111101110;
assign LUT_1[46769] = 32'b00000000000000000011000001101010;
assign LUT_1[46770] = 32'b00000000000000000101011101111111;
assign LUT_1[46771] = 32'b11111111111111111110101111111011;
assign LUT_1[46772] = 32'b00000000000000010001101001000101;
assign LUT_1[46773] = 32'b00000000000000001010111011000001;
assign LUT_1[46774] = 32'b00000000000000001101010111010110;
assign LUT_1[46775] = 32'b00000000000000000110101001010010;
assign LUT_1[46776] = 32'b00000000000000001000111101100011;
assign LUT_1[46777] = 32'b00000000000000000010001111011111;
assign LUT_1[46778] = 32'b00000000000000000100101011110100;
assign LUT_1[46779] = 32'b11111111111111111101111101110000;
assign LUT_1[46780] = 32'b00000000000000010000110110111010;
assign LUT_1[46781] = 32'b00000000000000001010001000110110;
assign LUT_1[46782] = 32'b00000000000000001100100101001011;
assign LUT_1[46783] = 32'b00000000000000000101110111000111;
assign LUT_1[46784] = 32'b00000000000000001000110110110101;
assign LUT_1[46785] = 32'b00000000000000000010001000110001;
assign LUT_1[46786] = 32'b00000000000000000100100101000110;
assign LUT_1[46787] = 32'b11111111111111111101110111000010;
assign LUT_1[46788] = 32'b00000000000000010000110000001100;
assign LUT_1[46789] = 32'b00000000000000001010000010001000;
assign LUT_1[46790] = 32'b00000000000000001100011110011101;
assign LUT_1[46791] = 32'b00000000000000000101110000011001;
assign LUT_1[46792] = 32'b00000000000000001000000100101010;
assign LUT_1[46793] = 32'b00000000000000000001010110100110;
assign LUT_1[46794] = 32'b00000000000000000011110010111011;
assign LUT_1[46795] = 32'b11111111111111111101000100110111;
assign LUT_1[46796] = 32'b00000000000000001111111110000001;
assign LUT_1[46797] = 32'b00000000000000001001001111111101;
assign LUT_1[46798] = 32'b00000000000000001011101100010010;
assign LUT_1[46799] = 32'b00000000000000000100111110001110;
assign LUT_1[46800] = 32'b00000000000000001010110010010111;
assign LUT_1[46801] = 32'b00000000000000000100000100010011;
assign LUT_1[46802] = 32'b00000000000000000110100000101000;
assign LUT_1[46803] = 32'b11111111111111111111110010100100;
assign LUT_1[46804] = 32'b00000000000000010010101011101110;
assign LUT_1[46805] = 32'b00000000000000001011111101101010;
assign LUT_1[46806] = 32'b00000000000000001110011001111111;
assign LUT_1[46807] = 32'b00000000000000000111101011111011;
assign LUT_1[46808] = 32'b00000000000000001010000000001100;
assign LUT_1[46809] = 32'b00000000000000000011010010001000;
assign LUT_1[46810] = 32'b00000000000000000101101110011101;
assign LUT_1[46811] = 32'b11111111111111111111000000011001;
assign LUT_1[46812] = 32'b00000000000000010001111001100011;
assign LUT_1[46813] = 32'b00000000000000001011001011011111;
assign LUT_1[46814] = 32'b00000000000000001101100111110100;
assign LUT_1[46815] = 32'b00000000000000000110111001110000;
assign LUT_1[46816] = 32'b00000000000000001001110001110100;
assign LUT_1[46817] = 32'b00000000000000000011000011110000;
assign LUT_1[46818] = 32'b00000000000000000101100000000101;
assign LUT_1[46819] = 32'b11111111111111111110110010000001;
assign LUT_1[46820] = 32'b00000000000000010001101011001011;
assign LUT_1[46821] = 32'b00000000000000001010111101000111;
assign LUT_1[46822] = 32'b00000000000000001101011001011100;
assign LUT_1[46823] = 32'b00000000000000000110101011011000;
assign LUT_1[46824] = 32'b00000000000000001000111111101001;
assign LUT_1[46825] = 32'b00000000000000000010010001100101;
assign LUT_1[46826] = 32'b00000000000000000100101101111010;
assign LUT_1[46827] = 32'b11111111111111111101111111110110;
assign LUT_1[46828] = 32'b00000000000000010000111001000000;
assign LUT_1[46829] = 32'b00000000000000001010001010111100;
assign LUT_1[46830] = 32'b00000000000000001100100111010001;
assign LUT_1[46831] = 32'b00000000000000000101111001001101;
assign LUT_1[46832] = 32'b00000000000000001011101101010110;
assign LUT_1[46833] = 32'b00000000000000000100111111010010;
assign LUT_1[46834] = 32'b00000000000000000111011011100111;
assign LUT_1[46835] = 32'b00000000000000000000101101100011;
assign LUT_1[46836] = 32'b00000000000000010011100110101101;
assign LUT_1[46837] = 32'b00000000000000001100111000101001;
assign LUT_1[46838] = 32'b00000000000000001111010100111110;
assign LUT_1[46839] = 32'b00000000000000001000100110111010;
assign LUT_1[46840] = 32'b00000000000000001010111011001011;
assign LUT_1[46841] = 32'b00000000000000000100001101000111;
assign LUT_1[46842] = 32'b00000000000000000110101001011100;
assign LUT_1[46843] = 32'b11111111111111111111111011011000;
assign LUT_1[46844] = 32'b00000000000000010010110100100010;
assign LUT_1[46845] = 32'b00000000000000001100000110011110;
assign LUT_1[46846] = 32'b00000000000000001110100010110011;
assign LUT_1[46847] = 32'b00000000000000000111110100101111;
assign LUT_1[46848] = 32'b00000000000000000001101101010110;
assign LUT_1[46849] = 32'b11111111111111111010111111010010;
assign LUT_1[46850] = 32'b11111111111111111101011011100111;
assign LUT_1[46851] = 32'b11111111111111110110101101100011;
assign LUT_1[46852] = 32'b00000000000000001001100110101101;
assign LUT_1[46853] = 32'b00000000000000000010111000101001;
assign LUT_1[46854] = 32'b00000000000000000101010100111110;
assign LUT_1[46855] = 32'b11111111111111111110100110111010;
assign LUT_1[46856] = 32'b00000000000000000000111011001011;
assign LUT_1[46857] = 32'b11111111111111111010001101000111;
assign LUT_1[46858] = 32'b11111111111111111100101001011100;
assign LUT_1[46859] = 32'b11111111111111110101111011011000;
assign LUT_1[46860] = 32'b00000000000000001000110100100010;
assign LUT_1[46861] = 32'b00000000000000000010000110011110;
assign LUT_1[46862] = 32'b00000000000000000100100010110011;
assign LUT_1[46863] = 32'b11111111111111111101110100101111;
assign LUT_1[46864] = 32'b00000000000000000011101000111000;
assign LUT_1[46865] = 32'b11111111111111111100111010110100;
assign LUT_1[46866] = 32'b11111111111111111111010111001001;
assign LUT_1[46867] = 32'b11111111111111111000101001000101;
assign LUT_1[46868] = 32'b00000000000000001011100010001111;
assign LUT_1[46869] = 32'b00000000000000000100110100001011;
assign LUT_1[46870] = 32'b00000000000000000111010000100000;
assign LUT_1[46871] = 32'b00000000000000000000100010011100;
assign LUT_1[46872] = 32'b00000000000000000010110110101101;
assign LUT_1[46873] = 32'b11111111111111111100001000101001;
assign LUT_1[46874] = 32'b11111111111111111110100100111110;
assign LUT_1[46875] = 32'b11111111111111110111110110111010;
assign LUT_1[46876] = 32'b00000000000000001010110000000100;
assign LUT_1[46877] = 32'b00000000000000000100000010000000;
assign LUT_1[46878] = 32'b00000000000000000110011110010101;
assign LUT_1[46879] = 32'b11111111111111111111110000010001;
assign LUT_1[46880] = 32'b00000000000000000010101000010101;
assign LUT_1[46881] = 32'b11111111111111111011111010010001;
assign LUT_1[46882] = 32'b11111111111111111110010110100110;
assign LUT_1[46883] = 32'b11111111111111110111101000100010;
assign LUT_1[46884] = 32'b00000000000000001010100001101100;
assign LUT_1[46885] = 32'b00000000000000000011110011101000;
assign LUT_1[46886] = 32'b00000000000000000110001111111101;
assign LUT_1[46887] = 32'b11111111111111111111100001111001;
assign LUT_1[46888] = 32'b00000000000000000001110110001010;
assign LUT_1[46889] = 32'b11111111111111111011001000000110;
assign LUT_1[46890] = 32'b11111111111111111101100100011011;
assign LUT_1[46891] = 32'b11111111111111110110110110010111;
assign LUT_1[46892] = 32'b00000000000000001001101111100001;
assign LUT_1[46893] = 32'b00000000000000000011000001011101;
assign LUT_1[46894] = 32'b00000000000000000101011101110010;
assign LUT_1[46895] = 32'b11111111111111111110101111101110;
assign LUT_1[46896] = 32'b00000000000000000100100011110111;
assign LUT_1[46897] = 32'b11111111111111111101110101110011;
assign LUT_1[46898] = 32'b00000000000000000000010010001000;
assign LUT_1[46899] = 32'b11111111111111111001100100000100;
assign LUT_1[46900] = 32'b00000000000000001100011101001110;
assign LUT_1[46901] = 32'b00000000000000000101101111001010;
assign LUT_1[46902] = 32'b00000000000000001000001011011111;
assign LUT_1[46903] = 32'b00000000000000000001011101011011;
assign LUT_1[46904] = 32'b00000000000000000011110001101100;
assign LUT_1[46905] = 32'b11111111111111111101000011101000;
assign LUT_1[46906] = 32'b11111111111111111111011111111101;
assign LUT_1[46907] = 32'b11111111111111111000110001111001;
assign LUT_1[46908] = 32'b00000000000000001011101011000011;
assign LUT_1[46909] = 32'b00000000000000000100111100111111;
assign LUT_1[46910] = 32'b00000000000000000111011001010100;
assign LUT_1[46911] = 32'b00000000000000000000101011010000;
assign LUT_1[46912] = 32'b00000000000000000011101010111110;
assign LUT_1[46913] = 32'b11111111111111111100111100111010;
assign LUT_1[46914] = 32'b11111111111111111111011001001111;
assign LUT_1[46915] = 32'b11111111111111111000101011001011;
assign LUT_1[46916] = 32'b00000000000000001011100100010101;
assign LUT_1[46917] = 32'b00000000000000000100110110010001;
assign LUT_1[46918] = 32'b00000000000000000111010010100110;
assign LUT_1[46919] = 32'b00000000000000000000100100100010;
assign LUT_1[46920] = 32'b00000000000000000010111000110011;
assign LUT_1[46921] = 32'b11111111111111111100001010101111;
assign LUT_1[46922] = 32'b11111111111111111110100111000100;
assign LUT_1[46923] = 32'b11111111111111110111111001000000;
assign LUT_1[46924] = 32'b00000000000000001010110010001010;
assign LUT_1[46925] = 32'b00000000000000000100000100000110;
assign LUT_1[46926] = 32'b00000000000000000110100000011011;
assign LUT_1[46927] = 32'b11111111111111111111110010010111;
assign LUT_1[46928] = 32'b00000000000000000101100110100000;
assign LUT_1[46929] = 32'b11111111111111111110111000011100;
assign LUT_1[46930] = 32'b00000000000000000001010100110001;
assign LUT_1[46931] = 32'b11111111111111111010100110101101;
assign LUT_1[46932] = 32'b00000000000000001101011111110111;
assign LUT_1[46933] = 32'b00000000000000000110110001110011;
assign LUT_1[46934] = 32'b00000000000000001001001110001000;
assign LUT_1[46935] = 32'b00000000000000000010100000000100;
assign LUT_1[46936] = 32'b00000000000000000100110100010101;
assign LUT_1[46937] = 32'b11111111111111111110000110010001;
assign LUT_1[46938] = 32'b00000000000000000000100010100110;
assign LUT_1[46939] = 32'b11111111111111111001110100100010;
assign LUT_1[46940] = 32'b00000000000000001100101101101100;
assign LUT_1[46941] = 32'b00000000000000000101111111101000;
assign LUT_1[46942] = 32'b00000000000000001000011011111101;
assign LUT_1[46943] = 32'b00000000000000000001101101111001;
assign LUT_1[46944] = 32'b00000000000000000100100101111101;
assign LUT_1[46945] = 32'b11111111111111111101110111111001;
assign LUT_1[46946] = 32'b00000000000000000000010100001110;
assign LUT_1[46947] = 32'b11111111111111111001100110001010;
assign LUT_1[46948] = 32'b00000000000000001100011111010100;
assign LUT_1[46949] = 32'b00000000000000000101110001010000;
assign LUT_1[46950] = 32'b00000000000000001000001101100101;
assign LUT_1[46951] = 32'b00000000000000000001011111100001;
assign LUT_1[46952] = 32'b00000000000000000011110011110010;
assign LUT_1[46953] = 32'b11111111111111111101000101101110;
assign LUT_1[46954] = 32'b11111111111111111111100010000011;
assign LUT_1[46955] = 32'b11111111111111111000110011111111;
assign LUT_1[46956] = 32'b00000000000000001011101101001001;
assign LUT_1[46957] = 32'b00000000000000000100111111000101;
assign LUT_1[46958] = 32'b00000000000000000111011011011010;
assign LUT_1[46959] = 32'b00000000000000000000101101010110;
assign LUT_1[46960] = 32'b00000000000000000110100001011111;
assign LUT_1[46961] = 32'b11111111111111111111110011011011;
assign LUT_1[46962] = 32'b00000000000000000010001111110000;
assign LUT_1[46963] = 32'b11111111111111111011100001101100;
assign LUT_1[46964] = 32'b00000000000000001110011010110110;
assign LUT_1[46965] = 32'b00000000000000000111101100110010;
assign LUT_1[46966] = 32'b00000000000000001010001001000111;
assign LUT_1[46967] = 32'b00000000000000000011011011000011;
assign LUT_1[46968] = 32'b00000000000000000101101111010100;
assign LUT_1[46969] = 32'b11111111111111111111000001010000;
assign LUT_1[46970] = 32'b00000000000000000001011101100101;
assign LUT_1[46971] = 32'b11111111111111111010101111100001;
assign LUT_1[46972] = 32'b00000000000000001101101000101011;
assign LUT_1[46973] = 32'b00000000000000000110111010100111;
assign LUT_1[46974] = 32'b00000000000000001001010110111100;
assign LUT_1[46975] = 32'b00000000000000000010101000111000;
assign LUT_1[46976] = 32'b00000000000000000100101101011001;
assign LUT_1[46977] = 32'b11111111111111111101111111010101;
assign LUT_1[46978] = 32'b00000000000000000000011011101010;
assign LUT_1[46979] = 32'b11111111111111111001101101100110;
assign LUT_1[46980] = 32'b00000000000000001100100110110000;
assign LUT_1[46981] = 32'b00000000000000000101111000101100;
assign LUT_1[46982] = 32'b00000000000000001000010101000001;
assign LUT_1[46983] = 32'b00000000000000000001100110111101;
assign LUT_1[46984] = 32'b00000000000000000011111011001110;
assign LUT_1[46985] = 32'b11111111111111111101001101001010;
assign LUT_1[46986] = 32'b11111111111111111111101001011111;
assign LUT_1[46987] = 32'b11111111111111111000111011011011;
assign LUT_1[46988] = 32'b00000000000000001011110100100101;
assign LUT_1[46989] = 32'b00000000000000000101000110100001;
assign LUT_1[46990] = 32'b00000000000000000111100010110110;
assign LUT_1[46991] = 32'b00000000000000000000110100110010;
assign LUT_1[46992] = 32'b00000000000000000110101000111011;
assign LUT_1[46993] = 32'b11111111111111111111111010110111;
assign LUT_1[46994] = 32'b00000000000000000010010111001100;
assign LUT_1[46995] = 32'b11111111111111111011101001001000;
assign LUT_1[46996] = 32'b00000000000000001110100010010010;
assign LUT_1[46997] = 32'b00000000000000000111110100001110;
assign LUT_1[46998] = 32'b00000000000000001010010000100011;
assign LUT_1[46999] = 32'b00000000000000000011100010011111;
assign LUT_1[47000] = 32'b00000000000000000101110110110000;
assign LUT_1[47001] = 32'b11111111111111111111001000101100;
assign LUT_1[47002] = 32'b00000000000000000001100101000001;
assign LUT_1[47003] = 32'b11111111111111111010110110111101;
assign LUT_1[47004] = 32'b00000000000000001101110000000111;
assign LUT_1[47005] = 32'b00000000000000000111000010000011;
assign LUT_1[47006] = 32'b00000000000000001001011110011000;
assign LUT_1[47007] = 32'b00000000000000000010110000010100;
assign LUT_1[47008] = 32'b00000000000000000101101000011000;
assign LUT_1[47009] = 32'b11111111111111111110111010010100;
assign LUT_1[47010] = 32'b00000000000000000001010110101001;
assign LUT_1[47011] = 32'b11111111111111111010101000100101;
assign LUT_1[47012] = 32'b00000000000000001101100001101111;
assign LUT_1[47013] = 32'b00000000000000000110110011101011;
assign LUT_1[47014] = 32'b00000000000000001001010000000000;
assign LUT_1[47015] = 32'b00000000000000000010100001111100;
assign LUT_1[47016] = 32'b00000000000000000100110110001101;
assign LUT_1[47017] = 32'b11111111111111111110001000001001;
assign LUT_1[47018] = 32'b00000000000000000000100100011110;
assign LUT_1[47019] = 32'b11111111111111111001110110011010;
assign LUT_1[47020] = 32'b00000000000000001100101111100100;
assign LUT_1[47021] = 32'b00000000000000000110000001100000;
assign LUT_1[47022] = 32'b00000000000000001000011101110101;
assign LUT_1[47023] = 32'b00000000000000000001101111110001;
assign LUT_1[47024] = 32'b00000000000000000111100011111010;
assign LUT_1[47025] = 32'b00000000000000000000110101110110;
assign LUT_1[47026] = 32'b00000000000000000011010010001011;
assign LUT_1[47027] = 32'b11111111111111111100100100000111;
assign LUT_1[47028] = 32'b00000000000000001111011101010001;
assign LUT_1[47029] = 32'b00000000000000001000101111001101;
assign LUT_1[47030] = 32'b00000000000000001011001011100010;
assign LUT_1[47031] = 32'b00000000000000000100011101011110;
assign LUT_1[47032] = 32'b00000000000000000110110001101111;
assign LUT_1[47033] = 32'b00000000000000000000000011101011;
assign LUT_1[47034] = 32'b00000000000000000010100000000000;
assign LUT_1[47035] = 32'b11111111111111111011110001111100;
assign LUT_1[47036] = 32'b00000000000000001110101011000110;
assign LUT_1[47037] = 32'b00000000000000000111111101000010;
assign LUT_1[47038] = 32'b00000000000000001010011001010111;
assign LUT_1[47039] = 32'b00000000000000000011101011010011;
assign LUT_1[47040] = 32'b00000000000000000110101011000001;
assign LUT_1[47041] = 32'b11111111111111111111111100111101;
assign LUT_1[47042] = 32'b00000000000000000010011001010010;
assign LUT_1[47043] = 32'b11111111111111111011101011001110;
assign LUT_1[47044] = 32'b00000000000000001110100100011000;
assign LUT_1[47045] = 32'b00000000000000000111110110010100;
assign LUT_1[47046] = 32'b00000000000000001010010010101001;
assign LUT_1[47047] = 32'b00000000000000000011100100100101;
assign LUT_1[47048] = 32'b00000000000000000101111000110110;
assign LUT_1[47049] = 32'b11111111111111111111001010110010;
assign LUT_1[47050] = 32'b00000000000000000001100111000111;
assign LUT_1[47051] = 32'b11111111111111111010111001000011;
assign LUT_1[47052] = 32'b00000000000000001101110010001101;
assign LUT_1[47053] = 32'b00000000000000000111000100001001;
assign LUT_1[47054] = 32'b00000000000000001001100000011110;
assign LUT_1[47055] = 32'b00000000000000000010110010011010;
assign LUT_1[47056] = 32'b00000000000000001000100110100011;
assign LUT_1[47057] = 32'b00000000000000000001111000011111;
assign LUT_1[47058] = 32'b00000000000000000100010100110100;
assign LUT_1[47059] = 32'b11111111111111111101100110110000;
assign LUT_1[47060] = 32'b00000000000000010000011111111010;
assign LUT_1[47061] = 32'b00000000000000001001110001110110;
assign LUT_1[47062] = 32'b00000000000000001100001110001011;
assign LUT_1[47063] = 32'b00000000000000000101100000000111;
assign LUT_1[47064] = 32'b00000000000000000111110100011000;
assign LUT_1[47065] = 32'b00000000000000000001000110010100;
assign LUT_1[47066] = 32'b00000000000000000011100010101001;
assign LUT_1[47067] = 32'b11111111111111111100110100100101;
assign LUT_1[47068] = 32'b00000000000000001111101101101111;
assign LUT_1[47069] = 32'b00000000000000001000111111101011;
assign LUT_1[47070] = 32'b00000000000000001011011100000000;
assign LUT_1[47071] = 32'b00000000000000000100101101111100;
assign LUT_1[47072] = 32'b00000000000000000111100110000000;
assign LUT_1[47073] = 32'b00000000000000000000110111111100;
assign LUT_1[47074] = 32'b00000000000000000011010100010001;
assign LUT_1[47075] = 32'b11111111111111111100100110001101;
assign LUT_1[47076] = 32'b00000000000000001111011111010111;
assign LUT_1[47077] = 32'b00000000000000001000110001010011;
assign LUT_1[47078] = 32'b00000000000000001011001101101000;
assign LUT_1[47079] = 32'b00000000000000000100011111100100;
assign LUT_1[47080] = 32'b00000000000000000110110011110101;
assign LUT_1[47081] = 32'b00000000000000000000000101110001;
assign LUT_1[47082] = 32'b00000000000000000010100010000110;
assign LUT_1[47083] = 32'b11111111111111111011110100000010;
assign LUT_1[47084] = 32'b00000000000000001110101101001100;
assign LUT_1[47085] = 32'b00000000000000000111111111001000;
assign LUT_1[47086] = 32'b00000000000000001010011011011101;
assign LUT_1[47087] = 32'b00000000000000000011101101011001;
assign LUT_1[47088] = 32'b00000000000000001001100001100010;
assign LUT_1[47089] = 32'b00000000000000000010110011011110;
assign LUT_1[47090] = 32'b00000000000000000101001111110011;
assign LUT_1[47091] = 32'b11111111111111111110100001101111;
assign LUT_1[47092] = 32'b00000000000000010001011010111001;
assign LUT_1[47093] = 32'b00000000000000001010101100110101;
assign LUT_1[47094] = 32'b00000000000000001101001001001010;
assign LUT_1[47095] = 32'b00000000000000000110011011000110;
assign LUT_1[47096] = 32'b00000000000000001000101111010111;
assign LUT_1[47097] = 32'b00000000000000000010000001010011;
assign LUT_1[47098] = 32'b00000000000000000100011101101000;
assign LUT_1[47099] = 32'b11111111111111111101101111100100;
assign LUT_1[47100] = 32'b00000000000000010000101000101110;
assign LUT_1[47101] = 32'b00000000000000001001111010101010;
assign LUT_1[47102] = 32'b00000000000000001100010110111111;
assign LUT_1[47103] = 32'b00000000000000000101101000111011;
assign LUT_1[47104] = 32'b00000000000000000100110101111000;
assign LUT_1[47105] = 32'b11111111111111111110000111110100;
assign LUT_1[47106] = 32'b00000000000000000000100100001001;
assign LUT_1[47107] = 32'b11111111111111111001110110000101;
assign LUT_1[47108] = 32'b00000000000000001100101111001111;
assign LUT_1[47109] = 32'b00000000000000000110000001001011;
assign LUT_1[47110] = 32'b00000000000000001000011101100000;
assign LUT_1[47111] = 32'b00000000000000000001101111011100;
assign LUT_1[47112] = 32'b00000000000000000100000011101101;
assign LUT_1[47113] = 32'b11111111111111111101010101101001;
assign LUT_1[47114] = 32'b11111111111111111111110001111110;
assign LUT_1[47115] = 32'b11111111111111111001000011111010;
assign LUT_1[47116] = 32'b00000000000000001011111101000100;
assign LUT_1[47117] = 32'b00000000000000000101001111000000;
assign LUT_1[47118] = 32'b00000000000000000111101011010101;
assign LUT_1[47119] = 32'b00000000000000000000111101010001;
assign LUT_1[47120] = 32'b00000000000000000110110001011010;
assign LUT_1[47121] = 32'b00000000000000000000000011010110;
assign LUT_1[47122] = 32'b00000000000000000010011111101011;
assign LUT_1[47123] = 32'b11111111111111111011110001100111;
assign LUT_1[47124] = 32'b00000000000000001110101010110001;
assign LUT_1[47125] = 32'b00000000000000000111111100101101;
assign LUT_1[47126] = 32'b00000000000000001010011001000010;
assign LUT_1[47127] = 32'b00000000000000000011101010111110;
assign LUT_1[47128] = 32'b00000000000000000101111111001111;
assign LUT_1[47129] = 32'b11111111111111111111010001001011;
assign LUT_1[47130] = 32'b00000000000000000001101101100000;
assign LUT_1[47131] = 32'b11111111111111111010111111011100;
assign LUT_1[47132] = 32'b00000000000000001101111000100110;
assign LUT_1[47133] = 32'b00000000000000000111001010100010;
assign LUT_1[47134] = 32'b00000000000000001001100110110111;
assign LUT_1[47135] = 32'b00000000000000000010111000110011;
assign LUT_1[47136] = 32'b00000000000000000101110000110111;
assign LUT_1[47137] = 32'b11111111111111111111000010110011;
assign LUT_1[47138] = 32'b00000000000000000001011111001000;
assign LUT_1[47139] = 32'b11111111111111111010110001000100;
assign LUT_1[47140] = 32'b00000000000000001101101010001110;
assign LUT_1[47141] = 32'b00000000000000000110111100001010;
assign LUT_1[47142] = 32'b00000000000000001001011000011111;
assign LUT_1[47143] = 32'b00000000000000000010101010011011;
assign LUT_1[47144] = 32'b00000000000000000100111110101100;
assign LUT_1[47145] = 32'b11111111111111111110010000101000;
assign LUT_1[47146] = 32'b00000000000000000000101100111101;
assign LUT_1[47147] = 32'b11111111111111111001111110111001;
assign LUT_1[47148] = 32'b00000000000000001100111000000011;
assign LUT_1[47149] = 32'b00000000000000000110001001111111;
assign LUT_1[47150] = 32'b00000000000000001000100110010100;
assign LUT_1[47151] = 32'b00000000000000000001111000010000;
assign LUT_1[47152] = 32'b00000000000000000111101100011001;
assign LUT_1[47153] = 32'b00000000000000000000111110010101;
assign LUT_1[47154] = 32'b00000000000000000011011010101010;
assign LUT_1[47155] = 32'b11111111111111111100101100100110;
assign LUT_1[47156] = 32'b00000000000000001111100101110000;
assign LUT_1[47157] = 32'b00000000000000001000110111101100;
assign LUT_1[47158] = 32'b00000000000000001011010100000001;
assign LUT_1[47159] = 32'b00000000000000000100100101111101;
assign LUT_1[47160] = 32'b00000000000000000110111010001110;
assign LUT_1[47161] = 32'b00000000000000000000001100001010;
assign LUT_1[47162] = 32'b00000000000000000010101000011111;
assign LUT_1[47163] = 32'b11111111111111111011111010011011;
assign LUT_1[47164] = 32'b00000000000000001110110011100101;
assign LUT_1[47165] = 32'b00000000000000001000000101100001;
assign LUT_1[47166] = 32'b00000000000000001010100001110110;
assign LUT_1[47167] = 32'b00000000000000000011110011110010;
assign LUT_1[47168] = 32'b00000000000000000110110011100000;
assign LUT_1[47169] = 32'b00000000000000000000000101011100;
assign LUT_1[47170] = 32'b00000000000000000010100001110001;
assign LUT_1[47171] = 32'b11111111111111111011110011101101;
assign LUT_1[47172] = 32'b00000000000000001110101100110111;
assign LUT_1[47173] = 32'b00000000000000000111111110110011;
assign LUT_1[47174] = 32'b00000000000000001010011011001000;
assign LUT_1[47175] = 32'b00000000000000000011101101000100;
assign LUT_1[47176] = 32'b00000000000000000110000001010101;
assign LUT_1[47177] = 32'b11111111111111111111010011010001;
assign LUT_1[47178] = 32'b00000000000000000001101111100110;
assign LUT_1[47179] = 32'b11111111111111111011000001100010;
assign LUT_1[47180] = 32'b00000000000000001101111010101100;
assign LUT_1[47181] = 32'b00000000000000000111001100101000;
assign LUT_1[47182] = 32'b00000000000000001001101000111101;
assign LUT_1[47183] = 32'b00000000000000000010111010111001;
assign LUT_1[47184] = 32'b00000000000000001000101111000010;
assign LUT_1[47185] = 32'b00000000000000000010000000111110;
assign LUT_1[47186] = 32'b00000000000000000100011101010011;
assign LUT_1[47187] = 32'b11111111111111111101101111001111;
assign LUT_1[47188] = 32'b00000000000000010000101000011001;
assign LUT_1[47189] = 32'b00000000000000001001111010010101;
assign LUT_1[47190] = 32'b00000000000000001100010110101010;
assign LUT_1[47191] = 32'b00000000000000000101101000100110;
assign LUT_1[47192] = 32'b00000000000000000111111100110111;
assign LUT_1[47193] = 32'b00000000000000000001001110110011;
assign LUT_1[47194] = 32'b00000000000000000011101011001000;
assign LUT_1[47195] = 32'b11111111111111111100111101000100;
assign LUT_1[47196] = 32'b00000000000000001111110110001110;
assign LUT_1[47197] = 32'b00000000000000001001001000001010;
assign LUT_1[47198] = 32'b00000000000000001011100100011111;
assign LUT_1[47199] = 32'b00000000000000000100110110011011;
assign LUT_1[47200] = 32'b00000000000000000111101110011111;
assign LUT_1[47201] = 32'b00000000000000000001000000011011;
assign LUT_1[47202] = 32'b00000000000000000011011100110000;
assign LUT_1[47203] = 32'b11111111111111111100101110101100;
assign LUT_1[47204] = 32'b00000000000000001111100111110110;
assign LUT_1[47205] = 32'b00000000000000001000111001110010;
assign LUT_1[47206] = 32'b00000000000000001011010110000111;
assign LUT_1[47207] = 32'b00000000000000000100101000000011;
assign LUT_1[47208] = 32'b00000000000000000110111100010100;
assign LUT_1[47209] = 32'b00000000000000000000001110010000;
assign LUT_1[47210] = 32'b00000000000000000010101010100101;
assign LUT_1[47211] = 32'b11111111111111111011111100100001;
assign LUT_1[47212] = 32'b00000000000000001110110101101011;
assign LUT_1[47213] = 32'b00000000000000001000000111100111;
assign LUT_1[47214] = 32'b00000000000000001010100011111100;
assign LUT_1[47215] = 32'b00000000000000000011110101111000;
assign LUT_1[47216] = 32'b00000000000000001001101010000001;
assign LUT_1[47217] = 32'b00000000000000000010111011111101;
assign LUT_1[47218] = 32'b00000000000000000101011000010010;
assign LUT_1[47219] = 32'b11111111111111111110101010001110;
assign LUT_1[47220] = 32'b00000000000000010001100011011000;
assign LUT_1[47221] = 32'b00000000000000001010110101010100;
assign LUT_1[47222] = 32'b00000000000000001101010001101001;
assign LUT_1[47223] = 32'b00000000000000000110100011100101;
assign LUT_1[47224] = 32'b00000000000000001000110111110110;
assign LUT_1[47225] = 32'b00000000000000000010001001110010;
assign LUT_1[47226] = 32'b00000000000000000100100110000111;
assign LUT_1[47227] = 32'b11111111111111111101111000000011;
assign LUT_1[47228] = 32'b00000000000000010000110001001101;
assign LUT_1[47229] = 32'b00000000000000001010000011001001;
assign LUT_1[47230] = 32'b00000000000000001100011111011110;
assign LUT_1[47231] = 32'b00000000000000000101110001011010;
assign LUT_1[47232] = 32'b00000000000000000111110101111011;
assign LUT_1[47233] = 32'b00000000000000000001000111110111;
assign LUT_1[47234] = 32'b00000000000000000011100100001100;
assign LUT_1[47235] = 32'b11111111111111111100110110001000;
assign LUT_1[47236] = 32'b00000000000000001111101111010010;
assign LUT_1[47237] = 32'b00000000000000001001000001001110;
assign LUT_1[47238] = 32'b00000000000000001011011101100011;
assign LUT_1[47239] = 32'b00000000000000000100101111011111;
assign LUT_1[47240] = 32'b00000000000000000111000011110000;
assign LUT_1[47241] = 32'b00000000000000000000010101101100;
assign LUT_1[47242] = 32'b00000000000000000010110010000001;
assign LUT_1[47243] = 32'b11111111111111111100000011111101;
assign LUT_1[47244] = 32'b00000000000000001110111101000111;
assign LUT_1[47245] = 32'b00000000000000001000001111000011;
assign LUT_1[47246] = 32'b00000000000000001010101011011000;
assign LUT_1[47247] = 32'b00000000000000000011111101010100;
assign LUT_1[47248] = 32'b00000000000000001001110001011101;
assign LUT_1[47249] = 32'b00000000000000000011000011011001;
assign LUT_1[47250] = 32'b00000000000000000101011111101110;
assign LUT_1[47251] = 32'b11111111111111111110110001101010;
assign LUT_1[47252] = 32'b00000000000000010001101010110100;
assign LUT_1[47253] = 32'b00000000000000001010111100110000;
assign LUT_1[47254] = 32'b00000000000000001101011001000101;
assign LUT_1[47255] = 32'b00000000000000000110101011000001;
assign LUT_1[47256] = 32'b00000000000000001000111111010010;
assign LUT_1[47257] = 32'b00000000000000000010010001001110;
assign LUT_1[47258] = 32'b00000000000000000100101101100011;
assign LUT_1[47259] = 32'b11111111111111111101111111011111;
assign LUT_1[47260] = 32'b00000000000000010000111000101001;
assign LUT_1[47261] = 32'b00000000000000001010001010100101;
assign LUT_1[47262] = 32'b00000000000000001100100110111010;
assign LUT_1[47263] = 32'b00000000000000000101111000110110;
assign LUT_1[47264] = 32'b00000000000000001000110000111010;
assign LUT_1[47265] = 32'b00000000000000000010000010110110;
assign LUT_1[47266] = 32'b00000000000000000100011111001011;
assign LUT_1[47267] = 32'b11111111111111111101110001000111;
assign LUT_1[47268] = 32'b00000000000000010000101010010001;
assign LUT_1[47269] = 32'b00000000000000001001111100001101;
assign LUT_1[47270] = 32'b00000000000000001100011000100010;
assign LUT_1[47271] = 32'b00000000000000000101101010011110;
assign LUT_1[47272] = 32'b00000000000000000111111110101111;
assign LUT_1[47273] = 32'b00000000000000000001010000101011;
assign LUT_1[47274] = 32'b00000000000000000011101101000000;
assign LUT_1[47275] = 32'b11111111111111111100111110111100;
assign LUT_1[47276] = 32'b00000000000000001111111000000110;
assign LUT_1[47277] = 32'b00000000000000001001001010000010;
assign LUT_1[47278] = 32'b00000000000000001011100110010111;
assign LUT_1[47279] = 32'b00000000000000000100111000010011;
assign LUT_1[47280] = 32'b00000000000000001010101100011100;
assign LUT_1[47281] = 32'b00000000000000000011111110011000;
assign LUT_1[47282] = 32'b00000000000000000110011010101101;
assign LUT_1[47283] = 32'b11111111111111111111101100101001;
assign LUT_1[47284] = 32'b00000000000000010010100101110011;
assign LUT_1[47285] = 32'b00000000000000001011110111101111;
assign LUT_1[47286] = 32'b00000000000000001110010100000100;
assign LUT_1[47287] = 32'b00000000000000000111100110000000;
assign LUT_1[47288] = 32'b00000000000000001001111010010001;
assign LUT_1[47289] = 32'b00000000000000000011001100001101;
assign LUT_1[47290] = 32'b00000000000000000101101000100010;
assign LUT_1[47291] = 32'b11111111111111111110111010011110;
assign LUT_1[47292] = 32'b00000000000000010001110011101000;
assign LUT_1[47293] = 32'b00000000000000001011000101100100;
assign LUT_1[47294] = 32'b00000000000000001101100001111001;
assign LUT_1[47295] = 32'b00000000000000000110110011110101;
assign LUT_1[47296] = 32'b00000000000000001001110011100011;
assign LUT_1[47297] = 32'b00000000000000000011000101011111;
assign LUT_1[47298] = 32'b00000000000000000101100001110100;
assign LUT_1[47299] = 32'b11111111111111111110110011110000;
assign LUT_1[47300] = 32'b00000000000000010001101100111010;
assign LUT_1[47301] = 32'b00000000000000001010111110110110;
assign LUT_1[47302] = 32'b00000000000000001101011011001011;
assign LUT_1[47303] = 32'b00000000000000000110101101000111;
assign LUT_1[47304] = 32'b00000000000000001001000001011000;
assign LUT_1[47305] = 32'b00000000000000000010010011010100;
assign LUT_1[47306] = 32'b00000000000000000100101111101001;
assign LUT_1[47307] = 32'b11111111111111111110000001100101;
assign LUT_1[47308] = 32'b00000000000000010000111010101111;
assign LUT_1[47309] = 32'b00000000000000001010001100101011;
assign LUT_1[47310] = 32'b00000000000000001100101001000000;
assign LUT_1[47311] = 32'b00000000000000000101111010111100;
assign LUT_1[47312] = 32'b00000000000000001011101111000101;
assign LUT_1[47313] = 32'b00000000000000000101000001000001;
assign LUT_1[47314] = 32'b00000000000000000111011101010110;
assign LUT_1[47315] = 32'b00000000000000000000101111010010;
assign LUT_1[47316] = 32'b00000000000000010011101000011100;
assign LUT_1[47317] = 32'b00000000000000001100111010011000;
assign LUT_1[47318] = 32'b00000000000000001111010110101101;
assign LUT_1[47319] = 32'b00000000000000001000101000101001;
assign LUT_1[47320] = 32'b00000000000000001010111100111010;
assign LUT_1[47321] = 32'b00000000000000000100001110110110;
assign LUT_1[47322] = 32'b00000000000000000110101011001011;
assign LUT_1[47323] = 32'b11111111111111111111111101000111;
assign LUT_1[47324] = 32'b00000000000000010010110110010001;
assign LUT_1[47325] = 32'b00000000000000001100001000001101;
assign LUT_1[47326] = 32'b00000000000000001110100100100010;
assign LUT_1[47327] = 32'b00000000000000000111110110011110;
assign LUT_1[47328] = 32'b00000000000000001010101110100010;
assign LUT_1[47329] = 32'b00000000000000000100000000011110;
assign LUT_1[47330] = 32'b00000000000000000110011100110011;
assign LUT_1[47331] = 32'b11111111111111111111101110101111;
assign LUT_1[47332] = 32'b00000000000000010010100111111001;
assign LUT_1[47333] = 32'b00000000000000001011111001110101;
assign LUT_1[47334] = 32'b00000000000000001110010110001010;
assign LUT_1[47335] = 32'b00000000000000000111101000000110;
assign LUT_1[47336] = 32'b00000000000000001001111100010111;
assign LUT_1[47337] = 32'b00000000000000000011001110010011;
assign LUT_1[47338] = 32'b00000000000000000101101010101000;
assign LUT_1[47339] = 32'b11111111111111111110111100100100;
assign LUT_1[47340] = 32'b00000000000000010001110101101110;
assign LUT_1[47341] = 32'b00000000000000001011000111101010;
assign LUT_1[47342] = 32'b00000000000000001101100011111111;
assign LUT_1[47343] = 32'b00000000000000000110110101111011;
assign LUT_1[47344] = 32'b00000000000000001100101010000100;
assign LUT_1[47345] = 32'b00000000000000000101111100000000;
assign LUT_1[47346] = 32'b00000000000000001000011000010101;
assign LUT_1[47347] = 32'b00000000000000000001101010010001;
assign LUT_1[47348] = 32'b00000000000000010100100011011011;
assign LUT_1[47349] = 32'b00000000000000001101110101010111;
assign LUT_1[47350] = 32'b00000000000000010000010001101100;
assign LUT_1[47351] = 32'b00000000000000001001100011101000;
assign LUT_1[47352] = 32'b00000000000000001011110111111001;
assign LUT_1[47353] = 32'b00000000000000000101001001110101;
assign LUT_1[47354] = 32'b00000000000000000111100110001010;
assign LUT_1[47355] = 32'b00000000000000000000111000000110;
assign LUT_1[47356] = 32'b00000000000000010011110001010000;
assign LUT_1[47357] = 32'b00000000000000001101000011001100;
assign LUT_1[47358] = 32'b00000000000000001111011111100001;
assign LUT_1[47359] = 32'b00000000000000001000110001011101;
assign LUT_1[47360] = 32'b00000000000000000010101010000100;
assign LUT_1[47361] = 32'b11111111111111111011111100000000;
assign LUT_1[47362] = 32'b11111111111111111110011000010101;
assign LUT_1[47363] = 32'b11111111111111110111101010010001;
assign LUT_1[47364] = 32'b00000000000000001010100011011011;
assign LUT_1[47365] = 32'b00000000000000000011110101010111;
assign LUT_1[47366] = 32'b00000000000000000110010001101100;
assign LUT_1[47367] = 32'b11111111111111111111100011101000;
assign LUT_1[47368] = 32'b00000000000000000001110111111001;
assign LUT_1[47369] = 32'b11111111111111111011001001110101;
assign LUT_1[47370] = 32'b11111111111111111101100110001010;
assign LUT_1[47371] = 32'b11111111111111110110111000000110;
assign LUT_1[47372] = 32'b00000000000000001001110001010000;
assign LUT_1[47373] = 32'b00000000000000000011000011001100;
assign LUT_1[47374] = 32'b00000000000000000101011111100001;
assign LUT_1[47375] = 32'b11111111111111111110110001011101;
assign LUT_1[47376] = 32'b00000000000000000100100101100110;
assign LUT_1[47377] = 32'b11111111111111111101110111100010;
assign LUT_1[47378] = 32'b00000000000000000000010011110111;
assign LUT_1[47379] = 32'b11111111111111111001100101110011;
assign LUT_1[47380] = 32'b00000000000000001100011110111101;
assign LUT_1[47381] = 32'b00000000000000000101110000111001;
assign LUT_1[47382] = 32'b00000000000000001000001101001110;
assign LUT_1[47383] = 32'b00000000000000000001011111001010;
assign LUT_1[47384] = 32'b00000000000000000011110011011011;
assign LUT_1[47385] = 32'b11111111111111111101000101010111;
assign LUT_1[47386] = 32'b11111111111111111111100001101100;
assign LUT_1[47387] = 32'b11111111111111111000110011101000;
assign LUT_1[47388] = 32'b00000000000000001011101100110010;
assign LUT_1[47389] = 32'b00000000000000000100111110101110;
assign LUT_1[47390] = 32'b00000000000000000111011011000011;
assign LUT_1[47391] = 32'b00000000000000000000101100111111;
assign LUT_1[47392] = 32'b00000000000000000011100101000011;
assign LUT_1[47393] = 32'b11111111111111111100110110111111;
assign LUT_1[47394] = 32'b11111111111111111111010011010100;
assign LUT_1[47395] = 32'b11111111111111111000100101010000;
assign LUT_1[47396] = 32'b00000000000000001011011110011010;
assign LUT_1[47397] = 32'b00000000000000000100110000010110;
assign LUT_1[47398] = 32'b00000000000000000111001100101011;
assign LUT_1[47399] = 32'b00000000000000000000011110100111;
assign LUT_1[47400] = 32'b00000000000000000010110010111000;
assign LUT_1[47401] = 32'b11111111111111111100000100110100;
assign LUT_1[47402] = 32'b11111111111111111110100001001001;
assign LUT_1[47403] = 32'b11111111111111110111110011000101;
assign LUT_1[47404] = 32'b00000000000000001010101100001111;
assign LUT_1[47405] = 32'b00000000000000000011111110001011;
assign LUT_1[47406] = 32'b00000000000000000110011010100000;
assign LUT_1[47407] = 32'b11111111111111111111101100011100;
assign LUT_1[47408] = 32'b00000000000000000101100000100101;
assign LUT_1[47409] = 32'b11111111111111111110110010100001;
assign LUT_1[47410] = 32'b00000000000000000001001110110110;
assign LUT_1[47411] = 32'b11111111111111111010100000110010;
assign LUT_1[47412] = 32'b00000000000000001101011001111100;
assign LUT_1[47413] = 32'b00000000000000000110101011111000;
assign LUT_1[47414] = 32'b00000000000000001001001000001101;
assign LUT_1[47415] = 32'b00000000000000000010011010001001;
assign LUT_1[47416] = 32'b00000000000000000100101110011010;
assign LUT_1[47417] = 32'b11111111111111111110000000010110;
assign LUT_1[47418] = 32'b00000000000000000000011100101011;
assign LUT_1[47419] = 32'b11111111111111111001101110100111;
assign LUT_1[47420] = 32'b00000000000000001100100111110001;
assign LUT_1[47421] = 32'b00000000000000000101111001101101;
assign LUT_1[47422] = 32'b00000000000000001000010110000010;
assign LUT_1[47423] = 32'b00000000000000000001100111111110;
assign LUT_1[47424] = 32'b00000000000000000100100111101100;
assign LUT_1[47425] = 32'b11111111111111111101111001101000;
assign LUT_1[47426] = 32'b00000000000000000000010101111101;
assign LUT_1[47427] = 32'b11111111111111111001100111111001;
assign LUT_1[47428] = 32'b00000000000000001100100001000011;
assign LUT_1[47429] = 32'b00000000000000000101110010111111;
assign LUT_1[47430] = 32'b00000000000000001000001111010100;
assign LUT_1[47431] = 32'b00000000000000000001100001010000;
assign LUT_1[47432] = 32'b00000000000000000011110101100001;
assign LUT_1[47433] = 32'b11111111111111111101000111011101;
assign LUT_1[47434] = 32'b11111111111111111111100011110010;
assign LUT_1[47435] = 32'b11111111111111111000110101101110;
assign LUT_1[47436] = 32'b00000000000000001011101110111000;
assign LUT_1[47437] = 32'b00000000000000000101000000110100;
assign LUT_1[47438] = 32'b00000000000000000111011101001001;
assign LUT_1[47439] = 32'b00000000000000000000101111000101;
assign LUT_1[47440] = 32'b00000000000000000110100011001110;
assign LUT_1[47441] = 32'b11111111111111111111110101001010;
assign LUT_1[47442] = 32'b00000000000000000010010001011111;
assign LUT_1[47443] = 32'b11111111111111111011100011011011;
assign LUT_1[47444] = 32'b00000000000000001110011100100101;
assign LUT_1[47445] = 32'b00000000000000000111101110100001;
assign LUT_1[47446] = 32'b00000000000000001010001010110110;
assign LUT_1[47447] = 32'b00000000000000000011011100110010;
assign LUT_1[47448] = 32'b00000000000000000101110001000011;
assign LUT_1[47449] = 32'b11111111111111111111000010111111;
assign LUT_1[47450] = 32'b00000000000000000001011111010100;
assign LUT_1[47451] = 32'b11111111111111111010110001010000;
assign LUT_1[47452] = 32'b00000000000000001101101010011010;
assign LUT_1[47453] = 32'b00000000000000000110111100010110;
assign LUT_1[47454] = 32'b00000000000000001001011000101011;
assign LUT_1[47455] = 32'b00000000000000000010101010100111;
assign LUT_1[47456] = 32'b00000000000000000101100010101011;
assign LUT_1[47457] = 32'b11111111111111111110110100100111;
assign LUT_1[47458] = 32'b00000000000000000001010000111100;
assign LUT_1[47459] = 32'b11111111111111111010100010111000;
assign LUT_1[47460] = 32'b00000000000000001101011100000010;
assign LUT_1[47461] = 32'b00000000000000000110101101111110;
assign LUT_1[47462] = 32'b00000000000000001001001010010011;
assign LUT_1[47463] = 32'b00000000000000000010011100001111;
assign LUT_1[47464] = 32'b00000000000000000100110000100000;
assign LUT_1[47465] = 32'b11111111111111111110000010011100;
assign LUT_1[47466] = 32'b00000000000000000000011110110001;
assign LUT_1[47467] = 32'b11111111111111111001110000101101;
assign LUT_1[47468] = 32'b00000000000000001100101001110111;
assign LUT_1[47469] = 32'b00000000000000000101111011110011;
assign LUT_1[47470] = 32'b00000000000000001000011000001000;
assign LUT_1[47471] = 32'b00000000000000000001101010000100;
assign LUT_1[47472] = 32'b00000000000000000111011110001101;
assign LUT_1[47473] = 32'b00000000000000000000110000001001;
assign LUT_1[47474] = 32'b00000000000000000011001100011110;
assign LUT_1[47475] = 32'b11111111111111111100011110011010;
assign LUT_1[47476] = 32'b00000000000000001111010111100100;
assign LUT_1[47477] = 32'b00000000000000001000101001100000;
assign LUT_1[47478] = 32'b00000000000000001011000101110101;
assign LUT_1[47479] = 32'b00000000000000000100010111110001;
assign LUT_1[47480] = 32'b00000000000000000110101100000010;
assign LUT_1[47481] = 32'b11111111111111111111111101111110;
assign LUT_1[47482] = 32'b00000000000000000010011010010011;
assign LUT_1[47483] = 32'b11111111111111111011101100001111;
assign LUT_1[47484] = 32'b00000000000000001110100101011001;
assign LUT_1[47485] = 32'b00000000000000000111110111010101;
assign LUT_1[47486] = 32'b00000000000000001010010011101010;
assign LUT_1[47487] = 32'b00000000000000000011100101100110;
assign LUT_1[47488] = 32'b00000000000000000101101010000111;
assign LUT_1[47489] = 32'b11111111111111111110111100000011;
assign LUT_1[47490] = 32'b00000000000000000001011000011000;
assign LUT_1[47491] = 32'b11111111111111111010101010010100;
assign LUT_1[47492] = 32'b00000000000000001101100011011110;
assign LUT_1[47493] = 32'b00000000000000000110110101011010;
assign LUT_1[47494] = 32'b00000000000000001001010001101111;
assign LUT_1[47495] = 32'b00000000000000000010100011101011;
assign LUT_1[47496] = 32'b00000000000000000100110111111100;
assign LUT_1[47497] = 32'b11111111111111111110001001111000;
assign LUT_1[47498] = 32'b00000000000000000000100110001101;
assign LUT_1[47499] = 32'b11111111111111111001111000001001;
assign LUT_1[47500] = 32'b00000000000000001100110001010011;
assign LUT_1[47501] = 32'b00000000000000000110000011001111;
assign LUT_1[47502] = 32'b00000000000000001000011111100100;
assign LUT_1[47503] = 32'b00000000000000000001110001100000;
assign LUT_1[47504] = 32'b00000000000000000111100101101001;
assign LUT_1[47505] = 32'b00000000000000000000110111100101;
assign LUT_1[47506] = 32'b00000000000000000011010011111010;
assign LUT_1[47507] = 32'b11111111111111111100100101110110;
assign LUT_1[47508] = 32'b00000000000000001111011111000000;
assign LUT_1[47509] = 32'b00000000000000001000110000111100;
assign LUT_1[47510] = 32'b00000000000000001011001101010001;
assign LUT_1[47511] = 32'b00000000000000000100011111001101;
assign LUT_1[47512] = 32'b00000000000000000110110011011110;
assign LUT_1[47513] = 32'b00000000000000000000000101011010;
assign LUT_1[47514] = 32'b00000000000000000010100001101111;
assign LUT_1[47515] = 32'b11111111111111111011110011101011;
assign LUT_1[47516] = 32'b00000000000000001110101100110101;
assign LUT_1[47517] = 32'b00000000000000000111111110110001;
assign LUT_1[47518] = 32'b00000000000000001010011011000110;
assign LUT_1[47519] = 32'b00000000000000000011101101000010;
assign LUT_1[47520] = 32'b00000000000000000110100101000110;
assign LUT_1[47521] = 32'b11111111111111111111110111000010;
assign LUT_1[47522] = 32'b00000000000000000010010011010111;
assign LUT_1[47523] = 32'b11111111111111111011100101010011;
assign LUT_1[47524] = 32'b00000000000000001110011110011101;
assign LUT_1[47525] = 32'b00000000000000000111110000011001;
assign LUT_1[47526] = 32'b00000000000000001010001100101110;
assign LUT_1[47527] = 32'b00000000000000000011011110101010;
assign LUT_1[47528] = 32'b00000000000000000101110010111011;
assign LUT_1[47529] = 32'b11111111111111111111000100110111;
assign LUT_1[47530] = 32'b00000000000000000001100001001100;
assign LUT_1[47531] = 32'b11111111111111111010110011001000;
assign LUT_1[47532] = 32'b00000000000000001101101100010010;
assign LUT_1[47533] = 32'b00000000000000000110111110001110;
assign LUT_1[47534] = 32'b00000000000000001001011010100011;
assign LUT_1[47535] = 32'b00000000000000000010101100011111;
assign LUT_1[47536] = 32'b00000000000000001000100000101000;
assign LUT_1[47537] = 32'b00000000000000000001110010100100;
assign LUT_1[47538] = 32'b00000000000000000100001110111001;
assign LUT_1[47539] = 32'b11111111111111111101100000110101;
assign LUT_1[47540] = 32'b00000000000000010000011001111111;
assign LUT_1[47541] = 32'b00000000000000001001101011111011;
assign LUT_1[47542] = 32'b00000000000000001100001000010000;
assign LUT_1[47543] = 32'b00000000000000000101011010001100;
assign LUT_1[47544] = 32'b00000000000000000111101110011101;
assign LUT_1[47545] = 32'b00000000000000000001000000011001;
assign LUT_1[47546] = 32'b00000000000000000011011100101110;
assign LUT_1[47547] = 32'b11111111111111111100101110101010;
assign LUT_1[47548] = 32'b00000000000000001111100111110100;
assign LUT_1[47549] = 32'b00000000000000001000111001110000;
assign LUT_1[47550] = 32'b00000000000000001011010110000101;
assign LUT_1[47551] = 32'b00000000000000000100101000000001;
assign LUT_1[47552] = 32'b00000000000000000111100111101111;
assign LUT_1[47553] = 32'b00000000000000000000111001101011;
assign LUT_1[47554] = 32'b00000000000000000011010110000000;
assign LUT_1[47555] = 32'b11111111111111111100100111111100;
assign LUT_1[47556] = 32'b00000000000000001111100001000110;
assign LUT_1[47557] = 32'b00000000000000001000110011000010;
assign LUT_1[47558] = 32'b00000000000000001011001111010111;
assign LUT_1[47559] = 32'b00000000000000000100100001010011;
assign LUT_1[47560] = 32'b00000000000000000110110101100100;
assign LUT_1[47561] = 32'b00000000000000000000000111100000;
assign LUT_1[47562] = 32'b00000000000000000010100011110101;
assign LUT_1[47563] = 32'b11111111111111111011110101110001;
assign LUT_1[47564] = 32'b00000000000000001110101110111011;
assign LUT_1[47565] = 32'b00000000000000001000000000110111;
assign LUT_1[47566] = 32'b00000000000000001010011101001100;
assign LUT_1[47567] = 32'b00000000000000000011101111001000;
assign LUT_1[47568] = 32'b00000000000000001001100011010001;
assign LUT_1[47569] = 32'b00000000000000000010110101001101;
assign LUT_1[47570] = 32'b00000000000000000101010001100010;
assign LUT_1[47571] = 32'b11111111111111111110100011011110;
assign LUT_1[47572] = 32'b00000000000000010001011100101000;
assign LUT_1[47573] = 32'b00000000000000001010101110100100;
assign LUT_1[47574] = 32'b00000000000000001101001010111001;
assign LUT_1[47575] = 32'b00000000000000000110011100110101;
assign LUT_1[47576] = 32'b00000000000000001000110001000110;
assign LUT_1[47577] = 32'b00000000000000000010000011000010;
assign LUT_1[47578] = 32'b00000000000000000100011111010111;
assign LUT_1[47579] = 32'b11111111111111111101110001010011;
assign LUT_1[47580] = 32'b00000000000000010000101010011101;
assign LUT_1[47581] = 32'b00000000000000001001111100011001;
assign LUT_1[47582] = 32'b00000000000000001100011000101110;
assign LUT_1[47583] = 32'b00000000000000000101101010101010;
assign LUT_1[47584] = 32'b00000000000000001000100010101110;
assign LUT_1[47585] = 32'b00000000000000000001110100101010;
assign LUT_1[47586] = 32'b00000000000000000100010000111111;
assign LUT_1[47587] = 32'b11111111111111111101100010111011;
assign LUT_1[47588] = 32'b00000000000000010000011100000101;
assign LUT_1[47589] = 32'b00000000000000001001101110000001;
assign LUT_1[47590] = 32'b00000000000000001100001010010110;
assign LUT_1[47591] = 32'b00000000000000000101011100010010;
assign LUT_1[47592] = 32'b00000000000000000111110000100011;
assign LUT_1[47593] = 32'b00000000000000000001000010011111;
assign LUT_1[47594] = 32'b00000000000000000011011110110100;
assign LUT_1[47595] = 32'b11111111111111111100110000110000;
assign LUT_1[47596] = 32'b00000000000000001111101001111010;
assign LUT_1[47597] = 32'b00000000000000001000111011110110;
assign LUT_1[47598] = 32'b00000000000000001011011000001011;
assign LUT_1[47599] = 32'b00000000000000000100101010000111;
assign LUT_1[47600] = 32'b00000000000000001010011110010000;
assign LUT_1[47601] = 32'b00000000000000000011110000001100;
assign LUT_1[47602] = 32'b00000000000000000110001100100001;
assign LUT_1[47603] = 32'b11111111111111111111011110011101;
assign LUT_1[47604] = 32'b00000000000000010010010111100111;
assign LUT_1[47605] = 32'b00000000000000001011101001100011;
assign LUT_1[47606] = 32'b00000000000000001110000101111000;
assign LUT_1[47607] = 32'b00000000000000000111010111110100;
assign LUT_1[47608] = 32'b00000000000000001001101100000101;
assign LUT_1[47609] = 32'b00000000000000000010111110000001;
assign LUT_1[47610] = 32'b00000000000000000101011010010110;
assign LUT_1[47611] = 32'b11111111111111111110101100010010;
assign LUT_1[47612] = 32'b00000000000000010001100101011100;
assign LUT_1[47613] = 32'b00000000000000001010110111011000;
assign LUT_1[47614] = 32'b00000000000000001101010011101101;
assign LUT_1[47615] = 32'b00000000000000000110100101101001;
assign LUT_1[47616] = 32'b11111111111111111110100100010101;
assign LUT_1[47617] = 32'b11111111111111110111110110010001;
assign LUT_1[47618] = 32'b11111111111111111010010010100110;
assign LUT_1[47619] = 32'b11111111111111110011100100100010;
assign LUT_1[47620] = 32'b00000000000000000110011101101100;
assign LUT_1[47621] = 32'b11111111111111111111101111101000;
assign LUT_1[47622] = 32'b00000000000000000010001011111101;
assign LUT_1[47623] = 32'b11111111111111111011011101111001;
assign LUT_1[47624] = 32'b11111111111111111101110010001010;
assign LUT_1[47625] = 32'b11111111111111110111000100000110;
assign LUT_1[47626] = 32'b11111111111111111001100000011011;
assign LUT_1[47627] = 32'b11111111111111110010110010010111;
assign LUT_1[47628] = 32'b00000000000000000101101011100001;
assign LUT_1[47629] = 32'b11111111111111111110111101011101;
assign LUT_1[47630] = 32'b00000000000000000001011001110010;
assign LUT_1[47631] = 32'b11111111111111111010101011101110;
assign LUT_1[47632] = 32'b00000000000000000000011111110111;
assign LUT_1[47633] = 32'b11111111111111111001110001110011;
assign LUT_1[47634] = 32'b11111111111111111100001110001000;
assign LUT_1[47635] = 32'b11111111111111110101100000000100;
assign LUT_1[47636] = 32'b00000000000000001000011001001110;
assign LUT_1[47637] = 32'b00000000000000000001101011001010;
assign LUT_1[47638] = 32'b00000000000000000100000111011111;
assign LUT_1[47639] = 32'b11111111111111111101011001011011;
assign LUT_1[47640] = 32'b11111111111111111111101101101100;
assign LUT_1[47641] = 32'b11111111111111111000111111101000;
assign LUT_1[47642] = 32'b11111111111111111011011011111101;
assign LUT_1[47643] = 32'b11111111111111110100101101111001;
assign LUT_1[47644] = 32'b00000000000000000111100111000011;
assign LUT_1[47645] = 32'b00000000000000000000111000111111;
assign LUT_1[47646] = 32'b00000000000000000011010101010100;
assign LUT_1[47647] = 32'b11111111111111111100100111010000;
assign LUT_1[47648] = 32'b11111111111111111111011111010100;
assign LUT_1[47649] = 32'b11111111111111111000110001010000;
assign LUT_1[47650] = 32'b11111111111111111011001101100101;
assign LUT_1[47651] = 32'b11111111111111110100011111100001;
assign LUT_1[47652] = 32'b00000000000000000111011000101011;
assign LUT_1[47653] = 32'b00000000000000000000101010100111;
assign LUT_1[47654] = 32'b00000000000000000011000110111100;
assign LUT_1[47655] = 32'b11111111111111111100011000111000;
assign LUT_1[47656] = 32'b11111111111111111110101101001001;
assign LUT_1[47657] = 32'b11111111111111110111111111000101;
assign LUT_1[47658] = 32'b11111111111111111010011011011010;
assign LUT_1[47659] = 32'b11111111111111110011101101010110;
assign LUT_1[47660] = 32'b00000000000000000110100110100000;
assign LUT_1[47661] = 32'b11111111111111111111111000011100;
assign LUT_1[47662] = 32'b00000000000000000010010100110001;
assign LUT_1[47663] = 32'b11111111111111111011100110101101;
assign LUT_1[47664] = 32'b00000000000000000001011010110110;
assign LUT_1[47665] = 32'b11111111111111111010101100110010;
assign LUT_1[47666] = 32'b11111111111111111101001001000111;
assign LUT_1[47667] = 32'b11111111111111110110011011000011;
assign LUT_1[47668] = 32'b00000000000000001001010100001101;
assign LUT_1[47669] = 32'b00000000000000000010100110001001;
assign LUT_1[47670] = 32'b00000000000000000101000010011110;
assign LUT_1[47671] = 32'b11111111111111111110010100011010;
assign LUT_1[47672] = 32'b00000000000000000000101000101011;
assign LUT_1[47673] = 32'b11111111111111111001111010100111;
assign LUT_1[47674] = 32'b11111111111111111100010110111100;
assign LUT_1[47675] = 32'b11111111111111110101101000111000;
assign LUT_1[47676] = 32'b00000000000000001000100010000010;
assign LUT_1[47677] = 32'b00000000000000000001110011111110;
assign LUT_1[47678] = 32'b00000000000000000100010000010011;
assign LUT_1[47679] = 32'b11111111111111111101100010001111;
assign LUT_1[47680] = 32'b00000000000000000000100001111101;
assign LUT_1[47681] = 32'b11111111111111111001110011111001;
assign LUT_1[47682] = 32'b11111111111111111100010000001110;
assign LUT_1[47683] = 32'b11111111111111110101100010001010;
assign LUT_1[47684] = 32'b00000000000000001000011011010100;
assign LUT_1[47685] = 32'b00000000000000000001101101010000;
assign LUT_1[47686] = 32'b00000000000000000100001001100101;
assign LUT_1[47687] = 32'b11111111111111111101011011100001;
assign LUT_1[47688] = 32'b11111111111111111111101111110010;
assign LUT_1[47689] = 32'b11111111111111111001000001101110;
assign LUT_1[47690] = 32'b11111111111111111011011110000011;
assign LUT_1[47691] = 32'b11111111111111110100101111111111;
assign LUT_1[47692] = 32'b00000000000000000111101001001001;
assign LUT_1[47693] = 32'b00000000000000000000111011000101;
assign LUT_1[47694] = 32'b00000000000000000011010111011010;
assign LUT_1[47695] = 32'b11111111111111111100101001010110;
assign LUT_1[47696] = 32'b00000000000000000010011101011111;
assign LUT_1[47697] = 32'b11111111111111111011101111011011;
assign LUT_1[47698] = 32'b11111111111111111110001011110000;
assign LUT_1[47699] = 32'b11111111111111110111011101101100;
assign LUT_1[47700] = 32'b00000000000000001010010110110110;
assign LUT_1[47701] = 32'b00000000000000000011101000110010;
assign LUT_1[47702] = 32'b00000000000000000110000101000111;
assign LUT_1[47703] = 32'b11111111111111111111010111000011;
assign LUT_1[47704] = 32'b00000000000000000001101011010100;
assign LUT_1[47705] = 32'b11111111111111111010111101010000;
assign LUT_1[47706] = 32'b11111111111111111101011001100101;
assign LUT_1[47707] = 32'b11111111111111110110101011100001;
assign LUT_1[47708] = 32'b00000000000000001001100100101011;
assign LUT_1[47709] = 32'b00000000000000000010110110100111;
assign LUT_1[47710] = 32'b00000000000000000101010010111100;
assign LUT_1[47711] = 32'b11111111111111111110100100111000;
assign LUT_1[47712] = 32'b00000000000000000001011100111100;
assign LUT_1[47713] = 32'b11111111111111111010101110111000;
assign LUT_1[47714] = 32'b11111111111111111101001011001101;
assign LUT_1[47715] = 32'b11111111111111110110011101001001;
assign LUT_1[47716] = 32'b00000000000000001001010110010011;
assign LUT_1[47717] = 32'b00000000000000000010101000001111;
assign LUT_1[47718] = 32'b00000000000000000101000100100100;
assign LUT_1[47719] = 32'b11111111111111111110010110100000;
assign LUT_1[47720] = 32'b00000000000000000000101010110001;
assign LUT_1[47721] = 32'b11111111111111111001111100101101;
assign LUT_1[47722] = 32'b11111111111111111100011001000010;
assign LUT_1[47723] = 32'b11111111111111110101101010111110;
assign LUT_1[47724] = 32'b00000000000000001000100100001000;
assign LUT_1[47725] = 32'b00000000000000000001110110000100;
assign LUT_1[47726] = 32'b00000000000000000100010010011001;
assign LUT_1[47727] = 32'b11111111111111111101100100010101;
assign LUT_1[47728] = 32'b00000000000000000011011000011110;
assign LUT_1[47729] = 32'b11111111111111111100101010011010;
assign LUT_1[47730] = 32'b11111111111111111111000110101111;
assign LUT_1[47731] = 32'b11111111111111111000011000101011;
assign LUT_1[47732] = 32'b00000000000000001011010001110101;
assign LUT_1[47733] = 32'b00000000000000000100100011110001;
assign LUT_1[47734] = 32'b00000000000000000111000000000110;
assign LUT_1[47735] = 32'b00000000000000000000010010000010;
assign LUT_1[47736] = 32'b00000000000000000010100110010011;
assign LUT_1[47737] = 32'b11111111111111111011111000001111;
assign LUT_1[47738] = 32'b11111111111111111110010100100100;
assign LUT_1[47739] = 32'b11111111111111110111100110100000;
assign LUT_1[47740] = 32'b00000000000000001010011111101010;
assign LUT_1[47741] = 32'b00000000000000000011110001100110;
assign LUT_1[47742] = 32'b00000000000000000110001101111011;
assign LUT_1[47743] = 32'b11111111111111111111011111110111;
assign LUT_1[47744] = 32'b00000000000000000001100100011000;
assign LUT_1[47745] = 32'b11111111111111111010110110010100;
assign LUT_1[47746] = 32'b11111111111111111101010010101001;
assign LUT_1[47747] = 32'b11111111111111110110100100100101;
assign LUT_1[47748] = 32'b00000000000000001001011101101111;
assign LUT_1[47749] = 32'b00000000000000000010101111101011;
assign LUT_1[47750] = 32'b00000000000000000101001100000000;
assign LUT_1[47751] = 32'b11111111111111111110011101111100;
assign LUT_1[47752] = 32'b00000000000000000000110010001101;
assign LUT_1[47753] = 32'b11111111111111111010000100001001;
assign LUT_1[47754] = 32'b11111111111111111100100000011110;
assign LUT_1[47755] = 32'b11111111111111110101110010011010;
assign LUT_1[47756] = 32'b00000000000000001000101011100100;
assign LUT_1[47757] = 32'b00000000000000000001111101100000;
assign LUT_1[47758] = 32'b00000000000000000100011001110101;
assign LUT_1[47759] = 32'b11111111111111111101101011110001;
assign LUT_1[47760] = 32'b00000000000000000011011111111010;
assign LUT_1[47761] = 32'b11111111111111111100110001110110;
assign LUT_1[47762] = 32'b11111111111111111111001110001011;
assign LUT_1[47763] = 32'b11111111111111111000100000000111;
assign LUT_1[47764] = 32'b00000000000000001011011001010001;
assign LUT_1[47765] = 32'b00000000000000000100101011001101;
assign LUT_1[47766] = 32'b00000000000000000111000111100010;
assign LUT_1[47767] = 32'b00000000000000000000011001011110;
assign LUT_1[47768] = 32'b00000000000000000010101101101111;
assign LUT_1[47769] = 32'b11111111111111111011111111101011;
assign LUT_1[47770] = 32'b11111111111111111110011100000000;
assign LUT_1[47771] = 32'b11111111111111110111101101111100;
assign LUT_1[47772] = 32'b00000000000000001010100111000110;
assign LUT_1[47773] = 32'b00000000000000000011111001000010;
assign LUT_1[47774] = 32'b00000000000000000110010101010111;
assign LUT_1[47775] = 32'b11111111111111111111100111010011;
assign LUT_1[47776] = 32'b00000000000000000010011111010111;
assign LUT_1[47777] = 32'b11111111111111111011110001010011;
assign LUT_1[47778] = 32'b11111111111111111110001101101000;
assign LUT_1[47779] = 32'b11111111111111110111011111100100;
assign LUT_1[47780] = 32'b00000000000000001010011000101110;
assign LUT_1[47781] = 32'b00000000000000000011101010101010;
assign LUT_1[47782] = 32'b00000000000000000110000110111111;
assign LUT_1[47783] = 32'b11111111111111111111011000111011;
assign LUT_1[47784] = 32'b00000000000000000001101101001100;
assign LUT_1[47785] = 32'b11111111111111111010111111001000;
assign LUT_1[47786] = 32'b11111111111111111101011011011101;
assign LUT_1[47787] = 32'b11111111111111110110101101011001;
assign LUT_1[47788] = 32'b00000000000000001001100110100011;
assign LUT_1[47789] = 32'b00000000000000000010111000011111;
assign LUT_1[47790] = 32'b00000000000000000101010100110100;
assign LUT_1[47791] = 32'b11111111111111111110100110110000;
assign LUT_1[47792] = 32'b00000000000000000100011010111001;
assign LUT_1[47793] = 32'b11111111111111111101101100110101;
assign LUT_1[47794] = 32'b00000000000000000000001001001010;
assign LUT_1[47795] = 32'b11111111111111111001011011000110;
assign LUT_1[47796] = 32'b00000000000000001100010100010000;
assign LUT_1[47797] = 32'b00000000000000000101100110001100;
assign LUT_1[47798] = 32'b00000000000000001000000010100001;
assign LUT_1[47799] = 32'b00000000000000000001010100011101;
assign LUT_1[47800] = 32'b00000000000000000011101000101110;
assign LUT_1[47801] = 32'b11111111111111111100111010101010;
assign LUT_1[47802] = 32'b11111111111111111111010110111111;
assign LUT_1[47803] = 32'b11111111111111111000101000111011;
assign LUT_1[47804] = 32'b00000000000000001011100010000101;
assign LUT_1[47805] = 32'b00000000000000000100110100000001;
assign LUT_1[47806] = 32'b00000000000000000111010000010110;
assign LUT_1[47807] = 32'b00000000000000000000100010010010;
assign LUT_1[47808] = 32'b00000000000000000011100010000000;
assign LUT_1[47809] = 32'b11111111111111111100110011111100;
assign LUT_1[47810] = 32'b11111111111111111111010000010001;
assign LUT_1[47811] = 32'b11111111111111111000100010001101;
assign LUT_1[47812] = 32'b00000000000000001011011011010111;
assign LUT_1[47813] = 32'b00000000000000000100101101010011;
assign LUT_1[47814] = 32'b00000000000000000111001001101000;
assign LUT_1[47815] = 32'b00000000000000000000011011100100;
assign LUT_1[47816] = 32'b00000000000000000010101111110101;
assign LUT_1[47817] = 32'b11111111111111111100000001110001;
assign LUT_1[47818] = 32'b11111111111111111110011110000110;
assign LUT_1[47819] = 32'b11111111111111110111110000000010;
assign LUT_1[47820] = 32'b00000000000000001010101001001100;
assign LUT_1[47821] = 32'b00000000000000000011111011001000;
assign LUT_1[47822] = 32'b00000000000000000110010111011101;
assign LUT_1[47823] = 32'b11111111111111111111101001011001;
assign LUT_1[47824] = 32'b00000000000000000101011101100010;
assign LUT_1[47825] = 32'b11111111111111111110101111011110;
assign LUT_1[47826] = 32'b00000000000000000001001011110011;
assign LUT_1[47827] = 32'b11111111111111111010011101101111;
assign LUT_1[47828] = 32'b00000000000000001101010110111001;
assign LUT_1[47829] = 32'b00000000000000000110101000110101;
assign LUT_1[47830] = 32'b00000000000000001001000101001010;
assign LUT_1[47831] = 32'b00000000000000000010010111000110;
assign LUT_1[47832] = 32'b00000000000000000100101011010111;
assign LUT_1[47833] = 32'b11111111111111111101111101010011;
assign LUT_1[47834] = 32'b00000000000000000000011001101000;
assign LUT_1[47835] = 32'b11111111111111111001101011100100;
assign LUT_1[47836] = 32'b00000000000000001100100100101110;
assign LUT_1[47837] = 32'b00000000000000000101110110101010;
assign LUT_1[47838] = 32'b00000000000000001000010010111111;
assign LUT_1[47839] = 32'b00000000000000000001100100111011;
assign LUT_1[47840] = 32'b00000000000000000100011100111111;
assign LUT_1[47841] = 32'b11111111111111111101101110111011;
assign LUT_1[47842] = 32'b00000000000000000000001011010000;
assign LUT_1[47843] = 32'b11111111111111111001011101001100;
assign LUT_1[47844] = 32'b00000000000000001100010110010110;
assign LUT_1[47845] = 32'b00000000000000000101101000010010;
assign LUT_1[47846] = 32'b00000000000000001000000100100111;
assign LUT_1[47847] = 32'b00000000000000000001010110100011;
assign LUT_1[47848] = 32'b00000000000000000011101010110100;
assign LUT_1[47849] = 32'b11111111111111111100111100110000;
assign LUT_1[47850] = 32'b11111111111111111111011001000101;
assign LUT_1[47851] = 32'b11111111111111111000101011000001;
assign LUT_1[47852] = 32'b00000000000000001011100100001011;
assign LUT_1[47853] = 32'b00000000000000000100110110000111;
assign LUT_1[47854] = 32'b00000000000000000111010010011100;
assign LUT_1[47855] = 32'b00000000000000000000100100011000;
assign LUT_1[47856] = 32'b00000000000000000110011000100001;
assign LUT_1[47857] = 32'b11111111111111111111101010011101;
assign LUT_1[47858] = 32'b00000000000000000010000110110010;
assign LUT_1[47859] = 32'b11111111111111111011011000101110;
assign LUT_1[47860] = 32'b00000000000000001110010001111000;
assign LUT_1[47861] = 32'b00000000000000000111100011110100;
assign LUT_1[47862] = 32'b00000000000000001010000000001001;
assign LUT_1[47863] = 32'b00000000000000000011010010000101;
assign LUT_1[47864] = 32'b00000000000000000101100110010110;
assign LUT_1[47865] = 32'b11111111111111111110111000010010;
assign LUT_1[47866] = 32'b00000000000000000001010100100111;
assign LUT_1[47867] = 32'b11111111111111111010100110100011;
assign LUT_1[47868] = 32'b00000000000000001101011111101101;
assign LUT_1[47869] = 32'b00000000000000000110110001101001;
assign LUT_1[47870] = 32'b00000000000000001001001101111110;
assign LUT_1[47871] = 32'b00000000000000000010011111111010;
assign LUT_1[47872] = 32'b11111111111111111100011000100001;
assign LUT_1[47873] = 32'b11111111111111110101101010011101;
assign LUT_1[47874] = 32'b11111111111111111000000110110010;
assign LUT_1[47875] = 32'b11111111111111110001011000101110;
assign LUT_1[47876] = 32'b00000000000000000100010001111000;
assign LUT_1[47877] = 32'b11111111111111111101100011110100;
assign LUT_1[47878] = 32'b00000000000000000000000000001001;
assign LUT_1[47879] = 32'b11111111111111111001010010000101;
assign LUT_1[47880] = 32'b11111111111111111011100110010110;
assign LUT_1[47881] = 32'b11111111111111110100111000010010;
assign LUT_1[47882] = 32'b11111111111111110111010100100111;
assign LUT_1[47883] = 32'b11111111111111110000100110100011;
assign LUT_1[47884] = 32'b00000000000000000011011111101101;
assign LUT_1[47885] = 32'b11111111111111111100110001101001;
assign LUT_1[47886] = 32'b11111111111111111111001101111110;
assign LUT_1[47887] = 32'b11111111111111111000011111111010;
assign LUT_1[47888] = 32'b11111111111111111110010100000011;
assign LUT_1[47889] = 32'b11111111111111110111100101111111;
assign LUT_1[47890] = 32'b11111111111111111010000010010100;
assign LUT_1[47891] = 32'b11111111111111110011010100010000;
assign LUT_1[47892] = 32'b00000000000000000110001101011010;
assign LUT_1[47893] = 32'b11111111111111111111011111010110;
assign LUT_1[47894] = 32'b00000000000000000001111011101011;
assign LUT_1[47895] = 32'b11111111111111111011001101100111;
assign LUT_1[47896] = 32'b11111111111111111101100001111000;
assign LUT_1[47897] = 32'b11111111111111110110110011110100;
assign LUT_1[47898] = 32'b11111111111111111001010000001001;
assign LUT_1[47899] = 32'b11111111111111110010100010000101;
assign LUT_1[47900] = 32'b00000000000000000101011011001111;
assign LUT_1[47901] = 32'b11111111111111111110101101001011;
assign LUT_1[47902] = 32'b00000000000000000001001001100000;
assign LUT_1[47903] = 32'b11111111111111111010011011011100;
assign LUT_1[47904] = 32'b11111111111111111101010011100000;
assign LUT_1[47905] = 32'b11111111111111110110100101011100;
assign LUT_1[47906] = 32'b11111111111111111001000001110001;
assign LUT_1[47907] = 32'b11111111111111110010010011101101;
assign LUT_1[47908] = 32'b00000000000000000101001100110111;
assign LUT_1[47909] = 32'b11111111111111111110011110110011;
assign LUT_1[47910] = 32'b00000000000000000000111011001000;
assign LUT_1[47911] = 32'b11111111111111111010001101000100;
assign LUT_1[47912] = 32'b11111111111111111100100001010101;
assign LUT_1[47913] = 32'b11111111111111110101110011010001;
assign LUT_1[47914] = 32'b11111111111111111000001111100110;
assign LUT_1[47915] = 32'b11111111111111110001100001100010;
assign LUT_1[47916] = 32'b00000000000000000100011010101100;
assign LUT_1[47917] = 32'b11111111111111111101101100101000;
assign LUT_1[47918] = 32'b00000000000000000000001000111101;
assign LUT_1[47919] = 32'b11111111111111111001011010111001;
assign LUT_1[47920] = 32'b11111111111111111111001111000010;
assign LUT_1[47921] = 32'b11111111111111111000100000111110;
assign LUT_1[47922] = 32'b11111111111111111010111101010011;
assign LUT_1[47923] = 32'b11111111111111110100001111001111;
assign LUT_1[47924] = 32'b00000000000000000111001000011001;
assign LUT_1[47925] = 32'b00000000000000000000011010010101;
assign LUT_1[47926] = 32'b00000000000000000010110110101010;
assign LUT_1[47927] = 32'b11111111111111111100001000100110;
assign LUT_1[47928] = 32'b11111111111111111110011100110111;
assign LUT_1[47929] = 32'b11111111111111110111101110110011;
assign LUT_1[47930] = 32'b11111111111111111010001011001000;
assign LUT_1[47931] = 32'b11111111111111110011011101000100;
assign LUT_1[47932] = 32'b00000000000000000110010110001110;
assign LUT_1[47933] = 32'b11111111111111111111101000001010;
assign LUT_1[47934] = 32'b00000000000000000010000100011111;
assign LUT_1[47935] = 32'b11111111111111111011010110011011;
assign LUT_1[47936] = 32'b11111111111111111110010110001001;
assign LUT_1[47937] = 32'b11111111111111110111101000000101;
assign LUT_1[47938] = 32'b11111111111111111010000100011010;
assign LUT_1[47939] = 32'b11111111111111110011010110010110;
assign LUT_1[47940] = 32'b00000000000000000110001111100000;
assign LUT_1[47941] = 32'b11111111111111111111100001011100;
assign LUT_1[47942] = 32'b00000000000000000001111101110001;
assign LUT_1[47943] = 32'b11111111111111111011001111101101;
assign LUT_1[47944] = 32'b11111111111111111101100011111110;
assign LUT_1[47945] = 32'b11111111111111110110110101111010;
assign LUT_1[47946] = 32'b11111111111111111001010010001111;
assign LUT_1[47947] = 32'b11111111111111110010100100001011;
assign LUT_1[47948] = 32'b00000000000000000101011101010101;
assign LUT_1[47949] = 32'b11111111111111111110101111010001;
assign LUT_1[47950] = 32'b00000000000000000001001011100110;
assign LUT_1[47951] = 32'b11111111111111111010011101100010;
assign LUT_1[47952] = 32'b00000000000000000000010001101011;
assign LUT_1[47953] = 32'b11111111111111111001100011100111;
assign LUT_1[47954] = 32'b11111111111111111011111111111100;
assign LUT_1[47955] = 32'b11111111111111110101010001111000;
assign LUT_1[47956] = 32'b00000000000000001000001011000010;
assign LUT_1[47957] = 32'b00000000000000000001011100111110;
assign LUT_1[47958] = 32'b00000000000000000011111001010011;
assign LUT_1[47959] = 32'b11111111111111111101001011001111;
assign LUT_1[47960] = 32'b11111111111111111111011111100000;
assign LUT_1[47961] = 32'b11111111111111111000110001011100;
assign LUT_1[47962] = 32'b11111111111111111011001101110001;
assign LUT_1[47963] = 32'b11111111111111110100011111101101;
assign LUT_1[47964] = 32'b00000000000000000111011000110111;
assign LUT_1[47965] = 32'b00000000000000000000101010110011;
assign LUT_1[47966] = 32'b00000000000000000011000111001000;
assign LUT_1[47967] = 32'b11111111111111111100011001000100;
assign LUT_1[47968] = 32'b11111111111111111111010001001000;
assign LUT_1[47969] = 32'b11111111111111111000100011000100;
assign LUT_1[47970] = 32'b11111111111111111010111111011001;
assign LUT_1[47971] = 32'b11111111111111110100010001010101;
assign LUT_1[47972] = 32'b00000000000000000111001010011111;
assign LUT_1[47973] = 32'b00000000000000000000011100011011;
assign LUT_1[47974] = 32'b00000000000000000010111000110000;
assign LUT_1[47975] = 32'b11111111111111111100001010101100;
assign LUT_1[47976] = 32'b11111111111111111110011110111101;
assign LUT_1[47977] = 32'b11111111111111110111110000111001;
assign LUT_1[47978] = 32'b11111111111111111010001101001110;
assign LUT_1[47979] = 32'b11111111111111110011011111001010;
assign LUT_1[47980] = 32'b00000000000000000110011000010100;
assign LUT_1[47981] = 32'b11111111111111111111101010010000;
assign LUT_1[47982] = 32'b00000000000000000010000110100101;
assign LUT_1[47983] = 32'b11111111111111111011011000100001;
assign LUT_1[47984] = 32'b00000000000000000001001100101010;
assign LUT_1[47985] = 32'b11111111111111111010011110100110;
assign LUT_1[47986] = 32'b11111111111111111100111010111011;
assign LUT_1[47987] = 32'b11111111111111110110001100110111;
assign LUT_1[47988] = 32'b00000000000000001001000110000001;
assign LUT_1[47989] = 32'b00000000000000000010010111111101;
assign LUT_1[47990] = 32'b00000000000000000100110100010010;
assign LUT_1[47991] = 32'b11111111111111111110000110001110;
assign LUT_1[47992] = 32'b00000000000000000000011010011111;
assign LUT_1[47993] = 32'b11111111111111111001101100011011;
assign LUT_1[47994] = 32'b11111111111111111100001000110000;
assign LUT_1[47995] = 32'b11111111111111110101011010101100;
assign LUT_1[47996] = 32'b00000000000000001000010011110110;
assign LUT_1[47997] = 32'b00000000000000000001100101110010;
assign LUT_1[47998] = 32'b00000000000000000100000010000111;
assign LUT_1[47999] = 32'b11111111111111111101010100000011;
assign LUT_1[48000] = 32'b11111111111111111111011000100100;
assign LUT_1[48001] = 32'b11111111111111111000101010100000;
assign LUT_1[48002] = 32'b11111111111111111011000110110101;
assign LUT_1[48003] = 32'b11111111111111110100011000110001;
assign LUT_1[48004] = 32'b00000000000000000111010001111011;
assign LUT_1[48005] = 32'b00000000000000000000100011110111;
assign LUT_1[48006] = 32'b00000000000000000011000000001100;
assign LUT_1[48007] = 32'b11111111111111111100010010001000;
assign LUT_1[48008] = 32'b11111111111111111110100110011001;
assign LUT_1[48009] = 32'b11111111111111110111111000010101;
assign LUT_1[48010] = 32'b11111111111111111010010100101010;
assign LUT_1[48011] = 32'b11111111111111110011100110100110;
assign LUT_1[48012] = 32'b00000000000000000110011111110000;
assign LUT_1[48013] = 32'b11111111111111111111110001101100;
assign LUT_1[48014] = 32'b00000000000000000010001110000001;
assign LUT_1[48015] = 32'b11111111111111111011011111111101;
assign LUT_1[48016] = 32'b00000000000000000001010100000110;
assign LUT_1[48017] = 32'b11111111111111111010100110000010;
assign LUT_1[48018] = 32'b11111111111111111101000010010111;
assign LUT_1[48019] = 32'b11111111111111110110010100010011;
assign LUT_1[48020] = 32'b00000000000000001001001101011101;
assign LUT_1[48021] = 32'b00000000000000000010011111011001;
assign LUT_1[48022] = 32'b00000000000000000100111011101110;
assign LUT_1[48023] = 32'b11111111111111111110001101101010;
assign LUT_1[48024] = 32'b00000000000000000000100001111011;
assign LUT_1[48025] = 32'b11111111111111111001110011110111;
assign LUT_1[48026] = 32'b11111111111111111100010000001100;
assign LUT_1[48027] = 32'b11111111111111110101100010001000;
assign LUT_1[48028] = 32'b00000000000000001000011011010010;
assign LUT_1[48029] = 32'b00000000000000000001101101001110;
assign LUT_1[48030] = 32'b00000000000000000100001001100011;
assign LUT_1[48031] = 32'b11111111111111111101011011011111;
assign LUT_1[48032] = 32'b00000000000000000000010011100011;
assign LUT_1[48033] = 32'b11111111111111111001100101011111;
assign LUT_1[48034] = 32'b11111111111111111100000001110100;
assign LUT_1[48035] = 32'b11111111111111110101010011110000;
assign LUT_1[48036] = 32'b00000000000000001000001100111010;
assign LUT_1[48037] = 32'b00000000000000000001011110110110;
assign LUT_1[48038] = 32'b00000000000000000011111011001011;
assign LUT_1[48039] = 32'b11111111111111111101001101000111;
assign LUT_1[48040] = 32'b11111111111111111111100001011000;
assign LUT_1[48041] = 32'b11111111111111111000110011010100;
assign LUT_1[48042] = 32'b11111111111111111011001111101001;
assign LUT_1[48043] = 32'b11111111111111110100100001100101;
assign LUT_1[48044] = 32'b00000000000000000111011010101111;
assign LUT_1[48045] = 32'b00000000000000000000101100101011;
assign LUT_1[48046] = 32'b00000000000000000011001001000000;
assign LUT_1[48047] = 32'b11111111111111111100011010111100;
assign LUT_1[48048] = 32'b00000000000000000010001111000101;
assign LUT_1[48049] = 32'b11111111111111111011100001000001;
assign LUT_1[48050] = 32'b11111111111111111101111101010110;
assign LUT_1[48051] = 32'b11111111111111110111001111010010;
assign LUT_1[48052] = 32'b00000000000000001010001000011100;
assign LUT_1[48053] = 32'b00000000000000000011011010011000;
assign LUT_1[48054] = 32'b00000000000000000101110110101101;
assign LUT_1[48055] = 32'b11111111111111111111001000101001;
assign LUT_1[48056] = 32'b00000000000000000001011100111010;
assign LUT_1[48057] = 32'b11111111111111111010101110110110;
assign LUT_1[48058] = 32'b11111111111111111101001011001011;
assign LUT_1[48059] = 32'b11111111111111110110011101000111;
assign LUT_1[48060] = 32'b00000000000000001001010110010001;
assign LUT_1[48061] = 32'b00000000000000000010101000001101;
assign LUT_1[48062] = 32'b00000000000000000101000100100010;
assign LUT_1[48063] = 32'b11111111111111111110010110011110;
assign LUT_1[48064] = 32'b00000000000000000001010110001100;
assign LUT_1[48065] = 32'b11111111111111111010101000001000;
assign LUT_1[48066] = 32'b11111111111111111101000100011101;
assign LUT_1[48067] = 32'b11111111111111110110010110011001;
assign LUT_1[48068] = 32'b00000000000000001001001111100011;
assign LUT_1[48069] = 32'b00000000000000000010100001011111;
assign LUT_1[48070] = 32'b00000000000000000100111101110100;
assign LUT_1[48071] = 32'b11111111111111111110001111110000;
assign LUT_1[48072] = 32'b00000000000000000000100100000001;
assign LUT_1[48073] = 32'b11111111111111111001110101111101;
assign LUT_1[48074] = 32'b11111111111111111100010010010010;
assign LUT_1[48075] = 32'b11111111111111110101100100001110;
assign LUT_1[48076] = 32'b00000000000000001000011101011000;
assign LUT_1[48077] = 32'b00000000000000000001101111010100;
assign LUT_1[48078] = 32'b00000000000000000100001011101001;
assign LUT_1[48079] = 32'b11111111111111111101011101100101;
assign LUT_1[48080] = 32'b00000000000000000011010001101110;
assign LUT_1[48081] = 32'b11111111111111111100100011101010;
assign LUT_1[48082] = 32'b11111111111111111110111111111111;
assign LUT_1[48083] = 32'b11111111111111111000010001111011;
assign LUT_1[48084] = 32'b00000000000000001011001011000101;
assign LUT_1[48085] = 32'b00000000000000000100011101000001;
assign LUT_1[48086] = 32'b00000000000000000110111001010110;
assign LUT_1[48087] = 32'b00000000000000000000001011010010;
assign LUT_1[48088] = 32'b00000000000000000010011111100011;
assign LUT_1[48089] = 32'b11111111111111111011110001011111;
assign LUT_1[48090] = 32'b11111111111111111110001101110100;
assign LUT_1[48091] = 32'b11111111111111110111011111110000;
assign LUT_1[48092] = 32'b00000000000000001010011000111010;
assign LUT_1[48093] = 32'b00000000000000000011101010110110;
assign LUT_1[48094] = 32'b00000000000000000110000111001011;
assign LUT_1[48095] = 32'b11111111111111111111011001000111;
assign LUT_1[48096] = 32'b00000000000000000010010001001011;
assign LUT_1[48097] = 32'b11111111111111111011100011000111;
assign LUT_1[48098] = 32'b11111111111111111101111111011100;
assign LUT_1[48099] = 32'b11111111111111110111010001011000;
assign LUT_1[48100] = 32'b00000000000000001010001010100010;
assign LUT_1[48101] = 32'b00000000000000000011011100011110;
assign LUT_1[48102] = 32'b00000000000000000101111000110011;
assign LUT_1[48103] = 32'b11111111111111111111001010101111;
assign LUT_1[48104] = 32'b00000000000000000001011111000000;
assign LUT_1[48105] = 32'b11111111111111111010110000111100;
assign LUT_1[48106] = 32'b11111111111111111101001101010001;
assign LUT_1[48107] = 32'b11111111111111110110011111001101;
assign LUT_1[48108] = 32'b00000000000000001001011000010111;
assign LUT_1[48109] = 32'b00000000000000000010101010010011;
assign LUT_1[48110] = 32'b00000000000000000101000110101000;
assign LUT_1[48111] = 32'b11111111111111111110011000100100;
assign LUT_1[48112] = 32'b00000000000000000100001100101101;
assign LUT_1[48113] = 32'b11111111111111111101011110101001;
assign LUT_1[48114] = 32'b11111111111111111111111010111110;
assign LUT_1[48115] = 32'b11111111111111111001001100111010;
assign LUT_1[48116] = 32'b00000000000000001100000110000100;
assign LUT_1[48117] = 32'b00000000000000000101011000000000;
assign LUT_1[48118] = 32'b00000000000000000111110100010101;
assign LUT_1[48119] = 32'b00000000000000000001000110010001;
assign LUT_1[48120] = 32'b00000000000000000011011010100010;
assign LUT_1[48121] = 32'b11111111111111111100101100011110;
assign LUT_1[48122] = 32'b11111111111111111111001000110011;
assign LUT_1[48123] = 32'b11111111111111111000011010101111;
assign LUT_1[48124] = 32'b00000000000000001011010011111001;
assign LUT_1[48125] = 32'b00000000000000000100100101110101;
assign LUT_1[48126] = 32'b00000000000000000111000010001010;
assign LUT_1[48127] = 32'b00000000000000000000010100000110;
assign LUT_1[48128] = 32'b00000000000000001011001100101000;
assign LUT_1[48129] = 32'b00000000000000000100011110100100;
assign LUT_1[48130] = 32'b00000000000000000110111010111001;
assign LUT_1[48131] = 32'b00000000000000000000001100110101;
assign LUT_1[48132] = 32'b00000000000000010011000101111111;
assign LUT_1[48133] = 32'b00000000000000001100010111111011;
assign LUT_1[48134] = 32'b00000000000000001110110100010000;
assign LUT_1[48135] = 32'b00000000000000001000000110001100;
assign LUT_1[48136] = 32'b00000000000000001010011010011101;
assign LUT_1[48137] = 32'b00000000000000000011101100011001;
assign LUT_1[48138] = 32'b00000000000000000110001000101110;
assign LUT_1[48139] = 32'b11111111111111111111011010101010;
assign LUT_1[48140] = 32'b00000000000000010010010011110100;
assign LUT_1[48141] = 32'b00000000000000001011100101110000;
assign LUT_1[48142] = 32'b00000000000000001110000010000101;
assign LUT_1[48143] = 32'b00000000000000000111010100000001;
assign LUT_1[48144] = 32'b00000000000000001101001000001010;
assign LUT_1[48145] = 32'b00000000000000000110011010000110;
assign LUT_1[48146] = 32'b00000000000000001000110110011011;
assign LUT_1[48147] = 32'b00000000000000000010001000010111;
assign LUT_1[48148] = 32'b00000000000000010101000001100001;
assign LUT_1[48149] = 32'b00000000000000001110010011011101;
assign LUT_1[48150] = 32'b00000000000000010000101111110010;
assign LUT_1[48151] = 32'b00000000000000001010000001101110;
assign LUT_1[48152] = 32'b00000000000000001100010101111111;
assign LUT_1[48153] = 32'b00000000000000000101100111111011;
assign LUT_1[48154] = 32'b00000000000000001000000100010000;
assign LUT_1[48155] = 32'b00000000000000000001010110001100;
assign LUT_1[48156] = 32'b00000000000000010100001111010110;
assign LUT_1[48157] = 32'b00000000000000001101100001010010;
assign LUT_1[48158] = 32'b00000000000000001111111101100111;
assign LUT_1[48159] = 32'b00000000000000001001001111100011;
assign LUT_1[48160] = 32'b00000000000000001100000111100111;
assign LUT_1[48161] = 32'b00000000000000000101011001100011;
assign LUT_1[48162] = 32'b00000000000000000111110101111000;
assign LUT_1[48163] = 32'b00000000000000000001000111110100;
assign LUT_1[48164] = 32'b00000000000000010100000000111110;
assign LUT_1[48165] = 32'b00000000000000001101010010111010;
assign LUT_1[48166] = 32'b00000000000000001111101111001111;
assign LUT_1[48167] = 32'b00000000000000001001000001001011;
assign LUT_1[48168] = 32'b00000000000000001011010101011100;
assign LUT_1[48169] = 32'b00000000000000000100100111011000;
assign LUT_1[48170] = 32'b00000000000000000111000011101101;
assign LUT_1[48171] = 32'b00000000000000000000010101101001;
assign LUT_1[48172] = 32'b00000000000000010011001110110011;
assign LUT_1[48173] = 32'b00000000000000001100100000101111;
assign LUT_1[48174] = 32'b00000000000000001110111101000100;
assign LUT_1[48175] = 32'b00000000000000001000001111000000;
assign LUT_1[48176] = 32'b00000000000000001110000011001001;
assign LUT_1[48177] = 32'b00000000000000000111010101000101;
assign LUT_1[48178] = 32'b00000000000000001001110001011010;
assign LUT_1[48179] = 32'b00000000000000000011000011010110;
assign LUT_1[48180] = 32'b00000000000000010101111100100000;
assign LUT_1[48181] = 32'b00000000000000001111001110011100;
assign LUT_1[48182] = 32'b00000000000000010001101010110001;
assign LUT_1[48183] = 32'b00000000000000001010111100101101;
assign LUT_1[48184] = 32'b00000000000000001101010000111110;
assign LUT_1[48185] = 32'b00000000000000000110100010111010;
assign LUT_1[48186] = 32'b00000000000000001000111111001111;
assign LUT_1[48187] = 32'b00000000000000000010010001001011;
assign LUT_1[48188] = 32'b00000000000000010101001010010101;
assign LUT_1[48189] = 32'b00000000000000001110011100010001;
assign LUT_1[48190] = 32'b00000000000000010000111000100110;
assign LUT_1[48191] = 32'b00000000000000001010001010100010;
assign LUT_1[48192] = 32'b00000000000000001101001010010000;
assign LUT_1[48193] = 32'b00000000000000000110011100001100;
assign LUT_1[48194] = 32'b00000000000000001000111000100001;
assign LUT_1[48195] = 32'b00000000000000000010001010011101;
assign LUT_1[48196] = 32'b00000000000000010101000011100111;
assign LUT_1[48197] = 32'b00000000000000001110010101100011;
assign LUT_1[48198] = 32'b00000000000000010000110001111000;
assign LUT_1[48199] = 32'b00000000000000001010000011110100;
assign LUT_1[48200] = 32'b00000000000000001100011000000101;
assign LUT_1[48201] = 32'b00000000000000000101101010000001;
assign LUT_1[48202] = 32'b00000000000000001000000110010110;
assign LUT_1[48203] = 32'b00000000000000000001011000010010;
assign LUT_1[48204] = 32'b00000000000000010100010001011100;
assign LUT_1[48205] = 32'b00000000000000001101100011011000;
assign LUT_1[48206] = 32'b00000000000000001111111111101101;
assign LUT_1[48207] = 32'b00000000000000001001010001101001;
assign LUT_1[48208] = 32'b00000000000000001111000101110010;
assign LUT_1[48209] = 32'b00000000000000001000010111101110;
assign LUT_1[48210] = 32'b00000000000000001010110100000011;
assign LUT_1[48211] = 32'b00000000000000000100000101111111;
assign LUT_1[48212] = 32'b00000000000000010110111111001001;
assign LUT_1[48213] = 32'b00000000000000010000010001000101;
assign LUT_1[48214] = 32'b00000000000000010010101101011010;
assign LUT_1[48215] = 32'b00000000000000001011111111010110;
assign LUT_1[48216] = 32'b00000000000000001110010011100111;
assign LUT_1[48217] = 32'b00000000000000000111100101100011;
assign LUT_1[48218] = 32'b00000000000000001010000001111000;
assign LUT_1[48219] = 32'b00000000000000000011010011110100;
assign LUT_1[48220] = 32'b00000000000000010110001100111110;
assign LUT_1[48221] = 32'b00000000000000001111011110111010;
assign LUT_1[48222] = 32'b00000000000000010001111011001111;
assign LUT_1[48223] = 32'b00000000000000001011001101001011;
assign LUT_1[48224] = 32'b00000000000000001110000101001111;
assign LUT_1[48225] = 32'b00000000000000000111010111001011;
assign LUT_1[48226] = 32'b00000000000000001001110011100000;
assign LUT_1[48227] = 32'b00000000000000000011000101011100;
assign LUT_1[48228] = 32'b00000000000000010101111110100110;
assign LUT_1[48229] = 32'b00000000000000001111010000100010;
assign LUT_1[48230] = 32'b00000000000000010001101100110111;
assign LUT_1[48231] = 32'b00000000000000001010111110110011;
assign LUT_1[48232] = 32'b00000000000000001101010011000100;
assign LUT_1[48233] = 32'b00000000000000000110100101000000;
assign LUT_1[48234] = 32'b00000000000000001001000001010101;
assign LUT_1[48235] = 32'b00000000000000000010010011010001;
assign LUT_1[48236] = 32'b00000000000000010101001100011011;
assign LUT_1[48237] = 32'b00000000000000001110011110010111;
assign LUT_1[48238] = 32'b00000000000000010000111010101100;
assign LUT_1[48239] = 32'b00000000000000001010001100101000;
assign LUT_1[48240] = 32'b00000000000000010000000000110001;
assign LUT_1[48241] = 32'b00000000000000001001010010101101;
assign LUT_1[48242] = 32'b00000000000000001011101111000010;
assign LUT_1[48243] = 32'b00000000000000000101000000111110;
assign LUT_1[48244] = 32'b00000000000000010111111010001000;
assign LUT_1[48245] = 32'b00000000000000010001001100000100;
assign LUT_1[48246] = 32'b00000000000000010011101000011001;
assign LUT_1[48247] = 32'b00000000000000001100111010010101;
assign LUT_1[48248] = 32'b00000000000000001111001110100110;
assign LUT_1[48249] = 32'b00000000000000001000100000100010;
assign LUT_1[48250] = 32'b00000000000000001010111100110111;
assign LUT_1[48251] = 32'b00000000000000000100001110110011;
assign LUT_1[48252] = 32'b00000000000000010111000111111101;
assign LUT_1[48253] = 32'b00000000000000010000011001111001;
assign LUT_1[48254] = 32'b00000000000000010010110110001110;
assign LUT_1[48255] = 32'b00000000000000001100001000001010;
assign LUT_1[48256] = 32'b00000000000000001110001100101011;
assign LUT_1[48257] = 32'b00000000000000000111011110100111;
assign LUT_1[48258] = 32'b00000000000000001001111010111100;
assign LUT_1[48259] = 32'b00000000000000000011001100111000;
assign LUT_1[48260] = 32'b00000000000000010110000110000010;
assign LUT_1[48261] = 32'b00000000000000001111010111111110;
assign LUT_1[48262] = 32'b00000000000000010001110100010011;
assign LUT_1[48263] = 32'b00000000000000001011000110001111;
assign LUT_1[48264] = 32'b00000000000000001101011010100000;
assign LUT_1[48265] = 32'b00000000000000000110101100011100;
assign LUT_1[48266] = 32'b00000000000000001001001000110001;
assign LUT_1[48267] = 32'b00000000000000000010011010101101;
assign LUT_1[48268] = 32'b00000000000000010101010011110111;
assign LUT_1[48269] = 32'b00000000000000001110100101110011;
assign LUT_1[48270] = 32'b00000000000000010001000010001000;
assign LUT_1[48271] = 32'b00000000000000001010010100000100;
assign LUT_1[48272] = 32'b00000000000000010000001000001101;
assign LUT_1[48273] = 32'b00000000000000001001011010001001;
assign LUT_1[48274] = 32'b00000000000000001011110110011110;
assign LUT_1[48275] = 32'b00000000000000000101001000011010;
assign LUT_1[48276] = 32'b00000000000000011000000001100100;
assign LUT_1[48277] = 32'b00000000000000010001010011100000;
assign LUT_1[48278] = 32'b00000000000000010011101111110101;
assign LUT_1[48279] = 32'b00000000000000001101000001110001;
assign LUT_1[48280] = 32'b00000000000000001111010110000010;
assign LUT_1[48281] = 32'b00000000000000001000100111111110;
assign LUT_1[48282] = 32'b00000000000000001011000100010011;
assign LUT_1[48283] = 32'b00000000000000000100010110001111;
assign LUT_1[48284] = 32'b00000000000000010111001111011001;
assign LUT_1[48285] = 32'b00000000000000010000100001010101;
assign LUT_1[48286] = 32'b00000000000000010010111101101010;
assign LUT_1[48287] = 32'b00000000000000001100001111100110;
assign LUT_1[48288] = 32'b00000000000000001111000111101010;
assign LUT_1[48289] = 32'b00000000000000001000011001100110;
assign LUT_1[48290] = 32'b00000000000000001010110101111011;
assign LUT_1[48291] = 32'b00000000000000000100000111110111;
assign LUT_1[48292] = 32'b00000000000000010111000001000001;
assign LUT_1[48293] = 32'b00000000000000010000010010111101;
assign LUT_1[48294] = 32'b00000000000000010010101111010010;
assign LUT_1[48295] = 32'b00000000000000001100000001001110;
assign LUT_1[48296] = 32'b00000000000000001110010101011111;
assign LUT_1[48297] = 32'b00000000000000000111100111011011;
assign LUT_1[48298] = 32'b00000000000000001010000011110000;
assign LUT_1[48299] = 32'b00000000000000000011010101101100;
assign LUT_1[48300] = 32'b00000000000000010110001110110110;
assign LUT_1[48301] = 32'b00000000000000001111100000110010;
assign LUT_1[48302] = 32'b00000000000000010001111101000111;
assign LUT_1[48303] = 32'b00000000000000001011001111000011;
assign LUT_1[48304] = 32'b00000000000000010001000011001100;
assign LUT_1[48305] = 32'b00000000000000001010010101001000;
assign LUT_1[48306] = 32'b00000000000000001100110001011101;
assign LUT_1[48307] = 32'b00000000000000000110000011011001;
assign LUT_1[48308] = 32'b00000000000000011000111100100011;
assign LUT_1[48309] = 32'b00000000000000010010001110011111;
assign LUT_1[48310] = 32'b00000000000000010100101010110100;
assign LUT_1[48311] = 32'b00000000000000001101111100110000;
assign LUT_1[48312] = 32'b00000000000000010000010001000001;
assign LUT_1[48313] = 32'b00000000000000001001100010111101;
assign LUT_1[48314] = 32'b00000000000000001011111111010010;
assign LUT_1[48315] = 32'b00000000000000000101010001001110;
assign LUT_1[48316] = 32'b00000000000000011000001010011000;
assign LUT_1[48317] = 32'b00000000000000010001011100010100;
assign LUT_1[48318] = 32'b00000000000000010011111000101001;
assign LUT_1[48319] = 32'b00000000000000001101001010100101;
assign LUT_1[48320] = 32'b00000000000000010000001010010011;
assign LUT_1[48321] = 32'b00000000000000001001011100001111;
assign LUT_1[48322] = 32'b00000000000000001011111000100100;
assign LUT_1[48323] = 32'b00000000000000000101001010100000;
assign LUT_1[48324] = 32'b00000000000000011000000011101010;
assign LUT_1[48325] = 32'b00000000000000010001010101100110;
assign LUT_1[48326] = 32'b00000000000000010011110001111011;
assign LUT_1[48327] = 32'b00000000000000001101000011110111;
assign LUT_1[48328] = 32'b00000000000000001111011000001000;
assign LUT_1[48329] = 32'b00000000000000001000101010000100;
assign LUT_1[48330] = 32'b00000000000000001011000110011001;
assign LUT_1[48331] = 32'b00000000000000000100011000010101;
assign LUT_1[48332] = 32'b00000000000000010111010001011111;
assign LUT_1[48333] = 32'b00000000000000010000100011011011;
assign LUT_1[48334] = 32'b00000000000000010010111111110000;
assign LUT_1[48335] = 32'b00000000000000001100010001101100;
assign LUT_1[48336] = 32'b00000000000000010010000101110101;
assign LUT_1[48337] = 32'b00000000000000001011010111110001;
assign LUT_1[48338] = 32'b00000000000000001101110100000110;
assign LUT_1[48339] = 32'b00000000000000000111000110000010;
assign LUT_1[48340] = 32'b00000000000000011001111111001100;
assign LUT_1[48341] = 32'b00000000000000010011010001001000;
assign LUT_1[48342] = 32'b00000000000000010101101101011101;
assign LUT_1[48343] = 32'b00000000000000001110111111011001;
assign LUT_1[48344] = 32'b00000000000000010001010011101010;
assign LUT_1[48345] = 32'b00000000000000001010100101100110;
assign LUT_1[48346] = 32'b00000000000000001101000001111011;
assign LUT_1[48347] = 32'b00000000000000000110010011110111;
assign LUT_1[48348] = 32'b00000000000000011001001101000001;
assign LUT_1[48349] = 32'b00000000000000010010011110111101;
assign LUT_1[48350] = 32'b00000000000000010100111011010010;
assign LUT_1[48351] = 32'b00000000000000001110001101001110;
assign LUT_1[48352] = 32'b00000000000000010001000101010010;
assign LUT_1[48353] = 32'b00000000000000001010010111001110;
assign LUT_1[48354] = 32'b00000000000000001100110011100011;
assign LUT_1[48355] = 32'b00000000000000000110000101011111;
assign LUT_1[48356] = 32'b00000000000000011000111110101001;
assign LUT_1[48357] = 32'b00000000000000010010010000100101;
assign LUT_1[48358] = 32'b00000000000000010100101100111010;
assign LUT_1[48359] = 32'b00000000000000001101111110110110;
assign LUT_1[48360] = 32'b00000000000000010000010011000111;
assign LUT_1[48361] = 32'b00000000000000001001100101000011;
assign LUT_1[48362] = 32'b00000000000000001100000001011000;
assign LUT_1[48363] = 32'b00000000000000000101010011010100;
assign LUT_1[48364] = 32'b00000000000000011000001100011110;
assign LUT_1[48365] = 32'b00000000000000010001011110011010;
assign LUT_1[48366] = 32'b00000000000000010011111010101111;
assign LUT_1[48367] = 32'b00000000000000001101001100101011;
assign LUT_1[48368] = 32'b00000000000000010011000000110100;
assign LUT_1[48369] = 32'b00000000000000001100010010110000;
assign LUT_1[48370] = 32'b00000000000000001110101111000101;
assign LUT_1[48371] = 32'b00000000000000001000000001000001;
assign LUT_1[48372] = 32'b00000000000000011010111010001011;
assign LUT_1[48373] = 32'b00000000000000010100001100000111;
assign LUT_1[48374] = 32'b00000000000000010110101000011100;
assign LUT_1[48375] = 32'b00000000000000001111111010011000;
assign LUT_1[48376] = 32'b00000000000000010010001110101001;
assign LUT_1[48377] = 32'b00000000000000001011100000100101;
assign LUT_1[48378] = 32'b00000000000000001101111100111010;
assign LUT_1[48379] = 32'b00000000000000000111001110110110;
assign LUT_1[48380] = 32'b00000000000000011010001000000000;
assign LUT_1[48381] = 32'b00000000000000010011011001111100;
assign LUT_1[48382] = 32'b00000000000000010101110110010001;
assign LUT_1[48383] = 32'b00000000000000001111001000001101;
assign LUT_1[48384] = 32'b00000000000000001001000000110100;
assign LUT_1[48385] = 32'b00000000000000000010010010110000;
assign LUT_1[48386] = 32'b00000000000000000100101111000101;
assign LUT_1[48387] = 32'b11111111111111111110000001000001;
assign LUT_1[48388] = 32'b00000000000000010000111010001011;
assign LUT_1[48389] = 32'b00000000000000001010001100000111;
assign LUT_1[48390] = 32'b00000000000000001100101000011100;
assign LUT_1[48391] = 32'b00000000000000000101111010011000;
assign LUT_1[48392] = 32'b00000000000000001000001110101001;
assign LUT_1[48393] = 32'b00000000000000000001100000100101;
assign LUT_1[48394] = 32'b00000000000000000011111100111010;
assign LUT_1[48395] = 32'b11111111111111111101001110110110;
assign LUT_1[48396] = 32'b00000000000000010000001000000000;
assign LUT_1[48397] = 32'b00000000000000001001011001111100;
assign LUT_1[48398] = 32'b00000000000000001011110110010001;
assign LUT_1[48399] = 32'b00000000000000000101001000001101;
assign LUT_1[48400] = 32'b00000000000000001010111100010110;
assign LUT_1[48401] = 32'b00000000000000000100001110010010;
assign LUT_1[48402] = 32'b00000000000000000110101010100111;
assign LUT_1[48403] = 32'b11111111111111111111111100100011;
assign LUT_1[48404] = 32'b00000000000000010010110101101101;
assign LUT_1[48405] = 32'b00000000000000001100000111101001;
assign LUT_1[48406] = 32'b00000000000000001110100011111110;
assign LUT_1[48407] = 32'b00000000000000000111110101111010;
assign LUT_1[48408] = 32'b00000000000000001010001010001011;
assign LUT_1[48409] = 32'b00000000000000000011011100000111;
assign LUT_1[48410] = 32'b00000000000000000101111000011100;
assign LUT_1[48411] = 32'b11111111111111111111001010011000;
assign LUT_1[48412] = 32'b00000000000000010010000011100010;
assign LUT_1[48413] = 32'b00000000000000001011010101011110;
assign LUT_1[48414] = 32'b00000000000000001101110001110011;
assign LUT_1[48415] = 32'b00000000000000000111000011101111;
assign LUT_1[48416] = 32'b00000000000000001001111011110011;
assign LUT_1[48417] = 32'b00000000000000000011001101101111;
assign LUT_1[48418] = 32'b00000000000000000101101010000100;
assign LUT_1[48419] = 32'b11111111111111111110111100000000;
assign LUT_1[48420] = 32'b00000000000000010001110101001010;
assign LUT_1[48421] = 32'b00000000000000001011000111000110;
assign LUT_1[48422] = 32'b00000000000000001101100011011011;
assign LUT_1[48423] = 32'b00000000000000000110110101010111;
assign LUT_1[48424] = 32'b00000000000000001001001001101000;
assign LUT_1[48425] = 32'b00000000000000000010011011100100;
assign LUT_1[48426] = 32'b00000000000000000100110111111001;
assign LUT_1[48427] = 32'b11111111111111111110001001110101;
assign LUT_1[48428] = 32'b00000000000000010001000010111111;
assign LUT_1[48429] = 32'b00000000000000001010010100111011;
assign LUT_1[48430] = 32'b00000000000000001100110001010000;
assign LUT_1[48431] = 32'b00000000000000000110000011001100;
assign LUT_1[48432] = 32'b00000000000000001011110111010101;
assign LUT_1[48433] = 32'b00000000000000000101001001010001;
assign LUT_1[48434] = 32'b00000000000000000111100101100110;
assign LUT_1[48435] = 32'b00000000000000000000110111100010;
assign LUT_1[48436] = 32'b00000000000000010011110000101100;
assign LUT_1[48437] = 32'b00000000000000001101000010101000;
assign LUT_1[48438] = 32'b00000000000000001111011110111101;
assign LUT_1[48439] = 32'b00000000000000001000110000111001;
assign LUT_1[48440] = 32'b00000000000000001011000101001010;
assign LUT_1[48441] = 32'b00000000000000000100010111000110;
assign LUT_1[48442] = 32'b00000000000000000110110011011011;
assign LUT_1[48443] = 32'b00000000000000000000000101010111;
assign LUT_1[48444] = 32'b00000000000000010010111110100001;
assign LUT_1[48445] = 32'b00000000000000001100010000011101;
assign LUT_1[48446] = 32'b00000000000000001110101100110010;
assign LUT_1[48447] = 32'b00000000000000000111111110101110;
assign LUT_1[48448] = 32'b00000000000000001010111110011100;
assign LUT_1[48449] = 32'b00000000000000000100010000011000;
assign LUT_1[48450] = 32'b00000000000000000110101100101101;
assign LUT_1[48451] = 32'b11111111111111111111111110101001;
assign LUT_1[48452] = 32'b00000000000000010010110111110011;
assign LUT_1[48453] = 32'b00000000000000001100001001101111;
assign LUT_1[48454] = 32'b00000000000000001110100110000100;
assign LUT_1[48455] = 32'b00000000000000000111111000000000;
assign LUT_1[48456] = 32'b00000000000000001010001100010001;
assign LUT_1[48457] = 32'b00000000000000000011011110001101;
assign LUT_1[48458] = 32'b00000000000000000101111010100010;
assign LUT_1[48459] = 32'b11111111111111111111001100011110;
assign LUT_1[48460] = 32'b00000000000000010010000101101000;
assign LUT_1[48461] = 32'b00000000000000001011010111100100;
assign LUT_1[48462] = 32'b00000000000000001101110011111001;
assign LUT_1[48463] = 32'b00000000000000000111000101110101;
assign LUT_1[48464] = 32'b00000000000000001100111001111110;
assign LUT_1[48465] = 32'b00000000000000000110001011111010;
assign LUT_1[48466] = 32'b00000000000000001000101000001111;
assign LUT_1[48467] = 32'b00000000000000000001111010001011;
assign LUT_1[48468] = 32'b00000000000000010100110011010101;
assign LUT_1[48469] = 32'b00000000000000001110000101010001;
assign LUT_1[48470] = 32'b00000000000000010000100001100110;
assign LUT_1[48471] = 32'b00000000000000001001110011100010;
assign LUT_1[48472] = 32'b00000000000000001100000111110011;
assign LUT_1[48473] = 32'b00000000000000000101011001101111;
assign LUT_1[48474] = 32'b00000000000000000111110110000100;
assign LUT_1[48475] = 32'b00000000000000000001001000000000;
assign LUT_1[48476] = 32'b00000000000000010100000001001010;
assign LUT_1[48477] = 32'b00000000000000001101010011000110;
assign LUT_1[48478] = 32'b00000000000000001111101111011011;
assign LUT_1[48479] = 32'b00000000000000001001000001010111;
assign LUT_1[48480] = 32'b00000000000000001011111001011011;
assign LUT_1[48481] = 32'b00000000000000000101001011010111;
assign LUT_1[48482] = 32'b00000000000000000111100111101100;
assign LUT_1[48483] = 32'b00000000000000000000111001101000;
assign LUT_1[48484] = 32'b00000000000000010011110010110010;
assign LUT_1[48485] = 32'b00000000000000001101000100101110;
assign LUT_1[48486] = 32'b00000000000000001111100001000011;
assign LUT_1[48487] = 32'b00000000000000001000110010111111;
assign LUT_1[48488] = 32'b00000000000000001011000111010000;
assign LUT_1[48489] = 32'b00000000000000000100011001001100;
assign LUT_1[48490] = 32'b00000000000000000110110101100001;
assign LUT_1[48491] = 32'b00000000000000000000000111011101;
assign LUT_1[48492] = 32'b00000000000000010011000000100111;
assign LUT_1[48493] = 32'b00000000000000001100010010100011;
assign LUT_1[48494] = 32'b00000000000000001110101110111000;
assign LUT_1[48495] = 32'b00000000000000001000000000110100;
assign LUT_1[48496] = 32'b00000000000000001101110100111101;
assign LUT_1[48497] = 32'b00000000000000000111000110111001;
assign LUT_1[48498] = 32'b00000000000000001001100011001110;
assign LUT_1[48499] = 32'b00000000000000000010110101001010;
assign LUT_1[48500] = 32'b00000000000000010101101110010100;
assign LUT_1[48501] = 32'b00000000000000001111000000010000;
assign LUT_1[48502] = 32'b00000000000000010001011100100101;
assign LUT_1[48503] = 32'b00000000000000001010101110100001;
assign LUT_1[48504] = 32'b00000000000000001101000010110010;
assign LUT_1[48505] = 32'b00000000000000000110010100101110;
assign LUT_1[48506] = 32'b00000000000000001000110001000011;
assign LUT_1[48507] = 32'b00000000000000000010000010111111;
assign LUT_1[48508] = 32'b00000000000000010100111100001001;
assign LUT_1[48509] = 32'b00000000000000001110001110000101;
assign LUT_1[48510] = 32'b00000000000000010000101010011010;
assign LUT_1[48511] = 32'b00000000000000001001111100010110;
assign LUT_1[48512] = 32'b00000000000000001100000000110111;
assign LUT_1[48513] = 32'b00000000000000000101010010110011;
assign LUT_1[48514] = 32'b00000000000000000111101111001000;
assign LUT_1[48515] = 32'b00000000000000000001000001000100;
assign LUT_1[48516] = 32'b00000000000000010011111010001110;
assign LUT_1[48517] = 32'b00000000000000001101001100001010;
assign LUT_1[48518] = 32'b00000000000000001111101000011111;
assign LUT_1[48519] = 32'b00000000000000001000111010011011;
assign LUT_1[48520] = 32'b00000000000000001011001110101100;
assign LUT_1[48521] = 32'b00000000000000000100100000101000;
assign LUT_1[48522] = 32'b00000000000000000110111100111101;
assign LUT_1[48523] = 32'b00000000000000000000001110111001;
assign LUT_1[48524] = 32'b00000000000000010011001000000011;
assign LUT_1[48525] = 32'b00000000000000001100011001111111;
assign LUT_1[48526] = 32'b00000000000000001110110110010100;
assign LUT_1[48527] = 32'b00000000000000001000001000010000;
assign LUT_1[48528] = 32'b00000000000000001101111100011001;
assign LUT_1[48529] = 32'b00000000000000000111001110010101;
assign LUT_1[48530] = 32'b00000000000000001001101010101010;
assign LUT_1[48531] = 32'b00000000000000000010111100100110;
assign LUT_1[48532] = 32'b00000000000000010101110101110000;
assign LUT_1[48533] = 32'b00000000000000001111000111101100;
assign LUT_1[48534] = 32'b00000000000000010001100100000001;
assign LUT_1[48535] = 32'b00000000000000001010110101111101;
assign LUT_1[48536] = 32'b00000000000000001101001010001110;
assign LUT_1[48537] = 32'b00000000000000000110011100001010;
assign LUT_1[48538] = 32'b00000000000000001000111000011111;
assign LUT_1[48539] = 32'b00000000000000000010001010011011;
assign LUT_1[48540] = 32'b00000000000000010101000011100101;
assign LUT_1[48541] = 32'b00000000000000001110010101100001;
assign LUT_1[48542] = 32'b00000000000000010000110001110110;
assign LUT_1[48543] = 32'b00000000000000001010000011110010;
assign LUT_1[48544] = 32'b00000000000000001100111011110110;
assign LUT_1[48545] = 32'b00000000000000000110001101110010;
assign LUT_1[48546] = 32'b00000000000000001000101010000111;
assign LUT_1[48547] = 32'b00000000000000000001111100000011;
assign LUT_1[48548] = 32'b00000000000000010100110101001101;
assign LUT_1[48549] = 32'b00000000000000001110000111001001;
assign LUT_1[48550] = 32'b00000000000000010000100011011110;
assign LUT_1[48551] = 32'b00000000000000001001110101011010;
assign LUT_1[48552] = 32'b00000000000000001100001001101011;
assign LUT_1[48553] = 32'b00000000000000000101011011100111;
assign LUT_1[48554] = 32'b00000000000000000111110111111100;
assign LUT_1[48555] = 32'b00000000000000000001001001111000;
assign LUT_1[48556] = 32'b00000000000000010100000011000010;
assign LUT_1[48557] = 32'b00000000000000001101010100111110;
assign LUT_1[48558] = 32'b00000000000000001111110001010011;
assign LUT_1[48559] = 32'b00000000000000001001000011001111;
assign LUT_1[48560] = 32'b00000000000000001110110111011000;
assign LUT_1[48561] = 32'b00000000000000001000001001010100;
assign LUT_1[48562] = 32'b00000000000000001010100101101001;
assign LUT_1[48563] = 32'b00000000000000000011110111100101;
assign LUT_1[48564] = 32'b00000000000000010110110000101111;
assign LUT_1[48565] = 32'b00000000000000010000000010101011;
assign LUT_1[48566] = 32'b00000000000000010010011111000000;
assign LUT_1[48567] = 32'b00000000000000001011110000111100;
assign LUT_1[48568] = 32'b00000000000000001110000101001101;
assign LUT_1[48569] = 32'b00000000000000000111010111001001;
assign LUT_1[48570] = 32'b00000000000000001001110011011110;
assign LUT_1[48571] = 32'b00000000000000000011000101011010;
assign LUT_1[48572] = 32'b00000000000000010101111110100100;
assign LUT_1[48573] = 32'b00000000000000001111010000100000;
assign LUT_1[48574] = 32'b00000000000000010001101100110101;
assign LUT_1[48575] = 32'b00000000000000001010111110110001;
assign LUT_1[48576] = 32'b00000000000000001101111110011111;
assign LUT_1[48577] = 32'b00000000000000000111010000011011;
assign LUT_1[48578] = 32'b00000000000000001001101100110000;
assign LUT_1[48579] = 32'b00000000000000000010111110101100;
assign LUT_1[48580] = 32'b00000000000000010101110111110110;
assign LUT_1[48581] = 32'b00000000000000001111001001110010;
assign LUT_1[48582] = 32'b00000000000000010001100110000111;
assign LUT_1[48583] = 32'b00000000000000001010111000000011;
assign LUT_1[48584] = 32'b00000000000000001101001100010100;
assign LUT_1[48585] = 32'b00000000000000000110011110010000;
assign LUT_1[48586] = 32'b00000000000000001000111010100101;
assign LUT_1[48587] = 32'b00000000000000000010001100100001;
assign LUT_1[48588] = 32'b00000000000000010101000101101011;
assign LUT_1[48589] = 32'b00000000000000001110010111100111;
assign LUT_1[48590] = 32'b00000000000000010000110011111100;
assign LUT_1[48591] = 32'b00000000000000001010000101111000;
assign LUT_1[48592] = 32'b00000000000000001111111010000001;
assign LUT_1[48593] = 32'b00000000000000001001001011111101;
assign LUT_1[48594] = 32'b00000000000000001011101000010010;
assign LUT_1[48595] = 32'b00000000000000000100111010001110;
assign LUT_1[48596] = 32'b00000000000000010111110011011000;
assign LUT_1[48597] = 32'b00000000000000010001000101010100;
assign LUT_1[48598] = 32'b00000000000000010011100001101001;
assign LUT_1[48599] = 32'b00000000000000001100110011100101;
assign LUT_1[48600] = 32'b00000000000000001111000111110110;
assign LUT_1[48601] = 32'b00000000000000001000011001110010;
assign LUT_1[48602] = 32'b00000000000000001010110110000111;
assign LUT_1[48603] = 32'b00000000000000000100001000000011;
assign LUT_1[48604] = 32'b00000000000000010111000001001101;
assign LUT_1[48605] = 32'b00000000000000010000010011001001;
assign LUT_1[48606] = 32'b00000000000000010010101111011110;
assign LUT_1[48607] = 32'b00000000000000001100000001011010;
assign LUT_1[48608] = 32'b00000000000000001110111001011110;
assign LUT_1[48609] = 32'b00000000000000001000001011011010;
assign LUT_1[48610] = 32'b00000000000000001010100111101111;
assign LUT_1[48611] = 32'b00000000000000000011111001101011;
assign LUT_1[48612] = 32'b00000000000000010110110010110101;
assign LUT_1[48613] = 32'b00000000000000010000000100110001;
assign LUT_1[48614] = 32'b00000000000000010010100001000110;
assign LUT_1[48615] = 32'b00000000000000001011110011000010;
assign LUT_1[48616] = 32'b00000000000000001110000111010011;
assign LUT_1[48617] = 32'b00000000000000000111011001001111;
assign LUT_1[48618] = 32'b00000000000000001001110101100100;
assign LUT_1[48619] = 32'b00000000000000000011000111100000;
assign LUT_1[48620] = 32'b00000000000000010110000000101010;
assign LUT_1[48621] = 32'b00000000000000001111010010100110;
assign LUT_1[48622] = 32'b00000000000000010001101110111011;
assign LUT_1[48623] = 32'b00000000000000001011000000110111;
assign LUT_1[48624] = 32'b00000000000000010000110101000000;
assign LUT_1[48625] = 32'b00000000000000001010000110111100;
assign LUT_1[48626] = 32'b00000000000000001100100011010001;
assign LUT_1[48627] = 32'b00000000000000000101110101001101;
assign LUT_1[48628] = 32'b00000000000000011000101110010111;
assign LUT_1[48629] = 32'b00000000000000010010000000010011;
assign LUT_1[48630] = 32'b00000000000000010100011100101000;
assign LUT_1[48631] = 32'b00000000000000001101101110100100;
assign LUT_1[48632] = 32'b00000000000000010000000010110101;
assign LUT_1[48633] = 32'b00000000000000001001010100110001;
assign LUT_1[48634] = 32'b00000000000000001011110001000110;
assign LUT_1[48635] = 32'b00000000000000000101000011000010;
assign LUT_1[48636] = 32'b00000000000000010111111100001100;
assign LUT_1[48637] = 32'b00000000000000010001001110001000;
assign LUT_1[48638] = 32'b00000000000000010011101010011101;
assign LUT_1[48639] = 32'b00000000000000001100111100011001;
assign LUT_1[48640] = 32'b00000000000000000100111011000101;
assign LUT_1[48641] = 32'b11111111111111111110001101000001;
assign LUT_1[48642] = 32'b00000000000000000000101001010110;
assign LUT_1[48643] = 32'b11111111111111111001111011010010;
assign LUT_1[48644] = 32'b00000000000000001100110100011100;
assign LUT_1[48645] = 32'b00000000000000000110000110011000;
assign LUT_1[48646] = 32'b00000000000000001000100010101101;
assign LUT_1[48647] = 32'b00000000000000000001110100101001;
assign LUT_1[48648] = 32'b00000000000000000100001000111010;
assign LUT_1[48649] = 32'b11111111111111111101011010110110;
assign LUT_1[48650] = 32'b11111111111111111111110111001011;
assign LUT_1[48651] = 32'b11111111111111111001001001000111;
assign LUT_1[48652] = 32'b00000000000000001100000010010001;
assign LUT_1[48653] = 32'b00000000000000000101010100001101;
assign LUT_1[48654] = 32'b00000000000000000111110000100010;
assign LUT_1[48655] = 32'b00000000000000000001000010011110;
assign LUT_1[48656] = 32'b00000000000000000110110110100111;
assign LUT_1[48657] = 32'b00000000000000000000001000100011;
assign LUT_1[48658] = 32'b00000000000000000010100100111000;
assign LUT_1[48659] = 32'b11111111111111111011110110110100;
assign LUT_1[48660] = 32'b00000000000000001110101111111110;
assign LUT_1[48661] = 32'b00000000000000001000000001111010;
assign LUT_1[48662] = 32'b00000000000000001010011110001111;
assign LUT_1[48663] = 32'b00000000000000000011110000001011;
assign LUT_1[48664] = 32'b00000000000000000110000100011100;
assign LUT_1[48665] = 32'b11111111111111111111010110011000;
assign LUT_1[48666] = 32'b00000000000000000001110010101101;
assign LUT_1[48667] = 32'b11111111111111111011000100101001;
assign LUT_1[48668] = 32'b00000000000000001101111101110011;
assign LUT_1[48669] = 32'b00000000000000000111001111101111;
assign LUT_1[48670] = 32'b00000000000000001001101100000100;
assign LUT_1[48671] = 32'b00000000000000000010111110000000;
assign LUT_1[48672] = 32'b00000000000000000101110110000100;
assign LUT_1[48673] = 32'b11111111111111111111001000000000;
assign LUT_1[48674] = 32'b00000000000000000001100100010101;
assign LUT_1[48675] = 32'b11111111111111111010110110010001;
assign LUT_1[48676] = 32'b00000000000000001101101111011011;
assign LUT_1[48677] = 32'b00000000000000000111000001010111;
assign LUT_1[48678] = 32'b00000000000000001001011101101100;
assign LUT_1[48679] = 32'b00000000000000000010101111101000;
assign LUT_1[48680] = 32'b00000000000000000101000011111001;
assign LUT_1[48681] = 32'b11111111111111111110010101110101;
assign LUT_1[48682] = 32'b00000000000000000000110010001010;
assign LUT_1[48683] = 32'b11111111111111111010000100000110;
assign LUT_1[48684] = 32'b00000000000000001100111101010000;
assign LUT_1[48685] = 32'b00000000000000000110001111001100;
assign LUT_1[48686] = 32'b00000000000000001000101011100001;
assign LUT_1[48687] = 32'b00000000000000000001111101011101;
assign LUT_1[48688] = 32'b00000000000000000111110001100110;
assign LUT_1[48689] = 32'b00000000000000000001000011100010;
assign LUT_1[48690] = 32'b00000000000000000011011111110111;
assign LUT_1[48691] = 32'b11111111111111111100110001110011;
assign LUT_1[48692] = 32'b00000000000000001111101010111101;
assign LUT_1[48693] = 32'b00000000000000001000111100111001;
assign LUT_1[48694] = 32'b00000000000000001011011001001110;
assign LUT_1[48695] = 32'b00000000000000000100101011001010;
assign LUT_1[48696] = 32'b00000000000000000110111111011011;
assign LUT_1[48697] = 32'b00000000000000000000010001010111;
assign LUT_1[48698] = 32'b00000000000000000010101101101100;
assign LUT_1[48699] = 32'b11111111111111111011111111101000;
assign LUT_1[48700] = 32'b00000000000000001110111000110010;
assign LUT_1[48701] = 32'b00000000000000001000001010101110;
assign LUT_1[48702] = 32'b00000000000000001010100111000011;
assign LUT_1[48703] = 32'b00000000000000000011111000111111;
assign LUT_1[48704] = 32'b00000000000000000110111000101101;
assign LUT_1[48705] = 32'b00000000000000000000001010101001;
assign LUT_1[48706] = 32'b00000000000000000010100110111110;
assign LUT_1[48707] = 32'b11111111111111111011111000111010;
assign LUT_1[48708] = 32'b00000000000000001110110010000100;
assign LUT_1[48709] = 32'b00000000000000001000000100000000;
assign LUT_1[48710] = 32'b00000000000000001010100000010101;
assign LUT_1[48711] = 32'b00000000000000000011110010010001;
assign LUT_1[48712] = 32'b00000000000000000110000110100010;
assign LUT_1[48713] = 32'b11111111111111111111011000011110;
assign LUT_1[48714] = 32'b00000000000000000001110100110011;
assign LUT_1[48715] = 32'b11111111111111111011000110101111;
assign LUT_1[48716] = 32'b00000000000000001101111111111001;
assign LUT_1[48717] = 32'b00000000000000000111010001110101;
assign LUT_1[48718] = 32'b00000000000000001001101110001010;
assign LUT_1[48719] = 32'b00000000000000000011000000000110;
assign LUT_1[48720] = 32'b00000000000000001000110100001111;
assign LUT_1[48721] = 32'b00000000000000000010000110001011;
assign LUT_1[48722] = 32'b00000000000000000100100010100000;
assign LUT_1[48723] = 32'b11111111111111111101110100011100;
assign LUT_1[48724] = 32'b00000000000000010000101101100110;
assign LUT_1[48725] = 32'b00000000000000001001111111100010;
assign LUT_1[48726] = 32'b00000000000000001100011011110111;
assign LUT_1[48727] = 32'b00000000000000000101101101110011;
assign LUT_1[48728] = 32'b00000000000000001000000010000100;
assign LUT_1[48729] = 32'b00000000000000000001010100000000;
assign LUT_1[48730] = 32'b00000000000000000011110000010101;
assign LUT_1[48731] = 32'b11111111111111111101000010010001;
assign LUT_1[48732] = 32'b00000000000000001111111011011011;
assign LUT_1[48733] = 32'b00000000000000001001001101010111;
assign LUT_1[48734] = 32'b00000000000000001011101001101100;
assign LUT_1[48735] = 32'b00000000000000000100111011101000;
assign LUT_1[48736] = 32'b00000000000000000111110011101100;
assign LUT_1[48737] = 32'b00000000000000000001000101101000;
assign LUT_1[48738] = 32'b00000000000000000011100001111101;
assign LUT_1[48739] = 32'b11111111111111111100110011111001;
assign LUT_1[48740] = 32'b00000000000000001111101101000011;
assign LUT_1[48741] = 32'b00000000000000001000111110111111;
assign LUT_1[48742] = 32'b00000000000000001011011011010100;
assign LUT_1[48743] = 32'b00000000000000000100101101010000;
assign LUT_1[48744] = 32'b00000000000000000111000001100001;
assign LUT_1[48745] = 32'b00000000000000000000010011011101;
assign LUT_1[48746] = 32'b00000000000000000010101111110010;
assign LUT_1[48747] = 32'b11111111111111111100000001101110;
assign LUT_1[48748] = 32'b00000000000000001110111010111000;
assign LUT_1[48749] = 32'b00000000000000001000001100110100;
assign LUT_1[48750] = 32'b00000000000000001010101001001001;
assign LUT_1[48751] = 32'b00000000000000000011111011000101;
assign LUT_1[48752] = 32'b00000000000000001001101111001110;
assign LUT_1[48753] = 32'b00000000000000000011000001001010;
assign LUT_1[48754] = 32'b00000000000000000101011101011111;
assign LUT_1[48755] = 32'b11111111111111111110101111011011;
assign LUT_1[48756] = 32'b00000000000000010001101000100101;
assign LUT_1[48757] = 32'b00000000000000001010111010100001;
assign LUT_1[48758] = 32'b00000000000000001101010110110110;
assign LUT_1[48759] = 32'b00000000000000000110101000110010;
assign LUT_1[48760] = 32'b00000000000000001000111101000011;
assign LUT_1[48761] = 32'b00000000000000000010001110111111;
assign LUT_1[48762] = 32'b00000000000000000100101011010100;
assign LUT_1[48763] = 32'b11111111111111111101111101010000;
assign LUT_1[48764] = 32'b00000000000000010000110110011010;
assign LUT_1[48765] = 32'b00000000000000001010001000010110;
assign LUT_1[48766] = 32'b00000000000000001100100100101011;
assign LUT_1[48767] = 32'b00000000000000000101110110100111;
assign LUT_1[48768] = 32'b00000000000000000111111011001000;
assign LUT_1[48769] = 32'b00000000000000000001001101000100;
assign LUT_1[48770] = 32'b00000000000000000011101001011001;
assign LUT_1[48771] = 32'b11111111111111111100111011010101;
assign LUT_1[48772] = 32'b00000000000000001111110100011111;
assign LUT_1[48773] = 32'b00000000000000001001000110011011;
assign LUT_1[48774] = 32'b00000000000000001011100010110000;
assign LUT_1[48775] = 32'b00000000000000000100110100101100;
assign LUT_1[48776] = 32'b00000000000000000111001000111101;
assign LUT_1[48777] = 32'b00000000000000000000011010111001;
assign LUT_1[48778] = 32'b00000000000000000010110111001110;
assign LUT_1[48779] = 32'b11111111111111111100001001001010;
assign LUT_1[48780] = 32'b00000000000000001111000010010100;
assign LUT_1[48781] = 32'b00000000000000001000010100010000;
assign LUT_1[48782] = 32'b00000000000000001010110000100101;
assign LUT_1[48783] = 32'b00000000000000000100000010100001;
assign LUT_1[48784] = 32'b00000000000000001001110110101010;
assign LUT_1[48785] = 32'b00000000000000000011001000100110;
assign LUT_1[48786] = 32'b00000000000000000101100100111011;
assign LUT_1[48787] = 32'b11111111111111111110110110110111;
assign LUT_1[48788] = 32'b00000000000000010001110000000001;
assign LUT_1[48789] = 32'b00000000000000001011000001111101;
assign LUT_1[48790] = 32'b00000000000000001101011110010010;
assign LUT_1[48791] = 32'b00000000000000000110110000001110;
assign LUT_1[48792] = 32'b00000000000000001001000100011111;
assign LUT_1[48793] = 32'b00000000000000000010010110011011;
assign LUT_1[48794] = 32'b00000000000000000100110010110000;
assign LUT_1[48795] = 32'b11111111111111111110000100101100;
assign LUT_1[48796] = 32'b00000000000000010000111101110110;
assign LUT_1[48797] = 32'b00000000000000001010001111110010;
assign LUT_1[48798] = 32'b00000000000000001100101100000111;
assign LUT_1[48799] = 32'b00000000000000000101111110000011;
assign LUT_1[48800] = 32'b00000000000000001000110110000111;
assign LUT_1[48801] = 32'b00000000000000000010001000000011;
assign LUT_1[48802] = 32'b00000000000000000100100100011000;
assign LUT_1[48803] = 32'b11111111111111111101110110010100;
assign LUT_1[48804] = 32'b00000000000000010000101111011110;
assign LUT_1[48805] = 32'b00000000000000001010000001011010;
assign LUT_1[48806] = 32'b00000000000000001100011101101111;
assign LUT_1[48807] = 32'b00000000000000000101101111101011;
assign LUT_1[48808] = 32'b00000000000000001000000011111100;
assign LUT_1[48809] = 32'b00000000000000000001010101111000;
assign LUT_1[48810] = 32'b00000000000000000011110010001101;
assign LUT_1[48811] = 32'b11111111111111111101000100001001;
assign LUT_1[48812] = 32'b00000000000000001111111101010011;
assign LUT_1[48813] = 32'b00000000000000001001001111001111;
assign LUT_1[48814] = 32'b00000000000000001011101011100100;
assign LUT_1[48815] = 32'b00000000000000000100111101100000;
assign LUT_1[48816] = 32'b00000000000000001010110001101001;
assign LUT_1[48817] = 32'b00000000000000000100000011100101;
assign LUT_1[48818] = 32'b00000000000000000110011111111010;
assign LUT_1[48819] = 32'b11111111111111111111110001110110;
assign LUT_1[48820] = 32'b00000000000000010010101011000000;
assign LUT_1[48821] = 32'b00000000000000001011111100111100;
assign LUT_1[48822] = 32'b00000000000000001110011001010001;
assign LUT_1[48823] = 32'b00000000000000000111101011001101;
assign LUT_1[48824] = 32'b00000000000000001001111111011110;
assign LUT_1[48825] = 32'b00000000000000000011010001011010;
assign LUT_1[48826] = 32'b00000000000000000101101101101111;
assign LUT_1[48827] = 32'b11111111111111111110111111101011;
assign LUT_1[48828] = 32'b00000000000000010001111000110101;
assign LUT_1[48829] = 32'b00000000000000001011001010110001;
assign LUT_1[48830] = 32'b00000000000000001101100111000110;
assign LUT_1[48831] = 32'b00000000000000000110111001000010;
assign LUT_1[48832] = 32'b00000000000000001001111000110000;
assign LUT_1[48833] = 32'b00000000000000000011001010101100;
assign LUT_1[48834] = 32'b00000000000000000101100111000001;
assign LUT_1[48835] = 32'b11111111111111111110111000111101;
assign LUT_1[48836] = 32'b00000000000000010001110010000111;
assign LUT_1[48837] = 32'b00000000000000001011000100000011;
assign LUT_1[48838] = 32'b00000000000000001101100000011000;
assign LUT_1[48839] = 32'b00000000000000000110110010010100;
assign LUT_1[48840] = 32'b00000000000000001001000110100101;
assign LUT_1[48841] = 32'b00000000000000000010011000100001;
assign LUT_1[48842] = 32'b00000000000000000100110100110110;
assign LUT_1[48843] = 32'b11111111111111111110000110110010;
assign LUT_1[48844] = 32'b00000000000000010000111111111100;
assign LUT_1[48845] = 32'b00000000000000001010010001111000;
assign LUT_1[48846] = 32'b00000000000000001100101110001101;
assign LUT_1[48847] = 32'b00000000000000000110000000001001;
assign LUT_1[48848] = 32'b00000000000000001011110100010010;
assign LUT_1[48849] = 32'b00000000000000000101000110001110;
assign LUT_1[48850] = 32'b00000000000000000111100010100011;
assign LUT_1[48851] = 32'b00000000000000000000110100011111;
assign LUT_1[48852] = 32'b00000000000000010011101101101001;
assign LUT_1[48853] = 32'b00000000000000001100111111100101;
assign LUT_1[48854] = 32'b00000000000000001111011011111010;
assign LUT_1[48855] = 32'b00000000000000001000101101110110;
assign LUT_1[48856] = 32'b00000000000000001011000010000111;
assign LUT_1[48857] = 32'b00000000000000000100010100000011;
assign LUT_1[48858] = 32'b00000000000000000110110000011000;
assign LUT_1[48859] = 32'b00000000000000000000000010010100;
assign LUT_1[48860] = 32'b00000000000000010010111011011110;
assign LUT_1[48861] = 32'b00000000000000001100001101011010;
assign LUT_1[48862] = 32'b00000000000000001110101001101111;
assign LUT_1[48863] = 32'b00000000000000000111111011101011;
assign LUT_1[48864] = 32'b00000000000000001010110011101111;
assign LUT_1[48865] = 32'b00000000000000000100000101101011;
assign LUT_1[48866] = 32'b00000000000000000110100010000000;
assign LUT_1[48867] = 32'b11111111111111111111110011111100;
assign LUT_1[48868] = 32'b00000000000000010010101101000110;
assign LUT_1[48869] = 32'b00000000000000001011111111000010;
assign LUT_1[48870] = 32'b00000000000000001110011011010111;
assign LUT_1[48871] = 32'b00000000000000000111101101010011;
assign LUT_1[48872] = 32'b00000000000000001010000001100100;
assign LUT_1[48873] = 32'b00000000000000000011010011100000;
assign LUT_1[48874] = 32'b00000000000000000101101111110101;
assign LUT_1[48875] = 32'b11111111111111111111000001110001;
assign LUT_1[48876] = 32'b00000000000000010001111010111011;
assign LUT_1[48877] = 32'b00000000000000001011001100110111;
assign LUT_1[48878] = 32'b00000000000000001101101001001100;
assign LUT_1[48879] = 32'b00000000000000000110111011001000;
assign LUT_1[48880] = 32'b00000000000000001100101111010001;
assign LUT_1[48881] = 32'b00000000000000000110000001001101;
assign LUT_1[48882] = 32'b00000000000000001000011101100010;
assign LUT_1[48883] = 32'b00000000000000000001101111011110;
assign LUT_1[48884] = 32'b00000000000000010100101000101000;
assign LUT_1[48885] = 32'b00000000000000001101111010100100;
assign LUT_1[48886] = 32'b00000000000000010000010110111001;
assign LUT_1[48887] = 32'b00000000000000001001101000110101;
assign LUT_1[48888] = 32'b00000000000000001011111101000110;
assign LUT_1[48889] = 32'b00000000000000000101001111000010;
assign LUT_1[48890] = 32'b00000000000000000111101011010111;
assign LUT_1[48891] = 32'b00000000000000000000111101010011;
assign LUT_1[48892] = 32'b00000000000000010011110110011101;
assign LUT_1[48893] = 32'b00000000000000001101001000011001;
assign LUT_1[48894] = 32'b00000000000000001111100100101110;
assign LUT_1[48895] = 32'b00000000000000001000110110101010;
assign LUT_1[48896] = 32'b00000000000000000010101111010001;
assign LUT_1[48897] = 32'b11111111111111111100000001001101;
assign LUT_1[48898] = 32'b11111111111111111110011101100010;
assign LUT_1[48899] = 32'b11111111111111110111101111011110;
assign LUT_1[48900] = 32'b00000000000000001010101000101000;
assign LUT_1[48901] = 32'b00000000000000000011111010100100;
assign LUT_1[48902] = 32'b00000000000000000110010110111001;
assign LUT_1[48903] = 32'b11111111111111111111101000110101;
assign LUT_1[48904] = 32'b00000000000000000001111101000110;
assign LUT_1[48905] = 32'b11111111111111111011001111000010;
assign LUT_1[48906] = 32'b11111111111111111101101011010111;
assign LUT_1[48907] = 32'b11111111111111110110111101010011;
assign LUT_1[48908] = 32'b00000000000000001001110110011101;
assign LUT_1[48909] = 32'b00000000000000000011001000011001;
assign LUT_1[48910] = 32'b00000000000000000101100100101110;
assign LUT_1[48911] = 32'b11111111111111111110110110101010;
assign LUT_1[48912] = 32'b00000000000000000100101010110011;
assign LUT_1[48913] = 32'b11111111111111111101111100101111;
assign LUT_1[48914] = 32'b00000000000000000000011001000100;
assign LUT_1[48915] = 32'b11111111111111111001101011000000;
assign LUT_1[48916] = 32'b00000000000000001100100100001010;
assign LUT_1[48917] = 32'b00000000000000000101110110000110;
assign LUT_1[48918] = 32'b00000000000000001000010010011011;
assign LUT_1[48919] = 32'b00000000000000000001100100010111;
assign LUT_1[48920] = 32'b00000000000000000011111000101000;
assign LUT_1[48921] = 32'b11111111111111111101001010100100;
assign LUT_1[48922] = 32'b11111111111111111111100110111001;
assign LUT_1[48923] = 32'b11111111111111111000111000110101;
assign LUT_1[48924] = 32'b00000000000000001011110001111111;
assign LUT_1[48925] = 32'b00000000000000000101000011111011;
assign LUT_1[48926] = 32'b00000000000000000111100000010000;
assign LUT_1[48927] = 32'b00000000000000000000110010001100;
assign LUT_1[48928] = 32'b00000000000000000011101010010000;
assign LUT_1[48929] = 32'b11111111111111111100111100001100;
assign LUT_1[48930] = 32'b11111111111111111111011000100001;
assign LUT_1[48931] = 32'b11111111111111111000101010011101;
assign LUT_1[48932] = 32'b00000000000000001011100011100111;
assign LUT_1[48933] = 32'b00000000000000000100110101100011;
assign LUT_1[48934] = 32'b00000000000000000111010001111000;
assign LUT_1[48935] = 32'b00000000000000000000100011110100;
assign LUT_1[48936] = 32'b00000000000000000010111000000101;
assign LUT_1[48937] = 32'b11111111111111111100001010000001;
assign LUT_1[48938] = 32'b11111111111111111110100110010110;
assign LUT_1[48939] = 32'b11111111111111110111111000010010;
assign LUT_1[48940] = 32'b00000000000000001010110001011100;
assign LUT_1[48941] = 32'b00000000000000000100000011011000;
assign LUT_1[48942] = 32'b00000000000000000110011111101101;
assign LUT_1[48943] = 32'b11111111111111111111110001101001;
assign LUT_1[48944] = 32'b00000000000000000101100101110010;
assign LUT_1[48945] = 32'b11111111111111111110110111101110;
assign LUT_1[48946] = 32'b00000000000000000001010100000011;
assign LUT_1[48947] = 32'b11111111111111111010100101111111;
assign LUT_1[48948] = 32'b00000000000000001101011111001001;
assign LUT_1[48949] = 32'b00000000000000000110110001000101;
assign LUT_1[48950] = 32'b00000000000000001001001101011010;
assign LUT_1[48951] = 32'b00000000000000000010011111010110;
assign LUT_1[48952] = 32'b00000000000000000100110011100111;
assign LUT_1[48953] = 32'b11111111111111111110000101100011;
assign LUT_1[48954] = 32'b00000000000000000000100001111000;
assign LUT_1[48955] = 32'b11111111111111111001110011110100;
assign LUT_1[48956] = 32'b00000000000000001100101100111110;
assign LUT_1[48957] = 32'b00000000000000000101111110111010;
assign LUT_1[48958] = 32'b00000000000000001000011011001111;
assign LUT_1[48959] = 32'b00000000000000000001101101001011;
assign LUT_1[48960] = 32'b00000000000000000100101100111001;
assign LUT_1[48961] = 32'b11111111111111111101111110110101;
assign LUT_1[48962] = 32'b00000000000000000000011011001010;
assign LUT_1[48963] = 32'b11111111111111111001101101000110;
assign LUT_1[48964] = 32'b00000000000000001100100110010000;
assign LUT_1[48965] = 32'b00000000000000000101111000001100;
assign LUT_1[48966] = 32'b00000000000000001000010100100001;
assign LUT_1[48967] = 32'b00000000000000000001100110011101;
assign LUT_1[48968] = 32'b00000000000000000011111010101110;
assign LUT_1[48969] = 32'b11111111111111111101001100101010;
assign LUT_1[48970] = 32'b11111111111111111111101000111111;
assign LUT_1[48971] = 32'b11111111111111111000111010111011;
assign LUT_1[48972] = 32'b00000000000000001011110100000101;
assign LUT_1[48973] = 32'b00000000000000000101000110000001;
assign LUT_1[48974] = 32'b00000000000000000111100010010110;
assign LUT_1[48975] = 32'b00000000000000000000110100010010;
assign LUT_1[48976] = 32'b00000000000000000110101000011011;
assign LUT_1[48977] = 32'b11111111111111111111111010010111;
assign LUT_1[48978] = 32'b00000000000000000010010110101100;
assign LUT_1[48979] = 32'b11111111111111111011101000101000;
assign LUT_1[48980] = 32'b00000000000000001110100001110010;
assign LUT_1[48981] = 32'b00000000000000000111110011101110;
assign LUT_1[48982] = 32'b00000000000000001010010000000011;
assign LUT_1[48983] = 32'b00000000000000000011100001111111;
assign LUT_1[48984] = 32'b00000000000000000101110110010000;
assign LUT_1[48985] = 32'b11111111111111111111001000001100;
assign LUT_1[48986] = 32'b00000000000000000001100100100001;
assign LUT_1[48987] = 32'b11111111111111111010110110011101;
assign LUT_1[48988] = 32'b00000000000000001101101111100111;
assign LUT_1[48989] = 32'b00000000000000000111000001100011;
assign LUT_1[48990] = 32'b00000000000000001001011101111000;
assign LUT_1[48991] = 32'b00000000000000000010101111110100;
assign LUT_1[48992] = 32'b00000000000000000101100111111000;
assign LUT_1[48993] = 32'b11111111111111111110111001110100;
assign LUT_1[48994] = 32'b00000000000000000001010110001001;
assign LUT_1[48995] = 32'b11111111111111111010101000000101;
assign LUT_1[48996] = 32'b00000000000000001101100001001111;
assign LUT_1[48997] = 32'b00000000000000000110110011001011;
assign LUT_1[48998] = 32'b00000000000000001001001111100000;
assign LUT_1[48999] = 32'b00000000000000000010100001011100;
assign LUT_1[49000] = 32'b00000000000000000100110101101101;
assign LUT_1[49001] = 32'b11111111111111111110000111101001;
assign LUT_1[49002] = 32'b00000000000000000000100011111110;
assign LUT_1[49003] = 32'b11111111111111111001110101111010;
assign LUT_1[49004] = 32'b00000000000000001100101111000100;
assign LUT_1[49005] = 32'b00000000000000000110000001000000;
assign LUT_1[49006] = 32'b00000000000000001000011101010101;
assign LUT_1[49007] = 32'b00000000000000000001101111010001;
assign LUT_1[49008] = 32'b00000000000000000111100011011010;
assign LUT_1[49009] = 32'b00000000000000000000110101010110;
assign LUT_1[49010] = 32'b00000000000000000011010001101011;
assign LUT_1[49011] = 32'b11111111111111111100100011100111;
assign LUT_1[49012] = 32'b00000000000000001111011100110001;
assign LUT_1[49013] = 32'b00000000000000001000101110101101;
assign LUT_1[49014] = 32'b00000000000000001011001011000010;
assign LUT_1[49015] = 32'b00000000000000000100011100111110;
assign LUT_1[49016] = 32'b00000000000000000110110001001111;
assign LUT_1[49017] = 32'b00000000000000000000000011001011;
assign LUT_1[49018] = 32'b00000000000000000010011111100000;
assign LUT_1[49019] = 32'b11111111111111111011110001011100;
assign LUT_1[49020] = 32'b00000000000000001110101010100110;
assign LUT_1[49021] = 32'b00000000000000000111111100100010;
assign LUT_1[49022] = 32'b00000000000000001010011000110111;
assign LUT_1[49023] = 32'b00000000000000000011101010110011;
assign LUT_1[49024] = 32'b00000000000000000101101111010100;
assign LUT_1[49025] = 32'b11111111111111111111000001010000;
assign LUT_1[49026] = 32'b00000000000000000001011101100101;
assign LUT_1[49027] = 32'b11111111111111111010101111100001;
assign LUT_1[49028] = 32'b00000000000000001101101000101011;
assign LUT_1[49029] = 32'b00000000000000000110111010100111;
assign LUT_1[49030] = 32'b00000000000000001001010110111100;
assign LUT_1[49031] = 32'b00000000000000000010101000111000;
assign LUT_1[49032] = 32'b00000000000000000100111101001001;
assign LUT_1[49033] = 32'b11111111111111111110001111000101;
assign LUT_1[49034] = 32'b00000000000000000000101011011010;
assign LUT_1[49035] = 32'b11111111111111111001111101010110;
assign LUT_1[49036] = 32'b00000000000000001100110110100000;
assign LUT_1[49037] = 32'b00000000000000000110001000011100;
assign LUT_1[49038] = 32'b00000000000000001000100100110001;
assign LUT_1[49039] = 32'b00000000000000000001110110101101;
assign LUT_1[49040] = 32'b00000000000000000111101010110110;
assign LUT_1[49041] = 32'b00000000000000000000111100110010;
assign LUT_1[49042] = 32'b00000000000000000011011001000111;
assign LUT_1[49043] = 32'b11111111111111111100101011000011;
assign LUT_1[49044] = 32'b00000000000000001111100100001101;
assign LUT_1[49045] = 32'b00000000000000001000110110001001;
assign LUT_1[49046] = 32'b00000000000000001011010010011110;
assign LUT_1[49047] = 32'b00000000000000000100100100011010;
assign LUT_1[49048] = 32'b00000000000000000110111000101011;
assign LUT_1[49049] = 32'b00000000000000000000001010100111;
assign LUT_1[49050] = 32'b00000000000000000010100110111100;
assign LUT_1[49051] = 32'b11111111111111111011111000111000;
assign LUT_1[49052] = 32'b00000000000000001110110010000010;
assign LUT_1[49053] = 32'b00000000000000001000000011111110;
assign LUT_1[49054] = 32'b00000000000000001010100000010011;
assign LUT_1[49055] = 32'b00000000000000000011110010001111;
assign LUT_1[49056] = 32'b00000000000000000110101010010011;
assign LUT_1[49057] = 32'b11111111111111111111111100001111;
assign LUT_1[49058] = 32'b00000000000000000010011000100100;
assign LUT_1[49059] = 32'b11111111111111111011101010100000;
assign LUT_1[49060] = 32'b00000000000000001110100011101010;
assign LUT_1[49061] = 32'b00000000000000000111110101100110;
assign LUT_1[49062] = 32'b00000000000000001010010001111011;
assign LUT_1[49063] = 32'b00000000000000000011100011110111;
assign LUT_1[49064] = 32'b00000000000000000101111000001000;
assign LUT_1[49065] = 32'b11111111111111111111001010000100;
assign LUT_1[49066] = 32'b00000000000000000001100110011001;
assign LUT_1[49067] = 32'b11111111111111111010111000010101;
assign LUT_1[49068] = 32'b00000000000000001101110001011111;
assign LUT_1[49069] = 32'b00000000000000000111000011011011;
assign LUT_1[49070] = 32'b00000000000000001001011111110000;
assign LUT_1[49071] = 32'b00000000000000000010110001101100;
assign LUT_1[49072] = 32'b00000000000000001000100101110101;
assign LUT_1[49073] = 32'b00000000000000000001110111110001;
assign LUT_1[49074] = 32'b00000000000000000100010100000110;
assign LUT_1[49075] = 32'b11111111111111111101100110000010;
assign LUT_1[49076] = 32'b00000000000000010000011111001100;
assign LUT_1[49077] = 32'b00000000000000001001110001001000;
assign LUT_1[49078] = 32'b00000000000000001100001101011101;
assign LUT_1[49079] = 32'b00000000000000000101011111011001;
assign LUT_1[49080] = 32'b00000000000000000111110011101010;
assign LUT_1[49081] = 32'b00000000000000000001000101100110;
assign LUT_1[49082] = 32'b00000000000000000011100001111011;
assign LUT_1[49083] = 32'b11111111111111111100110011110111;
assign LUT_1[49084] = 32'b00000000000000001111101101000001;
assign LUT_1[49085] = 32'b00000000000000001000111110111101;
assign LUT_1[49086] = 32'b00000000000000001011011011010010;
assign LUT_1[49087] = 32'b00000000000000000100101101001110;
assign LUT_1[49088] = 32'b00000000000000000111101100111100;
assign LUT_1[49089] = 32'b00000000000000000000111110111000;
assign LUT_1[49090] = 32'b00000000000000000011011011001101;
assign LUT_1[49091] = 32'b11111111111111111100101101001001;
assign LUT_1[49092] = 32'b00000000000000001111100110010011;
assign LUT_1[49093] = 32'b00000000000000001000111000001111;
assign LUT_1[49094] = 32'b00000000000000001011010100100100;
assign LUT_1[49095] = 32'b00000000000000000100100110100000;
assign LUT_1[49096] = 32'b00000000000000000110111010110001;
assign LUT_1[49097] = 32'b00000000000000000000001100101101;
assign LUT_1[49098] = 32'b00000000000000000010101001000010;
assign LUT_1[49099] = 32'b11111111111111111011111010111110;
assign LUT_1[49100] = 32'b00000000000000001110110100001000;
assign LUT_1[49101] = 32'b00000000000000001000000110000100;
assign LUT_1[49102] = 32'b00000000000000001010100010011001;
assign LUT_1[49103] = 32'b00000000000000000011110100010101;
assign LUT_1[49104] = 32'b00000000000000001001101000011110;
assign LUT_1[49105] = 32'b00000000000000000010111010011010;
assign LUT_1[49106] = 32'b00000000000000000101010110101111;
assign LUT_1[49107] = 32'b11111111111111111110101000101011;
assign LUT_1[49108] = 32'b00000000000000010001100001110101;
assign LUT_1[49109] = 32'b00000000000000001010110011110001;
assign LUT_1[49110] = 32'b00000000000000001101010000000110;
assign LUT_1[49111] = 32'b00000000000000000110100010000010;
assign LUT_1[49112] = 32'b00000000000000001000110110010011;
assign LUT_1[49113] = 32'b00000000000000000010001000001111;
assign LUT_1[49114] = 32'b00000000000000000100100100100100;
assign LUT_1[49115] = 32'b11111111111111111101110110100000;
assign LUT_1[49116] = 32'b00000000000000010000101111101010;
assign LUT_1[49117] = 32'b00000000000000001010000001100110;
assign LUT_1[49118] = 32'b00000000000000001100011101111011;
assign LUT_1[49119] = 32'b00000000000000000101101111110111;
assign LUT_1[49120] = 32'b00000000000000001000100111111011;
assign LUT_1[49121] = 32'b00000000000000000001111001110111;
assign LUT_1[49122] = 32'b00000000000000000100010110001100;
assign LUT_1[49123] = 32'b11111111111111111101101000001000;
assign LUT_1[49124] = 32'b00000000000000010000100001010010;
assign LUT_1[49125] = 32'b00000000000000001001110011001110;
assign LUT_1[49126] = 32'b00000000000000001100001111100011;
assign LUT_1[49127] = 32'b00000000000000000101100001011111;
assign LUT_1[49128] = 32'b00000000000000000111110101110000;
assign LUT_1[49129] = 32'b00000000000000000001000111101100;
assign LUT_1[49130] = 32'b00000000000000000011100100000001;
assign LUT_1[49131] = 32'b11111111111111111100110101111101;
assign LUT_1[49132] = 32'b00000000000000001111101111000111;
assign LUT_1[49133] = 32'b00000000000000001001000001000011;
assign LUT_1[49134] = 32'b00000000000000001011011101011000;
assign LUT_1[49135] = 32'b00000000000000000100101111010100;
assign LUT_1[49136] = 32'b00000000000000001010100011011101;
assign LUT_1[49137] = 32'b00000000000000000011110101011001;
assign LUT_1[49138] = 32'b00000000000000000110010001101110;
assign LUT_1[49139] = 32'b11111111111111111111100011101010;
assign LUT_1[49140] = 32'b00000000000000010010011100110100;
assign LUT_1[49141] = 32'b00000000000000001011101110110000;
assign LUT_1[49142] = 32'b00000000000000001110001011000101;
assign LUT_1[49143] = 32'b00000000000000000111011101000001;
assign LUT_1[49144] = 32'b00000000000000001001110001010010;
assign LUT_1[49145] = 32'b00000000000000000011000011001110;
assign LUT_1[49146] = 32'b00000000000000000101011111100011;
assign LUT_1[49147] = 32'b11111111111111111110110001011111;
assign LUT_1[49148] = 32'b00000000000000010001101010101001;
assign LUT_1[49149] = 32'b00000000000000001010111100100101;
assign LUT_1[49150] = 32'b00000000000000001101011000111010;
assign LUT_1[49151] = 32'b00000000000000000110101010110110;
assign LUT_1[49152] = 32'b11111111111111111111001010010001;
assign LUT_1[49153] = 32'b11111111111111111000011100001101;
assign LUT_1[49154] = 32'b11111111111111111010111000100010;
assign LUT_1[49155] = 32'b11111111111111110100001010011110;
assign LUT_1[49156] = 32'b00000000000000000111000011101000;
assign LUT_1[49157] = 32'b00000000000000000000010101100100;
assign LUT_1[49158] = 32'b00000000000000000010110001111001;
assign LUT_1[49159] = 32'b11111111111111111100000011110101;
assign LUT_1[49160] = 32'b11111111111111111110011000000110;
assign LUT_1[49161] = 32'b11111111111111110111101010000010;
assign LUT_1[49162] = 32'b11111111111111111010000110010111;
assign LUT_1[49163] = 32'b11111111111111110011011000010011;
assign LUT_1[49164] = 32'b00000000000000000110010001011101;
assign LUT_1[49165] = 32'b11111111111111111111100011011001;
assign LUT_1[49166] = 32'b00000000000000000001111111101110;
assign LUT_1[49167] = 32'b11111111111111111011010001101010;
assign LUT_1[49168] = 32'b00000000000000000001000101110011;
assign LUT_1[49169] = 32'b11111111111111111010010111101111;
assign LUT_1[49170] = 32'b11111111111111111100110100000100;
assign LUT_1[49171] = 32'b11111111111111110110000110000000;
assign LUT_1[49172] = 32'b00000000000000001000111111001010;
assign LUT_1[49173] = 32'b00000000000000000010010001000110;
assign LUT_1[49174] = 32'b00000000000000000100101101011011;
assign LUT_1[49175] = 32'b11111111111111111101111111010111;
assign LUT_1[49176] = 32'b00000000000000000000010011101000;
assign LUT_1[49177] = 32'b11111111111111111001100101100100;
assign LUT_1[49178] = 32'b11111111111111111100000001111001;
assign LUT_1[49179] = 32'b11111111111111110101010011110101;
assign LUT_1[49180] = 32'b00000000000000001000001100111111;
assign LUT_1[49181] = 32'b00000000000000000001011110111011;
assign LUT_1[49182] = 32'b00000000000000000011111011010000;
assign LUT_1[49183] = 32'b11111111111111111101001101001100;
assign LUT_1[49184] = 32'b00000000000000000000000101010000;
assign LUT_1[49185] = 32'b11111111111111111001010111001100;
assign LUT_1[49186] = 32'b11111111111111111011110011100001;
assign LUT_1[49187] = 32'b11111111111111110101000101011101;
assign LUT_1[49188] = 32'b00000000000000000111111110100111;
assign LUT_1[49189] = 32'b00000000000000000001010000100011;
assign LUT_1[49190] = 32'b00000000000000000011101100111000;
assign LUT_1[49191] = 32'b11111111111111111100111110110100;
assign LUT_1[49192] = 32'b11111111111111111111010011000101;
assign LUT_1[49193] = 32'b11111111111111111000100101000001;
assign LUT_1[49194] = 32'b11111111111111111011000001010110;
assign LUT_1[49195] = 32'b11111111111111110100010011010010;
assign LUT_1[49196] = 32'b00000000000000000111001100011100;
assign LUT_1[49197] = 32'b00000000000000000000011110011000;
assign LUT_1[49198] = 32'b00000000000000000010111010101101;
assign LUT_1[49199] = 32'b11111111111111111100001100101001;
assign LUT_1[49200] = 32'b00000000000000000010000000110010;
assign LUT_1[49201] = 32'b11111111111111111011010010101110;
assign LUT_1[49202] = 32'b11111111111111111101101111000011;
assign LUT_1[49203] = 32'b11111111111111110111000000111111;
assign LUT_1[49204] = 32'b00000000000000001001111010001001;
assign LUT_1[49205] = 32'b00000000000000000011001100000101;
assign LUT_1[49206] = 32'b00000000000000000101101000011010;
assign LUT_1[49207] = 32'b11111111111111111110111010010110;
assign LUT_1[49208] = 32'b00000000000000000001001110100111;
assign LUT_1[49209] = 32'b11111111111111111010100000100011;
assign LUT_1[49210] = 32'b11111111111111111100111100111000;
assign LUT_1[49211] = 32'b11111111111111110110001110110100;
assign LUT_1[49212] = 32'b00000000000000001001000111111110;
assign LUT_1[49213] = 32'b00000000000000000010011001111010;
assign LUT_1[49214] = 32'b00000000000000000100110110001111;
assign LUT_1[49215] = 32'b11111111111111111110001000001011;
assign LUT_1[49216] = 32'b00000000000000000001000111111001;
assign LUT_1[49217] = 32'b11111111111111111010011001110101;
assign LUT_1[49218] = 32'b11111111111111111100110110001010;
assign LUT_1[49219] = 32'b11111111111111110110001000000110;
assign LUT_1[49220] = 32'b00000000000000001001000001010000;
assign LUT_1[49221] = 32'b00000000000000000010010011001100;
assign LUT_1[49222] = 32'b00000000000000000100101111100001;
assign LUT_1[49223] = 32'b11111111111111111110000001011101;
assign LUT_1[49224] = 32'b00000000000000000000010101101110;
assign LUT_1[49225] = 32'b11111111111111111001100111101010;
assign LUT_1[49226] = 32'b11111111111111111100000011111111;
assign LUT_1[49227] = 32'b11111111111111110101010101111011;
assign LUT_1[49228] = 32'b00000000000000001000001111000101;
assign LUT_1[49229] = 32'b00000000000000000001100001000001;
assign LUT_1[49230] = 32'b00000000000000000011111101010110;
assign LUT_1[49231] = 32'b11111111111111111101001111010010;
assign LUT_1[49232] = 32'b00000000000000000011000011011011;
assign LUT_1[49233] = 32'b11111111111111111100010101010111;
assign LUT_1[49234] = 32'b11111111111111111110110001101100;
assign LUT_1[49235] = 32'b11111111111111111000000011101000;
assign LUT_1[49236] = 32'b00000000000000001010111100110010;
assign LUT_1[49237] = 32'b00000000000000000100001110101110;
assign LUT_1[49238] = 32'b00000000000000000110101011000011;
assign LUT_1[49239] = 32'b11111111111111111111111100111111;
assign LUT_1[49240] = 32'b00000000000000000010010001010000;
assign LUT_1[49241] = 32'b11111111111111111011100011001100;
assign LUT_1[49242] = 32'b11111111111111111101111111100001;
assign LUT_1[49243] = 32'b11111111111111110111010001011101;
assign LUT_1[49244] = 32'b00000000000000001010001010100111;
assign LUT_1[49245] = 32'b00000000000000000011011100100011;
assign LUT_1[49246] = 32'b00000000000000000101111000111000;
assign LUT_1[49247] = 32'b11111111111111111111001010110100;
assign LUT_1[49248] = 32'b00000000000000000010000010111000;
assign LUT_1[49249] = 32'b11111111111111111011010100110100;
assign LUT_1[49250] = 32'b11111111111111111101110001001001;
assign LUT_1[49251] = 32'b11111111111111110111000011000101;
assign LUT_1[49252] = 32'b00000000000000001001111100001111;
assign LUT_1[49253] = 32'b00000000000000000011001110001011;
assign LUT_1[49254] = 32'b00000000000000000101101010100000;
assign LUT_1[49255] = 32'b11111111111111111110111100011100;
assign LUT_1[49256] = 32'b00000000000000000001010000101101;
assign LUT_1[49257] = 32'b11111111111111111010100010101001;
assign LUT_1[49258] = 32'b11111111111111111100111110111110;
assign LUT_1[49259] = 32'b11111111111111110110010000111010;
assign LUT_1[49260] = 32'b00000000000000001001001010000100;
assign LUT_1[49261] = 32'b00000000000000000010011100000000;
assign LUT_1[49262] = 32'b00000000000000000100111000010101;
assign LUT_1[49263] = 32'b11111111111111111110001010010001;
assign LUT_1[49264] = 32'b00000000000000000011111110011010;
assign LUT_1[49265] = 32'b11111111111111111101010000010110;
assign LUT_1[49266] = 32'b11111111111111111111101100101011;
assign LUT_1[49267] = 32'b11111111111111111000111110100111;
assign LUT_1[49268] = 32'b00000000000000001011110111110001;
assign LUT_1[49269] = 32'b00000000000000000101001001101101;
assign LUT_1[49270] = 32'b00000000000000000111100110000010;
assign LUT_1[49271] = 32'b00000000000000000000110111111110;
assign LUT_1[49272] = 32'b00000000000000000011001100001111;
assign LUT_1[49273] = 32'b11111111111111111100011110001011;
assign LUT_1[49274] = 32'b11111111111111111110111010100000;
assign LUT_1[49275] = 32'b11111111111111111000001100011100;
assign LUT_1[49276] = 32'b00000000000000001011000101100110;
assign LUT_1[49277] = 32'b00000000000000000100010111100010;
assign LUT_1[49278] = 32'b00000000000000000110110011110111;
assign LUT_1[49279] = 32'b00000000000000000000000101110011;
assign LUT_1[49280] = 32'b00000000000000000010001010010100;
assign LUT_1[49281] = 32'b11111111111111111011011100010000;
assign LUT_1[49282] = 32'b11111111111111111101111000100101;
assign LUT_1[49283] = 32'b11111111111111110111001010100001;
assign LUT_1[49284] = 32'b00000000000000001010000011101011;
assign LUT_1[49285] = 32'b00000000000000000011010101100111;
assign LUT_1[49286] = 32'b00000000000000000101110001111100;
assign LUT_1[49287] = 32'b11111111111111111111000011111000;
assign LUT_1[49288] = 32'b00000000000000000001011000001001;
assign LUT_1[49289] = 32'b11111111111111111010101010000101;
assign LUT_1[49290] = 32'b11111111111111111101000110011010;
assign LUT_1[49291] = 32'b11111111111111110110011000010110;
assign LUT_1[49292] = 32'b00000000000000001001010001100000;
assign LUT_1[49293] = 32'b00000000000000000010100011011100;
assign LUT_1[49294] = 32'b00000000000000000100111111110001;
assign LUT_1[49295] = 32'b11111111111111111110010001101101;
assign LUT_1[49296] = 32'b00000000000000000100000101110110;
assign LUT_1[49297] = 32'b11111111111111111101010111110010;
assign LUT_1[49298] = 32'b11111111111111111111110100000111;
assign LUT_1[49299] = 32'b11111111111111111001000110000011;
assign LUT_1[49300] = 32'b00000000000000001011111111001101;
assign LUT_1[49301] = 32'b00000000000000000101010001001001;
assign LUT_1[49302] = 32'b00000000000000000111101101011110;
assign LUT_1[49303] = 32'b00000000000000000000111111011010;
assign LUT_1[49304] = 32'b00000000000000000011010011101011;
assign LUT_1[49305] = 32'b11111111111111111100100101100111;
assign LUT_1[49306] = 32'b11111111111111111111000001111100;
assign LUT_1[49307] = 32'b11111111111111111000010011111000;
assign LUT_1[49308] = 32'b00000000000000001011001101000010;
assign LUT_1[49309] = 32'b00000000000000000100011110111110;
assign LUT_1[49310] = 32'b00000000000000000110111011010011;
assign LUT_1[49311] = 32'b00000000000000000000001101001111;
assign LUT_1[49312] = 32'b00000000000000000011000101010011;
assign LUT_1[49313] = 32'b11111111111111111100010111001111;
assign LUT_1[49314] = 32'b11111111111111111110110011100100;
assign LUT_1[49315] = 32'b11111111111111111000000101100000;
assign LUT_1[49316] = 32'b00000000000000001010111110101010;
assign LUT_1[49317] = 32'b00000000000000000100010000100110;
assign LUT_1[49318] = 32'b00000000000000000110101100111011;
assign LUT_1[49319] = 32'b11111111111111111111111110110111;
assign LUT_1[49320] = 32'b00000000000000000010010011001000;
assign LUT_1[49321] = 32'b11111111111111111011100101000100;
assign LUT_1[49322] = 32'b11111111111111111110000001011001;
assign LUT_1[49323] = 32'b11111111111111110111010011010101;
assign LUT_1[49324] = 32'b00000000000000001010001100011111;
assign LUT_1[49325] = 32'b00000000000000000011011110011011;
assign LUT_1[49326] = 32'b00000000000000000101111010110000;
assign LUT_1[49327] = 32'b11111111111111111111001100101100;
assign LUT_1[49328] = 32'b00000000000000000101000000110101;
assign LUT_1[49329] = 32'b11111111111111111110010010110001;
assign LUT_1[49330] = 32'b00000000000000000000101111000110;
assign LUT_1[49331] = 32'b11111111111111111010000001000010;
assign LUT_1[49332] = 32'b00000000000000001100111010001100;
assign LUT_1[49333] = 32'b00000000000000000110001100001000;
assign LUT_1[49334] = 32'b00000000000000001000101000011101;
assign LUT_1[49335] = 32'b00000000000000000001111010011001;
assign LUT_1[49336] = 32'b00000000000000000100001110101010;
assign LUT_1[49337] = 32'b11111111111111111101100000100110;
assign LUT_1[49338] = 32'b11111111111111111111111100111011;
assign LUT_1[49339] = 32'b11111111111111111001001110110111;
assign LUT_1[49340] = 32'b00000000000000001100001000000001;
assign LUT_1[49341] = 32'b00000000000000000101011001111101;
assign LUT_1[49342] = 32'b00000000000000000111110110010010;
assign LUT_1[49343] = 32'b00000000000000000001001000001110;
assign LUT_1[49344] = 32'b00000000000000000100000111111100;
assign LUT_1[49345] = 32'b11111111111111111101011001111000;
assign LUT_1[49346] = 32'b11111111111111111111110110001101;
assign LUT_1[49347] = 32'b11111111111111111001001000001001;
assign LUT_1[49348] = 32'b00000000000000001100000001010011;
assign LUT_1[49349] = 32'b00000000000000000101010011001111;
assign LUT_1[49350] = 32'b00000000000000000111101111100100;
assign LUT_1[49351] = 32'b00000000000000000001000001100000;
assign LUT_1[49352] = 32'b00000000000000000011010101110001;
assign LUT_1[49353] = 32'b11111111111111111100100111101101;
assign LUT_1[49354] = 32'b11111111111111111111000100000010;
assign LUT_1[49355] = 32'b11111111111111111000010101111110;
assign LUT_1[49356] = 32'b00000000000000001011001111001000;
assign LUT_1[49357] = 32'b00000000000000000100100001000100;
assign LUT_1[49358] = 32'b00000000000000000110111101011001;
assign LUT_1[49359] = 32'b00000000000000000000001111010101;
assign LUT_1[49360] = 32'b00000000000000000110000011011110;
assign LUT_1[49361] = 32'b11111111111111111111010101011010;
assign LUT_1[49362] = 32'b00000000000000000001110001101111;
assign LUT_1[49363] = 32'b11111111111111111011000011101011;
assign LUT_1[49364] = 32'b00000000000000001101111100110101;
assign LUT_1[49365] = 32'b00000000000000000111001110110001;
assign LUT_1[49366] = 32'b00000000000000001001101011000110;
assign LUT_1[49367] = 32'b00000000000000000010111101000010;
assign LUT_1[49368] = 32'b00000000000000000101010001010011;
assign LUT_1[49369] = 32'b11111111111111111110100011001111;
assign LUT_1[49370] = 32'b00000000000000000000111111100100;
assign LUT_1[49371] = 32'b11111111111111111010010001100000;
assign LUT_1[49372] = 32'b00000000000000001101001010101010;
assign LUT_1[49373] = 32'b00000000000000000110011100100110;
assign LUT_1[49374] = 32'b00000000000000001000111000111011;
assign LUT_1[49375] = 32'b00000000000000000010001010110111;
assign LUT_1[49376] = 32'b00000000000000000101000010111011;
assign LUT_1[49377] = 32'b11111111111111111110010100110111;
assign LUT_1[49378] = 32'b00000000000000000000110001001100;
assign LUT_1[49379] = 32'b11111111111111111010000011001000;
assign LUT_1[49380] = 32'b00000000000000001100111100010010;
assign LUT_1[49381] = 32'b00000000000000000110001110001110;
assign LUT_1[49382] = 32'b00000000000000001000101010100011;
assign LUT_1[49383] = 32'b00000000000000000001111100011111;
assign LUT_1[49384] = 32'b00000000000000000100010000110000;
assign LUT_1[49385] = 32'b11111111111111111101100010101100;
assign LUT_1[49386] = 32'b11111111111111111111111111000001;
assign LUT_1[49387] = 32'b11111111111111111001010000111101;
assign LUT_1[49388] = 32'b00000000000000001100001010000111;
assign LUT_1[49389] = 32'b00000000000000000101011100000011;
assign LUT_1[49390] = 32'b00000000000000000111111000011000;
assign LUT_1[49391] = 32'b00000000000000000001001010010100;
assign LUT_1[49392] = 32'b00000000000000000110111110011101;
assign LUT_1[49393] = 32'b00000000000000000000010000011001;
assign LUT_1[49394] = 32'b00000000000000000010101100101110;
assign LUT_1[49395] = 32'b11111111111111111011111110101010;
assign LUT_1[49396] = 32'b00000000000000001110110111110100;
assign LUT_1[49397] = 32'b00000000000000001000001001110000;
assign LUT_1[49398] = 32'b00000000000000001010100110000101;
assign LUT_1[49399] = 32'b00000000000000000011111000000001;
assign LUT_1[49400] = 32'b00000000000000000110001100010010;
assign LUT_1[49401] = 32'b11111111111111111111011110001110;
assign LUT_1[49402] = 32'b00000000000000000001111010100011;
assign LUT_1[49403] = 32'b11111111111111111011001100011111;
assign LUT_1[49404] = 32'b00000000000000001110000101101001;
assign LUT_1[49405] = 32'b00000000000000000111010111100101;
assign LUT_1[49406] = 32'b00000000000000001001110011111010;
assign LUT_1[49407] = 32'b00000000000000000011000101110110;
assign LUT_1[49408] = 32'b11111111111111111100111110011101;
assign LUT_1[49409] = 32'b11111111111111110110010000011001;
assign LUT_1[49410] = 32'b11111111111111111000101100101110;
assign LUT_1[49411] = 32'b11111111111111110001111110101010;
assign LUT_1[49412] = 32'b00000000000000000100110111110100;
assign LUT_1[49413] = 32'b11111111111111111110001001110000;
assign LUT_1[49414] = 32'b00000000000000000000100110000101;
assign LUT_1[49415] = 32'b11111111111111111001111000000001;
assign LUT_1[49416] = 32'b11111111111111111100001100010010;
assign LUT_1[49417] = 32'b11111111111111110101011110001110;
assign LUT_1[49418] = 32'b11111111111111110111111010100011;
assign LUT_1[49419] = 32'b11111111111111110001001100011111;
assign LUT_1[49420] = 32'b00000000000000000100000101101001;
assign LUT_1[49421] = 32'b11111111111111111101010111100101;
assign LUT_1[49422] = 32'b11111111111111111111110011111010;
assign LUT_1[49423] = 32'b11111111111111111001000101110110;
assign LUT_1[49424] = 32'b11111111111111111110111001111111;
assign LUT_1[49425] = 32'b11111111111111111000001011111011;
assign LUT_1[49426] = 32'b11111111111111111010101000010000;
assign LUT_1[49427] = 32'b11111111111111110011111010001100;
assign LUT_1[49428] = 32'b00000000000000000110110011010110;
assign LUT_1[49429] = 32'b00000000000000000000000101010010;
assign LUT_1[49430] = 32'b00000000000000000010100001100111;
assign LUT_1[49431] = 32'b11111111111111111011110011100011;
assign LUT_1[49432] = 32'b11111111111111111110000111110100;
assign LUT_1[49433] = 32'b11111111111111110111011001110000;
assign LUT_1[49434] = 32'b11111111111111111001110110000101;
assign LUT_1[49435] = 32'b11111111111111110011001000000001;
assign LUT_1[49436] = 32'b00000000000000000110000001001011;
assign LUT_1[49437] = 32'b11111111111111111111010011000111;
assign LUT_1[49438] = 32'b00000000000000000001101111011100;
assign LUT_1[49439] = 32'b11111111111111111011000001011000;
assign LUT_1[49440] = 32'b11111111111111111101111001011100;
assign LUT_1[49441] = 32'b11111111111111110111001011011000;
assign LUT_1[49442] = 32'b11111111111111111001100111101101;
assign LUT_1[49443] = 32'b11111111111111110010111001101001;
assign LUT_1[49444] = 32'b00000000000000000101110010110011;
assign LUT_1[49445] = 32'b11111111111111111111000100101111;
assign LUT_1[49446] = 32'b00000000000000000001100001000100;
assign LUT_1[49447] = 32'b11111111111111111010110011000000;
assign LUT_1[49448] = 32'b11111111111111111101000111010001;
assign LUT_1[49449] = 32'b11111111111111110110011001001101;
assign LUT_1[49450] = 32'b11111111111111111000110101100010;
assign LUT_1[49451] = 32'b11111111111111110010000111011110;
assign LUT_1[49452] = 32'b00000000000000000101000000101000;
assign LUT_1[49453] = 32'b11111111111111111110010010100100;
assign LUT_1[49454] = 32'b00000000000000000000101110111001;
assign LUT_1[49455] = 32'b11111111111111111010000000110101;
assign LUT_1[49456] = 32'b11111111111111111111110100111110;
assign LUT_1[49457] = 32'b11111111111111111001000110111010;
assign LUT_1[49458] = 32'b11111111111111111011100011001111;
assign LUT_1[49459] = 32'b11111111111111110100110101001011;
assign LUT_1[49460] = 32'b00000000000000000111101110010101;
assign LUT_1[49461] = 32'b00000000000000000001000000010001;
assign LUT_1[49462] = 32'b00000000000000000011011100100110;
assign LUT_1[49463] = 32'b11111111111111111100101110100010;
assign LUT_1[49464] = 32'b11111111111111111111000010110011;
assign LUT_1[49465] = 32'b11111111111111111000010100101111;
assign LUT_1[49466] = 32'b11111111111111111010110001000100;
assign LUT_1[49467] = 32'b11111111111111110100000011000000;
assign LUT_1[49468] = 32'b00000000000000000110111100001010;
assign LUT_1[49469] = 32'b00000000000000000000001110000110;
assign LUT_1[49470] = 32'b00000000000000000010101010011011;
assign LUT_1[49471] = 32'b11111111111111111011111100010111;
assign LUT_1[49472] = 32'b11111111111111111110111100000101;
assign LUT_1[49473] = 32'b11111111111111111000001110000001;
assign LUT_1[49474] = 32'b11111111111111111010101010010110;
assign LUT_1[49475] = 32'b11111111111111110011111100010010;
assign LUT_1[49476] = 32'b00000000000000000110110101011100;
assign LUT_1[49477] = 32'b00000000000000000000000111011000;
assign LUT_1[49478] = 32'b00000000000000000010100011101101;
assign LUT_1[49479] = 32'b11111111111111111011110101101001;
assign LUT_1[49480] = 32'b11111111111111111110001001111010;
assign LUT_1[49481] = 32'b11111111111111110111011011110110;
assign LUT_1[49482] = 32'b11111111111111111001111000001011;
assign LUT_1[49483] = 32'b11111111111111110011001010000111;
assign LUT_1[49484] = 32'b00000000000000000110000011010001;
assign LUT_1[49485] = 32'b11111111111111111111010101001101;
assign LUT_1[49486] = 32'b00000000000000000001110001100010;
assign LUT_1[49487] = 32'b11111111111111111011000011011110;
assign LUT_1[49488] = 32'b00000000000000000000110111100111;
assign LUT_1[49489] = 32'b11111111111111111010001001100011;
assign LUT_1[49490] = 32'b11111111111111111100100101111000;
assign LUT_1[49491] = 32'b11111111111111110101110111110100;
assign LUT_1[49492] = 32'b00000000000000001000110000111110;
assign LUT_1[49493] = 32'b00000000000000000010000010111010;
assign LUT_1[49494] = 32'b00000000000000000100011111001111;
assign LUT_1[49495] = 32'b11111111111111111101110001001011;
assign LUT_1[49496] = 32'b00000000000000000000000101011100;
assign LUT_1[49497] = 32'b11111111111111111001010111011000;
assign LUT_1[49498] = 32'b11111111111111111011110011101101;
assign LUT_1[49499] = 32'b11111111111111110101000101101001;
assign LUT_1[49500] = 32'b00000000000000000111111110110011;
assign LUT_1[49501] = 32'b00000000000000000001010000101111;
assign LUT_1[49502] = 32'b00000000000000000011101101000100;
assign LUT_1[49503] = 32'b11111111111111111100111111000000;
assign LUT_1[49504] = 32'b11111111111111111111110111000100;
assign LUT_1[49505] = 32'b11111111111111111001001001000000;
assign LUT_1[49506] = 32'b11111111111111111011100101010101;
assign LUT_1[49507] = 32'b11111111111111110100110111010001;
assign LUT_1[49508] = 32'b00000000000000000111110000011011;
assign LUT_1[49509] = 32'b00000000000000000001000010010111;
assign LUT_1[49510] = 32'b00000000000000000011011110101100;
assign LUT_1[49511] = 32'b11111111111111111100110000101000;
assign LUT_1[49512] = 32'b11111111111111111111000100111001;
assign LUT_1[49513] = 32'b11111111111111111000010110110101;
assign LUT_1[49514] = 32'b11111111111111111010110011001010;
assign LUT_1[49515] = 32'b11111111111111110100000101000110;
assign LUT_1[49516] = 32'b00000000000000000110111110010000;
assign LUT_1[49517] = 32'b00000000000000000000010000001100;
assign LUT_1[49518] = 32'b00000000000000000010101100100001;
assign LUT_1[49519] = 32'b11111111111111111011111110011101;
assign LUT_1[49520] = 32'b00000000000000000001110010100110;
assign LUT_1[49521] = 32'b11111111111111111011000100100010;
assign LUT_1[49522] = 32'b11111111111111111101100000110111;
assign LUT_1[49523] = 32'b11111111111111110110110010110011;
assign LUT_1[49524] = 32'b00000000000000001001101011111101;
assign LUT_1[49525] = 32'b00000000000000000010111101111001;
assign LUT_1[49526] = 32'b00000000000000000101011010001110;
assign LUT_1[49527] = 32'b11111111111111111110101100001010;
assign LUT_1[49528] = 32'b00000000000000000001000000011011;
assign LUT_1[49529] = 32'b11111111111111111010010010010111;
assign LUT_1[49530] = 32'b11111111111111111100101110101100;
assign LUT_1[49531] = 32'b11111111111111110110000000101000;
assign LUT_1[49532] = 32'b00000000000000001000111001110010;
assign LUT_1[49533] = 32'b00000000000000000010001011101110;
assign LUT_1[49534] = 32'b00000000000000000100101000000011;
assign LUT_1[49535] = 32'b11111111111111111101111001111111;
assign LUT_1[49536] = 32'b11111111111111111111111110100000;
assign LUT_1[49537] = 32'b11111111111111111001010000011100;
assign LUT_1[49538] = 32'b11111111111111111011101100110001;
assign LUT_1[49539] = 32'b11111111111111110100111110101101;
assign LUT_1[49540] = 32'b00000000000000000111110111110111;
assign LUT_1[49541] = 32'b00000000000000000001001001110011;
assign LUT_1[49542] = 32'b00000000000000000011100110001000;
assign LUT_1[49543] = 32'b11111111111111111100111000000100;
assign LUT_1[49544] = 32'b11111111111111111111001100010101;
assign LUT_1[49545] = 32'b11111111111111111000011110010001;
assign LUT_1[49546] = 32'b11111111111111111010111010100110;
assign LUT_1[49547] = 32'b11111111111111110100001100100010;
assign LUT_1[49548] = 32'b00000000000000000111000101101100;
assign LUT_1[49549] = 32'b00000000000000000000010111101000;
assign LUT_1[49550] = 32'b00000000000000000010110011111101;
assign LUT_1[49551] = 32'b11111111111111111100000101111001;
assign LUT_1[49552] = 32'b00000000000000000001111010000010;
assign LUT_1[49553] = 32'b11111111111111111011001011111110;
assign LUT_1[49554] = 32'b11111111111111111101101000010011;
assign LUT_1[49555] = 32'b11111111111111110110111010001111;
assign LUT_1[49556] = 32'b00000000000000001001110011011001;
assign LUT_1[49557] = 32'b00000000000000000011000101010101;
assign LUT_1[49558] = 32'b00000000000000000101100001101010;
assign LUT_1[49559] = 32'b11111111111111111110110011100110;
assign LUT_1[49560] = 32'b00000000000000000001000111110111;
assign LUT_1[49561] = 32'b11111111111111111010011001110011;
assign LUT_1[49562] = 32'b11111111111111111100110110001000;
assign LUT_1[49563] = 32'b11111111111111110110001000000100;
assign LUT_1[49564] = 32'b00000000000000001001000001001110;
assign LUT_1[49565] = 32'b00000000000000000010010011001010;
assign LUT_1[49566] = 32'b00000000000000000100101111011111;
assign LUT_1[49567] = 32'b11111111111111111110000001011011;
assign LUT_1[49568] = 32'b00000000000000000000111001011111;
assign LUT_1[49569] = 32'b11111111111111111010001011011011;
assign LUT_1[49570] = 32'b11111111111111111100100111110000;
assign LUT_1[49571] = 32'b11111111111111110101111001101100;
assign LUT_1[49572] = 32'b00000000000000001000110010110110;
assign LUT_1[49573] = 32'b00000000000000000010000100110010;
assign LUT_1[49574] = 32'b00000000000000000100100001000111;
assign LUT_1[49575] = 32'b11111111111111111101110011000011;
assign LUT_1[49576] = 32'b00000000000000000000000111010100;
assign LUT_1[49577] = 32'b11111111111111111001011001010000;
assign LUT_1[49578] = 32'b11111111111111111011110101100101;
assign LUT_1[49579] = 32'b11111111111111110101000111100001;
assign LUT_1[49580] = 32'b00000000000000001000000000101011;
assign LUT_1[49581] = 32'b00000000000000000001010010100111;
assign LUT_1[49582] = 32'b00000000000000000011101110111100;
assign LUT_1[49583] = 32'b11111111111111111101000000111000;
assign LUT_1[49584] = 32'b00000000000000000010110101000001;
assign LUT_1[49585] = 32'b11111111111111111100000110111101;
assign LUT_1[49586] = 32'b11111111111111111110100011010010;
assign LUT_1[49587] = 32'b11111111111111110111110101001110;
assign LUT_1[49588] = 32'b00000000000000001010101110011000;
assign LUT_1[49589] = 32'b00000000000000000100000000010100;
assign LUT_1[49590] = 32'b00000000000000000110011100101001;
assign LUT_1[49591] = 32'b11111111111111111111101110100101;
assign LUT_1[49592] = 32'b00000000000000000010000010110110;
assign LUT_1[49593] = 32'b11111111111111111011010100110010;
assign LUT_1[49594] = 32'b11111111111111111101110001000111;
assign LUT_1[49595] = 32'b11111111111111110111000011000011;
assign LUT_1[49596] = 32'b00000000000000001001111100001101;
assign LUT_1[49597] = 32'b00000000000000000011001110001001;
assign LUT_1[49598] = 32'b00000000000000000101101010011110;
assign LUT_1[49599] = 32'b11111111111111111110111100011010;
assign LUT_1[49600] = 32'b00000000000000000001111100001000;
assign LUT_1[49601] = 32'b11111111111111111011001110000100;
assign LUT_1[49602] = 32'b11111111111111111101101010011001;
assign LUT_1[49603] = 32'b11111111111111110110111100010101;
assign LUT_1[49604] = 32'b00000000000000001001110101011111;
assign LUT_1[49605] = 32'b00000000000000000011000111011011;
assign LUT_1[49606] = 32'b00000000000000000101100011110000;
assign LUT_1[49607] = 32'b11111111111111111110110101101100;
assign LUT_1[49608] = 32'b00000000000000000001001001111101;
assign LUT_1[49609] = 32'b11111111111111111010011011111001;
assign LUT_1[49610] = 32'b11111111111111111100111000001110;
assign LUT_1[49611] = 32'b11111111111111110110001010001010;
assign LUT_1[49612] = 32'b00000000000000001001000011010100;
assign LUT_1[49613] = 32'b00000000000000000010010101010000;
assign LUT_1[49614] = 32'b00000000000000000100110001100101;
assign LUT_1[49615] = 32'b11111111111111111110000011100001;
assign LUT_1[49616] = 32'b00000000000000000011110111101010;
assign LUT_1[49617] = 32'b11111111111111111101001001100110;
assign LUT_1[49618] = 32'b11111111111111111111100101111011;
assign LUT_1[49619] = 32'b11111111111111111000110111110111;
assign LUT_1[49620] = 32'b00000000000000001011110001000001;
assign LUT_1[49621] = 32'b00000000000000000101000010111101;
assign LUT_1[49622] = 32'b00000000000000000111011111010010;
assign LUT_1[49623] = 32'b00000000000000000000110001001110;
assign LUT_1[49624] = 32'b00000000000000000011000101011111;
assign LUT_1[49625] = 32'b11111111111111111100010111011011;
assign LUT_1[49626] = 32'b11111111111111111110110011110000;
assign LUT_1[49627] = 32'b11111111111111111000000101101100;
assign LUT_1[49628] = 32'b00000000000000001010111110110110;
assign LUT_1[49629] = 32'b00000000000000000100010000110010;
assign LUT_1[49630] = 32'b00000000000000000110101101000111;
assign LUT_1[49631] = 32'b11111111111111111111111111000011;
assign LUT_1[49632] = 32'b00000000000000000010110111000111;
assign LUT_1[49633] = 32'b11111111111111111100001001000011;
assign LUT_1[49634] = 32'b11111111111111111110100101011000;
assign LUT_1[49635] = 32'b11111111111111110111110111010100;
assign LUT_1[49636] = 32'b00000000000000001010110000011110;
assign LUT_1[49637] = 32'b00000000000000000100000010011010;
assign LUT_1[49638] = 32'b00000000000000000110011110101111;
assign LUT_1[49639] = 32'b11111111111111111111110000101011;
assign LUT_1[49640] = 32'b00000000000000000010000100111100;
assign LUT_1[49641] = 32'b11111111111111111011010110111000;
assign LUT_1[49642] = 32'b11111111111111111101110011001101;
assign LUT_1[49643] = 32'b11111111111111110111000101001001;
assign LUT_1[49644] = 32'b00000000000000001001111110010011;
assign LUT_1[49645] = 32'b00000000000000000011010000001111;
assign LUT_1[49646] = 32'b00000000000000000101101100100100;
assign LUT_1[49647] = 32'b11111111111111111110111110100000;
assign LUT_1[49648] = 32'b00000000000000000100110010101001;
assign LUT_1[49649] = 32'b11111111111111111110000100100101;
assign LUT_1[49650] = 32'b00000000000000000000100000111010;
assign LUT_1[49651] = 32'b11111111111111111001110010110110;
assign LUT_1[49652] = 32'b00000000000000001100101100000000;
assign LUT_1[49653] = 32'b00000000000000000101111101111100;
assign LUT_1[49654] = 32'b00000000000000001000011010010001;
assign LUT_1[49655] = 32'b00000000000000000001101100001101;
assign LUT_1[49656] = 32'b00000000000000000100000000011110;
assign LUT_1[49657] = 32'b11111111111111111101010010011010;
assign LUT_1[49658] = 32'b11111111111111111111101110101111;
assign LUT_1[49659] = 32'b11111111111111111001000000101011;
assign LUT_1[49660] = 32'b00000000000000001011111001110101;
assign LUT_1[49661] = 32'b00000000000000000101001011110001;
assign LUT_1[49662] = 32'b00000000000000000111101000000110;
assign LUT_1[49663] = 32'b00000000000000000000111010000010;
assign LUT_1[49664] = 32'b11111111111111111000111000101110;
assign LUT_1[49665] = 32'b11111111111111110010001010101010;
assign LUT_1[49666] = 32'b11111111111111110100100110111111;
assign LUT_1[49667] = 32'b11111111111111101101111000111011;
assign LUT_1[49668] = 32'b00000000000000000000110010000101;
assign LUT_1[49669] = 32'b11111111111111111010000100000001;
assign LUT_1[49670] = 32'b11111111111111111100100000010110;
assign LUT_1[49671] = 32'b11111111111111110101110010010010;
assign LUT_1[49672] = 32'b11111111111111111000000110100011;
assign LUT_1[49673] = 32'b11111111111111110001011000011111;
assign LUT_1[49674] = 32'b11111111111111110011110100110100;
assign LUT_1[49675] = 32'b11111111111111101101000110110000;
assign LUT_1[49676] = 32'b11111111111111111111111111111010;
assign LUT_1[49677] = 32'b11111111111111111001010001110110;
assign LUT_1[49678] = 32'b11111111111111111011101110001011;
assign LUT_1[49679] = 32'b11111111111111110101000000000111;
assign LUT_1[49680] = 32'b11111111111111111010110100010000;
assign LUT_1[49681] = 32'b11111111111111110100000110001100;
assign LUT_1[49682] = 32'b11111111111111110110100010100001;
assign LUT_1[49683] = 32'b11111111111111101111110100011101;
assign LUT_1[49684] = 32'b00000000000000000010101101100111;
assign LUT_1[49685] = 32'b11111111111111111011111111100011;
assign LUT_1[49686] = 32'b11111111111111111110011011111000;
assign LUT_1[49687] = 32'b11111111111111110111101101110100;
assign LUT_1[49688] = 32'b11111111111111111010000010000101;
assign LUT_1[49689] = 32'b11111111111111110011010100000001;
assign LUT_1[49690] = 32'b11111111111111110101110000010110;
assign LUT_1[49691] = 32'b11111111111111101111000010010010;
assign LUT_1[49692] = 32'b00000000000000000001111011011100;
assign LUT_1[49693] = 32'b11111111111111111011001101011000;
assign LUT_1[49694] = 32'b11111111111111111101101001101101;
assign LUT_1[49695] = 32'b11111111111111110110111011101001;
assign LUT_1[49696] = 32'b11111111111111111001110011101101;
assign LUT_1[49697] = 32'b11111111111111110011000101101001;
assign LUT_1[49698] = 32'b11111111111111110101100001111110;
assign LUT_1[49699] = 32'b11111111111111101110110011111010;
assign LUT_1[49700] = 32'b00000000000000000001101101000100;
assign LUT_1[49701] = 32'b11111111111111111010111111000000;
assign LUT_1[49702] = 32'b11111111111111111101011011010101;
assign LUT_1[49703] = 32'b11111111111111110110101101010001;
assign LUT_1[49704] = 32'b11111111111111111001000001100010;
assign LUT_1[49705] = 32'b11111111111111110010010011011110;
assign LUT_1[49706] = 32'b11111111111111110100101111110011;
assign LUT_1[49707] = 32'b11111111111111101110000001101111;
assign LUT_1[49708] = 32'b00000000000000000000111010111001;
assign LUT_1[49709] = 32'b11111111111111111010001100110101;
assign LUT_1[49710] = 32'b11111111111111111100101001001010;
assign LUT_1[49711] = 32'b11111111111111110101111011000110;
assign LUT_1[49712] = 32'b11111111111111111011101111001111;
assign LUT_1[49713] = 32'b11111111111111110101000001001011;
assign LUT_1[49714] = 32'b11111111111111110111011101100000;
assign LUT_1[49715] = 32'b11111111111111110000101111011100;
assign LUT_1[49716] = 32'b00000000000000000011101000100110;
assign LUT_1[49717] = 32'b11111111111111111100111010100010;
assign LUT_1[49718] = 32'b11111111111111111111010110110111;
assign LUT_1[49719] = 32'b11111111111111111000101000110011;
assign LUT_1[49720] = 32'b11111111111111111010111101000100;
assign LUT_1[49721] = 32'b11111111111111110100001111000000;
assign LUT_1[49722] = 32'b11111111111111110110101011010101;
assign LUT_1[49723] = 32'b11111111111111101111111101010001;
assign LUT_1[49724] = 32'b00000000000000000010110110011011;
assign LUT_1[49725] = 32'b11111111111111111100001000010111;
assign LUT_1[49726] = 32'b11111111111111111110100100101100;
assign LUT_1[49727] = 32'b11111111111111110111110110101000;
assign LUT_1[49728] = 32'b11111111111111111010110110010110;
assign LUT_1[49729] = 32'b11111111111111110100001000010010;
assign LUT_1[49730] = 32'b11111111111111110110100100100111;
assign LUT_1[49731] = 32'b11111111111111101111110110100011;
assign LUT_1[49732] = 32'b00000000000000000010101111101101;
assign LUT_1[49733] = 32'b11111111111111111100000001101001;
assign LUT_1[49734] = 32'b11111111111111111110011101111110;
assign LUT_1[49735] = 32'b11111111111111110111101111111010;
assign LUT_1[49736] = 32'b11111111111111111010000100001011;
assign LUT_1[49737] = 32'b11111111111111110011010110000111;
assign LUT_1[49738] = 32'b11111111111111110101110010011100;
assign LUT_1[49739] = 32'b11111111111111101111000100011000;
assign LUT_1[49740] = 32'b00000000000000000001111101100010;
assign LUT_1[49741] = 32'b11111111111111111011001111011110;
assign LUT_1[49742] = 32'b11111111111111111101101011110011;
assign LUT_1[49743] = 32'b11111111111111110110111101101111;
assign LUT_1[49744] = 32'b11111111111111111100110001111000;
assign LUT_1[49745] = 32'b11111111111111110110000011110100;
assign LUT_1[49746] = 32'b11111111111111111000100000001001;
assign LUT_1[49747] = 32'b11111111111111110001110010000101;
assign LUT_1[49748] = 32'b00000000000000000100101011001111;
assign LUT_1[49749] = 32'b11111111111111111101111101001011;
assign LUT_1[49750] = 32'b00000000000000000000011001100000;
assign LUT_1[49751] = 32'b11111111111111111001101011011100;
assign LUT_1[49752] = 32'b11111111111111111011111111101101;
assign LUT_1[49753] = 32'b11111111111111110101010001101001;
assign LUT_1[49754] = 32'b11111111111111110111101101111110;
assign LUT_1[49755] = 32'b11111111111111110000111111111010;
assign LUT_1[49756] = 32'b00000000000000000011111001000100;
assign LUT_1[49757] = 32'b11111111111111111101001011000000;
assign LUT_1[49758] = 32'b11111111111111111111100111010101;
assign LUT_1[49759] = 32'b11111111111111111000111001010001;
assign LUT_1[49760] = 32'b11111111111111111011110001010101;
assign LUT_1[49761] = 32'b11111111111111110101000011010001;
assign LUT_1[49762] = 32'b11111111111111110111011111100110;
assign LUT_1[49763] = 32'b11111111111111110000110001100010;
assign LUT_1[49764] = 32'b00000000000000000011101010101100;
assign LUT_1[49765] = 32'b11111111111111111100111100101000;
assign LUT_1[49766] = 32'b11111111111111111111011000111101;
assign LUT_1[49767] = 32'b11111111111111111000101010111001;
assign LUT_1[49768] = 32'b11111111111111111010111111001010;
assign LUT_1[49769] = 32'b11111111111111110100010001000110;
assign LUT_1[49770] = 32'b11111111111111110110101101011011;
assign LUT_1[49771] = 32'b11111111111111101111111111010111;
assign LUT_1[49772] = 32'b00000000000000000010111000100001;
assign LUT_1[49773] = 32'b11111111111111111100001010011101;
assign LUT_1[49774] = 32'b11111111111111111110100110110010;
assign LUT_1[49775] = 32'b11111111111111110111111000101110;
assign LUT_1[49776] = 32'b11111111111111111101101100110111;
assign LUT_1[49777] = 32'b11111111111111110110111110110011;
assign LUT_1[49778] = 32'b11111111111111111001011011001000;
assign LUT_1[49779] = 32'b11111111111111110010101101000100;
assign LUT_1[49780] = 32'b00000000000000000101100110001110;
assign LUT_1[49781] = 32'b11111111111111111110111000001010;
assign LUT_1[49782] = 32'b00000000000000000001010100011111;
assign LUT_1[49783] = 32'b11111111111111111010100110011011;
assign LUT_1[49784] = 32'b11111111111111111100111010101100;
assign LUT_1[49785] = 32'b11111111111111110110001100101000;
assign LUT_1[49786] = 32'b11111111111111111000101000111101;
assign LUT_1[49787] = 32'b11111111111111110001111010111001;
assign LUT_1[49788] = 32'b00000000000000000100110100000011;
assign LUT_1[49789] = 32'b11111111111111111110000101111111;
assign LUT_1[49790] = 32'b00000000000000000000100010010100;
assign LUT_1[49791] = 32'b11111111111111111001110100010000;
assign LUT_1[49792] = 32'b11111111111111111011111000110001;
assign LUT_1[49793] = 32'b11111111111111110101001010101101;
assign LUT_1[49794] = 32'b11111111111111110111100111000010;
assign LUT_1[49795] = 32'b11111111111111110000111000111110;
assign LUT_1[49796] = 32'b00000000000000000011110010001000;
assign LUT_1[49797] = 32'b11111111111111111101000100000100;
assign LUT_1[49798] = 32'b11111111111111111111100000011001;
assign LUT_1[49799] = 32'b11111111111111111000110010010101;
assign LUT_1[49800] = 32'b11111111111111111011000110100110;
assign LUT_1[49801] = 32'b11111111111111110100011000100010;
assign LUT_1[49802] = 32'b11111111111111110110110100110111;
assign LUT_1[49803] = 32'b11111111111111110000000110110011;
assign LUT_1[49804] = 32'b00000000000000000010111111111101;
assign LUT_1[49805] = 32'b11111111111111111100010001111001;
assign LUT_1[49806] = 32'b11111111111111111110101110001110;
assign LUT_1[49807] = 32'b11111111111111111000000000001010;
assign LUT_1[49808] = 32'b11111111111111111101110100010011;
assign LUT_1[49809] = 32'b11111111111111110111000110001111;
assign LUT_1[49810] = 32'b11111111111111111001100010100100;
assign LUT_1[49811] = 32'b11111111111111110010110100100000;
assign LUT_1[49812] = 32'b00000000000000000101101101101010;
assign LUT_1[49813] = 32'b11111111111111111110111111100110;
assign LUT_1[49814] = 32'b00000000000000000001011011111011;
assign LUT_1[49815] = 32'b11111111111111111010101101110111;
assign LUT_1[49816] = 32'b11111111111111111101000010001000;
assign LUT_1[49817] = 32'b11111111111111110110010100000100;
assign LUT_1[49818] = 32'b11111111111111111000110000011001;
assign LUT_1[49819] = 32'b11111111111111110010000010010101;
assign LUT_1[49820] = 32'b00000000000000000100111011011111;
assign LUT_1[49821] = 32'b11111111111111111110001101011011;
assign LUT_1[49822] = 32'b00000000000000000000101001110000;
assign LUT_1[49823] = 32'b11111111111111111001111011101100;
assign LUT_1[49824] = 32'b11111111111111111100110011110000;
assign LUT_1[49825] = 32'b11111111111111110110000101101100;
assign LUT_1[49826] = 32'b11111111111111111000100010000001;
assign LUT_1[49827] = 32'b11111111111111110001110011111101;
assign LUT_1[49828] = 32'b00000000000000000100101101000111;
assign LUT_1[49829] = 32'b11111111111111111101111111000011;
assign LUT_1[49830] = 32'b00000000000000000000011011011000;
assign LUT_1[49831] = 32'b11111111111111111001101101010100;
assign LUT_1[49832] = 32'b11111111111111111100000001100101;
assign LUT_1[49833] = 32'b11111111111111110101010011100001;
assign LUT_1[49834] = 32'b11111111111111110111101111110110;
assign LUT_1[49835] = 32'b11111111111111110001000001110010;
assign LUT_1[49836] = 32'b00000000000000000011111010111100;
assign LUT_1[49837] = 32'b11111111111111111101001100111000;
assign LUT_1[49838] = 32'b11111111111111111111101001001101;
assign LUT_1[49839] = 32'b11111111111111111000111011001001;
assign LUT_1[49840] = 32'b11111111111111111110101111010010;
assign LUT_1[49841] = 32'b11111111111111111000000001001110;
assign LUT_1[49842] = 32'b11111111111111111010011101100011;
assign LUT_1[49843] = 32'b11111111111111110011101111011111;
assign LUT_1[49844] = 32'b00000000000000000110101000101001;
assign LUT_1[49845] = 32'b11111111111111111111111010100101;
assign LUT_1[49846] = 32'b00000000000000000010010110111010;
assign LUT_1[49847] = 32'b11111111111111111011101000110110;
assign LUT_1[49848] = 32'b11111111111111111101111101000111;
assign LUT_1[49849] = 32'b11111111111111110111001111000011;
assign LUT_1[49850] = 32'b11111111111111111001101011011000;
assign LUT_1[49851] = 32'b11111111111111110010111101010100;
assign LUT_1[49852] = 32'b00000000000000000101110110011110;
assign LUT_1[49853] = 32'b11111111111111111111001000011010;
assign LUT_1[49854] = 32'b00000000000000000001100100101111;
assign LUT_1[49855] = 32'b11111111111111111010110110101011;
assign LUT_1[49856] = 32'b11111111111111111101110110011001;
assign LUT_1[49857] = 32'b11111111111111110111001000010101;
assign LUT_1[49858] = 32'b11111111111111111001100100101010;
assign LUT_1[49859] = 32'b11111111111111110010110110100110;
assign LUT_1[49860] = 32'b00000000000000000101101111110000;
assign LUT_1[49861] = 32'b11111111111111111111000001101100;
assign LUT_1[49862] = 32'b00000000000000000001011110000001;
assign LUT_1[49863] = 32'b11111111111111111010101111111101;
assign LUT_1[49864] = 32'b11111111111111111101000100001110;
assign LUT_1[49865] = 32'b11111111111111110110010110001010;
assign LUT_1[49866] = 32'b11111111111111111000110010011111;
assign LUT_1[49867] = 32'b11111111111111110010000100011011;
assign LUT_1[49868] = 32'b00000000000000000100111101100101;
assign LUT_1[49869] = 32'b11111111111111111110001111100001;
assign LUT_1[49870] = 32'b00000000000000000000101011110110;
assign LUT_1[49871] = 32'b11111111111111111001111101110010;
assign LUT_1[49872] = 32'b11111111111111111111110001111011;
assign LUT_1[49873] = 32'b11111111111111111001000011110111;
assign LUT_1[49874] = 32'b11111111111111111011100000001100;
assign LUT_1[49875] = 32'b11111111111111110100110010001000;
assign LUT_1[49876] = 32'b00000000000000000111101011010010;
assign LUT_1[49877] = 32'b00000000000000000000111101001110;
assign LUT_1[49878] = 32'b00000000000000000011011001100011;
assign LUT_1[49879] = 32'b11111111111111111100101011011111;
assign LUT_1[49880] = 32'b11111111111111111110111111110000;
assign LUT_1[49881] = 32'b11111111111111111000010001101100;
assign LUT_1[49882] = 32'b11111111111111111010101110000001;
assign LUT_1[49883] = 32'b11111111111111110011111111111101;
assign LUT_1[49884] = 32'b00000000000000000110111001000111;
assign LUT_1[49885] = 32'b00000000000000000000001011000011;
assign LUT_1[49886] = 32'b00000000000000000010100111011000;
assign LUT_1[49887] = 32'b11111111111111111011111001010100;
assign LUT_1[49888] = 32'b11111111111111111110110001011000;
assign LUT_1[49889] = 32'b11111111111111111000000011010100;
assign LUT_1[49890] = 32'b11111111111111111010011111101001;
assign LUT_1[49891] = 32'b11111111111111110011110001100101;
assign LUT_1[49892] = 32'b00000000000000000110101010101111;
assign LUT_1[49893] = 32'b11111111111111111111111100101011;
assign LUT_1[49894] = 32'b00000000000000000010011001000000;
assign LUT_1[49895] = 32'b11111111111111111011101010111100;
assign LUT_1[49896] = 32'b11111111111111111101111111001101;
assign LUT_1[49897] = 32'b11111111111111110111010001001001;
assign LUT_1[49898] = 32'b11111111111111111001101101011110;
assign LUT_1[49899] = 32'b11111111111111110010111111011010;
assign LUT_1[49900] = 32'b00000000000000000101111000100100;
assign LUT_1[49901] = 32'b11111111111111111111001010100000;
assign LUT_1[49902] = 32'b00000000000000000001100110110101;
assign LUT_1[49903] = 32'b11111111111111111010111000110001;
assign LUT_1[49904] = 32'b00000000000000000000101100111010;
assign LUT_1[49905] = 32'b11111111111111111001111110110110;
assign LUT_1[49906] = 32'b11111111111111111100011011001011;
assign LUT_1[49907] = 32'b11111111111111110101101101000111;
assign LUT_1[49908] = 32'b00000000000000001000100110010001;
assign LUT_1[49909] = 32'b00000000000000000001111000001101;
assign LUT_1[49910] = 32'b00000000000000000100010100100010;
assign LUT_1[49911] = 32'b11111111111111111101100110011110;
assign LUT_1[49912] = 32'b11111111111111111111111010101111;
assign LUT_1[49913] = 32'b11111111111111111001001100101011;
assign LUT_1[49914] = 32'b11111111111111111011101001000000;
assign LUT_1[49915] = 32'b11111111111111110100111010111100;
assign LUT_1[49916] = 32'b00000000000000000111110100000110;
assign LUT_1[49917] = 32'b00000000000000000001000110000010;
assign LUT_1[49918] = 32'b00000000000000000011100010010111;
assign LUT_1[49919] = 32'b11111111111111111100110100010011;
assign LUT_1[49920] = 32'b11111111111111110110101100111010;
assign LUT_1[49921] = 32'b11111111111111101111111110110110;
assign LUT_1[49922] = 32'b11111111111111110010011011001011;
assign LUT_1[49923] = 32'b11111111111111101011101101000111;
assign LUT_1[49924] = 32'b11111111111111111110100110010001;
assign LUT_1[49925] = 32'b11111111111111110111111000001101;
assign LUT_1[49926] = 32'b11111111111111111010010100100010;
assign LUT_1[49927] = 32'b11111111111111110011100110011110;
assign LUT_1[49928] = 32'b11111111111111110101111010101111;
assign LUT_1[49929] = 32'b11111111111111101111001100101011;
assign LUT_1[49930] = 32'b11111111111111110001101001000000;
assign LUT_1[49931] = 32'b11111111111111101010111010111100;
assign LUT_1[49932] = 32'b11111111111111111101110100000110;
assign LUT_1[49933] = 32'b11111111111111110111000110000010;
assign LUT_1[49934] = 32'b11111111111111111001100010010111;
assign LUT_1[49935] = 32'b11111111111111110010110100010011;
assign LUT_1[49936] = 32'b11111111111111111000101000011100;
assign LUT_1[49937] = 32'b11111111111111110001111010011000;
assign LUT_1[49938] = 32'b11111111111111110100010110101101;
assign LUT_1[49939] = 32'b11111111111111101101101000101001;
assign LUT_1[49940] = 32'b00000000000000000000100001110011;
assign LUT_1[49941] = 32'b11111111111111111001110011101111;
assign LUT_1[49942] = 32'b11111111111111111100010000000100;
assign LUT_1[49943] = 32'b11111111111111110101100010000000;
assign LUT_1[49944] = 32'b11111111111111110111110110010001;
assign LUT_1[49945] = 32'b11111111111111110001001000001101;
assign LUT_1[49946] = 32'b11111111111111110011100100100010;
assign LUT_1[49947] = 32'b11111111111111101100110110011110;
assign LUT_1[49948] = 32'b11111111111111111111101111101000;
assign LUT_1[49949] = 32'b11111111111111111001000001100100;
assign LUT_1[49950] = 32'b11111111111111111011011101111001;
assign LUT_1[49951] = 32'b11111111111111110100101111110101;
assign LUT_1[49952] = 32'b11111111111111110111100111111001;
assign LUT_1[49953] = 32'b11111111111111110000111001110101;
assign LUT_1[49954] = 32'b11111111111111110011010110001010;
assign LUT_1[49955] = 32'b11111111111111101100101000000110;
assign LUT_1[49956] = 32'b11111111111111111111100001010000;
assign LUT_1[49957] = 32'b11111111111111111000110011001100;
assign LUT_1[49958] = 32'b11111111111111111011001111100001;
assign LUT_1[49959] = 32'b11111111111111110100100001011101;
assign LUT_1[49960] = 32'b11111111111111110110110101101110;
assign LUT_1[49961] = 32'b11111111111111110000000111101010;
assign LUT_1[49962] = 32'b11111111111111110010100011111111;
assign LUT_1[49963] = 32'b11111111111111101011110101111011;
assign LUT_1[49964] = 32'b11111111111111111110101111000101;
assign LUT_1[49965] = 32'b11111111111111111000000001000001;
assign LUT_1[49966] = 32'b11111111111111111010011101010110;
assign LUT_1[49967] = 32'b11111111111111110011101111010010;
assign LUT_1[49968] = 32'b11111111111111111001100011011011;
assign LUT_1[49969] = 32'b11111111111111110010110101010111;
assign LUT_1[49970] = 32'b11111111111111110101010001101100;
assign LUT_1[49971] = 32'b11111111111111101110100011101000;
assign LUT_1[49972] = 32'b00000000000000000001011100110010;
assign LUT_1[49973] = 32'b11111111111111111010101110101110;
assign LUT_1[49974] = 32'b11111111111111111101001011000011;
assign LUT_1[49975] = 32'b11111111111111110110011100111111;
assign LUT_1[49976] = 32'b11111111111111111000110001010000;
assign LUT_1[49977] = 32'b11111111111111110010000011001100;
assign LUT_1[49978] = 32'b11111111111111110100011111100001;
assign LUT_1[49979] = 32'b11111111111111101101110001011101;
assign LUT_1[49980] = 32'b00000000000000000000101010100111;
assign LUT_1[49981] = 32'b11111111111111111001111100100011;
assign LUT_1[49982] = 32'b11111111111111111100011000111000;
assign LUT_1[49983] = 32'b11111111111111110101101010110100;
assign LUT_1[49984] = 32'b11111111111111111000101010100010;
assign LUT_1[49985] = 32'b11111111111111110001111100011110;
assign LUT_1[49986] = 32'b11111111111111110100011000110011;
assign LUT_1[49987] = 32'b11111111111111101101101010101111;
assign LUT_1[49988] = 32'b00000000000000000000100011111001;
assign LUT_1[49989] = 32'b11111111111111111001110101110101;
assign LUT_1[49990] = 32'b11111111111111111100010010001010;
assign LUT_1[49991] = 32'b11111111111111110101100100000110;
assign LUT_1[49992] = 32'b11111111111111110111111000010111;
assign LUT_1[49993] = 32'b11111111111111110001001010010011;
assign LUT_1[49994] = 32'b11111111111111110011100110101000;
assign LUT_1[49995] = 32'b11111111111111101100111000100100;
assign LUT_1[49996] = 32'b11111111111111111111110001101110;
assign LUT_1[49997] = 32'b11111111111111111001000011101010;
assign LUT_1[49998] = 32'b11111111111111111011011111111111;
assign LUT_1[49999] = 32'b11111111111111110100110001111011;
assign LUT_1[50000] = 32'b11111111111111111010100110000100;
assign LUT_1[50001] = 32'b11111111111111110011111000000000;
assign LUT_1[50002] = 32'b11111111111111110110010100010101;
assign LUT_1[50003] = 32'b11111111111111101111100110010001;
assign LUT_1[50004] = 32'b00000000000000000010011111011011;
assign LUT_1[50005] = 32'b11111111111111111011110001010111;
assign LUT_1[50006] = 32'b11111111111111111110001101101100;
assign LUT_1[50007] = 32'b11111111111111110111011111101000;
assign LUT_1[50008] = 32'b11111111111111111001110011111001;
assign LUT_1[50009] = 32'b11111111111111110011000101110101;
assign LUT_1[50010] = 32'b11111111111111110101100010001010;
assign LUT_1[50011] = 32'b11111111111111101110110100000110;
assign LUT_1[50012] = 32'b00000000000000000001101101010000;
assign LUT_1[50013] = 32'b11111111111111111010111111001100;
assign LUT_1[50014] = 32'b11111111111111111101011011100001;
assign LUT_1[50015] = 32'b11111111111111110110101101011101;
assign LUT_1[50016] = 32'b11111111111111111001100101100001;
assign LUT_1[50017] = 32'b11111111111111110010110111011101;
assign LUT_1[50018] = 32'b11111111111111110101010011110010;
assign LUT_1[50019] = 32'b11111111111111101110100101101110;
assign LUT_1[50020] = 32'b00000000000000000001011110111000;
assign LUT_1[50021] = 32'b11111111111111111010110000110100;
assign LUT_1[50022] = 32'b11111111111111111101001101001001;
assign LUT_1[50023] = 32'b11111111111111110110011111000101;
assign LUT_1[50024] = 32'b11111111111111111000110011010110;
assign LUT_1[50025] = 32'b11111111111111110010000101010010;
assign LUT_1[50026] = 32'b11111111111111110100100001100111;
assign LUT_1[50027] = 32'b11111111111111101101110011100011;
assign LUT_1[50028] = 32'b00000000000000000000101100101101;
assign LUT_1[50029] = 32'b11111111111111111001111110101001;
assign LUT_1[50030] = 32'b11111111111111111100011010111110;
assign LUT_1[50031] = 32'b11111111111111110101101100111010;
assign LUT_1[50032] = 32'b11111111111111111011100001000011;
assign LUT_1[50033] = 32'b11111111111111110100110010111111;
assign LUT_1[50034] = 32'b11111111111111110111001111010100;
assign LUT_1[50035] = 32'b11111111111111110000100001010000;
assign LUT_1[50036] = 32'b00000000000000000011011010011010;
assign LUT_1[50037] = 32'b11111111111111111100101100010110;
assign LUT_1[50038] = 32'b11111111111111111111001000101011;
assign LUT_1[50039] = 32'b11111111111111111000011010100111;
assign LUT_1[50040] = 32'b11111111111111111010101110111000;
assign LUT_1[50041] = 32'b11111111111111110100000000110100;
assign LUT_1[50042] = 32'b11111111111111110110011101001001;
assign LUT_1[50043] = 32'b11111111111111101111101111000101;
assign LUT_1[50044] = 32'b00000000000000000010101000001111;
assign LUT_1[50045] = 32'b11111111111111111011111010001011;
assign LUT_1[50046] = 32'b11111111111111111110010110100000;
assign LUT_1[50047] = 32'b11111111111111110111101000011100;
assign LUT_1[50048] = 32'b11111111111111111001101100111101;
assign LUT_1[50049] = 32'b11111111111111110010111110111001;
assign LUT_1[50050] = 32'b11111111111111110101011011001110;
assign LUT_1[50051] = 32'b11111111111111101110101101001010;
assign LUT_1[50052] = 32'b00000000000000000001100110010100;
assign LUT_1[50053] = 32'b11111111111111111010111000010000;
assign LUT_1[50054] = 32'b11111111111111111101010100100101;
assign LUT_1[50055] = 32'b11111111111111110110100110100001;
assign LUT_1[50056] = 32'b11111111111111111000111010110010;
assign LUT_1[50057] = 32'b11111111111111110010001100101110;
assign LUT_1[50058] = 32'b11111111111111110100101001000011;
assign LUT_1[50059] = 32'b11111111111111101101111010111111;
assign LUT_1[50060] = 32'b00000000000000000000110100001001;
assign LUT_1[50061] = 32'b11111111111111111010000110000101;
assign LUT_1[50062] = 32'b11111111111111111100100010011010;
assign LUT_1[50063] = 32'b11111111111111110101110100010110;
assign LUT_1[50064] = 32'b11111111111111111011101000011111;
assign LUT_1[50065] = 32'b11111111111111110100111010011011;
assign LUT_1[50066] = 32'b11111111111111110111010110110000;
assign LUT_1[50067] = 32'b11111111111111110000101000101100;
assign LUT_1[50068] = 32'b00000000000000000011100001110110;
assign LUT_1[50069] = 32'b11111111111111111100110011110010;
assign LUT_1[50070] = 32'b11111111111111111111010000000111;
assign LUT_1[50071] = 32'b11111111111111111000100010000011;
assign LUT_1[50072] = 32'b11111111111111111010110110010100;
assign LUT_1[50073] = 32'b11111111111111110100001000010000;
assign LUT_1[50074] = 32'b11111111111111110110100100100101;
assign LUT_1[50075] = 32'b11111111111111101111110110100001;
assign LUT_1[50076] = 32'b00000000000000000010101111101011;
assign LUT_1[50077] = 32'b11111111111111111100000001100111;
assign LUT_1[50078] = 32'b11111111111111111110011101111100;
assign LUT_1[50079] = 32'b11111111111111110111101111111000;
assign LUT_1[50080] = 32'b11111111111111111010100111111100;
assign LUT_1[50081] = 32'b11111111111111110011111001111000;
assign LUT_1[50082] = 32'b11111111111111110110010110001101;
assign LUT_1[50083] = 32'b11111111111111101111101000001001;
assign LUT_1[50084] = 32'b00000000000000000010100001010011;
assign LUT_1[50085] = 32'b11111111111111111011110011001111;
assign LUT_1[50086] = 32'b11111111111111111110001111100100;
assign LUT_1[50087] = 32'b11111111111111110111100001100000;
assign LUT_1[50088] = 32'b11111111111111111001110101110001;
assign LUT_1[50089] = 32'b11111111111111110011000111101101;
assign LUT_1[50090] = 32'b11111111111111110101100100000010;
assign LUT_1[50091] = 32'b11111111111111101110110101111110;
assign LUT_1[50092] = 32'b00000000000000000001101111001000;
assign LUT_1[50093] = 32'b11111111111111111011000001000100;
assign LUT_1[50094] = 32'b11111111111111111101011101011001;
assign LUT_1[50095] = 32'b11111111111111110110101111010101;
assign LUT_1[50096] = 32'b11111111111111111100100011011110;
assign LUT_1[50097] = 32'b11111111111111110101110101011010;
assign LUT_1[50098] = 32'b11111111111111111000010001101111;
assign LUT_1[50099] = 32'b11111111111111110001100011101011;
assign LUT_1[50100] = 32'b00000000000000000100011100110101;
assign LUT_1[50101] = 32'b11111111111111111101101110110001;
assign LUT_1[50102] = 32'b00000000000000000000001011000110;
assign LUT_1[50103] = 32'b11111111111111111001011101000010;
assign LUT_1[50104] = 32'b11111111111111111011110001010011;
assign LUT_1[50105] = 32'b11111111111111110101000011001111;
assign LUT_1[50106] = 32'b11111111111111110111011111100100;
assign LUT_1[50107] = 32'b11111111111111110000110001100000;
assign LUT_1[50108] = 32'b00000000000000000011101010101010;
assign LUT_1[50109] = 32'b11111111111111111100111100100110;
assign LUT_1[50110] = 32'b11111111111111111111011000111011;
assign LUT_1[50111] = 32'b11111111111111111000101010110111;
assign LUT_1[50112] = 32'b11111111111111111011101010100101;
assign LUT_1[50113] = 32'b11111111111111110100111100100001;
assign LUT_1[50114] = 32'b11111111111111110111011000110110;
assign LUT_1[50115] = 32'b11111111111111110000101010110010;
assign LUT_1[50116] = 32'b00000000000000000011100011111100;
assign LUT_1[50117] = 32'b11111111111111111100110101111000;
assign LUT_1[50118] = 32'b11111111111111111111010010001101;
assign LUT_1[50119] = 32'b11111111111111111000100100001001;
assign LUT_1[50120] = 32'b11111111111111111010111000011010;
assign LUT_1[50121] = 32'b11111111111111110100001010010110;
assign LUT_1[50122] = 32'b11111111111111110110100110101011;
assign LUT_1[50123] = 32'b11111111111111101111111000100111;
assign LUT_1[50124] = 32'b00000000000000000010110001110001;
assign LUT_1[50125] = 32'b11111111111111111100000011101101;
assign LUT_1[50126] = 32'b11111111111111111110100000000010;
assign LUT_1[50127] = 32'b11111111111111110111110001111110;
assign LUT_1[50128] = 32'b11111111111111111101100110000111;
assign LUT_1[50129] = 32'b11111111111111110110111000000011;
assign LUT_1[50130] = 32'b11111111111111111001010100011000;
assign LUT_1[50131] = 32'b11111111111111110010100110010100;
assign LUT_1[50132] = 32'b00000000000000000101011111011110;
assign LUT_1[50133] = 32'b11111111111111111110110001011010;
assign LUT_1[50134] = 32'b00000000000000000001001101101111;
assign LUT_1[50135] = 32'b11111111111111111010011111101011;
assign LUT_1[50136] = 32'b11111111111111111100110011111100;
assign LUT_1[50137] = 32'b11111111111111110110000101111000;
assign LUT_1[50138] = 32'b11111111111111111000100010001101;
assign LUT_1[50139] = 32'b11111111111111110001110100001001;
assign LUT_1[50140] = 32'b00000000000000000100101101010011;
assign LUT_1[50141] = 32'b11111111111111111101111111001111;
assign LUT_1[50142] = 32'b00000000000000000000011011100100;
assign LUT_1[50143] = 32'b11111111111111111001101101100000;
assign LUT_1[50144] = 32'b11111111111111111100100101100100;
assign LUT_1[50145] = 32'b11111111111111110101110111100000;
assign LUT_1[50146] = 32'b11111111111111111000010011110101;
assign LUT_1[50147] = 32'b11111111111111110001100101110001;
assign LUT_1[50148] = 32'b00000000000000000100011110111011;
assign LUT_1[50149] = 32'b11111111111111111101110000110111;
assign LUT_1[50150] = 32'b00000000000000000000001101001100;
assign LUT_1[50151] = 32'b11111111111111111001011111001000;
assign LUT_1[50152] = 32'b11111111111111111011110011011001;
assign LUT_1[50153] = 32'b11111111111111110101000101010101;
assign LUT_1[50154] = 32'b11111111111111110111100001101010;
assign LUT_1[50155] = 32'b11111111111111110000110011100110;
assign LUT_1[50156] = 32'b00000000000000000011101100110000;
assign LUT_1[50157] = 32'b11111111111111111100111110101100;
assign LUT_1[50158] = 32'b11111111111111111111011011000001;
assign LUT_1[50159] = 32'b11111111111111111000101100111101;
assign LUT_1[50160] = 32'b11111111111111111110100001000110;
assign LUT_1[50161] = 32'b11111111111111110111110011000010;
assign LUT_1[50162] = 32'b11111111111111111010001111010111;
assign LUT_1[50163] = 32'b11111111111111110011100001010011;
assign LUT_1[50164] = 32'b00000000000000000110011010011101;
assign LUT_1[50165] = 32'b11111111111111111111101100011001;
assign LUT_1[50166] = 32'b00000000000000000010001000101110;
assign LUT_1[50167] = 32'b11111111111111111011011010101010;
assign LUT_1[50168] = 32'b11111111111111111101101110111011;
assign LUT_1[50169] = 32'b11111111111111110111000000110111;
assign LUT_1[50170] = 32'b11111111111111111001011101001100;
assign LUT_1[50171] = 32'b11111111111111110010101111001000;
assign LUT_1[50172] = 32'b00000000000000000101101000010010;
assign LUT_1[50173] = 32'b11111111111111111110111010001110;
assign LUT_1[50174] = 32'b00000000000000000001010110100011;
assign LUT_1[50175] = 32'b11111111111111111010101000011111;
assign LUT_1[50176] = 32'b00000000000000000101100001000001;
assign LUT_1[50177] = 32'b11111111111111111110110010111101;
assign LUT_1[50178] = 32'b00000000000000000001001111010010;
assign LUT_1[50179] = 32'b11111111111111111010100001001110;
assign LUT_1[50180] = 32'b00000000000000001101011010011000;
assign LUT_1[50181] = 32'b00000000000000000110101100010100;
assign LUT_1[50182] = 32'b00000000000000001001001000101001;
assign LUT_1[50183] = 32'b00000000000000000010011010100101;
assign LUT_1[50184] = 32'b00000000000000000100101110110110;
assign LUT_1[50185] = 32'b11111111111111111110000000110010;
assign LUT_1[50186] = 32'b00000000000000000000011101000111;
assign LUT_1[50187] = 32'b11111111111111111001101111000011;
assign LUT_1[50188] = 32'b00000000000000001100101000001101;
assign LUT_1[50189] = 32'b00000000000000000101111010001001;
assign LUT_1[50190] = 32'b00000000000000001000010110011110;
assign LUT_1[50191] = 32'b00000000000000000001101000011010;
assign LUT_1[50192] = 32'b00000000000000000111011100100011;
assign LUT_1[50193] = 32'b00000000000000000000101110011111;
assign LUT_1[50194] = 32'b00000000000000000011001010110100;
assign LUT_1[50195] = 32'b11111111111111111100011100110000;
assign LUT_1[50196] = 32'b00000000000000001111010101111010;
assign LUT_1[50197] = 32'b00000000000000001000100111110110;
assign LUT_1[50198] = 32'b00000000000000001011000100001011;
assign LUT_1[50199] = 32'b00000000000000000100010110000111;
assign LUT_1[50200] = 32'b00000000000000000110101010011000;
assign LUT_1[50201] = 32'b11111111111111111111111100010100;
assign LUT_1[50202] = 32'b00000000000000000010011000101001;
assign LUT_1[50203] = 32'b11111111111111111011101010100101;
assign LUT_1[50204] = 32'b00000000000000001110100011101111;
assign LUT_1[50205] = 32'b00000000000000000111110101101011;
assign LUT_1[50206] = 32'b00000000000000001010010010000000;
assign LUT_1[50207] = 32'b00000000000000000011100011111100;
assign LUT_1[50208] = 32'b00000000000000000110011100000000;
assign LUT_1[50209] = 32'b11111111111111111111101101111100;
assign LUT_1[50210] = 32'b00000000000000000010001010010001;
assign LUT_1[50211] = 32'b11111111111111111011011100001101;
assign LUT_1[50212] = 32'b00000000000000001110010101010111;
assign LUT_1[50213] = 32'b00000000000000000111100111010011;
assign LUT_1[50214] = 32'b00000000000000001010000011101000;
assign LUT_1[50215] = 32'b00000000000000000011010101100100;
assign LUT_1[50216] = 32'b00000000000000000101101001110101;
assign LUT_1[50217] = 32'b11111111111111111110111011110001;
assign LUT_1[50218] = 32'b00000000000000000001011000000110;
assign LUT_1[50219] = 32'b11111111111111111010101010000010;
assign LUT_1[50220] = 32'b00000000000000001101100011001100;
assign LUT_1[50221] = 32'b00000000000000000110110101001000;
assign LUT_1[50222] = 32'b00000000000000001001010001011101;
assign LUT_1[50223] = 32'b00000000000000000010100011011001;
assign LUT_1[50224] = 32'b00000000000000001000010111100010;
assign LUT_1[50225] = 32'b00000000000000000001101001011110;
assign LUT_1[50226] = 32'b00000000000000000100000101110011;
assign LUT_1[50227] = 32'b11111111111111111101010111101111;
assign LUT_1[50228] = 32'b00000000000000010000010000111001;
assign LUT_1[50229] = 32'b00000000000000001001100010110101;
assign LUT_1[50230] = 32'b00000000000000001011111111001010;
assign LUT_1[50231] = 32'b00000000000000000101010001000110;
assign LUT_1[50232] = 32'b00000000000000000111100101010111;
assign LUT_1[50233] = 32'b00000000000000000000110111010011;
assign LUT_1[50234] = 32'b00000000000000000011010011101000;
assign LUT_1[50235] = 32'b11111111111111111100100101100100;
assign LUT_1[50236] = 32'b00000000000000001111011110101110;
assign LUT_1[50237] = 32'b00000000000000001000110000101010;
assign LUT_1[50238] = 32'b00000000000000001011001100111111;
assign LUT_1[50239] = 32'b00000000000000000100011110111011;
assign LUT_1[50240] = 32'b00000000000000000111011110101001;
assign LUT_1[50241] = 32'b00000000000000000000110000100101;
assign LUT_1[50242] = 32'b00000000000000000011001100111010;
assign LUT_1[50243] = 32'b11111111111111111100011110110110;
assign LUT_1[50244] = 32'b00000000000000001111011000000000;
assign LUT_1[50245] = 32'b00000000000000001000101001111100;
assign LUT_1[50246] = 32'b00000000000000001011000110010001;
assign LUT_1[50247] = 32'b00000000000000000100011000001101;
assign LUT_1[50248] = 32'b00000000000000000110101100011110;
assign LUT_1[50249] = 32'b11111111111111111111111110011010;
assign LUT_1[50250] = 32'b00000000000000000010011010101111;
assign LUT_1[50251] = 32'b11111111111111111011101100101011;
assign LUT_1[50252] = 32'b00000000000000001110100101110101;
assign LUT_1[50253] = 32'b00000000000000000111110111110001;
assign LUT_1[50254] = 32'b00000000000000001010010100000110;
assign LUT_1[50255] = 32'b00000000000000000011100110000010;
assign LUT_1[50256] = 32'b00000000000000001001011010001011;
assign LUT_1[50257] = 32'b00000000000000000010101100000111;
assign LUT_1[50258] = 32'b00000000000000000101001000011100;
assign LUT_1[50259] = 32'b11111111111111111110011010011000;
assign LUT_1[50260] = 32'b00000000000000010001010011100010;
assign LUT_1[50261] = 32'b00000000000000001010100101011110;
assign LUT_1[50262] = 32'b00000000000000001101000001110011;
assign LUT_1[50263] = 32'b00000000000000000110010011101111;
assign LUT_1[50264] = 32'b00000000000000001000101000000000;
assign LUT_1[50265] = 32'b00000000000000000001111001111100;
assign LUT_1[50266] = 32'b00000000000000000100010110010001;
assign LUT_1[50267] = 32'b11111111111111111101101000001101;
assign LUT_1[50268] = 32'b00000000000000010000100001010111;
assign LUT_1[50269] = 32'b00000000000000001001110011010011;
assign LUT_1[50270] = 32'b00000000000000001100001111101000;
assign LUT_1[50271] = 32'b00000000000000000101100001100100;
assign LUT_1[50272] = 32'b00000000000000001000011001101000;
assign LUT_1[50273] = 32'b00000000000000000001101011100100;
assign LUT_1[50274] = 32'b00000000000000000100000111111001;
assign LUT_1[50275] = 32'b11111111111111111101011001110101;
assign LUT_1[50276] = 32'b00000000000000010000010010111111;
assign LUT_1[50277] = 32'b00000000000000001001100100111011;
assign LUT_1[50278] = 32'b00000000000000001100000001010000;
assign LUT_1[50279] = 32'b00000000000000000101010011001100;
assign LUT_1[50280] = 32'b00000000000000000111100111011101;
assign LUT_1[50281] = 32'b00000000000000000000111001011001;
assign LUT_1[50282] = 32'b00000000000000000011010101101110;
assign LUT_1[50283] = 32'b11111111111111111100100111101010;
assign LUT_1[50284] = 32'b00000000000000001111100000110100;
assign LUT_1[50285] = 32'b00000000000000001000110010110000;
assign LUT_1[50286] = 32'b00000000000000001011001111000101;
assign LUT_1[50287] = 32'b00000000000000000100100001000001;
assign LUT_1[50288] = 32'b00000000000000001010010101001010;
assign LUT_1[50289] = 32'b00000000000000000011100111000110;
assign LUT_1[50290] = 32'b00000000000000000110000011011011;
assign LUT_1[50291] = 32'b11111111111111111111010101010111;
assign LUT_1[50292] = 32'b00000000000000010010001110100001;
assign LUT_1[50293] = 32'b00000000000000001011100000011101;
assign LUT_1[50294] = 32'b00000000000000001101111100110010;
assign LUT_1[50295] = 32'b00000000000000000111001110101110;
assign LUT_1[50296] = 32'b00000000000000001001100010111111;
assign LUT_1[50297] = 32'b00000000000000000010110100111011;
assign LUT_1[50298] = 32'b00000000000000000101010001010000;
assign LUT_1[50299] = 32'b11111111111111111110100011001100;
assign LUT_1[50300] = 32'b00000000000000010001011100010110;
assign LUT_1[50301] = 32'b00000000000000001010101110010010;
assign LUT_1[50302] = 32'b00000000000000001101001010100111;
assign LUT_1[50303] = 32'b00000000000000000110011100100011;
assign LUT_1[50304] = 32'b00000000000000001000100001000100;
assign LUT_1[50305] = 32'b00000000000000000001110011000000;
assign LUT_1[50306] = 32'b00000000000000000100001111010101;
assign LUT_1[50307] = 32'b11111111111111111101100001010001;
assign LUT_1[50308] = 32'b00000000000000010000011010011011;
assign LUT_1[50309] = 32'b00000000000000001001101100010111;
assign LUT_1[50310] = 32'b00000000000000001100001000101100;
assign LUT_1[50311] = 32'b00000000000000000101011010101000;
assign LUT_1[50312] = 32'b00000000000000000111101110111001;
assign LUT_1[50313] = 32'b00000000000000000001000000110101;
assign LUT_1[50314] = 32'b00000000000000000011011101001010;
assign LUT_1[50315] = 32'b11111111111111111100101111000110;
assign LUT_1[50316] = 32'b00000000000000001111101000010000;
assign LUT_1[50317] = 32'b00000000000000001000111010001100;
assign LUT_1[50318] = 32'b00000000000000001011010110100001;
assign LUT_1[50319] = 32'b00000000000000000100101000011101;
assign LUT_1[50320] = 32'b00000000000000001010011100100110;
assign LUT_1[50321] = 32'b00000000000000000011101110100010;
assign LUT_1[50322] = 32'b00000000000000000110001010110111;
assign LUT_1[50323] = 32'b11111111111111111111011100110011;
assign LUT_1[50324] = 32'b00000000000000010010010101111101;
assign LUT_1[50325] = 32'b00000000000000001011100111111001;
assign LUT_1[50326] = 32'b00000000000000001110000100001110;
assign LUT_1[50327] = 32'b00000000000000000111010110001010;
assign LUT_1[50328] = 32'b00000000000000001001101010011011;
assign LUT_1[50329] = 32'b00000000000000000010111100010111;
assign LUT_1[50330] = 32'b00000000000000000101011000101100;
assign LUT_1[50331] = 32'b11111111111111111110101010101000;
assign LUT_1[50332] = 32'b00000000000000010001100011110010;
assign LUT_1[50333] = 32'b00000000000000001010110101101110;
assign LUT_1[50334] = 32'b00000000000000001101010010000011;
assign LUT_1[50335] = 32'b00000000000000000110100011111111;
assign LUT_1[50336] = 32'b00000000000000001001011100000011;
assign LUT_1[50337] = 32'b00000000000000000010101101111111;
assign LUT_1[50338] = 32'b00000000000000000101001010010100;
assign LUT_1[50339] = 32'b11111111111111111110011100010000;
assign LUT_1[50340] = 32'b00000000000000010001010101011010;
assign LUT_1[50341] = 32'b00000000000000001010100111010110;
assign LUT_1[50342] = 32'b00000000000000001101000011101011;
assign LUT_1[50343] = 32'b00000000000000000110010101100111;
assign LUT_1[50344] = 32'b00000000000000001000101001111000;
assign LUT_1[50345] = 32'b00000000000000000001111011110100;
assign LUT_1[50346] = 32'b00000000000000000100011000001001;
assign LUT_1[50347] = 32'b11111111111111111101101010000101;
assign LUT_1[50348] = 32'b00000000000000010000100011001111;
assign LUT_1[50349] = 32'b00000000000000001001110101001011;
assign LUT_1[50350] = 32'b00000000000000001100010001100000;
assign LUT_1[50351] = 32'b00000000000000000101100011011100;
assign LUT_1[50352] = 32'b00000000000000001011010111100101;
assign LUT_1[50353] = 32'b00000000000000000100101001100001;
assign LUT_1[50354] = 32'b00000000000000000111000101110110;
assign LUT_1[50355] = 32'b00000000000000000000010111110010;
assign LUT_1[50356] = 32'b00000000000000010011010000111100;
assign LUT_1[50357] = 32'b00000000000000001100100010111000;
assign LUT_1[50358] = 32'b00000000000000001110111111001101;
assign LUT_1[50359] = 32'b00000000000000001000010001001001;
assign LUT_1[50360] = 32'b00000000000000001010100101011010;
assign LUT_1[50361] = 32'b00000000000000000011110111010110;
assign LUT_1[50362] = 32'b00000000000000000110010011101011;
assign LUT_1[50363] = 32'b11111111111111111111100101100111;
assign LUT_1[50364] = 32'b00000000000000010010011110110001;
assign LUT_1[50365] = 32'b00000000000000001011110000101101;
assign LUT_1[50366] = 32'b00000000000000001110001101000010;
assign LUT_1[50367] = 32'b00000000000000000111011110111110;
assign LUT_1[50368] = 32'b00000000000000001010011110101100;
assign LUT_1[50369] = 32'b00000000000000000011110000101000;
assign LUT_1[50370] = 32'b00000000000000000110001100111101;
assign LUT_1[50371] = 32'b11111111111111111111011110111001;
assign LUT_1[50372] = 32'b00000000000000010010011000000011;
assign LUT_1[50373] = 32'b00000000000000001011101001111111;
assign LUT_1[50374] = 32'b00000000000000001110000110010100;
assign LUT_1[50375] = 32'b00000000000000000111011000010000;
assign LUT_1[50376] = 32'b00000000000000001001101100100001;
assign LUT_1[50377] = 32'b00000000000000000010111110011101;
assign LUT_1[50378] = 32'b00000000000000000101011010110010;
assign LUT_1[50379] = 32'b11111111111111111110101100101110;
assign LUT_1[50380] = 32'b00000000000000010001100101111000;
assign LUT_1[50381] = 32'b00000000000000001010110111110100;
assign LUT_1[50382] = 32'b00000000000000001101010100001001;
assign LUT_1[50383] = 32'b00000000000000000110100110000101;
assign LUT_1[50384] = 32'b00000000000000001100011010001110;
assign LUT_1[50385] = 32'b00000000000000000101101100001010;
assign LUT_1[50386] = 32'b00000000000000001000001000011111;
assign LUT_1[50387] = 32'b00000000000000000001011010011011;
assign LUT_1[50388] = 32'b00000000000000010100010011100101;
assign LUT_1[50389] = 32'b00000000000000001101100101100001;
assign LUT_1[50390] = 32'b00000000000000010000000001110110;
assign LUT_1[50391] = 32'b00000000000000001001010011110010;
assign LUT_1[50392] = 32'b00000000000000001011101000000011;
assign LUT_1[50393] = 32'b00000000000000000100111001111111;
assign LUT_1[50394] = 32'b00000000000000000111010110010100;
assign LUT_1[50395] = 32'b00000000000000000000101000010000;
assign LUT_1[50396] = 32'b00000000000000010011100001011010;
assign LUT_1[50397] = 32'b00000000000000001100110011010110;
assign LUT_1[50398] = 32'b00000000000000001111001111101011;
assign LUT_1[50399] = 32'b00000000000000001000100001100111;
assign LUT_1[50400] = 32'b00000000000000001011011001101011;
assign LUT_1[50401] = 32'b00000000000000000100101011100111;
assign LUT_1[50402] = 32'b00000000000000000111000111111100;
assign LUT_1[50403] = 32'b00000000000000000000011001111000;
assign LUT_1[50404] = 32'b00000000000000010011010011000010;
assign LUT_1[50405] = 32'b00000000000000001100100100111110;
assign LUT_1[50406] = 32'b00000000000000001111000001010011;
assign LUT_1[50407] = 32'b00000000000000001000010011001111;
assign LUT_1[50408] = 32'b00000000000000001010100111100000;
assign LUT_1[50409] = 32'b00000000000000000011111001011100;
assign LUT_1[50410] = 32'b00000000000000000110010101110001;
assign LUT_1[50411] = 32'b11111111111111111111100111101101;
assign LUT_1[50412] = 32'b00000000000000010010100000110111;
assign LUT_1[50413] = 32'b00000000000000001011110010110011;
assign LUT_1[50414] = 32'b00000000000000001110001111001000;
assign LUT_1[50415] = 32'b00000000000000000111100001000100;
assign LUT_1[50416] = 32'b00000000000000001101010101001101;
assign LUT_1[50417] = 32'b00000000000000000110100111001001;
assign LUT_1[50418] = 32'b00000000000000001001000011011110;
assign LUT_1[50419] = 32'b00000000000000000010010101011010;
assign LUT_1[50420] = 32'b00000000000000010101001110100100;
assign LUT_1[50421] = 32'b00000000000000001110100000100000;
assign LUT_1[50422] = 32'b00000000000000010000111100110101;
assign LUT_1[50423] = 32'b00000000000000001010001110110001;
assign LUT_1[50424] = 32'b00000000000000001100100011000010;
assign LUT_1[50425] = 32'b00000000000000000101110100111110;
assign LUT_1[50426] = 32'b00000000000000001000010001010011;
assign LUT_1[50427] = 32'b00000000000000000001100011001111;
assign LUT_1[50428] = 32'b00000000000000010100011100011001;
assign LUT_1[50429] = 32'b00000000000000001101101110010101;
assign LUT_1[50430] = 32'b00000000000000010000001010101010;
assign LUT_1[50431] = 32'b00000000000000001001011100100110;
assign LUT_1[50432] = 32'b00000000000000000011010101001101;
assign LUT_1[50433] = 32'b11111111111111111100100111001001;
assign LUT_1[50434] = 32'b11111111111111111111000011011110;
assign LUT_1[50435] = 32'b11111111111111111000010101011010;
assign LUT_1[50436] = 32'b00000000000000001011001110100100;
assign LUT_1[50437] = 32'b00000000000000000100100000100000;
assign LUT_1[50438] = 32'b00000000000000000110111100110101;
assign LUT_1[50439] = 32'b00000000000000000000001110110001;
assign LUT_1[50440] = 32'b00000000000000000010100011000010;
assign LUT_1[50441] = 32'b11111111111111111011110100111110;
assign LUT_1[50442] = 32'b11111111111111111110010001010011;
assign LUT_1[50443] = 32'b11111111111111110111100011001111;
assign LUT_1[50444] = 32'b00000000000000001010011100011001;
assign LUT_1[50445] = 32'b00000000000000000011101110010101;
assign LUT_1[50446] = 32'b00000000000000000110001010101010;
assign LUT_1[50447] = 32'b11111111111111111111011100100110;
assign LUT_1[50448] = 32'b00000000000000000101010000101111;
assign LUT_1[50449] = 32'b11111111111111111110100010101011;
assign LUT_1[50450] = 32'b00000000000000000000111111000000;
assign LUT_1[50451] = 32'b11111111111111111010010000111100;
assign LUT_1[50452] = 32'b00000000000000001101001010000110;
assign LUT_1[50453] = 32'b00000000000000000110011100000010;
assign LUT_1[50454] = 32'b00000000000000001000111000010111;
assign LUT_1[50455] = 32'b00000000000000000010001010010011;
assign LUT_1[50456] = 32'b00000000000000000100011110100100;
assign LUT_1[50457] = 32'b11111111111111111101110000100000;
assign LUT_1[50458] = 32'b00000000000000000000001100110101;
assign LUT_1[50459] = 32'b11111111111111111001011110110001;
assign LUT_1[50460] = 32'b00000000000000001100010111111011;
assign LUT_1[50461] = 32'b00000000000000000101101001110111;
assign LUT_1[50462] = 32'b00000000000000001000000110001100;
assign LUT_1[50463] = 32'b00000000000000000001011000001000;
assign LUT_1[50464] = 32'b00000000000000000100010000001100;
assign LUT_1[50465] = 32'b11111111111111111101100010001000;
assign LUT_1[50466] = 32'b11111111111111111111111110011101;
assign LUT_1[50467] = 32'b11111111111111111001010000011001;
assign LUT_1[50468] = 32'b00000000000000001100001001100011;
assign LUT_1[50469] = 32'b00000000000000000101011011011111;
assign LUT_1[50470] = 32'b00000000000000000111110111110100;
assign LUT_1[50471] = 32'b00000000000000000001001001110000;
assign LUT_1[50472] = 32'b00000000000000000011011110000001;
assign LUT_1[50473] = 32'b11111111111111111100101111111101;
assign LUT_1[50474] = 32'b11111111111111111111001100010010;
assign LUT_1[50475] = 32'b11111111111111111000011110001110;
assign LUT_1[50476] = 32'b00000000000000001011010111011000;
assign LUT_1[50477] = 32'b00000000000000000100101001010100;
assign LUT_1[50478] = 32'b00000000000000000111000101101001;
assign LUT_1[50479] = 32'b00000000000000000000010111100101;
assign LUT_1[50480] = 32'b00000000000000000110001011101110;
assign LUT_1[50481] = 32'b11111111111111111111011101101010;
assign LUT_1[50482] = 32'b00000000000000000001111001111111;
assign LUT_1[50483] = 32'b11111111111111111011001011111011;
assign LUT_1[50484] = 32'b00000000000000001110000101000101;
assign LUT_1[50485] = 32'b00000000000000000111010111000001;
assign LUT_1[50486] = 32'b00000000000000001001110011010110;
assign LUT_1[50487] = 32'b00000000000000000011000101010010;
assign LUT_1[50488] = 32'b00000000000000000101011001100011;
assign LUT_1[50489] = 32'b11111111111111111110101011011111;
assign LUT_1[50490] = 32'b00000000000000000001000111110100;
assign LUT_1[50491] = 32'b11111111111111111010011001110000;
assign LUT_1[50492] = 32'b00000000000000001101010010111010;
assign LUT_1[50493] = 32'b00000000000000000110100100110110;
assign LUT_1[50494] = 32'b00000000000000001001000001001011;
assign LUT_1[50495] = 32'b00000000000000000010010011000111;
assign LUT_1[50496] = 32'b00000000000000000101010010110101;
assign LUT_1[50497] = 32'b11111111111111111110100100110001;
assign LUT_1[50498] = 32'b00000000000000000001000001000110;
assign LUT_1[50499] = 32'b11111111111111111010010011000010;
assign LUT_1[50500] = 32'b00000000000000001101001100001100;
assign LUT_1[50501] = 32'b00000000000000000110011110001000;
assign LUT_1[50502] = 32'b00000000000000001000111010011101;
assign LUT_1[50503] = 32'b00000000000000000010001100011001;
assign LUT_1[50504] = 32'b00000000000000000100100000101010;
assign LUT_1[50505] = 32'b11111111111111111101110010100110;
assign LUT_1[50506] = 32'b00000000000000000000001110111011;
assign LUT_1[50507] = 32'b11111111111111111001100000110111;
assign LUT_1[50508] = 32'b00000000000000001100011010000001;
assign LUT_1[50509] = 32'b00000000000000000101101011111101;
assign LUT_1[50510] = 32'b00000000000000001000001000010010;
assign LUT_1[50511] = 32'b00000000000000000001011010001110;
assign LUT_1[50512] = 32'b00000000000000000111001110010111;
assign LUT_1[50513] = 32'b00000000000000000000100000010011;
assign LUT_1[50514] = 32'b00000000000000000010111100101000;
assign LUT_1[50515] = 32'b11111111111111111100001110100100;
assign LUT_1[50516] = 32'b00000000000000001111000111101110;
assign LUT_1[50517] = 32'b00000000000000001000011001101010;
assign LUT_1[50518] = 32'b00000000000000001010110101111111;
assign LUT_1[50519] = 32'b00000000000000000100000111111011;
assign LUT_1[50520] = 32'b00000000000000000110011100001100;
assign LUT_1[50521] = 32'b11111111111111111111101110001000;
assign LUT_1[50522] = 32'b00000000000000000010001010011101;
assign LUT_1[50523] = 32'b11111111111111111011011100011001;
assign LUT_1[50524] = 32'b00000000000000001110010101100011;
assign LUT_1[50525] = 32'b00000000000000000111100111011111;
assign LUT_1[50526] = 32'b00000000000000001010000011110100;
assign LUT_1[50527] = 32'b00000000000000000011010101110000;
assign LUT_1[50528] = 32'b00000000000000000110001101110100;
assign LUT_1[50529] = 32'b11111111111111111111011111110000;
assign LUT_1[50530] = 32'b00000000000000000001111100000101;
assign LUT_1[50531] = 32'b11111111111111111011001110000001;
assign LUT_1[50532] = 32'b00000000000000001110000111001011;
assign LUT_1[50533] = 32'b00000000000000000111011001000111;
assign LUT_1[50534] = 32'b00000000000000001001110101011100;
assign LUT_1[50535] = 32'b00000000000000000011000111011000;
assign LUT_1[50536] = 32'b00000000000000000101011011101001;
assign LUT_1[50537] = 32'b11111111111111111110101101100101;
assign LUT_1[50538] = 32'b00000000000000000001001001111010;
assign LUT_1[50539] = 32'b11111111111111111010011011110110;
assign LUT_1[50540] = 32'b00000000000000001101010101000000;
assign LUT_1[50541] = 32'b00000000000000000110100110111100;
assign LUT_1[50542] = 32'b00000000000000001001000011010001;
assign LUT_1[50543] = 32'b00000000000000000010010101001101;
assign LUT_1[50544] = 32'b00000000000000001000001001010110;
assign LUT_1[50545] = 32'b00000000000000000001011011010010;
assign LUT_1[50546] = 32'b00000000000000000011110111100111;
assign LUT_1[50547] = 32'b11111111111111111101001001100011;
assign LUT_1[50548] = 32'b00000000000000010000000010101101;
assign LUT_1[50549] = 32'b00000000000000001001010100101001;
assign LUT_1[50550] = 32'b00000000000000001011110000111110;
assign LUT_1[50551] = 32'b00000000000000000101000010111010;
assign LUT_1[50552] = 32'b00000000000000000111010111001011;
assign LUT_1[50553] = 32'b00000000000000000000101001000111;
assign LUT_1[50554] = 32'b00000000000000000011000101011100;
assign LUT_1[50555] = 32'b11111111111111111100010111011000;
assign LUT_1[50556] = 32'b00000000000000001111010000100010;
assign LUT_1[50557] = 32'b00000000000000001000100010011110;
assign LUT_1[50558] = 32'b00000000000000001010111110110011;
assign LUT_1[50559] = 32'b00000000000000000100010000101111;
assign LUT_1[50560] = 32'b00000000000000000110010101010000;
assign LUT_1[50561] = 32'b11111111111111111111100111001100;
assign LUT_1[50562] = 32'b00000000000000000010000011100001;
assign LUT_1[50563] = 32'b11111111111111111011010101011101;
assign LUT_1[50564] = 32'b00000000000000001110001110100111;
assign LUT_1[50565] = 32'b00000000000000000111100000100011;
assign LUT_1[50566] = 32'b00000000000000001001111100111000;
assign LUT_1[50567] = 32'b00000000000000000011001110110100;
assign LUT_1[50568] = 32'b00000000000000000101100011000101;
assign LUT_1[50569] = 32'b11111111111111111110110101000001;
assign LUT_1[50570] = 32'b00000000000000000001010001010110;
assign LUT_1[50571] = 32'b11111111111111111010100011010010;
assign LUT_1[50572] = 32'b00000000000000001101011100011100;
assign LUT_1[50573] = 32'b00000000000000000110101110011000;
assign LUT_1[50574] = 32'b00000000000000001001001010101101;
assign LUT_1[50575] = 32'b00000000000000000010011100101001;
assign LUT_1[50576] = 32'b00000000000000001000010000110010;
assign LUT_1[50577] = 32'b00000000000000000001100010101110;
assign LUT_1[50578] = 32'b00000000000000000011111111000011;
assign LUT_1[50579] = 32'b11111111111111111101010000111111;
assign LUT_1[50580] = 32'b00000000000000010000001010001001;
assign LUT_1[50581] = 32'b00000000000000001001011100000101;
assign LUT_1[50582] = 32'b00000000000000001011111000011010;
assign LUT_1[50583] = 32'b00000000000000000101001010010110;
assign LUT_1[50584] = 32'b00000000000000000111011110100111;
assign LUT_1[50585] = 32'b00000000000000000000110000100011;
assign LUT_1[50586] = 32'b00000000000000000011001100111000;
assign LUT_1[50587] = 32'b11111111111111111100011110110100;
assign LUT_1[50588] = 32'b00000000000000001111010111111110;
assign LUT_1[50589] = 32'b00000000000000001000101001111010;
assign LUT_1[50590] = 32'b00000000000000001011000110001111;
assign LUT_1[50591] = 32'b00000000000000000100011000001011;
assign LUT_1[50592] = 32'b00000000000000000111010000001111;
assign LUT_1[50593] = 32'b00000000000000000000100010001011;
assign LUT_1[50594] = 32'b00000000000000000010111110100000;
assign LUT_1[50595] = 32'b11111111111111111100010000011100;
assign LUT_1[50596] = 32'b00000000000000001111001001100110;
assign LUT_1[50597] = 32'b00000000000000001000011011100010;
assign LUT_1[50598] = 32'b00000000000000001010110111110111;
assign LUT_1[50599] = 32'b00000000000000000100001001110011;
assign LUT_1[50600] = 32'b00000000000000000110011110000100;
assign LUT_1[50601] = 32'b11111111111111111111110000000000;
assign LUT_1[50602] = 32'b00000000000000000010001100010101;
assign LUT_1[50603] = 32'b11111111111111111011011110010001;
assign LUT_1[50604] = 32'b00000000000000001110010111011011;
assign LUT_1[50605] = 32'b00000000000000000111101001010111;
assign LUT_1[50606] = 32'b00000000000000001010000101101100;
assign LUT_1[50607] = 32'b00000000000000000011010111101000;
assign LUT_1[50608] = 32'b00000000000000001001001011110001;
assign LUT_1[50609] = 32'b00000000000000000010011101101101;
assign LUT_1[50610] = 32'b00000000000000000100111010000010;
assign LUT_1[50611] = 32'b11111111111111111110001011111110;
assign LUT_1[50612] = 32'b00000000000000010001000101001000;
assign LUT_1[50613] = 32'b00000000000000001010010111000100;
assign LUT_1[50614] = 32'b00000000000000001100110011011001;
assign LUT_1[50615] = 32'b00000000000000000110000101010101;
assign LUT_1[50616] = 32'b00000000000000001000011001100110;
assign LUT_1[50617] = 32'b00000000000000000001101011100010;
assign LUT_1[50618] = 32'b00000000000000000100000111110111;
assign LUT_1[50619] = 32'b11111111111111111101011001110011;
assign LUT_1[50620] = 32'b00000000000000010000010010111101;
assign LUT_1[50621] = 32'b00000000000000001001100100111001;
assign LUT_1[50622] = 32'b00000000000000001100000001001110;
assign LUT_1[50623] = 32'b00000000000000000101010011001010;
assign LUT_1[50624] = 32'b00000000000000001000010010111000;
assign LUT_1[50625] = 32'b00000000000000000001100100110100;
assign LUT_1[50626] = 32'b00000000000000000100000001001001;
assign LUT_1[50627] = 32'b11111111111111111101010011000101;
assign LUT_1[50628] = 32'b00000000000000010000001100001111;
assign LUT_1[50629] = 32'b00000000000000001001011110001011;
assign LUT_1[50630] = 32'b00000000000000001011111010100000;
assign LUT_1[50631] = 32'b00000000000000000101001100011100;
assign LUT_1[50632] = 32'b00000000000000000111100000101101;
assign LUT_1[50633] = 32'b00000000000000000000110010101001;
assign LUT_1[50634] = 32'b00000000000000000011001110111110;
assign LUT_1[50635] = 32'b11111111111111111100100000111010;
assign LUT_1[50636] = 32'b00000000000000001111011010000100;
assign LUT_1[50637] = 32'b00000000000000001000101100000000;
assign LUT_1[50638] = 32'b00000000000000001011001000010101;
assign LUT_1[50639] = 32'b00000000000000000100011010010001;
assign LUT_1[50640] = 32'b00000000000000001010001110011010;
assign LUT_1[50641] = 32'b00000000000000000011100000010110;
assign LUT_1[50642] = 32'b00000000000000000101111100101011;
assign LUT_1[50643] = 32'b11111111111111111111001110100111;
assign LUT_1[50644] = 32'b00000000000000010010000111110001;
assign LUT_1[50645] = 32'b00000000000000001011011001101101;
assign LUT_1[50646] = 32'b00000000000000001101110110000010;
assign LUT_1[50647] = 32'b00000000000000000111000111111110;
assign LUT_1[50648] = 32'b00000000000000001001011100001111;
assign LUT_1[50649] = 32'b00000000000000000010101110001011;
assign LUT_1[50650] = 32'b00000000000000000101001010100000;
assign LUT_1[50651] = 32'b11111111111111111110011100011100;
assign LUT_1[50652] = 32'b00000000000000010001010101100110;
assign LUT_1[50653] = 32'b00000000000000001010100111100010;
assign LUT_1[50654] = 32'b00000000000000001101000011110111;
assign LUT_1[50655] = 32'b00000000000000000110010101110011;
assign LUT_1[50656] = 32'b00000000000000001001001101110111;
assign LUT_1[50657] = 32'b00000000000000000010011111110011;
assign LUT_1[50658] = 32'b00000000000000000100111100001000;
assign LUT_1[50659] = 32'b11111111111111111110001110000100;
assign LUT_1[50660] = 32'b00000000000000010001000111001110;
assign LUT_1[50661] = 32'b00000000000000001010011001001010;
assign LUT_1[50662] = 32'b00000000000000001100110101011111;
assign LUT_1[50663] = 32'b00000000000000000110000111011011;
assign LUT_1[50664] = 32'b00000000000000001000011011101100;
assign LUT_1[50665] = 32'b00000000000000000001101101101000;
assign LUT_1[50666] = 32'b00000000000000000100001001111101;
assign LUT_1[50667] = 32'b11111111111111111101011011111001;
assign LUT_1[50668] = 32'b00000000000000010000010101000011;
assign LUT_1[50669] = 32'b00000000000000001001100110111111;
assign LUT_1[50670] = 32'b00000000000000001100000011010100;
assign LUT_1[50671] = 32'b00000000000000000101010101010000;
assign LUT_1[50672] = 32'b00000000000000001011001001011001;
assign LUT_1[50673] = 32'b00000000000000000100011011010101;
assign LUT_1[50674] = 32'b00000000000000000110110111101010;
assign LUT_1[50675] = 32'b00000000000000000000001001100110;
assign LUT_1[50676] = 32'b00000000000000010011000010110000;
assign LUT_1[50677] = 32'b00000000000000001100010100101100;
assign LUT_1[50678] = 32'b00000000000000001110110001000001;
assign LUT_1[50679] = 32'b00000000000000001000000010111101;
assign LUT_1[50680] = 32'b00000000000000001010010111001110;
assign LUT_1[50681] = 32'b00000000000000000011101001001010;
assign LUT_1[50682] = 32'b00000000000000000110000101011111;
assign LUT_1[50683] = 32'b11111111111111111111010111011011;
assign LUT_1[50684] = 32'b00000000000000010010010000100101;
assign LUT_1[50685] = 32'b00000000000000001011100010100001;
assign LUT_1[50686] = 32'b00000000000000001101111110110110;
assign LUT_1[50687] = 32'b00000000000000000111010000110010;
assign LUT_1[50688] = 32'b11111111111111111111001111011110;
assign LUT_1[50689] = 32'b11111111111111111000100001011010;
assign LUT_1[50690] = 32'b11111111111111111010111101101111;
assign LUT_1[50691] = 32'b11111111111111110100001111101011;
assign LUT_1[50692] = 32'b00000000000000000111001000110101;
assign LUT_1[50693] = 32'b00000000000000000000011010110001;
assign LUT_1[50694] = 32'b00000000000000000010110111000110;
assign LUT_1[50695] = 32'b11111111111111111100001001000010;
assign LUT_1[50696] = 32'b11111111111111111110011101010011;
assign LUT_1[50697] = 32'b11111111111111110111101111001111;
assign LUT_1[50698] = 32'b11111111111111111010001011100100;
assign LUT_1[50699] = 32'b11111111111111110011011101100000;
assign LUT_1[50700] = 32'b00000000000000000110010110101010;
assign LUT_1[50701] = 32'b11111111111111111111101000100110;
assign LUT_1[50702] = 32'b00000000000000000010000100111011;
assign LUT_1[50703] = 32'b11111111111111111011010110110111;
assign LUT_1[50704] = 32'b00000000000000000001001011000000;
assign LUT_1[50705] = 32'b11111111111111111010011100111100;
assign LUT_1[50706] = 32'b11111111111111111100111001010001;
assign LUT_1[50707] = 32'b11111111111111110110001011001101;
assign LUT_1[50708] = 32'b00000000000000001001000100010111;
assign LUT_1[50709] = 32'b00000000000000000010010110010011;
assign LUT_1[50710] = 32'b00000000000000000100110010101000;
assign LUT_1[50711] = 32'b11111111111111111110000100100100;
assign LUT_1[50712] = 32'b00000000000000000000011000110101;
assign LUT_1[50713] = 32'b11111111111111111001101010110001;
assign LUT_1[50714] = 32'b11111111111111111100000111000110;
assign LUT_1[50715] = 32'b11111111111111110101011001000010;
assign LUT_1[50716] = 32'b00000000000000001000010010001100;
assign LUT_1[50717] = 32'b00000000000000000001100100001000;
assign LUT_1[50718] = 32'b00000000000000000100000000011101;
assign LUT_1[50719] = 32'b11111111111111111101010010011001;
assign LUT_1[50720] = 32'b00000000000000000000001010011101;
assign LUT_1[50721] = 32'b11111111111111111001011100011001;
assign LUT_1[50722] = 32'b11111111111111111011111000101110;
assign LUT_1[50723] = 32'b11111111111111110101001010101010;
assign LUT_1[50724] = 32'b00000000000000001000000011110100;
assign LUT_1[50725] = 32'b00000000000000000001010101110000;
assign LUT_1[50726] = 32'b00000000000000000011110010000101;
assign LUT_1[50727] = 32'b11111111111111111101000100000001;
assign LUT_1[50728] = 32'b11111111111111111111011000010010;
assign LUT_1[50729] = 32'b11111111111111111000101010001110;
assign LUT_1[50730] = 32'b11111111111111111011000110100011;
assign LUT_1[50731] = 32'b11111111111111110100011000011111;
assign LUT_1[50732] = 32'b00000000000000000111010001101001;
assign LUT_1[50733] = 32'b00000000000000000000100011100101;
assign LUT_1[50734] = 32'b00000000000000000010111111111010;
assign LUT_1[50735] = 32'b11111111111111111100010001110110;
assign LUT_1[50736] = 32'b00000000000000000010000101111111;
assign LUT_1[50737] = 32'b11111111111111111011010111111011;
assign LUT_1[50738] = 32'b11111111111111111101110100010000;
assign LUT_1[50739] = 32'b11111111111111110111000110001100;
assign LUT_1[50740] = 32'b00000000000000001001111111010110;
assign LUT_1[50741] = 32'b00000000000000000011010001010010;
assign LUT_1[50742] = 32'b00000000000000000101101101100111;
assign LUT_1[50743] = 32'b11111111111111111110111111100011;
assign LUT_1[50744] = 32'b00000000000000000001010011110100;
assign LUT_1[50745] = 32'b11111111111111111010100101110000;
assign LUT_1[50746] = 32'b11111111111111111101000010000101;
assign LUT_1[50747] = 32'b11111111111111110110010100000001;
assign LUT_1[50748] = 32'b00000000000000001001001101001011;
assign LUT_1[50749] = 32'b00000000000000000010011111000111;
assign LUT_1[50750] = 32'b00000000000000000100111011011100;
assign LUT_1[50751] = 32'b11111111111111111110001101011000;
assign LUT_1[50752] = 32'b00000000000000000001001101000110;
assign LUT_1[50753] = 32'b11111111111111111010011111000010;
assign LUT_1[50754] = 32'b11111111111111111100111011010111;
assign LUT_1[50755] = 32'b11111111111111110110001101010011;
assign LUT_1[50756] = 32'b00000000000000001001000110011101;
assign LUT_1[50757] = 32'b00000000000000000010011000011001;
assign LUT_1[50758] = 32'b00000000000000000100110100101110;
assign LUT_1[50759] = 32'b11111111111111111110000110101010;
assign LUT_1[50760] = 32'b00000000000000000000011010111011;
assign LUT_1[50761] = 32'b11111111111111111001101100110111;
assign LUT_1[50762] = 32'b11111111111111111100001001001100;
assign LUT_1[50763] = 32'b11111111111111110101011011001000;
assign LUT_1[50764] = 32'b00000000000000001000010100010010;
assign LUT_1[50765] = 32'b00000000000000000001100110001110;
assign LUT_1[50766] = 32'b00000000000000000100000010100011;
assign LUT_1[50767] = 32'b11111111111111111101010100011111;
assign LUT_1[50768] = 32'b00000000000000000011001000101000;
assign LUT_1[50769] = 32'b11111111111111111100011010100100;
assign LUT_1[50770] = 32'b11111111111111111110110110111001;
assign LUT_1[50771] = 32'b11111111111111111000001000110101;
assign LUT_1[50772] = 32'b00000000000000001011000001111111;
assign LUT_1[50773] = 32'b00000000000000000100010011111011;
assign LUT_1[50774] = 32'b00000000000000000110110000010000;
assign LUT_1[50775] = 32'b00000000000000000000000010001100;
assign LUT_1[50776] = 32'b00000000000000000010010110011101;
assign LUT_1[50777] = 32'b11111111111111111011101000011001;
assign LUT_1[50778] = 32'b11111111111111111110000100101110;
assign LUT_1[50779] = 32'b11111111111111110111010110101010;
assign LUT_1[50780] = 32'b00000000000000001010001111110100;
assign LUT_1[50781] = 32'b00000000000000000011100001110000;
assign LUT_1[50782] = 32'b00000000000000000101111110000101;
assign LUT_1[50783] = 32'b11111111111111111111010000000001;
assign LUT_1[50784] = 32'b00000000000000000010001000000101;
assign LUT_1[50785] = 32'b11111111111111111011011010000001;
assign LUT_1[50786] = 32'b11111111111111111101110110010110;
assign LUT_1[50787] = 32'b11111111111111110111001000010010;
assign LUT_1[50788] = 32'b00000000000000001010000001011100;
assign LUT_1[50789] = 32'b00000000000000000011010011011000;
assign LUT_1[50790] = 32'b00000000000000000101101111101101;
assign LUT_1[50791] = 32'b11111111111111111111000001101001;
assign LUT_1[50792] = 32'b00000000000000000001010101111010;
assign LUT_1[50793] = 32'b11111111111111111010100111110110;
assign LUT_1[50794] = 32'b11111111111111111101000100001011;
assign LUT_1[50795] = 32'b11111111111111110110010110000111;
assign LUT_1[50796] = 32'b00000000000000001001001111010001;
assign LUT_1[50797] = 32'b00000000000000000010100001001101;
assign LUT_1[50798] = 32'b00000000000000000100111101100010;
assign LUT_1[50799] = 32'b11111111111111111110001111011110;
assign LUT_1[50800] = 32'b00000000000000000100000011100111;
assign LUT_1[50801] = 32'b11111111111111111101010101100011;
assign LUT_1[50802] = 32'b11111111111111111111110001111000;
assign LUT_1[50803] = 32'b11111111111111111001000011110100;
assign LUT_1[50804] = 32'b00000000000000001011111100111110;
assign LUT_1[50805] = 32'b00000000000000000101001110111010;
assign LUT_1[50806] = 32'b00000000000000000111101011001111;
assign LUT_1[50807] = 32'b00000000000000000000111101001011;
assign LUT_1[50808] = 32'b00000000000000000011010001011100;
assign LUT_1[50809] = 32'b11111111111111111100100011011000;
assign LUT_1[50810] = 32'b11111111111111111110111111101101;
assign LUT_1[50811] = 32'b11111111111111111000010001101001;
assign LUT_1[50812] = 32'b00000000000000001011001010110011;
assign LUT_1[50813] = 32'b00000000000000000100011100101111;
assign LUT_1[50814] = 32'b00000000000000000110111001000100;
assign LUT_1[50815] = 32'b00000000000000000000001011000000;
assign LUT_1[50816] = 32'b00000000000000000010001111100001;
assign LUT_1[50817] = 32'b11111111111111111011100001011101;
assign LUT_1[50818] = 32'b11111111111111111101111101110010;
assign LUT_1[50819] = 32'b11111111111111110111001111101110;
assign LUT_1[50820] = 32'b00000000000000001010001000111000;
assign LUT_1[50821] = 32'b00000000000000000011011010110100;
assign LUT_1[50822] = 32'b00000000000000000101110111001001;
assign LUT_1[50823] = 32'b11111111111111111111001001000101;
assign LUT_1[50824] = 32'b00000000000000000001011101010110;
assign LUT_1[50825] = 32'b11111111111111111010101111010010;
assign LUT_1[50826] = 32'b11111111111111111101001011100111;
assign LUT_1[50827] = 32'b11111111111111110110011101100011;
assign LUT_1[50828] = 32'b00000000000000001001010110101101;
assign LUT_1[50829] = 32'b00000000000000000010101000101001;
assign LUT_1[50830] = 32'b00000000000000000101000100111110;
assign LUT_1[50831] = 32'b11111111111111111110010110111010;
assign LUT_1[50832] = 32'b00000000000000000100001011000011;
assign LUT_1[50833] = 32'b11111111111111111101011100111111;
assign LUT_1[50834] = 32'b11111111111111111111111001010100;
assign LUT_1[50835] = 32'b11111111111111111001001011010000;
assign LUT_1[50836] = 32'b00000000000000001100000100011010;
assign LUT_1[50837] = 32'b00000000000000000101010110010110;
assign LUT_1[50838] = 32'b00000000000000000111110010101011;
assign LUT_1[50839] = 32'b00000000000000000001000100100111;
assign LUT_1[50840] = 32'b00000000000000000011011000111000;
assign LUT_1[50841] = 32'b11111111111111111100101010110100;
assign LUT_1[50842] = 32'b11111111111111111111000111001001;
assign LUT_1[50843] = 32'b11111111111111111000011001000101;
assign LUT_1[50844] = 32'b00000000000000001011010010001111;
assign LUT_1[50845] = 32'b00000000000000000100100100001011;
assign LUT_1[50846] = 32'b00000000000000000111000000100000;
assign LUT_1[50847] = 32'b00000000000000000000010010011100;
assign LUT_1[50848] = 32'b00000000000000000011001010100000;
assign LUT_1[50849] = 32'b11111111111111111100011100011100;
assign LUT_1[50850] = 32'b11111111111111111110111000110001;
assign LUT_1[50851] = 32'b11111111111111111000001010101101;
assign LUT_1[50852] = 32'b00000000000000001011000011110111;
assign LUT_1[50853] = 32'b00000000000000000100010101110011;
assign LUT_1[50854] = 32'b00000000000000000110110010001000;
assign LUT_1[50855] = 32'b00000000000000000000000100000100;
assign LUT_1[50856] = 32'b00000000000000000010011000010101;
assign LUT_1[50857] = 32'b11111111111111111011101010010001;
assign LUT_1[50858] = 32'b11111111111111111110000110100110;
assign LUT_1[50859] = 32'b11111111111111110111011000100010;
assign LUT_1[50860] = 32'b00000000000000001010010001101100;
assign LUT_1[50861] = 32'b00000000000000000011100011101000;
assign LUT_1[50862] = 32'b00000000000000000101111111111101;
assign LUT_1[50863] = 32'b11111111111111111111010001111001;
assign LUT_1[50864] = 32'b00000000000000000101000110000010;
assign LUT_1[50865] = 32'b11111111111111111110010111111110;
assign LUT_1[50866] = 32'b00000000000000000000110100010011;
assign LUT_1[50867] = 32'b11111111111111111010000110001111;
assign LUT_1[50868] = 32'b00000000000000001100111111011001;
assign LUT_1[50869] = 32'b00000000000000000110010001010101;
assign LUT_1[50870] = 32'b00000000000000001000101101101010;
assign LUT_1[50871] = 32'b00000000000000000001111111100110;
assign LUT_1[50872] = 32'b00000000000000000100010011110111;
assign LUT_1[50873] = 32'b11111111111111111101100101110011;
assign LUT_1[50874] = 32'b00000000000000000000000010001000;
assign LUT_1[50875] = 32'b11111111111111111001010100000100;
assign LUT_1[50876] = 32'b00000000000000001100001101001110;
assign LUT_1[50877] = 32'b00000000000000000101011111001010;
assign LUT_1[50878] = 32'b00000000000000000111111011011111;
assign LUT_1[50879] = 32'b00000000000000000001001101011011;
assign LUT_1[50880] = 32'b00000000000000000100001101001001;
assign LUT_1[50881] = 32'b11111111111111111101011111000101;
assign LUT_1[50882] = 32'b11111111111111111111111011011010;
assign LUT_1[50883] = 32'b11111111111111111001001101010110;
assign LUT_1[50884] = 32'b00000000000000001100000110100000;
assign LUT_1[50885] = 32'b00000000000000000101011000011100;
assign LUT_1[50886] = 32'b00000000000000000111110100110001;
assign LUT_1[50887] = 32'b00000000000000000001000110101101;
assign LUT_1[50888] = 32'b00000000000000000011011010111110;
assign LUT_1[50889] = 32'b11111111111111111100101100111010;
assign LUT_1[50890] = 32'b11111111111111111111001001001111;
assign LUT_1[50891] = 32'b11111111111111111000011011001011;
assign LUT_1[50892] = 32'b00000000000000001011010100010101;
assign LUT_1[50893] = 32'b00000000000000000100100110010001;
assign LUT_1[50894] = 32'b00000000000000000111000010100110;
assign LUT_1[50895] = 32'b00000000000000000000010100100010;
assign LUT_1[50896] = 32'b00000000000000000110001000101011;
assign LUT_1[50897] = 32'b11111111111111111111011010100111;
assign LUT_1[50898] = 32'b00000000000000000001110110111100;
assign LUT_1[50899] = 32'b11111111111111111011001000111000;
assign LUT_1[50900] = 32'b00000000000000001110000010000010;
assign LUT_1[50901] = 32'b00000000000000000111010011111110;
assign LUT_1[50902] = 32'b00000000000000001001110000010011;
assign LUT_1[50903] = 32'b00000000000000000011000010001111;
assign LUT_1[50904] = 32'b00000000000000000101010110100000;
assign LUT_1[50905] = 32'b11111111111111111110101000011100;
assign LUT_1[50906] = 32'b00000000000000000001000100110001;
assign LUT_1[50907] = 32'b11111111111111111010010110101101;
assign LUT_1[50908] = 32'b00000000000000001101001111110111;
assign LUT_1[50909] = 32'b00000000000000000110100001110011;
assign LUT_1[50910] = 32'b00000000000000001000111110001000;
assign LUT_1[50911] = 32'b00000000000000000010010000000100;
assign LUT_1[50912] = 32'b00000000000000000101001000001000;
assign LUT_1[50913] = 32'b11111111111111111110011010000100;
assign LUT_1[50914] = 32'b00000000000000000000110110011001;
assign LUT_1[50915] = 32'b11111111111111111010001000010101;
assign LUT_1[50916] = 32'b00000000000000001101000001011111;
assign LUT_1[50917] = 32'b00000000000000000110010011011011;
assign LUT_1[50918] = 32'b00000000000000001000101111110000;
assign LUT_1[50919] = 32'b00000000000000000010000001101100;
assign LUT_1[50920] = 32'b00000000000000000100010101111101;
assign LUT_1[50921] = 32'b11111111111111111101100111111001;
assign LUT_1[50922] = 32'b00000000000000000000000100001110;
assign LUT_1[50923] = 32'b11111111111111111001010110001010;
assign LUT_1[50924] = 32'b00000000000000001100001111010100;
assign LUT_1[50925] = 32'b00000000000000000101100001010000;
assign LUT_1[50926] = 32'b00000000000000000111111101100101;
assign LUT_1[50927] = 32'b00000000000000000001001111100001;
assign LUT_1[50928] = 32'b00000000000000000111000011101010;
assign LUT_1[50929] = 32'b00000000000000000000010101100110;
assign LUT_1[50930] = 32'b00000000000000000010110001111011;
assign LUT_1[50931] = 32'b11111111111111111100000011110111;
assign LUT_1[50932] = 32'b00000000000000001110111101000001;
assign LUT_1[50933] = 32'b00000000000000001000001110111101;
assign LUT_1[50934] = 32'b00000000000000001010101011010010;
assign LUT_1[50935] = 32'b00000000000000000011111101001110;
assign LUT_1[50936] = 32'b00000000000000000110010001011111;
assign LUT_1[50937] = 32'b11111111111111111111100011011011;
assign LUT_1[50938] = 32'b00000000000000000001111111110000;
assign LUT_1[50939] = 32'b11111111111111111011010001101100;
assign LUT_1[50940] = 32'b00000000000000001110001010110110;
assign LUT_1[50941] = 32'b00000000000000000111011100110010;
assign LUT_1[50942] = 32'b00000000000000001001111001000111;
assign LUT_1[50943] = 32'b00000000000000000011001011000011;
assign LUT_1[50944] = 32'b11111111111111111101000011101010;
assign LUT_1[50945] = 32'b11111111111111110110010101100110;
assign LUT_1[50946] = 32'b11111111111111111000110001111011;
assign LUT_1[50947] = 32'b11111111111111110010000011110111;
assign LUT_1[50948] = 32'b00000000000000000100111101000001;
assign LUT_1[50949] = 32'b11111111111111111110001110111101;
assign LUT_1[50950] = 32'b00000000000000000000101011010010;
assign LUT_1[50951] = 32'b11111111111111111001111101001110;
assign LUT_1[50952] = 32'b11111111111111111100010001011111;
assign LUT_1[50953] = 32'b11111111111111110101100011011011;
assign LUT_1[50954] = 32'b11111111111111110111111111110000;
assign LUT_1[50955] = 32'b11111111111111110001010001101100;
assign LUT_1[50956] = 32'b00000000000000000100001010110110;
assign LUT_1[50957] = 32'b11111111111111111101011100110010;
assign LUT_1[50958] = 32'b11111111111111111111111001000111;
assign LUT_1[50959] = 32'b11111111111111111001001011000011;
assign LUT_1[50960] = 32'b11111111111111111110111111001100;
assign LUT_1[50961] = 32'b11111111111111111000010001001000;
assign LUT_1[50962] = 32'b11111111111111111010101101011101;
assign LUT_1[50963] = 32'b11111111111111110011111111011001;
assign LUT_1[50964] = 32'b00000000000000000110111000100011;
assign LUT_1[50965] = 32'b00000000000000000000001010011111;
assign LUT_1[50966] = 32'b00000000000000000010100110110100;
assign LUT_1[50967] = 32'b11111111111111111011111000110000;
assign LUT_1[50968] = 32'b11111111111111111110001101000001;
assign LUT_1[50969] = 32'b11111111111111110111011110111101;
assign LUT_1[50970] = 32'b11111111111111111001111011010010;
assign LUT_1[50971] = 32'b11111111111111110011001101001110;
assign LUT_1[50972] = 32'b00000000000000000110000110011000;
assign LUT_1[50973] = 32'b11111111111111111111011000010100;
assign LUT_1[50974] = 32'b00000000000000000001110100101001;
assign LUT_1[50975] = 32'b11111111111111111011000110100101;
assign LUT_1[50976] = 32'b11111111111111111101111110101001;
assign LUT_1[50977] = 32'b11111111111111110111010000100101;
assign LUT_1[50978] = 32'b11111111111111111001101100111010;
assign LUT_1[50979] = 32'b11111111111111110010111110110110;
assign LUT_1[50980] = 32'b00000000000000000101111000000000;
assign LUT_1[50981] = 32'b11111111111111111111001001111100;
assign LUT_1[50982] = 32'b00000000000000000001100110010001;
assign LUT_1[50983] = 32'b11111111111111111010111000001101;
assign LUT_1[50984] = 32'b11111111111111111101001100011110;
assign LUT_1[50985] = 32'b11111111111111110110011110011010;
assign LUT_1[50986] = 32'b11111111111111111000111010101111;
assign LUT_1[50987] = 32'b11111111111111110010001100101011;
assign LUT_1[50988] = 32'b00000000000000000101000101110101;
assign LUT_1[50989] = 32'b11111111111111111110010111110001;
assign LUT_1[50990] = 32'b00000000000000000000110100000110;
assign LUT_1[50991] = 32'b11111111111111111010000110000010;
assign LUT_1[50992] = 32'b11111111111111111111111010001011;
assign LUT_1[50993] = 32'b11111111111111111001001100000111;
assign LUT_1[50994] = 32'b11111111111111111011101000011100;
assign LUT_1[50995] = 32'b11111111111111110100111010011000;
assign LUT_1[50996] = 32'b00000000000000000111110011100010;
assign LUT_1[50997] = 32'b00000000000000000001000101011110;
assign LUT_1[50998] = 32'b00000000000000000011100001110011;
assign LUT_1[50999] = 32'b11111111111111111100110011101111;
assign LUT_1[51000] = 32'b11111111111111111111001000000000;
assign LUT_1[51001] = 32'b11111111111111111000011001111100;
assign LUT_1[51002] = 32'b11111111111111111010110110010001;
assign LUT_1[51003] = 32'b11111111111111110100001000001101;
assign LUT_1[51004] = 32'b00000000000000000111000001010111;
assign LUT_1[51005] = 32'b00000000000000000000010011010011;
assign LUT_1[51006] = 32'b00000000000000000010101111101000;
assign LUT_1[51007] = 32'b11111111111111111100000001100100;
assign LUT_1[51008] = 32'b11111111111111111111000001010010;
assign LUT_1[51009] = 32'b11111111111111111000010011001110;
assign LUT_1[51010] = 32'b11111111111111111010101111100011;
assign LUT_1[51011] = 32'b11111111111111110100000001011111;
assign LUT_1[51012] = 32'b00000000000000000110111010101001;
assign LUT_1[51013] = 32'b00000000000000000000001100100101;
assign LUT_1[51014] = 32'b00000000000000000010101000111010;
assign LUT_1[51015] = 32'b11111111111111111011111010110110;
assign LUT_1[51016] = 32'b11111111111111111110001111000111;
assign LUT_1[51017] = 32'b11111111111111110111100001000011;
assign LUT_1[51018] = 32'b11111111111111111001111101011000;
assign LUT_1[51019] = 32'b11111111111111110011001111010100;
assign LUT_1[51020] = 32'b00000000000000000110001000011110;
assign LUT_1[51021] = 32'b11111111111111111111011010011010;
assign LUT_1[51022] = 32'b00000000000000000001110110101111;
assign LUT_1[51023] = 32'b11111111111111111011001000101011;
assign LUT_1[51024] = 32'b00000000000000000000111100110100;
assign LUT_1[51025] = 32'b11111111111111111010001110110000;
assign LUT_1[51026] = 32'b11111111111111111100101011000101;
assign LUT_1[51027] = 32'b11111111111111110101111101000001;
assign LUT_1[51028] = 32'b00000000000000001000110110001011;
assign LUT_1[51029] = 32'b00000000000000000010001000000111;
assign LUT_1[51030] = 32'b00000000000000000100100100011100;
assign LUT_1[51031] = 32'b11111111111111111101110110011000;
assign LUT_1[51032] = 32'b00000000000000000000001010101001;
assign LUT_1[51033] = 32'b11111111111111111001011100100101;
assign LUT_1[51034] = 32'b11111111111111111011111000111010;
assign LUT_1[51035] = 32'b11111111111111110101001010110110;
assign LUT_1[51036] = 32'b00000000000000001000000100000000;
assign LUT_1[51037] = 32'b00000000000000000001010101111100;
assign LUT_1[51038] = 32'b00000000000000000011110010010001;
assign LUT_1[51039] = 32'b11111111111111111101000100001101;
assign LUT_1[51040] = 32'b11111111111111111111111100010001;
assign LUT_1[51041] = 32'b11111111111111111001001110001101;
assign LUT_1[51042] = 32'b11111111111111111011101010100010;
assign LUT_1[51043] = 32'b11111111111111110100111100011110;
assign LUT_1[51044] = 32'b00000000000000000111110101101000;
assign LUT_1[51045] = 32'b00000000000000000001000111100100;
assign LUT_1[51046] = 32'b00000000000000000011100011111001;
assign LUT_1[51047] = 32'b11111111111111111100110101110101;
assign LUT_1[51048] = 32'b11111111111111111111001010000110;
assign LUT_1[51049] = 32'b11111111111111111000011100000010;
assign LUT_1[51050] = 32'b11111111111111111010111000010111;
assign LUT_1[51051] = 32'b11111111111111110100001010010011;
assign LUT_1[51052] = 32'b00000000000000000111000011011101;
assign LUT_1[51053] = 32'b00000000000000000000010101011001;
assign LUT_1[51054] = 32'b00000000000000000010110001101110;
assign LUT_1[51055] = 32'b11111111111111111100000011101010;
assign LUT_1[51056] = 32'b00000000000000000001110111110011;
assign LUT_1[51057] = 32'b11111111111111111011001001101111;
assign LUT_1[51058] = 32'b11111111111111111101100110000100;
assign LUT_1[51059] = 32'b11111111111111110110111000000000;
assign LUT_1[51060] = 32'b00000000000000001001110001001010;
assign LUT_1[51061] = 32'b00000000000000000011000011000110;
assign LUT_1[51062] = 32'b00000000000000000101011111011011;
assign LUT_1[51063] = 32'b11111111111111111110110001010111;
assign LUT_1[51064] = 32'b00000000000000000001000101101000;
assign LUT_1[51065] = 32'b11111111111111111010010111100100;
assign LUT_1[51066] = 32'b11111111111111111100110011111001;
assign LUT_1[51067] = 32'b11111111111111110110000101110101;
assign LUT_1[51068] = 32'b00000000000000001000111110111111;
assign LUT_1[51069] = 32'b00000000000000000010010000111011;
assign LUT_1[51070] = 32'b00000000000000000100101101010000;
assign LUT_1[51071] = 32'b11111111111111111101111111001100;
assign LUT_1[51072] = 32'b00000000000000000000000011101101;
assign LUT_1[51073] = 32'b11111111111111111001010101101001;
assign LUT_1[51074] = 32'b11111111111111111011110001111110;
assign LUT_1[51075] = 32'b11111111111111110101000011111010;
assign LUT_1[51076] = 32'b00000000000000000111111101000100;
assign LUT_1[51077] = 32'b00000000000000000001001111000000;
assign LUT_1[51078] = 32'b00000000000000000011101011010101;
assign LUT_1[51079] = 32'b11111111111111111100111101010001;
assign LUT_1[51080] = 32'b11111111111111111111010001100010;
assign LUT_1[51081] = 32'b11111111111111111000100011011110;
assign LUT_1[51082] = 32'b11111111111111111010111111110011;
assign LUT_1[51083] = 32'b11111111111111110100010001101111;
assign LUT_1[51084] = 32'b00000000000000000111001010111001;
assign LUT_1[51085] = 32'b00000000000000000000011100110101;
assign LUT_1[51086] = 32'b00000000000000000010111001001010;
assign LUT_1[51087] = 32'b11111111111111111100001011000110;
assign LUT_1[51088] = 32'b00000000000000000001111111001111;
assign LUT_1[51089] = 32'b11111111111111111011010001001011;
assign LUT_1[51090] = 32'b11111111111111111101101101100000;
assign LUT_1[51091] = 32'b11111111111111110110111111011100;
assign LUT_1[51092] = 32'b00000000000000001001111000100110;
assign LUT_1[51093] = 32'b00000000000000000011001010100010;
assign LUT_1[51094] = 32'b00000000000000000101100110110111;
assign LUT_1[51095] = 32'b11111111111111111110111000110011;
assign LUT_1[51096] = 32'b00000000000000000001001101000100;
assign LUT_1[51097] = 32'b11111111111111111010011111000000;
assign LUT_1[51098] = 32'b11111111111111111100111011010101;
assign LUT_1[51099] = 32'b11111111111111110110001101010001;
assign LUT_1[51100] = 32'b00000000000000001001000110011011;
assign LUT_1[51101] = 32'b00000000000000000010011000010111;
assign LUT_1[51102] = 32'b00000000000000000100110100101100;
assign LUT_1[51103] = 32'b11111111111111111110000110101000;
assign LUT_1[51104] = 32'b00000000000000000000111110101100;
assign LUT_1[51105] = 32'b11111111111111111010010000101000;
assign LUT_1[51106] = 32'b11111111111111111100101100111101;
assign LUT_1[51107] = 32'b11111111111111110101111110111001;
assign LUT_1[51108] = 32'b00000000000000001000111000000011;
assign LUT_1[51109] = 32'b00000000000000000010001001111111;
assign LUT_1[51110] = 32'b00000000000000000100100110010100;
assign LUT_1[51111] = 32'b11111111111111111101111000010000;
assign LUT_1[51112] = 32'b00000000000000000000001100100001;
assign LUT_1[51113] = 32'b11111111111111111001011110011101;
assign LUT_1[51114] = 32'b11111111111111111011111010110010;
assign LUT_1[51115] = 32'b11111111111111110101001100101110;
assign LUT_1[51116] = 32'b00000000000000001000000101111000;
assign LUT_1[51117] = 32'b00000000000000000001010111110100;
assign LUT_1[51118] = 32'b00000000000000000011110100001001;
assign LUT_1[51119] = 32'b11111111111111111101000110000101;
assign LUT_1[51120] = 32'b00000000000000000010111010001110;
assign LUT_1[51121] = 32'b11111111111111111100001100001010;
assign LUT_1[51122] = 32'b11111111111111111110101000011111;
assign LUT_1[51123] = 32'b11111111111111110111111010011011;
assign LUT_1[51124] = 32'b00000000000000001010110011100101;
assign LUT_1[51125] = 32'b00000000000000000100000101100001;
assign LUT_1[51126] = 32'b00000000000000000110100001110110;
assign LUT_1[51127] = 32'b11111111111111111111110011110010;
assign LUT_1[51128] = 32'b00000000000000000010001000000011;
assign LUT_1[51129] = 32'b11111111111111111011011001111111;
assign LUT_1[51130] = 32'b11111111111111111101110110010100;
assign LUT_1[51131] = 32'b11111111111111110111001000010000;
assign LUT_1[51132] = 32'b00000000000000001010000001011010;
assign LUT_1[51133] = 32'b00000000000000000011010011010110;
assign LUT_1[51134] = 32'b00000000000000000101101111101011;
assign LUT_1[51135] = 32'b11111111111111111111000001100111;
assign LUT_1[51136] = 32'b00000000000000000010000001010101;
assign LUT_1[51137] = 32'b11111111111111111011010011010001;
assign LUT_1[51138] = 32'b11111111111111111101101111100110;
assign LUT_1[51139] = 32'b11111111111111110111000001100010;
assign LUT_1[51140] = 32'b00000000000000001001111010101100;
assign LUT_1[51141] = 32'b00000000000000000011001100101000;
assign LUT_1[51142] = 32'b00000000000000000101101000111101;
assign LUT_1[51143] = 32'b11111111111111111110111010111001;
assign LUT_1[51144] = 32'b00000000000000000001001111001010;
assign LUT_1[51145] = 32'b11111111111111111010100001000110;
assign LUT_1[51146] = 32'b11111111111111111100111101011011;
assign LUT_1[51147] = 32'b11111111111111110110001111010111;
assign LUT_1[51148] = 32'b00000000000000001001001000100001;
assign LUT_1[51149] = 32'b00000000000000000010011010011101;
assign LUT_1[51150] = 32'b00000000000000000100110110110010;
assign LUT_1[51151] = 32'b11111111111111111110001000101110;
assign LUT_1[51152] = 32'b00000000000000000011111100110111;
assign LUT_1[51153] = 32'b11111111111111111101001110110011;
assign LUT_1[51154] = 32'b11111111111111111111101011001000;
assign LUT_1[51155] = 32'b11111111111111111000111101000100;
assign LUT_1[51156] = 32'b00000000000000001011110110001110;
assign LUT_1[51157] = 32'b00000000000000000101001000001010;
assign LUT_1[51158] = 32'b00000000000000000111100100011111;
assign LUT_1[51159] = 32'b00000000000000000000110110011011;
assign LUT_1[51160] = 32'b00000000000000000011001010101100;
assign LUT_1[51161] = 32'b11111111111111111100011100101000;
assign LUT_1[51162] = 32'b11111111111111111110111000111101;
assign LUT_1[51163] = 32'b11111111111111111000001010111001;
assign LUT_1[51164] = 32'b00000000000000001011000100000011;
assign LUT_1[51165] = 32'b00000000000000000100010101111111;
assign LUT_1[51166] = 32'b00000000000000000110110010010100;
assign LUT_1[51167] = 32'b00000000000000000000000100010000;
assign LUT_1[51168] = 32'b00000000000000000010111100010100;
assign LUT_1[51169] = 32'b11111111111111111100001110010000;
assign LUT_1[51170] = 32'b11111111111111111110101010100101;
assign LUT_1[51171] = 32'b11111111111111110111111100100001;
assign LUT_1[51172] = 32'b00000000000000001010110101101011;
assign LUT_1[51173] = 32'b00000000000000000100000111100111;
assign LUT_1[51174] = 32'b00000000000000000110100011111100;
assign LUT_1[51175] = 32'b11111111111111111111110101111000;
assign LUT_1[51176] = 32'b00000000000000000010001010001001;
assign LUT_1[51177] = 32'b11111111111111111011011100000101;
assign LUT_1[51178] = 32'b11111111111111111101111000011010;
assign LUT_1[51179] = 32'b11111111111111110111001010010110;
assign LUT_1[51180] = 32'b00000000000000001010000011100000;
assign LUT_1[51181] = 32'b00000000000000000011010101011100;
assign LUT_1[51182] = 32'b00000000000000000101110001110001;
assign LUT_1[51183] = 32'b11111111111111111111000011101101;
assign LUT_1[51184] = 32'b00000000000000000100110111110110;
assign LUT_1[51185] = 32'b11111111111111111110001001110010;
assign LUT_1[51186] = 32'b00000000000000000000100110000111;
assign LUT_1[51187] = 32'b11111111111111111001111000000011;
assign LUT_1[51188] = 32'b00000000000000001100110001001101;
assign LUT_1[51189] = 32'b00000000000000000110000011001001;
assign LUT_1[51190] = 32'b00000000000000001000011111011110;
assign LUT_1[51191] = 32'b00000000000000000001110001011010;
assign LUT_1[51192] = 32'b00000000000000000100000101101011;
assign LUT_1[51193] = 32'b11111111111111111101010111100111;
assign LUT_1[51194] = 32'b11111111111111111111110011111100;
assign LUT_1[51195] = 32'b11111111111111111001000101111000;
assign LUT_1[51196] = 32'b00000000000000001011111111000010;
assign LUT_1[51197] = 32'b00000000000000000101010000111110;
assign LUT_1[51198] = 32'b00000000000000000111101101010011;
assign LUT_1[51199] = 32'b00000000000000000000111111001111;
assign LUT_1[51200] = 32'b00000000000000000000001100001100;
assign LUT_1[51201] = 32'b11111111111111111001011110001000;
assign LUT_1[51202] = 32'b11111111111111111011111010011101;
assign LUT_1[51203] = 32'b11111111111111110101001100011001;
assign LUT_1[51204] = 32'b00000000000000001000000101100011;
assign LUT_1[51205] = 32'b00000000000000000001010111011111;
assign LUT_1[51206] = 32'b00000000000000000011110011110100;
assign LUT_1[51207] = 32'b11111111111111111101000101110000;
assign LUT_1[51208] = 32'b11111111111111111111011010000001;
assign LUT_1[51209] = 32'b11111111111111111000101011111101;
assign LUT_1[51210] = 32'b11111111111111111011001000010010;
assign LUT_1[51211] = 32'b11111111111111110100011010001110;
assign LUT_1[51212] = 32'b00000000000000000111010011011000;
assign LUT_1[51213] = 32'b00000000000000000000100101010100;
assign LUT_1[51214] = 32'b00000000000000000011000001101001;
assign LUT_1[51215] = 32'b11111111111111111100010011100101;
assign LUT_1[51216] = 32'b00000000000000000010000111101110;
assign LUT_1[51217] = 32'b11111111111111111011011001101010;
assign LUT_1[51218] = 32'b11111111111111111101110101111111;
assign LUT_1[51219] = 32'b11111111111111110111000111111011;
assign LUT_1[51220] = 32'b00000000000000001010000001000101;
assign LUT_1[51221] = 32'b00000000000000000011010011000001;
assign LUT_1[51222] = 32'b00000000000000000101101111010110;
assign LUT_1[51223] = 32'b11111111111111111111000001010010;
assign LUT_1[51224] = 32'b00000000000000000001010101100011;
assign LUT_1[51225] = 32'b11111111111111111010100111011111;
assign LUT_1[51226] = 32'b11111111111111111101000011110100;
assign LUT_1[51227] = 32'b11111111111111110110010101110000;
assign LUT_1[51228] = 32'b00000000000000001001001110111010;
assign LUT_1[51229] = 32'b00000000000000000010100000110110;
assign LUT_1[51230] = 32'b00000000000000000100111101001011;
assign LUT_1[51231] = 32'b11111111111111111110001111000111;
assign LUT_1[51232] = 32'b00000000000000000001000111001011;
assign LUT_1[51233] = 32'b11111111111111111010011001000111;
assign LUT_1[51234] = 32'b11111111111111111100110101011100;
assign LUT_1[51235] = 32'b11111111111111110110000111011000;
assign LUT_1[51236] = 32'b00000000000000001001000000100010;
assign LUT_1[51237] = 32'b00000000000000000010010010011110;
assign LUT_1[51238] = 32'b00000000000000000100101110110011;
assign LUT_1[51239] = 32'b11111111111111111110000000101111;
assign LUT_1[51240] = 32'b00000000000000000000010101000000;
assign LUT_1[51241] = 32'b11111111111111111001100110111100;
assign LUT_1[51242] = 32'b11111111111111111100000011010001;
assign LUT_1[51243] = 32'b11111111111111110101010101001101;
assign LUT_1[51244] = 32'b00000000000000001000001110010111;
assign LUT_1[51245] = 32'b00000000000000000001100000010011;
assign LUT_1[51246] = 32'b00000000000000000011111100101000;
assign LUT_1[51247] = 32'b11111111111111111101001110100100;
assign LUT_1[51248] = 32'b00000000000000000011000010101101;
assign LUT_1[51249] = 32'b11111111111111111100010100101001;
assign LUT_1[51250] = 32'b11111111111111111110110000111110;
assign LUT_1[51251] = 32'b11111111111111111000000010111010;
assign LUT_1[51252] = 32'b00000000000000001010111100000100;
assign LUT_1[51253] = 32'b00000000000000000100001110000000;
assign LUT_1[51254] = 32'b00000000000000000110101010010101;
assign LUT_1[51255] = 32'b11111111111111111111111100010001;
assign LUT_1[51256] = 32'b00000000000000000010010000100010;
assign LUT_1[51257] = 32'b11111111111111111011100010011110;
assign LUT_1[51258] = 32'b11111111111111111101111110110011;
assign LUT_1[51259] = 32'b11111111111111110111010000101111;
assign LUT_1[51260] = 32'b00000000000000001010001001111001;
assign LUT_1[51261] = 32'b00000000000000000011011011110101;
assign LUT_1[51262] = 32'b00000000000000000101111000001010;
assign LUT_1[51263] = 32'b11111111111111111111001010000110;
assign LUT_1[51264] = 32'b00000000000000000010001001110100;
assign LUT_1[51265] = 32'b11111111111111111011011011110000;
assign LUT_1[51266] = 32'b11111111111111111101111000000101;
assign LUT_1[51267] = 32'b11111111111111110111001010000001;
assign LUT_1[51268] = 32'b00000000000000001010000011001011;
assign LUT_1[51269] = 32'b00000000000000000011010101000111;
assign LUT_1[51270] = 32'b00000000000000000101110001011100;
assign LUT_1[51271] = 32'b11111111111111111111000011011000;
assign LUT_1[51272] = 32'b00000000000000000001010111101001;
assign LUT_1[51273] = 32'b11111111111111111010101001100101;
assign LUT_1[51274] = 32'b11111111111111111101000101111010;
assign LUT_1[51275] = 32'b11111111111111110110010111110110;
assign LUT_1[51276] = 32'b00000000000000001001010001000000;
assign LUT_1[51277] = 32'b00000000000000000010100010111100;
assign LUT_1[51278] = 32'b00000000000000000100111111010001;
assign LUT_1[51279] = 32'b11111111111111111110010001001101;
assign LUT_1[51280] = 32'b00000000000000000100000101010110;
assign LUT_1[51281] = 32'b11111111111111111101010111010010;
assign LUT_1[51282] = 32'b11111111111111111111110011100111;
assign LUT_1[51283] = 32'b11111111111111111001000101100011;
assign LUT_1[51284] = 32'b00000000000000001011111110101101;
assign LUT_1[51285] = 32'b00000000000000000101010000101001;
assign LUT_1[51286] = 32'b00000000000000000111101100111110;
assign LUT_1[51287] = 32'b00000000000000000000111110111010;
assign LUT_1[51288] = 32'b00000000000000000011010011001011;
assign LUT_1[51289] = 32'b11111111111111111100100101000111;
assign LUT_1[51290] = 32'b11111111111111111111000001011100;
assign LUT_1[51291] = 32'b11111111111111111000010011011000;
assign LUT_1[51292] = 32'b00000000000000001011001100100010;
assign LUT_1[51293] = 32'b00000000000000000100011110011110;
assign LUT_1[51294] = 32'b00000000000000000110111010110011;
assign LUT_1[51295] = 32'b00000000000000000000001100101111;
assign LUT_1[51296] = 32'b00000000000000000011000100110011;
assign LUT_1[51297] = 32'b11111111111111111100010110101111;
assign LUT_1[51298] = 32'b11111111111111111110110011000100;
assign LUT_1[51299] = 32'b11111111111111111000000101000000;
assign LUT_1[51300] = 32'b00000000000000001010111110001010;
assign LUT_1[51301] = 32'b00000000000000000100010000000110;
assign LUT_1[51302] = 32'b00000000000000000110101100011011;
assign LUT_1[51303] = 32'b11111111111111111111111110010111;
assign LUT_1[51304] = 32'b00000000000000000010010010101000;
assign LUT_1[51305] = 32'b11111111111111111011100100100100;
assign LUT_1[51306] = 32'b11111111111111111110000000111001;
assign LUT_1[51307] = 32'b11111111111111110111010010110101;
assign LUT_1[51308] = 32'b00000000000000001010001011111111;
assign LUT_1[51309] = 32'b00000000000000000011011101111011;
assign LUT_1[51310] = 32'b00000000000000000101111010010000;
assign LUT_1[51311] = 32'b11111111111111111111001100001100;
assign LUT_1[51312] = 32'b00000000000000000101000000010101;
assign LUT_1[51313] = 32'b11111111111111111110010010010001;
assign LUT_1[51314] = 32'b00000000000000000000101110100110;
assign LUT_1[51315] = 32'b11111111111111111010000000100010;
assign LUT_1[51316] = 32'b00000000000000001100111001101100;
assign LUT_1[51317] = 32'b00000000000000000110001011101000;
assign LUT_1[51318] = 32'b00000000000000001000100111111101;
assign LUT_1[51319] = 32'b00000000000000000001111001111001;
assign LUT_1[51320] = 32'b00000000000000000100001110001010;
assign LUT_1[51321] = 32'b11111111111111111101100000000110;
assign LUT_1[51322] = 32'b11111111111111111111111100011011;
assign LUT_1[51323] = 32'b11111111111111111001001110010111;
assign LUT_1[51324] = 32'b00000000000000001100000111100001;
assign LUT_1[51325] = 32'b00000000000000000101011001011101;
assign LUT_1[51326] = 32'b00000000000000000111110101110010;
assign LUT_1[51327] = 32'b00000000000000000001000111101110;
assign LUT_1[51328] = 32'b00000000000000000011001100001111;
assign LUT_1[51329] = 32'b11111111111111111100011110001011;
assign LUT_1[51330] = 32'b11111111111111111110111010100000;
assign LUT_1[51331] = 32'b11111111111111111000001100011100;
assign LUT_1[51332] = 32'b00000000000000001011000101100110;
assign LUT_1[51333] = 32'b00000000000000000100010111100010;
assign LUT_1[51334] = 32'b00000000000000000110110011110111;
assign LUT_1[51335] = 32'b00000000000000000000000101110011;
assign LUT_1[51336] = 32'b00000000000000000010011010000100;
assign LUT_1[51337] = 32'b11111111111111111011101100000000;
assign LUT_1[51338] = 32'b11111111111111111110001000010101;
assign LUT_1[51339] = 32'b11111111111111110111011010010001;
assign LUT_1[51340] = 32'b00000000000000001010010011011011;
assign LUT_1[51341] = 32'b00000000000000000011100101010111;
assign LUT_1[51342] = 32'b00000000000000000110000001101100;
assign LUT_1[51343] = 32'b11111111111111111111010011101000;
assign LUT_1[51344] = 32'b00000000000000000101000111110001;
assign LUT_1[51345] = 32'b11111111111111111110011001101101;
assign LUT_1[51346] = 32'b00000000000000000000110110000010;
assign LUT_1[51347] = 32'b11111111111111111010000111111110;
assign LUT_1[51348] = 32'b00000000000000001101000001001000;
assign LUT_1[51349] = 32'b00000000000000000110010011000100;
assign LUT_1[51350] = 32'b00000000000000001000101111011001;
assign LUT_1[51351] = 32'b00000000000000000010000001010101;
assign LUT_1[51352] = 32'b00000000000000000100010101100110;
assign LUT_1[51353] = 32'b11111111111111111101100111100010;
assign LUT_1[51354] = 32'b00000000000000000000000011110111;
assign LUT_1[51355] = 32'b11111111111111111001010101110011;
assign LUT_1[51356] = 32'b00000000000000001100001110111101;
assign LUT_1[51357] = 32'b00000000000000000101100000111001;
assign LUT_1[51358] = 32'b00000000000000000111111101001110;
assign LUT_1[51359] = 32'b00000000000000000001001111001010;
assign LUT_1[51360] = 32'b00000000000000000100000111001110;
assign LUT_1[51361] = 32'b11111111111111111101011001001010;
assign LUT_1[51362] = 32'b11111111111111111111110101011111;
assign LUT_1[51363] = 32'b11111111111111111001000111011011;
assign LUT_1[51364] = 32'b00000000000000001100000000100101;
assign LUT_1[51365] = 32'b00000000000000000101010010100001;
assign LUT_1[51366] = 32'b00000000000000000111101110110110;
assign LUT_1[51367] = 32'b00000000000000000001000000110010;
assign LUT_1[51368] = 32'b00000000000000000011010101000011;
assign LUT_1[51369] = 32'b11111111111111111100100110111111;
assign LUT_1[51370] = 32'b11111111111111111111000011010100;
assign LUT_1[51371] = 32'b11111111111111111000010101010000;
assign LUT_1[51372] = 32'b00000000000000001011001110011010;
assign LUT_1[51373] = 32'b00000000000000000100100000010110;
assign LUT_1[51374] = 32'b00000000000000000110111100101011;
assign LUT_1[51375] = 32'b00000000000000000000001110100111;
assign LUT_1[51376] = 32'b00000000000000000110000010110000;
assign LUT_1[51377] = 32'b11111111111111111111010100101100;
assign LUT_1[51378] = 32'b00000000000000000001110001000001;
assign LUT_1[51379] = 32'b11111111111111111011000010111101;
assign LUT_1[51380] = 32'b00000000000000001101111100000111;
assign LUT_1[51381] = 32'b00000000000000000111001110000011;
assign LUT_1[51382] = 32'b00000000000000001001101010011000;
assign LUT_1[51383] = 32'b00000000000000000010111100010100;
assign LUT_1[51384] = 32'b00000000000000000101010000100101;
assign LUT_1[51385] = 32'b11111111111111111110100010100001;
assign LUT_1[51386] = 32'b00000000000000000000111110110110;
assign LUT_1[51387] = 32'b11111111111111111010010000110010;
assign LUT_1[51388] = 32'b00000000000000001101001001111100;
assign LUT_1[51389] = 32'b00000000000000000110011011111000;
assign LUT_1[51390] = 32'b00000000000000001000111000001101;
assign LUT_1[51391] = 32'b00000000000000000010001010001001;
assign LUT_1[51392] = 32'b00000000000000000101001001110111;
assign LUT_1[51393] = 32'b11111111111111111110011011110011;
assign LUT_1[51394] = 32'b00000000000000000000111000001000;
assign LUT_1[51395] = 32'b11111111111111111010001010000100;
assign LUT_1[51396] = 32'b00000000000000001101000011001110;
assign LUT_1[51397] = 32'b00000000000000000110010101001010;
assign LUT_1[51398] = 32'b00000000000000001000110001011111;
assign LUT_1[51399] = 32'b00000000000000000010000011011011;
assign LUT_1[51400] = 32'b00000000000000000100010111101100;
assign LUT_1[51401] = 32'b11111111111111111101101001101000;
assign LUT_1[51402] = 32'b00000000000000000000000101111101;
assign LUT_1[51403] = 32'b11111111111111111001010111111001;
assign LUT_1[51404] = 32'b00000000000000001100010001000011;
assign LUT_1[51405] = 32'b00000000000000000101100010111111;
assign LUT_1[51406] = 32'b00000000000000000111111111010100;
assign LUT_1[51407] = 32'b00000000000000000001010001010000;
assign LUT_1[51408] = 32'b00000000000000000111000101011001;
assign LUT_1[51409] = 32'b00000000000000000000010111010101;
assign LUT_1[51410] = 32'b00000000000000000010110011101010;
assign LUT_1[51411] = 32'b11111111111111111100000101100110;
assign LUT_1[51412] = 32'b00000000000000001110111110110000;
assign LUT_1[51413] = 32'b00000000000000001000010000101100;
assign LUT_1[51414] = 32'b00000000000000001010101101000001;
assign LUT_1[51415] = 32'b00000000000000000011111110111101;
assign LUT_1[51416] = 32'b00000000000000000110010011001110;
assign LUT_1[51417] = 32'b11111111111111111111100101001010;
assign LUT_1[51418] = 32'b00000000000000000010000001011111;
assign LUT_1[51419] = 32'b11111111111111111011010011011011;
assign LUT_1[51420] = 32'b00000000000000001110001100100101;
assign LUT_1[51421] = 32'b00000000000000000111011110100001;
assign LUT_1[51422] = 32'b00000000000000001001111010110110;
assign LUT_1[51423] = 32'b00000000000000000011001100110010;
assign LUT_1[51424] = 32'b00000000000000000110000100110110;
assign LUT_1[51425] = 32'b11111111111111111111010110110010;
assign LUT_1[51426] = 32'b00000000000000000001110011000111;
assign LUT_1[51427] = 32'b11111111111111111011000101000011;
assign LUT_1[51428] = 32'b00000000000000001101111110001101;
assign LUT_1[51429] = 32'b00000000000000000111010000001001;
assign LUT_1[51430] = 32'b00000000000000001001101100011110;
assign LUT_1[51431] = 32'b00000000000000000010111110011010;
assign LUT_1[51432] = 32'b00000000000000000101010010101011;
assign LUT_1[51433] = 32'b11111111111111111110100100100111;
assign LUT_1[51434] = 32'b00000000000000000001000000111100;
assign LUT_1[51435] = 32'b11111111111111111010010010111000;
assign LUT_1[51436] = 32'b00000000000000001101001100000010;
assign LUT_1[51437] = 32'b00000000000000000110011101111110;
assign LUT_1[51438] = 32'b00000000000000001000111010010011;
assign LUT_1[51439] = 32'b00000000000000000010001100001111;
assign LUT_1[51440] = 32'b00000000000000001000000000011000;
assign LUT_1[51441] = 32'b00000000000000000001010010010100;
assign LUT_1[51442] = 32'b00000000000000000011101110101001;
assign LUT_1[51443] = 32'b11111111111111111101000000100101;
assign LUT_1[51444] = 32'b00000000000000001111111001101111;
assign LUT_1[51445] = 32'b00000000000000001001001011101011;
assign LUT_1[51446] = 32'b00000000000000001011101000000000;
assign LUT_1[51447] = 32'b00000000000000000100111001111100;
assign LUT_1[51448] = 32'b00000000000000000111001110001101;
assign LUT_1[51449] = 32'b00000000000000000000100000001001;
assign LUT_1[51450] = 32'b00000000000000000010111100011110;
assign LUT_1[51451] = 32'b11111111111111111100001110011010;
assign LUT_1[51452] = 32'b00000000000000001111000111100100;
assign LUT_1[51453] = 32'b00000000000000001000011001100000;
assign LUT_1[51454] = 32'b00000000000000001010110101110101;
assign LUT_1[51455] = 32'b00000000000000000100000111110001;
assign LUT_1[51456] = 32'b11111111111111111110000000011000;
assign LUT_1[51457] = 32'b11111111111111110111010010010100;
assign LUT_1[51458] = 32'b11111111111111111001101110101001;
assign LUT_1[51459] = 32'b11111111111111110011000000100101;
assign LUT_1[51460] = 32'b00000000000000000101111001101111;
assign LUT_1[51461] = 32'b11111111111111111111001011101011;
assign LUT_1[51462] = 32'b00000000000000000001101000000000;
assign LUT_1[51463] = 32'b11111111111111111010111001111100;
assign LUT_1[51464] = 32'b11111111111111111101001110001101;
assign LUT_1[51465] = 32'b11111111111111110110100000001001;
assign LUT_1[51466] = 32'b11111111111111111000111100011110;
assign LUT_1[51467] = 32'b11111111111111110010001110011010;
assign LUT_1[51468] = 32'b00000000000000000101000111100100;
assign LUT_1[51469] = 32'b11111111111111111110011001100000;
assign LUT_1[51470] = 32'b00000000000000000000110101110101;
assign LUT_1[51471] = 32'b11111111111111111010000111110001;
assign LUT_1[51472] = 32'b11111111111111111111111011111010;
assign LUT_1[51473] = 32'b11111111111111111001001101110110;
assign LUT_1[51474] = 32'b11111111111111111011101010001011;
assign LUT_1[51475] = 32'b11111111111111110100111100000111;
assign LUT_1[51476] = 32'b00000000000000000111110101010001;
assign LUT_1[51477] = 32'b00000000000000000001000111001101;
assign LUT_1[51478] = 32'b00000000000000000011100011100010;
assign LUT_1[51479] = 32'b11111111111111111100110101011110;
assign LUT_1[51480] = 32'b11111111111111111111001001101111;
assign LUT_1[51481] = 32'b11111111111111111000011011101011;
assign LUT_1[51482] = 32'b11111111111111111010111000000000;
assign LUT_1[51483] = 32'b11111111111111110100001001111100;
assign LUT_1[51484] = 32'b00000000000000000111000011000110;
assign LUT_1[51485] = 32'b00000000000000000000010101000010;
assign LUT_1[51486] = 32'b00000000000000000010110001010111;
assign LUT_1[51487] = 32'b11111111111111111100000011010011;
assign LUT_1[51488] = 32'b11111111111111111110111011010111;
assign LUT_1[51489] = 32'b11111111111111111000001101010011;
assign LUT_1[51490] = 32'b11111111111111111010101001101000;
assign LUT_1[51491] = 32'b11111111111111110011111011100100;
assign LUT_1[51492] = 32'b00000000000000000110110100101110;
assign LUT_1[51493] = 32'b00000000000000000000000110101010;
assign LUT_1[51494] = 32'b00000000000000000010100010111111;
assign LUT_1[51495] = 32'b11111111111111111011110100111011;
assign LUT_1[51496] = 32'b11111111111111111110001001001100;
assign LUT_1[51497] = 32'b11111111111111110111011011001000;
assign LUT_1[51498] = 32'b11111111111111111001110111011101;
assign LUT_1[51499] = 32'b11111111111111110011001001011001;
assign LUT_1[51500] = 32'b00000000000000000110000010100011;
assign LUT_1[51501] = 32'b11111111111111111111010100011111;
assign LUT_1[51502] = 32'b00000000000000000001110000110100;
assign LUT_1[51503] = 32'b11111111111111111011000010110000;
assign LUT_1[51504] = 32'b00000000000000000000110110111001;
assign LUT_1[51505] = 32'b11111111111111111010001000110101;
assign LUT_1[51506] = 32'b11111111111111111100100101001010;
assign LUT_1[51507] = 32'b11111111111111110101110111000110;
assign LUT_1[51508] = 32'b00000000000000001000110000010000;
assign LUT_1[51509] = 32'b00000000000000000010000010001100;
assign LUT_1[51510] = 32'b00000000000000000100011110100001;
assign LUT_1[51511] = 32'b11111111111111111101110000011101;
assign LUT_1[51512] = 32'b00000000000000000000000100101110;
assign LUT_1[51513] = 32'b11111111111111111001010110101010;
assign LUT_1[51514] = 32'b11111111111111111011110010111111;
assign LUT_1[51515] = 32'b11111111111111110101000100111011;
assign LUT_1[51516] = 32'b00000000000000000111111110000101;
assign LUT_1[51517] = 32'b00000000000000000001010000000001;
assign LUT_1[51518] = 32'b00000000000000000011101100010110;
assign LUT_1[51519] = 32'b11111111111111111100111110010010;
assign LUT_1[51520] = 32'b11111111111111111111111110000000;
assign LUT_1[51521] = 32'b11111111111111111001001111111100;
assign LUT_1[51522] = 32'b11111111111111111011101100010001;
assign LUT_1[51523] = 32'b11111111111111110100111110001101;
assign LUT_1[51524] = 32'b00000000000000000111110111010111;
assign LUT_1[51525] = 32'b00000000000000000001001001010011;
assign LUT_1[51526] = 32'b00000000000000000011100101101000;
assign LUT_1[51527] = 32'b11111111111111111100110111100100;
assign LUT_1[51528] = 32'b11111111111111111111001011110101;
assign LUT_1[51529] = 32'b11111111111111111000011101110001;
assign LUT_1[51530] = 32'b11111111111111111010111010000110;
assign LUT_1[51531] = 32'b11111111111111110100001100000010;
assign LUT_1[51532] = 32'b00000000000000000111000101001100;
assign LUT_1[51533] = 32'b00000000000000000000010111001000;
assign LUT_1[51534] = 32'b00000000000000000010110011011101;
assign LUT_1[51535] = 32'b11111111111111111100000101011001;
assign LUT_1[51536] = 32'b00000000000000000001111001100010;
assign LUT_1[51537] = 32'b11111111111111111011001011011110;
assign LUT_1[51538] = 32'b11111111111111111101100111110011;
assign LUT_1[51539] = 32'b11111111111111110110111001101111;
assign LUT_1[51540] = 32'b00000000000000001001110010111001;
assign LUT_1[51541] = 32'b00000000000000000011000100110101;
assign LUT_1[51542] = 32'b00000000000000000101100001001010;
assign LUT_1[51543] = 32'b11111111111111111110110011000110;
assign LUT_1[51544] = 32'b00000000000000000001000111010111;
assign LUT_1[51545] = 32'b11111111111111111010011001010011;
assign LUT_1[51546] = 32'b11111111111111111100110101101000;
assign LUT_1[51547] = 32'b11111111111111110110000111100100;
assign LUT_1[51548] = 32'b00000000000000001001000000101110;
assign LUT_1[51549] = 32'b00000000000000000010010010101010;
assign LUT_1[51550] = 32'b00000000000000000100101110111111;
assign LUT_1[51551] = 32'b11111111111111111110000000111011;
assign LUT_1[51552] = 32'b00000000000000000000111000111111;
assign LUT_1[51553] = 32'b11111111111111111010001010111011;
assign LUT_1[51554] = 32'b11111111111111111100100111010000;
assign LUT_1[51555] = 32'b11111111111111110101111001001100;
assign LUT_1[51556] = 32'b00000000000000001000110010010110;
assign LUT_1[51557] = 32'b00000000000000000010000100010010;
assign LUT_1[51558] = 32'b00000000000000000100100000100111;
assign LUT_1[51559] = 32'b11111111111111111101110010100011;
assign LUT_1[51560] = 32'b00000000000000000000000110110100;
assign LUT_1[51561] = 32'b11111111111111111001011000110000;
assign LUT_1[51562] = 32'b11111111111111111011110101000101;
assign LUT_1[51563] = 32'b11111111111111110101000111000001;
assign LUT_1[51564] = 32'b00000000000000001000000000001011;
assign LUT_1[51565] = 32'b00000000000000000001010010000111;
assign LUT_1[51566] = 32'b00000000000000000011101110011100;
assign LUT_1[51567] = 32'b11111111111111111101000000011000;
assign LUT_1[51568] = 32'b00000000000000000010110100100001;
assign LUT_1[51569] = 32'b11111111111111111100000110011101;
assign LUT_1[51570] = 32'b11111111111111111110100010110010;
assign LUT_1[51571] = 32'b11111111111111110111110100101110;
assign LUT_1[51572] = 32'b00000000000000001010101101111000;
assign LUT_1[51573] = 32'b00000000000000000011111111110100;
assign LUT_1[51574] = 32'b00000000000000000110011100001001;
assign LUT_1[51575] = 32'b11111111111111111111101110000101;
assign LUT_1[51576] = 32'b00000000000000000010000010010110;
assign LUT_1[51577] = 32'b11111111111111111011010100010010;
assign LUT_1[51578] = 32'b11111111111111111101110000100111;
assign LUT_1[51579] = 32'b11111111111111110111000010100011;
assign LUT_1[51580] = 32'b00000000000000001001111011101101;
assign LUT_1[51581] = 32'b00000000000000000011001101101001;
assign LUT_1[51582] = 32'b00000000000000000101101001111110;
assign LUT_1[51583] = 32'b11111111111111111110111011111010;
assign LUT_1[51584] = 32'b00000000000000000001000000011011;
assign LUT_1[51585] = 32'b11111111111111111010010010010111;
assign LUT_1[51586] = 32'b11111111111111111100101110101100;
assign LUT_1[51587] = 32'b11111111111111110110000000101000;
assign LUT_1[51588] = 32'b00000000000000001000111001110010;
assign LUT_1[51589] = 32'b00000000000000000010001011101110;
assign LUT_1[51590] = 32'b00000000000000000100101000000011;
assign LUT_1[51591] = 32'b11111111111111111101111001111111;
assign LUT_1[51592] = 32'b00000000000000000000001110010000;
assign LUT_1[51593] = 32'b11111111111111111001100000001100;
assign LUT_1[51594] = 32'b11111111111111111011111100100001;
assign LUT_1[51595] = 32'b11111111111111110101001110011101;
assign LUT_1[51596] = 32'b00000000000000001000000111100111;
assign LUT_1[51597] = 32'b00000000000000000001011001100011;
assign LUT_1[51598] = 32'b00000000000000000011110101111000;
assign LUT_1[51599] = 32'b11111111111111111101000111110100;
assign LUT_1[51600] = 32'b00000000000000000010111011111101;
assign LUT_1[51601] = 32'b11111111111111111100001101111001;
assign LUT_1[51602] = 32'b11111111111111111110101010001110;
assign LUT_1[51603] = 32'b11111111111111110111111100001010;
assign LUT_1[51604] = 32'b00000000000000001010110101010100;
assign LUT_1[51605] = 32'b00000000000000000100000111010000;
assign LUT_1[51606] = 32'b00000000000000000110100011100101;
assign LUT_1[51607] = 32'b11111111111111111111110101100001;
assign LUT_1[51608] = 32'b00000000000000000010001001110010;
assign LUT_1[51609] = 32'b11111111111111111011011011101110;
assign LUT_1[51610] = 32'b11111111111111111101111000000011;
assign LUT_1[51611] = 32'b11111111111111110111001001111111;
assign LUT_1[51612] = 32'b00000000000000001010000011001001;
assign LUT_1[51613] = 32'b00000000000000000011010101000101;
assign LUT_1[51614] = 32'b00000000000000000101110001011010;
assign LUT_1[51615] = 32'b11111111111111111111000011010110;
assign LUT_1[51616] = 32'b00000000000000000001111011011010;
assign LUT_1[51617] = 32'b11111111111111111011001101010110;
assign LUT_1[51618] = 32'b11111111111111111101101001101011;
assign LUT_1[51619] = 32'b11111111111111110110111011100111;
assign LUT_1[51620] = 32'b00000000000000001001110100110001;
assign LUT_1[51621] = 32'b00000000000000000011000110101101;
assign LUT_1[51622] = 32'b00000000000000000101100011000010;
assign LUT_1[51623] = 32'b11111111111111111110110100111110;
assign LUT_1[51624] = 32'b00000000000000000001001001001111;
assign LUT_1[51625] = 32'b11111111111111111010011011001011;
assign LUT_1[51626] = 32'b11111111111111111100110111100000;
assign LUT_1[51627] = 32'b11111111111111110110001001011100;
assign LUT_1[51628] = 32'b00000000000000001001000010100110;
assign LUT_1[51629] = 32'b00000000000000000010010100100010;
assign LUT_1[51630] = 32'b00000000000000000100110000110111;
assign LUT_1[51631] = 32'b11111111111111111110000010110011;
assign LUT_1[51632] = 32'b00000000000000000011110110111100;
assign LUT_1[51633] = 32'b11111111111111111101001000111000;
assign LUT_1[51634] = 32'b11111111111111111111100101001101;
assign LUT_1[51635] = 32'b11111111111111111000110111001001;
assign LUT_1[51636] = 32'b00000000000000001011110000010011;
assign LUT_1[51637] = 32'b00000000000000000101000010001111;
assign LUT_1[51638] = 32'b00000000000000000111011110100100;
assign LUT_1[51639] = 32'b00000000000000000000110000100000;
assign LUT_1[51640] = 32'b00000000000000000011000100110001;
assign LUT_1[51641] = 32'b11111111111111111100010110101101;
assign LUT_1[51642] = 32'b11111111111111111110110011000010;
assign LUT_1[51643] = 32'b11111111111111111000000100111110;
assign LUT_1[51644] = 32'b00000000000000001010111110001000;
assign LUT_1[51645] = 32'b00000000000000000100010000000100;
assign LUT_1[51646] = 32'b00000000000000000110101100011001;
assign LUT_1[51647] = 32'b11111111111111111111111110010101;
assign LUT_1[51648] = 32'b00000000000000000010111110000011;
assign LUT_1[51649] = 32'b11111111111111111100001111111111;
assign LUT_1[51650] = 32'b11111111111111111110101100010100;
assign LUT_1[51651] = 32'b11111111111111110111111110010000;
assign LUT_1[51652] = 32'b00000000000000001010110111011010;
assign LUT_1[51653] = 32'b00000000000000000100001001010110;
assign LUT_1[51654] = 32'b00000000000000000110100101101011;
assign LUT_1[51655] = 32'b11111111111111111111110111100111;
assign LUT_1[51656] = 32'b00000000000000000010001011111000;
assign LUT_1[51657] = 32'b11111111111111111011011101110100;
assign LUT_1[51658] = 32'b11111111111111111101111010001001;
assign LUT_1[51659] = 32'b11111111111111110111001100000101;
assign LUT_1[51660] = 32'b00000000000000001010000101001111;
assign LUT_1[51661] = 32'b00000000000000000011010111001011;
assign LUT_1[51662] = 32'b00000000000000000101110011100000;
assign LUT_1[51663] = 32'b11111111111111111111000101011100;
assign LUT_1[51664] = 32'b00000000000000000100111001100101;
assign LUT_1[51665] = 32'b11111111111111111110001011100001;
assign LUT_1[51666] = 32'b00000000000000000000100111110110;
assign LUT_1[51667] = 32'b11111111111111111001111001110010;
assign LUT_1[51668] = 32'b00000000000000001100110010111100;
assign LUT_1[51669] = 32'b00000000000000000110000100111000;
assign LUT_1[51670] = 32'b00000000000000001000100001001101;
assign LUT_1[51671] = 32'b00000000000000000001110011001001;
assign LUT_1[51672] = 32'b00000000000000000100000111011010;
assign LUT_1[51673] = 32'b11111111111111111101011001010110;
assign LUT_1[51674] = 32'b11111111111111111111110101101011;
assign LUT_1[51675] = 32'b11111111111111111001000111100111;
assign LUT_1[51676] = 32'b00000000000000001100000000110001;
assign LUT_1[51677] = 32'b00000000000000000101010010101101;
assign LUT_1[51678] = 32'b00000000000000000111101111000010;
assign LUT_1[51679] = 32'b00000000000000000001000000111110;
assign LUT_1[51680] = 32'b00000000000000000011111001000010;
assign LUT_1[51681] = 32'b11111111111111111101001010111110;
assign LUT_1[51682] = 32'b11111111111111111111100111010011;
assign LUT_1[51683] = 32'b11111111111111111000111001001111;
assign LUT_1[51684] = 32'b00000000000000001011110010011001;
assign LUT_1[51685] = 32'b00000000000000000101000100010101;
assign LUT_1[51686] = 32'b00000000000000000111100000101010;
assign LUT_1[51687] = 32'b00000000000000000000110010100110;
assign LUT_1[51688] = 32'b00000000000000000011000110110111;
assign LUT_1[51689] = 32'b11111111111111111100011000110011;
assign LUT_1[51690] = 32'b11111111111111111110110101001000;
assign LUT_1[51691] = 32'b11111111111111111000000111000100;
assign LUT_1[51692] = 32'b00000000000000001011000000001110;
assign LUT_1[51693] = 32'b00000000000000000100010010001010;
assign LUT_1[51694] = 32'b00000000000000000110101110011111;
assign LUT_1[51695] = 32'b00000000000000000000000000011011;
assign LUT_1[51696] = 32'b00000000000000000101110100100100;
assign LUT_1[51697] = 32'b11111111111111111111000110100000;
assign LUT_1[51698] = 32'b00000000000000000001100010110101;
assign LUT_1[51699] = 32'b11111111111111111010110100110001;
assign LUT_1[51700] = 32'b00000000000000001101101101111011;
assign LUT_1[51701] = 32'b00000000000000000110111111110111;
assign LUT_1[51702] = 32'b00000000000000001001011100001100;
assign LUT_1[51703] = 32'b00000000000000000010101110001000;
assign LUT_1[51704] = 32'b00000000000000000101000010011001;
assign LUT_1[51705] = 32'b11111111111111111110010100010101;
assign LUT_1[51706] = 32'b00000000000000000000110000101010;
assign LUT_1[51707] = 32'b11111111111111111010000010100110;
assign LUT_1[51708] = 32'b00000000000000001100111011110000;
assign LUT_1[51709] = 32'b00000000000000000110001101101100;
assign LUT_1[51710] = 32'b00000000000000001000101010000001;
assign LUT_1[51711] = 32'b00000000000000000001111011111101;
assign LUT_1[51712] = 32'b11111111111111111001111010101001;
assign LUT_1[51713] = 32'b11111111111111110011001100100101;
assign LUT_1[51714] = 32'b11111111111111110101101000111010;
assign LUT_1[51715] = 32'b11111111111111101110111010110110;
assign LUT_1[51716] = 32'b00000000000000000001110100000000;
assign LUT_1[51717] = 32'b11111111111111111011000101111100;
assign LUT_1[51718] = 32'b11111111111111111101100010010001;
assign LUT_1[51719] = 32'b11111111111111110110110100001101;
assign LUT_1[51720] = 32'b11111111111111111001001000011110;
assign LUT_1[51721] = 32'b11111111111111110010011010011010;
assign LUT_1[51722] = 32'b11111111111111110100110110101111;
assign LUT_1[51723] = 32'b11111111111111101110001000101011;
assign LUT_1[51724] = 32'b00000000000000000001000001110101;
assign LUT_1[51725] = 32'b11111111111111111010010011110001;
assign LUT_1[51726] = 32'b11111111111111111100110000000110;
assign LUT_1[51727] = 32'b11111111111111110110000010000010;
assign LUT_1[51728] = 32'b11111111111111111011110110001011;
assign LUT_1[51729] = 32'b11111111111111110101001000000111;
assign LUT_1[51730] = 32'b11111111111111110111100100011100;
assign LUT_1[51731] = 32'b11111111111111110000110110011000;
assign LUT_1[51732] = 32'b00000000000000000011101111100010;
assign LUT_1[51733] = 32'b11111111111111111101000001011110;
assign LUT_1[51734] = 32'b11111111111111111111011101110011;
assign LUT_1[51735] = 32'b11111111111111111000101111101111;
assign LUT_1[51736] = 32'b11111111111111111011000100000000;
assign LUT_1[51737] = 32'b11111111111111110100010101111100;
assign LUT_1[51738] = 32'b11111111111111110110110010010001;
assign LUT_1[51739] = 32'b11111111111111110000000100001101;
assign LUT_1[51740] = 32'b00000000000000000010111101010111;
assign LUT_1[51741] = 32'b11111111111111111100001111010011;
assign LUT_1[51742] = 32'b11111111111111111110101011101000;
assign LUT_1[51743] = 32'b11111111111111110111111101100100;
assign LUT_1[51744] = 32'b11111111111111111010110101101000;
assign LUT_1[51745] = 32'b11111111111111110100000111100100;
assign LUT_1[51746] = 32'b11111111111111110110100011111001;
assign LUT_1[51747] = 32'b11111111111111101111110101110101;
assign LUT_1[51748] = 32'b00000000000000000010101110111111;
assign LUT_1[51749] = 32'b11111111111111111100000000111011;
assign LUT_1[51750] = 32'b11111111111111111110011101010000;
assign LUT_1[51751] = 32'b11111111111111110111101111001100;
assign LUT_1[51752] = 32'b11111111111111111010000011011101;
assign LUT_1[51753] = 32'b11111111111111110011010101011001;
assign LUT_1[51754] = 32'b11111111111111110101110001101110;
assign LUT_1[51755] = 32'b11111111111111101111000011101010;
assign LUT_1[51756] = 32'b00000000000000000001111100110100;
assign LUT_1[51757] = 32'b11111111111111111011001110110000;
assign LUT_1[51758] = 32'b11111111111111111101101011000101;
assign LUT_1[51759] = 32'b11111111111111110110111101000001;
assign LUT_1[51760] = 32'b11111111111111111100110001001010;
assign LUT_1[51761] = 32'b11111111111111110110000011000110;
assign LUT_1[51762] = 32'b11111111111111111000011111011011;
assign LUT_1[51763] = 32'b11111111111111110001110001010111;
assign LUT_1[51764] = 32'b00000000000000000100101010100001;
assign LUT_1[51765] = 32'b11111111111111111101111100011101;
assign LUT_1[51766] = 32'b00000000000000000000011000110010;
assign LUT_1[51767] = 32'b11111111111111111001101010101110;
assign LUT_1[51768] = 32'b11111111111111111011111110111111;
assign LUT_1[51769] = 32'b11111111111111110101010000111011;
assign LUT_1[51770] = 32'b11111111111111110111101101010000;
assign LUT_1[51771] = 32'b11111111111111110000111111001100;
assign LUT_1[51772] = 32'b00000000000000000011111000010110;
assign LUT_1[51773] = 32'b11111111111111111101001010010010;
assign LUT_1[51774] = 32'b11111111111111111111100110100111;
assign LUT_1[51775] = 32'b11111111111111111000111000100011;
assign LUT_1[51776] = 32'b11111111111111111011111000010001;
assign LUT_1[51777] = 32'b11111111111111110101001010001101;
assign LUT_1[51778] = 32'b11111111111111110111100110100010;
assign LUT_1[51779] = 32'b11111111111111110000111000011110;
assign LUT_1[51780] = 32'b00000000000000000011110001101000;
assign LUT_1[51781] = 32'b11111111111111111101000011100100;
assign LUT_1[51782] = 32'b11111111111111111111011111111001;
assign LUT_1[51783] = 32'b11111111111111111000110001110101;
assign LUT_1[51784] = 32'b11111111111111111011000110000110;
assign LUT_1[51785] = 32'b11111111111111110100011000000010;
assign LUT_1[51786] = 32'b11111111111111110110110100010111;
assign LUT_1[51787] = 32'b11111111111111110000000110010011;
assign LUT_1[51788] = 32'b00000000000000000010111111011101;
assign LUT_1[51789] = 32'b11111111111111111100010001011001;
assign LUT_1[51790] = 32'b11111111111111111110101101101110;
assign LUT_1[51791] = 32'b11111111111111110111111111101010;
assign LUT_1[51792] = 32'b11111111111111111101110011110011;
assign LUT_1[51793] = 32'b11111111111111110111000101101111;
assign LUT_1[51794] = 32'b11111111111111111001100010000100;
assign LUT_1[51795] = 32'b11111111111111110010110100000000;
assign LUT_1[51796] = 32'b00000000000000000101101101001010;
assign LUT_1[51797] = 32'b11111111111111111110111111000110;
assign LUT_1[51798] = 32'b00000000000000000001011011011011;
assign LUT_1[51799] = 32'b11111111111111111010101101010111;
assign LUT_1[51800] = 32'b11111111111111111101000001101000;
assign LUT_1[51801] = 32'b11111111111111110110010011100100;
assign LUT_1[51802] = 32'b11111111111111111000101111111001;
assign LUT_1[51803] = 32'b11111111111111110010000001110101;
assign LUT_1[51804] = 32'b00000000000000000100111010111111;
assign LUT_1[51805] = 32'b11111111111111111110001100111011;
assign LUT_1[51806] = 32'b00000000000000000000101001010000;
assign LUT_1[51807] = 32'b11111111111111111001111011001100;
assign LUT_1[51808] = 32'b11111111111111111100110011010000;
assign LUT_1[51809] = 32'b11111111111111110110000101001100;
assign LUT_1[51810] = 32'b11111111111111111000100001100001;
assign LUT_1[51811] = 32'b11111111111111110001110011011101;
assign LUT_1[51812] = 32'b00000000000000000100101100100111;
assign LUT_1[51813] = 32'b11111111111111111101111110100011;
assign LUT_1[51814] = 32'b00000000000000000000011010111000;
assign LUT_1[51815] = 32'b11111111111111111001101100110100;
assign LUT_1[51816] = 32'b11111111111111111100000001000101;
assign LUT_1[51817] = 32'b11111111111111110101010011000001;
assign LUT_1[51818] = 32'b11111111111111110111101111010110;
assign LUT_1[51819] = 32'b11111111111111110001000001010010;
assign LUT_1[51820] = 32'b00000000000000000011111010011100;
assign LUT_1[51821] = 32'b11111111111111111101001100011000;
assign LUT_1[51822] = 32'b11111111111111111111101000101101;
assign LUT_1[51823] = 32'b11111111111111111000111010101001;
assign LUT_1[51824] = 32'b11111111111111111110101110110010;
assign LUT_1[51825] = 32'b11111111111111111000000000101110;
assign LUT_1[51826] = 32'b11111111111111111010011101000011;
assign LUT_1[51827] = 32'b11111111111111110011101110111111;
assign LUT_1[51828] = 32'b00000000000000000110101000001001;
assign LUT_1[51829] = 32'b11111111111111111111111010000101;
assign LUT_1[51830] = 32'b00000000000000000010010110011010;
assign LUT_1[51831] = 32'b11111111111111111011101000010110;
assign LUT_1[51832] = 32'b11111111111111111101111100100111;
assign LUT_1[51833] = 32'b11111111111111110111001110100011;
assign LUT_1[51834] = 32'b11111111111111111001101010111000;
assign LUT_1[51835] = 32'b11111111111111110010111100110100;
assign LUT_1[51836] = 32'b00000000000000000101110101111110;
assign LUT_1[51837] = 32'b11111111111111111111000111111010;
assign LUT_1[51838] = 32'b00000000000000000001100100001111;
assign LUT_1[51839] = 32'b11111111111111111010110110001011;
assign LUT_1[51840] = 32'b11111111111111111100111010101100;
assign LUT_1[51841] = 32'b11111111111111110110001100101000;
assign LUT_1[51842] = 32'b11111111111111111000101000111101;
assign LUT_1[51843] = 32'b11111111111111110001111010111001;
assign LUT_1[51844] = 32'b00000000000000000100110100000011;
assign LUT_1[51845] = 32'b11111111111111111110000101111111;
assign LUT_1[51846] = 32'b00000000000000000000100010010100;
assign LUT_1[51847] = 32'b11111111111111111001110100010000;
assign LUT_1[51848] = 32'b11111111111111111100001000100001;
assign LUT_1[51849] = 32'b11111111111111110101011010011101;
assign LUT_1[51850] = 32'b11111111111111110111110110110010;
assign LUT_1[51851] = 32'b11111111111111110001001000101110;
assign LUT_1[51852] = 32'b00000000000000000100000001111000;
assign LUT_1[51853] = 32'b11111111111111111101010011110100;
assign LUT_1[51854] = 32'b11111111111111111111110000001001;
assign LUT_1[51855] = 32'b11111111111111111001000010000101;
assign LUT_1[51856] = 32'b11111111111111111110110110001110;
assign LUT_1[51857] = 32'b11111111111111111000001000001010;
assign LUT_1[51858] = 32'b11111111111111111010100100011111;
assign LUT_1[51859] = 32'b11111111111111110011110110011011;
assign LUT_1[51860] = 32'b00000000000000000110101111100101;
assign LUT_1[51861] = 32'b00000000000000000000000001100001;
assign LUT_1[51862] = 32'b00000000000000000010011101110110;
assign LUT_1[51863] = 32'b11111111111111111011101111110010;
assign LUT_1[51864] = 32'b11111111111111111110000100000011;
assign LUT_1[51865] = 32'b11111111111111110111010101111111;
assign LUT_1[51866] = 32'b11111111111111111001110010010100;
assign LUT_1[51867] = 32'b11111111111111110011000100010000;
assign LUT_1[51868] = 32'b00000000000000000101111101011010;
assign LUT_1[51869] = 32'b11111111111111111111001111010110;
assign LUT_1[51870] = 32'b00000000000000000001101011101011;
assign LUT_1[51871] = 32'b11111111111111111010111101100111;
assign LUT_1[51872] = 32'b11111111111111111101110101101011;
assign LUT_1[51873] = 32'b11111111111111110111000111100111;
assign LUT_1[51874] = 32'b11111111111111111001100011111100;
assign LUT_1[51875] = 32'b11111111111111110010110101111000;
assign LUT_1[51876] = 32'b00000000000000000101101111000010;
assign LUT_1[51877] = 32'b11111111111111111111000000111110;
assign LUT_1[51878] = 32'b00000000000000000001011101010011;
assign LUT_1[51879] = 32'b11111111111111111010101111001111;
assign LUT_1[51880] = 32'b11111111111111111101000011100000;
assign LUT_1[51881] = 32'b11111111111111110110010101011100;
assign LUT_1[51882] = 32'b11111111111111111000110001110001;
assign LUT_1[51883] = 32'b11111111111111110010000011101101;
assign LUT_1[51884] = 32'b00000000000000000100111100110111;
assign LUT_1[51885] = 32'b11111111111111111110001110110011;
assign LUT_1[51886] = 32'b00000000000000000000101011001000;
assign LUT_1[51887] = 32'b11111111111111111001111101000100;
assign LUT_1[51888] = 32'b11111111111111111111110001001101;
assign LUT_1[51889] = 32'b11111111111111111001000011001001;
assign LUT_1[51890] = 32'b11111111111111111011011111011110;
assign LUT_1[51891] = 32'b11111111111111110100110001011010;
assign LUT_1[51892] = 32'b00000000000000000111101010100100;
assign LUT_1[51893] = 32'b00000000000000000000111100100000;
assign LUT_1[51894] = 32'b00000000000000000011011000110101;
assign LUT_1[51895] = 32'b11111111111111111100101010110001;
assign LUT_1[51896] = 32'b11111111111111111110111111000010;
assign LUT_1[51897] = 32'b11111111111111111000010000111110;
assign LUT_1[51898] = 32'b11111111111111111010101101010011;
assign LUT_1[51899] = 32'b11111111111111110011111111001111;
assign LUT_1[51900] = 32'b00000000000000000110111000011001;
assign LUT_1[51901] = 32'b00000000000000000000001010010101;
assign LUT_1[51902] = 32'b00000000000000000010100110101010;
assign LUT_1[51903] = 32'b11111111111111111011111000100110;
assign LUT_1[51904] = 32'b11111111111111111110111000010100;
assign LUT_1[51905] = 32'b11111111111111111000001010010000;
assign LUT_1[51906] = 32'b11111111111111111010100110100101;
assign LUT_1[51907] = 32'b11111111111111110011111000100001;
assign LUT_1[51908] = 32'b00000000000000000110110001101011;
assign LUT_1[51909] = 32'b00000000000000000000000011100111;
assign LUT_1[51910] = 32'b00000000000000000010011111111100;
assign LUT_1[51911] = 32'b11111111111111111011110001111000;
assign LUT_1[51912] = 32'b11111111111111111110000110001001;
assign LUT_1[51913] = 32'b11111111111111110111011000000101;
assign LUT_1[51914] = 32'b11111111111111111001110100011010;
assign LUT_1[51915] = 32'b11111111111111110011000110010110;
assign LUT_1[51916] = 32'b00000000000000000101111111100000;
assign LUT_1[51917] = 32'b11111111111111111111010001011100;
assign LUT_1[51918] = 32'b00000000000000000001101101110001;
assign LUT_1[51919] = 32'b11111111111111111010111111101101;
assign LUT_1[51920] = 32'b00000000000000000000110011110110;
assign LUT_1[51921] = 32'b11111111111111111010000101110010;
assign LUT_1[51922] = 32'b11111111111111111100100010000111;
assign LUT_1[51923] = 32'b11111111111111110101110100000011;
assign LUT_1[51924] = 32'b00000000000000001000101101001101;
assign LUT_1[51925] = 32'b00000000000000000001111111001001;
assign LUT_1[51926] = 32'b00000000000000000100011011011110;
assign LUT_1[51927] = 32'b11111111111111111101101101011010;
assign LUT_1[51928] = 32'b00000000000000000000000001101011;
assign LUT_1[51929] = 32'b11111111111111111001010011100111;
assign LUT_1[51930] = 32'b11111111111111111011101111111100;
assign LUT_1[51931] = 32'b11111111111111110101000001111000;
assign LUT_1[51932] = 32'b00000000000000000111111011000010;
assign LUT_1[51933] = 32'b00000000000000000001001100111110;
assign LUT_1[51934] = 32'b00000000000000000011101001010011;
assign LUT_1[51935] = 32'b11111111111111111100111011001111;
assign LUT_1[51936] = 32'b11111111111111111111110011010011;
assign LUT_1[51937] = 32'b11111111111111111001000101001111;
assign LUT_1[51938] = 32'b11111111111111111011100001100100;
assign LUT_1[51939] = 32'b11111111111111110100110011100000;
assign LUT_1[51940] = 32'b00000000000000000111101100101010;
assign LUT_1[51941] = 32'b00000000000000000000111110100110;
assign LUT_1[51942] = 32'b00000000000000000011011010111011;
assign LUT_1[51943] = 32'b11111111111111111100101100110111;
assign LUT_1[51944] = 32'b11111111111111111111000001001000;
assign LUT_1[51945] = 32'b11111111111111111000010011000100;
assign LUT_1[51946] = 32'b11111111111111111010101111011001;
assign LUT_1[51947] = 32'b11111111111111110100000001010101;
assign LUT_1[51948] = 32'b00000000000000000110111010011111;
assign LUT_1[51949] = 32'b00000000000000000000001100011011;
assign LUT_1[51950] = 32'b00000000000000000010101000110000;
assign LUT_1[51951] = 32'b11111111111111111011111010101100;
assign LUT_1[51952] = 32'b00000000000000000001101110110101;
assign LUT_1[51953] = 32'b11111111111111111011000000110001;
assign LUT_1[51954] = 32'b11111111111111111101011101000110;
assign LUT_1[51955] = 32'b11111111111111110110101111000010;
assign LUT_1[51956] = 32'b00000000000000001001101000001100;
assign LUT_1[51957] = 32'b00000000000000000010111010001000;
assign LUT_1[51958] = 32'b00000000000000000101010110011101;
assign LUT_1[51959] = 32'b11111111111111111110101000011001;
assign LUT_1[51960] = 32'b00000000000000000000111100101010;
assign LUT_1[51961] = 32'b11111111111111111010001110100110;
assign LUT_1[51962] = 32'b11111111111111111100101010111011;
assign LUT_1[51963] = 32'b11111111111111110101111100110111;
assign LUT_1[51964] = 32'b00000000000000001000110110000001;
assign LUT_1[51965] = 32'b00000000000000000010000111111101;
assign LUT_1[51966] = 32'b00000000000000000100100100010010;
assign LUT_1[51967] = 32'b11111111111111111101110110001110;
assign LUT_1[51968] = 32'b11111111111111110111101110110101;
assign LUT_1[51969] = 32'b11111111111111110001000000110001;
assign LUT_1[51970] = 32'b11111111111111110011011101000110;
assign LUT_1[51971] = 32'b11111111111111101100101111000010;
assign LUT_1[51972] = 32'b11111111111111111111101000001100;
assign LUT_1[51973] = 32'b11111111111111111000111010001000;
assign LUT_1[51974] = 32'b11111111111111111011010110011101;
assign LUT_1[51975] = 32'b11111111111111110100101000011001;
assign LUT_1[51976] = 32'b11111111111111110110111100101010;
assign LUT_1[51977] = 32'b11111111111111110000001110100110;
assign LUT_1[51978] = 32'b11111111111111110010101010111011;
assign LUT_1[51979] = 32'b11111111111111101011111100110111;
assign LUT_1[51980] = 32'b11111111111111111110110110000001;
assign LUT_1[51981] = 32'b11111111111111111000000111111101;
assign LUT_1[51982] = 32'b11111111111111111010100100010010;
assign LUT_1[51983] = 32'b11111111111111110011110110001110;
assign LUT_1[51984] = 32'b11111111111111111001101010010111;
assign LUT_1[51985] = 32'b11111111111111110010111100010011;
assign LUT_1[51986] = 32'b11111111111111110101011000101000;
assign LUT_1[51987] = 32'b11111111111111101110101010100100;
assign LUT_1[51988] = 32'b00000000000000000001100011101110;
assign LUT_1[51989] = 32'b11111111111111111010110101101010;
assign LUT_1[51990] = 32'b11111111111111111101010001111111;
assign LUT_1[51991] = 32'b11111111111111110110100011111011;
assign LUT_1[51992] = 32'b11111111111111111000111000001100;
assign LUT_1[51993] = 32'b11111111111111110010001010001000;
assign LUT_1[51994] = 32'b11111111111111110100100110011101;
assign LUT_1[51995] = 32'b11111111111111101101111000011001;
assign LUT_1[51996] = 32'b00000000000000000000110001100011;
assign LUT_1[51997] = 32'b11111111111111111010000011011111;
assign LUT_1[51998] = 32'b11111111111111111100011111110100;
assign LUT_1[51999] = 32'b11111111111111110101110001110000;
assign LUT_1[52000] = 32'b11111111111111111000101001110100;
assign LUT_1[52001] = 32'b11111111111111110001111011110000;
assign LUT_1[52002] = 32'b11111111111111110100011000000101;
assign LUT_1[52003] = 32'b11111111111111101101101010000001;
assign LUT_1[52004] = 32'b00000000000000000000100011001011;
assign LUT_1[52005] = 32'b11111111111111111001110101000111;
assign LUT_1[52006] = 32'b11111111111111111100010001011100;
assign LUT_1[52007] = 32'b11111111111111110101100011011000;
assign LUT_1[52008] = 32'b11111111111111110111110111101001;
assign LUT_1[52009] = 32'b11111111111111110001001001100101;
assign LUT_1[52010] = 32'b11111111111111110011100101111010;
assign LUT_1[52011] = 32'b11111111111111101100110111110110;
assign LUT_1[52012] = 32'b11111111111111111111110001000000;
assign LUT_1[52013] = 32'b11111111111111111001000010111100;
assign LUT_1[52014] = 32'b11111111111111111011011111010001;
assign LUT_1[52015] = 32'b11111111111111110100110001001101;
assign LUT_1[52016] = 32'b11111111111111111010100101010110;
assign LUT_1[52017] = 32'b11111111111111110011110111010010;
assign LUT_1[52018] = 32'b11111111111111110110010011100111;
assign LUT_1[52019] = 32'b11111111111111101111100101100011;
assign LUT_1[52020] = 32'b00000000000000000010011110101101;
assign LUT_1[52021] = 32'b11111111111111111011110000101001;
assign LUT_1[52022] = 32'b11111111111111111110001100111110;
assign LUT_1[52023] = 32'b11111111111111110111011110111010;
assign LUT_1[52024] = 32'b11111111111111111001110011001011;
assign LUT_1[52025] = 32'b11111111111111110011000101000111;
assign LUT_1[52026] = 32'b11111111111111110101100001011100;
assign LUT_1[52027] = 32'b11111111111111101110110011011000;
assign LUT_1[52028] = 32'b00000000000000000001101100100010;
assign LUT_1[52029] = 32'b11111111111111111010111110011110;
assign LUT_1[52030] = 32'b11111111111111111101011010110011;
assign LUT_1[52031] = 32'b11111111111111110110101100101111;
assign LUT_1[52032] = 32'b11111111111111111001101100011101;
assign LUT_1[52033] = 32'b11111111111111110010111110011001;
assign LUT_1[52034] = 32'b11111111111111110101011010101110;
assign LUT_1[52035] = 32'b11111111111111101110101100101010;
assign LUT_1[52036] = 32'b00000000000000000001100101110100;
assign LUT_1[52037] = 32'b11111111111111111010110111110000;
assign LUT_1[52038] = 32'b11111111111111111101010100000101;
assign LUT_1[52039] = 32'b11111111111111110110100110000001;
assign LUT_1[52040] = 32'b11111111111111111000111010010010;
assign LUT_1[52041] = 32'b11111111111111110010001100001110;
assign LUT_1[52042] = 32'b11111111111111110100101000100011;
assign LUT_1[52043] = 32'b11111111111111101101111010011111;
assign LUT_1[52044] = 32'b00000000000000000000110011101001;
assign LUT_1[52045] = 32'b11111111111111111010000101100101;
assign LUT_1[52046] = 32'b11111111111111111100100001111010;
assign LUT_1[52047] = 32'b11111111111111110101110011110110;
assign LUT_1[52048] = 32'b11111111111111111011100111111111;
assign LUT_1[52049] = 32'b11111111111111110100111001111011;
assign LUT_1[52050] = 32'b11111111111111110111010110010000;
assign LUT_1[52051] = 32'b11111111111111110000101000001100;
assign LUT_1[52052] = 32'b00000000000000000011100001010110;
assign LUT_1[52053] = 32'b11111111111111111100110011010010;
assign LUT_1[52054] = 32'b11111111111111111111001111100111;
assign LUT_1[52055] = 32'b11111111111111111000100001100011;
assign LUT_1[52056] = 32'b11111111111111111010110101110100;
assign LUT_1[52057] = 32'b11111111111111110100000111110000;
assign LUT_1[52058] = 32'b11111111111111110110100100000101;
assign LUT_1[52059] = 32'b11111111111111101111110110000001;
assign LUT_1[52060] = 32'b00000000000000000010101111001011;
assign LUT_1[52061] = 32'b11111111111111111100000001000111;
assign LUT_1[52062] = 32'b11111111111111111110011101011100;
assign LUT_1[52063] = 32'b11111111111111110111101111011000;
assign LUT_1[52064] = 32'b11111111111111111010100111011100;
assign LUT_1[52065] = 32'b11111111111111110011111001011000;
assign LUT_1[52066] = 32'b11111111111111110110010101101101;
assign LUT_1[52067] = 32'b11111111111111101111100111101001;
assign LUT_1[52068] = 32'b00000000000000000010100000110011;
assign LUT_1[52069] = 32'b11111111111111111011110010101111;
assign LUT_1[52070] = 32'b11111111111111111110001111000100;
assign LUT_1[52071] = 32'b11111111111111110111100001000000;
assign LUT_1[52072] = 32'b11111111111111111001110101010001;
assign LUT_1[52073] = 32'b11111111111111110011000111001101;
assign LUT_1[52074] = 32'b11111111111111110101100011100010;
assign LUT_1[52075] = 32'b11111111111111101110110101011110;
assign LUT_1[52076] = 32'b00000000000000000001101110101000;
assign LUT_1[52077] = 32'b11111111111111111011000000100100;
assign LUT_1[52078] = 32'b11111111111111111101011100111001;
assign LUT_1[52079] = 32'b11111111111111110110101110110101;
assign LUT_1[52080] = 32'b11111111111111111100100010111110;
assign LUT_1[52081] = 32'b11111111111111110101110100111010;
assign LUT_1[52082] = 32'b11111111111111111000010001001111;
assign LUT_1[52083] = 32'b11111111111111110001100011001011;
assign LUT_1[52084] = 32'b00000000000000000100011100010101;
assign LUT_1[52085] = 32'b11111111111111111101101110010001;
assign LUT_1[52086] = 32'b00000000000000000000001010100110;
assign LUT_1[52087] = 32'b11111111111111111001011100100010;
assign LUT_1[52088] = 32'b11111111111111111011110000110011;
assign LUT_1[52089] = 32'b11111111111111110101000010101111;
assign LUT_1[52090] = 32'b11111111111111110111011111000100;
assign LUT_1[52091] = 32'b11111111111111110000110001000000;
assign LUT_1[52092] = 32'b00000000000000000011101010001010;
assign LUT_1[52093] = 32'b11111111111111111100111100000110;
assign LUT_1[52094] = 32'b11111111111111111111011000011011;
assign LUT_1[52095] = 32'b11111111111111111000101010010111;
assign LUT_1[52096] = 32'b11111111111111111010101110111000;
assign LUT_1[52097] = 32'b11111111111111110100000000110100;
assign LUT_1[52098] = 32'b11111111111111110110011101001001;
assign LUT_1[52099] = 32'b11111111111111101111101111000101;
assign LUT_1[52100] = 32'b00000000000000000010101000001111;
assign LUT_1[52101] = 32'b11111111111111111011111010001011;
assign LUT_1[52102] = 32'b11111111111111111110010110100000;
assign LUT_1[52103] = 32'b11111111111111110111101000011100;
assign LUT_1[52104] = 32'b11111111111111111001111100101101;
assign LUT_1[52105] = 32'b11111111111111110011001110101001;
assign LUT_1[52106] = 32'b11111111111111110101101010111110;
assign LUT_1[52107] = 32'b11111111111111101110111100111010;
assign LUT_1[52108] = 32'b00000000000000000001110110000100;
assign LUT_1[52109] = 32'b11111111111111111011001000000000;
assign LUT_1[52110] = 32'b11111111111111111101100100010101;
assign LUT_1[52111] = 32'b11111111111111110110110110010001;
assign LUT_1[52112] = 32'b11111111111111111100101010011010;
assign LUT_1[52113] = 32'b11111111111111110101111100010110;
assign LUT_1[52114] = 32'b11111111111111111000011000101011;
assign LUT_1[52115] = 32'b11111111111111110001101010100111;
assign LUT_1[52116] = 32'b00000000000000000100100011110001;
assign LUT_1[52117] = 32'b11111111111111111101110101101101;
assign LUT_1[52118] = 32'b00000000000000000000010010000010;
assign LUT_1[52119] = 32'b11111111111111111001100011111110;
assign LUT_1[52120] = 32'b11111111111111111011111000001111;
assign LUT_1[52121] = 32'b11111111111111110101001010001011;
assign LUT_1[52122] = 32'b11111111111111110111100110100000;
assign LUT_1[52123] = 32'b11111111111111110000111000011100;
assign LUT_1[52124] = 32'b00000000000000000011110001100110;
assign LUT_1[52125] = 32'b11111111111111111101000011100010;
assign LUT_1[52126] = 32'b11111111111111111111011111110111;
assign LUT_1[52127] = 32'b11111111111111111000110001110011;
assign LUT_1[52128] = 32'b11111111111111111011101001110111;
assign LUT_1[52129] = 32'b11111111111111110100111011110011;
assign LUT_1[52130] = 32'b11111111111111110111011000001000;
assign LUT_1[52131] = 32'b11111111111111110000101010000100;
assign LUT_1[52132] = 32'b00000000000000000011100011001110;
assign LUT_1[52133] = 32'b11111111111111111100110101001010;
assign LUT_1[52134] = 32'b11111111111111111111010001011111;
assign LUT_1[52135] = 32'b11111111111111111000100011011011;
assign LUT_1[52136] = 32'b11111111111111111010110111101100;
assign LUT_1[52137] = 32'b11111111111111110100001001101000;
assign LUT_1[52138] = 32'b11111111111111110110100101111101;
assign LUT_1[52139] = 32'b11111111111111101111110111111001;
assign LUT_1[52140] = 32'b00000000000000000010110001000011;
assign LUT_1[52141] = 32'b11111111111111111100000010111111;
assign LUT_1[52142] = 32'b11111111111111111110011111010100;
assign LUT_1[52143] = 32'b11111111111111110111110001010000;
assign LUT_1[52144] = 32'b11111111111111111101100101011001;
assign LUT_1[52145] = 32'b11111111111111110110110111010101;
assign LUT_1[52146] = 32'b11111111111111111001010011101010;
assign LUT_1[52147] = 32'b11111111111111110010100101100110;
assign LUT_1[52148] = 32'b00000000000000000101011110110000;
assign LUT_1[52149] = 32'b11111111111111111110110000101100;
assign LUT_1[52150] = 32'b00000000000000000001001101000001;
assign LUT_1[52151] = 32'b11111111111111111010011110111101;
assign LUT_1[52152] = 32'b11111111111111111100110011001110;
assign LUT_1[52153] = 32'b11111111111111110110000101001010;
assign LUT_1[52154] = 32'b11111111111111111000100001011111;
assign LUT_1[52155] = 32'b11111111111111110001110011011011;
assign LUT_1[52156] = 32'b00000000000000000100101100100101;
assign LUT_1[52157] = 32'b11111111111111111101111110100001;
assign LUT_1[52158] = 32'b00000000000000000000011010110110;
assign LUT_1[52159] = 32'b11111111111111111001101100110010;
assign LUT_1[52160] = 32'b11111111111111111100101100100000;
assign LUT_1[52161] = 32'b11111111111111110101111110011100;
assign LUT_1[52162] = 32'b11111111111111111000011010110001;
assign LUT_1[52163] = 32'b11111111111111110001101100101101;
assign LUT_1[52164] = 32'b00000000000000000100100101110111;
assign LUT_1[52165] = 32'b11111111111111111101110111110011;
assign LUT_1[52166] = 32'b00000000000000000000010100001000;
assign LUT_1[52167] = 32'b11111111111111111001100110000100;
assign LUT_1[52168] = 32'b11111111111111111011111010010101;
assign LUT_1[52169] = 32'b11111111111111110101001100010001;
assign LUT_1[52170] = 32'b11111111111111110111101000100110;
assign LUT_1[52171] = 32'b11111111111111110000111010100010;
assign LUT_1[52172] = 32'b00000000000000000011110011101100;
assign LUT_1[52173] = 32'b11111111111111111101000101101000;
assign LUT_1[52174] = 32'b11111111111111111111100001111101;
assign LUT_1[52175] = 32'b11111111111111111000110011111001;
assign LUT_1[52176] = 32'b11111111111111111110101000000010;
assign LUT_1[52177] = 32'b11111111111111110111111001111110;
assign LUT_1[52178] = 32'b11111111111111111010010110010011;
assign LUT_1[52179] = 32'b11111111111111110011101000001111;
assign LUT_1[52180] = 32'b00000000000000000110100001011001;
assign LUT_1[52181] = 32'b11111111111111111111110011010101;
assign LUT_1[52182] = 32'b00000000000000000010001111101010;
assign LUT_1[52183] = 32'b11111111111111111011100001100110;
assign LUT_1[52184] = 32'b11111111111111111101110101110111;
assign LUT_1[52185] = 32'b11111111111111110111000111110011;
assign LUT_1[52186] = 32'b11111111111111111001100100001000;
assign LUT_1[52187] = 32'b11111111111111110010110110000100;
assign LUT_1[52188] = 32'b00000000000000000101101111001110;
assign LUT_1[52189] = 32'b11111111111111111111000001001010;
assign LUT_1[52190] = 32'b00000000000000000001011101011111;
assign LUT_1[52191] = 32'b11111111111111111010101111011011;
assign LUT_1[52192] = 32'b11111111111111111101100111011111;
assign LUT_1[52193] = 32'b11111111111111110110111001011011;
assign LUT_1[52194] = 32'b11111111111111111001010101110000;
assign LUT_1[52195] = 32'b11111111111111110010100111101100;
assign LUT_1[52196] = 32'b00000000000000000101100000110110;
assign LUT_1[52197] = 32'b11111111111111111110110010110010;
assign LUT_1[52198] = 32'b00000000000000000001001111000111;
assign LUT_1[52199] = 32'b11111111111111111010100001000011;
assign LUT_1[52200] = 32'b11111111111111111100110101010100;
assign LUT_1[52201] = 32'b11111111111111110110000111010000;
assign LUT_1[52202] = 32'b11111111111111111000100011100101;
assign LUT_1[52203] = 32'b11111111111111110001110101100001;
assign LUT_1[52204] = 32'b00000000000000000100101110101011;
assign LUT_1[52205] = 32'b11111111111111111110000000100111;
assign LUT_1[52206] = 32'b00000000000000000000011100111100;
assign LUT_1[52207] = 32'b11111111111111111001101110111000;
assign LUT_1[52208] = 32'b11111111111111111111100011000001;
assign LUT_1[52209] = 32'b11111111111111111000110100111101;
assign LUT_1[52210] = 32'b11111111111111111011010001010010;
assign LUT_1[52211] = 32'b11111111111111110100100011001110;
assign LUT_1[52212] = 32'b00000000000000000111011100011000;
assign LUT_1[52213] = 32'b00000000000000000000101110010100;
assign LUT_1[52214] = 32'b00000000000000000011001010101001;
assign LUT_1[52215] = 32'b11111111111111111100011100100101;
assign LUT_1[52216] = 32'b11111111111111111110110000110110;
assign LUT_1[52217] = 32'b11111111111111111000000010110010;
assign LUT_1[52218] = 32'b11111111111111111010011111000111;
assign LUT_1[52219] = 32'b11111111111111110011110001000011;
assign LUT_1[52220] = 32'b00000000000000000110101010001101;
assign LUT_1[52221] = 32'b11111111111111111111111100001001;
assign LUT_1[52222] = 32'b00000000000000000010011000011110;
assign LUT_1[52223] = 32'b11111111111111111011101010011010;
assign LUT_1[52224] = 32'b00000000000000000110100010111100;
assign LUT_1[52225] = 32'b11111111111111111111110100111000;
assign LUT_1[52226] = 32'b00000000000000000010010001001101;
assign LUT_1[52227] = 32'b11111111111111111011100011001001;
assign LUT_1[52228] = 32'b00000000000000001110011100010011;
assign LUT_1[52229] = 32'b00000000000000000111101110001111;
assign LUT_1[52230] = 32'b00000000000000001010001010100100;
assign LUT_1[52231] = 32'b00000000000000000011011100100000;
assign LUT_1[52232] = 32'b00000000000000000101110000110001;
assign LUT_1[52233] = 32'b11111111111111111111000010101101;
assign LUT_1[52234] = 32'b00000000000000000001011111000010;
assign LUT_1[52235] = 32'b11111111111111111010110000111110;
assign LUT_1[52236] = 32'b00000000000000001101101010001000;
assign LUT_1[52237] = 32'b00000000000000000110111100000100;
assign LUT_1[52238] = 32'b00000000000000001001011000011001;
assign LUT_1[52239] = 32'b00000000000000000010101010010101;
assign LUT_1[52240] = 32'b00000000000000001000011110011110;
assign LUT_1[52241] = 32'b00000000000000000001110000011010;
assign LUT_1[52242] = 32'b00000000000000000100001100101111;
assign LUT_1[52243] = 32'b11111111111111111101011110101011;
assign LUT_1[52244] = 32'b00000000000000010000010111110101;
assign LUT_1[52245] = 32'b00000000000000001001101001110001;
assign LUT_1[52246] = 32'b00000000000000001100000110000110;
assign LUT_1[52247] = 32'b00000000000000000101011000000010;
assign LUT_1[52248] = 32'b00000000000000000111101100010011;
assign LUT_1[52249] = 32'b00000000000000000000111110001111;
assign LUT_1[52250] = 32'b00000000000000000011011010100100;
assign LUT_1[52251] = 32'b11111111111111111100101100100000;
assign LUT_1[52252] = 32'b00000000000000001111100101101010;
assign LUT_1[52253] = 32'b00000000000000001000110111100110;
assign LUT_1[52254] = 32'b00000000000000001011010011111011;
assign LUT_1[52255] = 32'b00000000000000000100100101110111;
assign LUT_1[52256] = 32'b00000000000000000111011101111011;
assign LUT_1[52257] = 32'b00000000000000000000101111110111;
assign LUT_1[52258] = 32'b00000000000000000011001100001100;
assign LUT_1[52259] = 32'b11111111111111111100011110001000;
assign LUT_1[52260] = 32'b00000000000000001111010111010010;
assign LUT_1[52261] = 32'b00000000000000001000101001001110;
assign LUT_1[52262] = 32'b00000000000000001011000101100011;
assign LUT_1[52263] = 32'b00000000000000000100010111011111;
assign LUT_1[52264] = 32'b00000000000000000110101011110000;
assign LUT_1[52265] = 32'b11111111111111111111111101101100;
assign LUT_1[52266] = 32'b00000000000000000010011010000001;
assign LUT_1[52267] = 32'b11111111111111111011101011111101;
assign LUT_1[52268] = 32'b00000000000000001110100101000111;
assign LUT_1[52269] = 32'b00000000000000000111110111000011;
assign LUT_1[52270] = 32'b00000000000000001010010011011000;
assign LUT_1[52271] = 32'b00000000000000000011100101010100;
assign LUT_1[52272] = 32'b00000000000000001001011001011101;
assign LUT_1[52273] = 32'b00000000000000000010101011011001;
assign LUT_1[52274] = 32'b00000000000000000101000111101110;
assign LUT_1[52275] = 32'b11111111111111111110011001101010;
assign LUT_1[52276] = 32'b00000000000000010001010010110100;
assign LUT_1[52277] = 32'b00000000000000001010100100110000;
assign LUT_1[52278] = 32'b00000000000000001101000001000101;
assign LUT_1[52279] = 32'b00000000000000000110010011000001;
assign LUT_1[52280] = 32'b00000000000000001000100111010010;
assign LUT_1[52281] = 32'b00000000000000000001111001001110;
assign LUT_1[52282] = 32'b00000000000000000100010101100011;
assign LUT_1[52283] = 32'b11111111111111111101100111011111;
assign LUT_1[52284] = 32'b00000000000000010000100000101001;
assign LUT_1[52285] = 32'b00000000000000001001110010100101;
assign LUT_1[52286] = 32'b00000000000000001100001110111010;
assign LUT_1[52287] = 32'b00000000000000000101100000110110;
assign LUT_1[52288] = 32'b00000000000000001000100000100100;
assign LUT_1[52289] = 32'b00000000000000000001110010100000;
assign LUT_1[52290] = 32'b00000000000000000100001110110101;
assign LUT_1[52291] = 32'b11111111111111111101100000110001;
assign LUT_1[52292] = 32'b00000000000000010000011001111011;
assign LUT_1[52293] = 32'b00000000000000001001101011110111;
assign LUT_1[52294] = 32'b00000000000000001100001000001100;
assign LUT_1[52295] = 32'b00000000000000000101011010001000;
assign LUT_1[52296] = 32'b00000000000000000111101110011001;
assign LUT_1[52297] = 32'b00000000000000000001000000010101;
assign LUT_1[52298] = 32'b00000000000000000011011100101010;
assign LUT_1[52299] = 32'b11111111111111111100101110100110;
assign LUT_1[52300] = 32'b00000000000000001111100111110000;
assign LUT_1[52301] = 32'b00000000000000001000111001101100;
assign LUT_1[52302] = 32'b00000000000000001011010110000001;
assign LUT_1[52303] = 32'b00000000000000000100100111111101;
assign LUT_1[52304] = 32'b00000000000000001010011100000110;
assign LUT_1[52305] = 32'b00000000000000000011101110000010;
assign LUT_1[52306] = 32'b00000000000000000110001010010111;
assign LUT_1[52307] = 32'b11111111111111111111011100010011;
assign LUT_1[52308] = 32'b00000000000000010010010101011101;
assign LUT_1[52309] = 32'b00000000000000001011100111011001;
assign LUT_1[52310] = 32'b00000000000000001110000011101110;
assign LUT_1[52311] = 32'b00000000000000000111010101101010;
assign LUT_1[52312] = 32'b00000000000000001001101001111011;
assign LUT_1[52313] = 32'b00000000000000000010111011110111;
assign LUT_1[52314] = 32'b00000000000000000101011000001100;
assign LUT_1[52315] = 32'b11111111111111111110101010001000;
assign LUT_1[52316] = 32'b00000000000000010001100011010010;
assign LUT_1[52317] = 32'b00000000000000001010110101001110;
assign LUT_1[52318] = 32'b00000000000000001101010001100011;
assign LUT_1[52319] = 32'b00000000000000000110100011011111;
assign LUT_1[52320] = 32'b00000000000000001001011011100011;
assign LUT_1[52321] = 32'b00000000000000000010101101011111;
assign LUT_1[52322] = 32'b00000000000000000101001001110100;
assign LUT_1[52323] = 32'b11111111111111111110011011110000;
assign LUT_1[52324] = 32'b00000000000000010001010100111010;
assign LUT_1[52325] = 32'b00000000000000001010100110110110;
assign LUT_1[52326] = 32'b00000000000000001101000011001011;
assign LUT_1[52327] = 32'b00000000000000000110010101000111;
assign LUT_1[52328] = 32'b00000000000000001000101001011000;
assign LUT_1[52329] = 32'b00000000000000000001111011010100;
assign LUT_1[52330] = 32'b00000000000000000100010111101001;
assign LUT_1[52331] = 32'b11111111111111111101101001100101;
assign LUT_1[52332] = 32'b00000000000000010000100010101111;
assign LUT_1[52333] = 32'b00000000000000001001110100101011;
assign LUT_1[52334] = 32'b00000000000000001100010001000000;
assign LUT_1[52335] = 32'b00000000000000000101100010111100;
assign LUT_1[52336] = 32'b00000000000000001011010111000101;
assign LUT_1[52337] = 32'b00000000000000000100101001000001;
assign LUT_1[52338] = 32'b00000000000000000111000101010110;
assign LUT_1[52339] = 32'b00000000000000000000010111010010;
assign LUT_1[52340] = 32'b00000000000000010011010000011100;
assign LUT_1[52341] = 32'b00000000000000001100100010011000;
assign LUT_1[52342] = 32'b00000000000000001110111110101101;
assign LUT_1[52343] = 32'b00000000000000001000010000101001;
assign LUT_1[52344] = 32'b00000000000000001010100100111010;
assign LUT_1[52345] = 32'b00000000000000000011110110110110;
assign LUT_1[52346] = 32'b00000000000000000110010011001011;
assign LUT_1[52347] = 32'b11111111111111111111100101000111;
assign LUT_1[52348] = 32'b00000000000000010010011110010001;
assign LUT_1[52349] = 32'b00000000000000001011110000001101;
assign LUT_1[52350] = 32'b00000000000000001110001100100010;
assign LUT_1[52351] = 32'b00000000000000000111011110011110;
assign LUT_1[52352] = 32'b00000000000000001001100010111111;
assign LUT_1[52353] = 32'b00000000000000000010110100111011;
assign LUT_1[52354] = 32'b00000000000000000101010001010000;
assign LUT_1[52355] = 32'b11111111111111111110100011001100;
assign LUT_1[52356] = 32'b00000000000000010001011100010110;
assign LUT_1[52357] = 32'b00000000000000001010101110010010;
assign LUT_1[52358] = 32'b00000000000000001101001010100111;
assign LUT_1[52359] = 32'b00000000000000000110011100100011;
assign LUT_1[52360] = 32'b00000000000000001000110000110100;
assign LUT_1[52361] = 32'b00000000000000000010000010110000;
assign LUT_1[52362] = 32'b00000000000000000100011111000101;
assign LUT_1[52363] = 32'b11111111111111111101110001000001;
assign LUT_1[52364] = 32'b00000000000000010000101010001011;
assign LUT_1[52365] = 32'b00000000000000001001111100000111;
assign LUT_1[52366] = 32'b00000000000000001100011000011100;
assign LUT_1[52367] = 32'b00000000000000000101101010011000;
assign LUT_1[52368] = 32'b00000000000000001011011110100001;
assign LUT_1[52369] = 32'b00000000000000000100110000011101;
assign LUT_1[52370] = 32'b00000000000000000111001100110010;
assign LUT_1[52371] = 32'b00000000000000000000011110101110;
assign LUT_1[52372] = 32'b00000000000000010011010111111000;
assign LUT_1[52373] = 32'b00000000000000001100101001110100;
assign LUT_1[52374] = 32'b00000000000000001111000110001001;
assign LUT_1[52375] = 32'b00000000000000001000011000000101;
assign LUT_1[52376] = 32'b00000000000000001010101100010110;
assign LUT_1[52377] = 32'b00000000000000000011111110010010;
assign LUT_1[52378] = 32'b00000000000000000110011010100111;
assign LUT_1[52379] = 32'b11111111111111111111101100100011;
assign LUT_1[52380] = 32'b00000000000000010010100101101101;
assign LUT_1[52381] = 32'b00000000000000001011110111101001;
assign LUT_1[52382] = 32'b00000000000000001110010011111110;
assign LUT_1[52383] = 32'b00000000000000000111100101111010;
assign LUT_1[52384] = 32'b00000000000000001010011101111110;
assign LUT_1[52385] = 32'b00000000000000000011101111111010;
assign LUT_1[52386] = 32'b00000000000000000110001100001111;
assign LUT_1[52387] = 32'b11111111111111111111011110001011;
assign LUT_1[52388] = 32'b00000000000000010010010111010101;
assign LUT_1[52389] = 32'b00000000000000001011101001010001;
assign LUT_1[52390] = 32'b00000000000000001110000101100110;
assign LUT_1[52391] = 32'b00000000000000000111010111100010;
assign LUT_1[52392] = 32'b00000000000000001001101011110011;
assign LUT_1[52393] = 32'b00000000000000000010111101101111;
assign LUT_1[52394] = 32'b00000000000000000101011010000100;
assign LUT_1[52395] = 32'b11111111111111111110101100000000;
assign LUT_1[52396] = 32'b00000000000000010001100101001010;
assign LUT_1[52397] = 32'b00000000000000001010110111000110;
assign LUT_1[52398] = 32'b00000000000000001101010011011011;
assign LUT_1[52399] = 32'b00000000000000000110100101010111;
assign LUT_1[52400] = 32'b00000000000000001100011001100000;
assign LUT_1[52401] = 32'b00000000000000000101101011011100;
assign LUT_1[52402] = 32'b00000000000000001000000111110001;
assign LUT_1[52403] = 32'b00000000000000000001011001101101;
assign LUT_1[52404] = 32'b00000000000000010100010010110111;
assign LUT_1[52405] = 32'b00000000000000001101100100110011;
assign LUT_1[52406] = 32'b00000000000000010000000001001000;
assign LUT_1[52407] = 32'b00000000000000001001010011000100;
assign LUT_1[52408] = 32'b00000000000000001011100111010101;
assign LUT_1[52409] = 32'b00000000000000000100111001010001;
assign LUT_1[52410] = 32'b00000000000000000111010101100110;
assign LUT_1[52411] = 32'b00000000000000000000100111100010;
assign LUT_1[52412] = 32'b00000000000000010011100000101100;
assign LUT_1[52413] = 32'b00000000000000001100110010101000;
assign LUT_1[52414] = 32'b00000000000000001111001110111101;
assign LUT_1[52415] = 32'b00000000000000001000100000111001;
assign LUT_1[52416] = 32'b00000000000000001011100000100111;
assign LUT_1[52417] = 32'b00000000000000000100110010100011;
assign LUT_1[52418] = 32'b00000000000000000111001110111000;
assign LUT_1[52419] = 32'b00000000000000000000100000110100;
assign LUT_1[52420] = 32'b00000000000000010011011001111110;
assign LUT_1[52421] = 32'b00000000000000001100101011111010;
assign LUT_1[52422] = 32'b00000000000000001111001000001111;
assign LUT_1[52423] = 32'b00000000000000001000011010001011;
assign LUT_1[52424] = 32'b00000000000000001010101110011100;
assign LUT_1[52425] = 32'b00000000000000000100000000011000;
assign LUT_1[52426] = 32'b00000000000000000110011100101101;
assign LUT_1[52427] = 32'b11111111111111111111101110101001;
assign LUT_1[52428] = 32'b00000000000000010010100111110011;
assign LUT_1[52429] = 32'b00000000000000001011111001101111;
assign LUT_1[52430] = 32'b00000000000000001110010110000100;
assign LUT_1[52431] = 32'b00000000000000000111101000000000;
assign LUT_1[52432] = 32'b00000000000000001101011100001001;
assign LUT_1[52433] = 32'b00000000000000000110101110000101;
assign LUT_1[52434] = 32'b00000000000000001001001010011010;
assign LUT_1[52435] = 32'b00000000000000000010011100010110;
assign LUT_1[52436] = 32'b00000000000000010101010101100000;
assign LUT_1[52437] = 32'b00000000000000001110100111011100;
assign LUT_1[52438] = 32'b00000000000000010001000011110001;
assign LUT_1[52439] = 32'b00000000000000001010010101101101;
assign LUT_1[52440] = 32'b00000000000000001100101001111110;
assign LUT_1[52441] = 32'b00000000000000000101111011111010;
assign LUT_1[52442] = 32'b00000000000000001000011000001111;
assign LUT_1[52443] = 32'b00000000000000000001101010001011;
assign LUT_1[52444] = 32'b00000000000000010100100011010101;
assign LUT_1[52445] = 32'b00000000000000001101110101010001;
assign LUT_1[52446] = 32'b00000000000000010000010001100110;
assign LUT_1[52447] = 32'b00000000000000001001100011100010;
assign LUT_1[52448] = 32'b00000000000000001100011011100110;
assign LUT_1[52449] = 32'b00000000000000000101101101100010;
assign LUT_1[52450] = 32'b00000000000000001000001001110111;
assign LUT_1[52451] = 32'b00000000000000000001011011110011;
assign LUT_1[52452] = 32'b00000000000000010100010100111101;
assign LUT_1[52453] = 32'b00000000000000001101100110111001;
assign LUT_1[52454] = 32'b00000000000000010000000011001110;
assign LUT_1[52455] = 32'b00000000000000001001010101001010;
assign LUT_1[52456] = 32'b00000000000000001011101001011011;
assign LUT_1[52457] = 32'b00000000000000000100111011010111;
assign LUT_1[52458] = 32'b00000000000000000111010111101100;
assign LUT_1[52459] = 32'b00000000000000000000101001101000;
assign LUT_1[52460] = 32'b00000000000000010011100010110010;
assign LUT_1[52461] = 32'b00000000000000001100110100101110;
assign LUT_1[52462] = 32'b00000000000000001111010001000011;
assign LUT_1[52463] = 32'b00000000000000001000100010111111;
assign LUT_1[52464] = 32'b00000000000000001110010111001000;
assign LUT_1[52465] = 32'b00000000000000000111101001000100;
assign LUT_1[52466] = 32'b00000000000000001010000101011001;
assign LUT_1[52467] = 32'b00000000000000000011010111010101;
assign LUT_1[52468] = 32'b00000000000000010110010000011111;
assign LUT_1[52469] = 32'b00000000000000001111100010011011;
assign LUT_1[52470] = 32'b00000000000000010001111110110000;
assign LUT_1[52471] = 32'b00000000000000001011010000101100;
assign LUT_1[52472] = 32'b00000000000000001101100100111101;
assign LUT_1[52473] = 32'b00000000000000000110110110111001;
assign LUT_1[52474] = 32'b00000000000000001001010011001110;
assign LUT_1[52475] = 32'b00000000000000000010100101001010;
assign LUT_1[52476] = 32'b00000000000000010101011110010100;
assign LUT_1[52477] = 32'b00000000000000001110110000010000;
assign LUT_1[52478] = 32'b00000000000000010001001100100101;
assign LUT_1[52479] = 32'b00000000000000001010011110100001;
assign LUT_1[52480] = 32'b00000000000000000100010111001000;
assign LUT_1[52481] = 32'b11111111111111111101101001000100;
assign LUT_1[52482] = 32'b00000000000000000000000101011001;
assign LUT_1[52483] = 32'b11111111111111111001010111010101;
assign LUT_1[52484] = 32'b00000000000000001100010000011111;
assign LUT_1[52485] = 32'b00000000000000000101100010011011;
assign LUT_1[52486] = 32'b00000000000000000111111110110000;
assign LUT_1[52487] = 32'b00000000000000000001010000101100;
assign LUT_1[52488] = 32'b00000000000000000011100100111101;
assign LUT_1[52489] = 32'b11111111111111111100110110111001;
assign LUT_1[52490] = 32'b11111111111111111111010011001110;
assign LUT_1[52491] = 32'b11111111111111111000100101001010;
assign LUT_1[52492] = 32'b00000000000000001011011110010100;
assign LUT_1[52493] = 32'b00000000000000000100110000010000;
assign LUT_1[52494] = 32'b00000000000000000111001100100101;
assign LUT_1[52495] = 32'b00000000000000000000011110100001;
assign LUT_1[52496] = 32'b00000000000000000110010010101010;
assign LUT_1[52497] = 32'b11111111111111111111100100100110;
assign LUT_1[52498] = 32'b00000000000000000010000000111011;
assign LUT_1[52499] = 32'b11111111111111111011010010110111;
assign LUT_1[52500] = 32'b00000000000000001110001100000001;
assign LUT_1[52501] = 32'b00000000000000000111011101111101;
assign LUT_1[52502] = 32'b00000000000000001001111010010010;
assign LUT_1[52503] = 32'b00000000000000000011001100001110;
assign LUT_1[52504] = 32'b00000000000000000101100000011111;
assign LUT_1[52505] = 32'b11111111111111111110110010011011;
assign LUT_1[52506] = 32'b00000000000000000001001110110000;
assign LUT_1[52507] = 32'b11111111111111111010100000101100;
assign LUT_1[52508] = 32'b00000000000000001101011001110110;
assign LUT_1[52509] = 32'b00000000000000000110101011110010;
assign LUT_1[52510] = 32'b00000000000000001001001000000111;
assign LUT_1[52511] = 32'b00000000000000000010011010000011;
assign LUT_1[52512] = 32'b00000000000000000101010010000111;
assign LUT_1[52513] = 32'b11111111111111111110100100000011;
assign LUT_1[52514] = 32'b00000000000000000001000000011000;
assign LUT_1[52515] = 32'b11111111111111111010010010010100;
assign LUT_1[52516] = 32'b00000000000000001101001011011110;
assign LUT_1[52517] = 32'b00000000000000000110011101011010;
assign LUT_1[52518] = 32'b00000000000000001000111001101111;
assign LUT_1[52519] = 32'b00000000000000000010001011101011;
assign LUT_1[52520] = 32'b00000000000000000100011111111100;
assign LUT_1[52521] = 32'b11111111111111111101110001111000;
assign LUT_1[52522] = 32'b00000000000000000000001110001101;
assign LUT_1[52523] = 32'b11111111111111111001100000001001;
assign LUT_1[52524] = 32'b00000000000000001100011001010011;
assign LUT_1[52525] = 32'b00000000000000000101101011001111;
assign LUT_1[52526] = 32'b00000000000000001000000111100100;
assign LUT_1[52527] = 32'b00000000000000000001011001100000;
assign LUT_1[52528] = 32'b00000000000000000111001101101001;
assign LUT_1[52529] = 32'b00000000000000000000011111100101;
assign LUT_1[52530] = 32'b00000000000000000010111011111010;
assign LUT_1[52531] = 32'b11111111111111111100001101110110;
assign LUT_1[52532] = 32'b00000000000000001111000111000000;
assign LUT_1[52533] = 32'b00000000000000001000011000111100;
assign LUT_1[52534] = 32'b00000000000000001010110101010001;
assign LUT_1[52535] = 32'b00000000000000000100000111001101;
assign LUT_1[52536] = 32'b00000000000000000110011011011110;
assign LUT_1[52537] = 32'b11111111111111111111101101011010;
assign LUT_1[52538] = 32'b00000000000000000010001001101111;
assign LUT_1[52539] = 32'b11111111111111111011011011101011;
assign LUT_1[52540] = 32'b00000000000000001110010100110101;
assign LUT_1[52541] = 32'b00000000000000000111100110110001;
assign LUT_1[52542] = 32'b00000000000000001010000011000110;
assign LUT_1[52543] = 32'b00000000000000000011010101000010;
assign LUT_1[52544] = 32'b00000000000000000110010100110000;
assign LUT_1[52545] = 32'b11111111111111111111100110101100;
assign LUT_1[52546] = 32'b00000000000000000010000011000001;
assign LUT_1[52547] = 32'b11111111111111111011010100111101;
assign LUT_1[52548] = 32'b00000000000000001110001110000111;
assign LUT_1[52549] = 32'b00000000000000000111100000000011;
assign LUT_1[52550] = 32'b00000000000000001001111100011000;
assign LUT_1[52551] = 32'b00000000000000000011001110010100;
assign LUT_1[52552] = 32'b00000000000000000101100010100101;
assign LUT_1[52553] = 32'b11111111111111111110110100100001;
assign LUT_1[52554] = 32'b00000000000000000001010000110110;
assign LUT_1[52555] = 32'b11111111111111111010100010110010;
assign LUT_1[52556] = 32'b00000000000000001101011011111100;
assign LUT_1[52557] = 32'b00000000000000000110101101111000;
assign LUT_1[52558] = 32'b00000000000000001001001010001101;
assign LUT_1[52559] = 32'b00000000000000000010011100001001;
assign LUT_1[52560] = 32'b00000000000000001000010000010010;
assign LUT_1[52561] = 32'b00000000000000000001100010001110;
assign LUT_1[52562] = 32'b00000000000000000011111110100011;
assign LUT_1[52563] = 32'b11111111111111111101010000011111;
assign LUT_1[52564] = 32'b00000000000000010000001001101001;
assign LUT_1[52565] = 32'b00000000000000001001011011100101;
assign LUT_1[52566] = 32'b00000000000000001011110111111010;
assign LUT_1[52567] = 32'b00000000000000000101001001110110;
assign LUT_1[52568] = 32'b00000000000000000111011110000111;
assign LUT_1[52569] = 32'b00000000000000000000110000000011;
assign LUT_1[52570] = 32'b00000000000000000011001100011000;
assign LUT_1[52571] = 32'b11111111111111111100011110010100;
assign LUT_1[52572] = 32'b00000000000000001111010111011110;
assign LUT_1[52573] = 32'b00000000000000001000101001011010;
assign LUT_1[52574] = 32'b00000000000000001011000101101111;
assign LUT_1[52575] = 32'b00000000000000000100010111101011;
assign LUT_1[52576] = 32'b00000000000000000111001111101111;
assign LUT_1[52577] = 32'b00000000000000000000100001101011;
assign LUT_1[52578] = 32'b00000000000000000010111110000000;
assign LUT_1[52579] = 32'b11111111111111111100001111111100;
assign LUT_1[52580] = 32'b00000000000000001111001001000110;
assign LUT_1[52581] = 32'b00000000000000001000011011000010;
assign LUT_1[52582] = 32'b00000000000000001010110111010111;
assign LUT_1[52583] = 32'b00000000000000000100001001010011;
assign LUT_1[52584] = 32'b00000000000000000110011101100100;
assign LUT_1[52585] = 32'b11111111111111111111101111100000;
assign LUT_1[52586] = 32'b00000000000000000010001011110101;
assign LUT_1[52587] = 32'b11111111111111111011011101110001;
assign LUT_1[52588] = 32'b00000000000000001110010110111011;
assign LUT_1[52589] = 32'b00000000000000000111101000110111;
assign LUT_1[52590] = 32'b00000000000000001010000101001100;
assign LUT_1[52591] = 32'b00000000000000000011010111001000;
assign LUT_1[52592] = 32'b00000000000000001001001011010001;
assign LUT_1[52593] = 32'b00000000000000000010011101001101;
assign LUT_1[52594] = 32'b00000000000000000100111001100010;
assign LUT_1[52595] = 32'b11111111111111111110001011011110;
assign LUT_1[52596] = 32'b00000000000000010001000100101000;
assign LUT_1[52597] = 32'b00000000000000001010010110100100;
assign LUT_1[52598] = 32'b00000000000000001100110010111001;
assign LUT_1[52599] = 32'b00000000000000000110000100110101;
assign LUT_1[52600] = 32'b00000000000000001000011001000110;
assign LUT_1[52601] = 32'b00000000000000000001101011000010;
assign LUT_1[52602] = 32'b00000000000000000100000111010111;
assign LUT_1[52603] = 32'b11111111111111111101011001010011;
assign LUT_1[52604] = 32'b00000000000000010000010010011101;
assign LUT_1[52605] = 32'b00000000000000001001100100011001;
assign LUT_1[52606] = 32'b00000000000000001100000000101110;
assign LUT_1[52607] = 32'b00000000000000000101010010101010;
assign LUT_1[52608] = 32'b00000000000000000111010111001011;
assign LUT_1[52609] = 32'b00000000000000000000101001000111;
assign LUT_1[52610] = 32'b00000000000000000011000101011100;
assign LUT_1[52611] = 32'b11111111111111111100010111011000;
assign LUT_1[52612] = 32'b00000000000000001111010000100010;
assign LUT_1[52613] = 32'b00000000000000001000100010011110;
assign LUT_1[52614] = 32'b00000000000000001010111110110011;
assign LUT_1[52615] = 32'b00000000000000000100010000101111;
assign LUT_1[52616] = 32'b00000000000000000110100101000000;
assign LUT_1[52617] = 32'b11111111111111111111110110111100;
assign LUT_1[52618] = 32'b00000000000000000010010011010001;
assign LUT_1[52619] = 32'b11111111111111111011100101001101;
assign LUT_1[52620] = 32'b00000000000000001110011110010111;
assign LUT_1[52621] = 32'b00000000000000000111110000010011;
assign LUT_1[52622] = 32'b00000000000000001010001100101000;
assign LUT_1[52623] = 32'b00000000000000000011011110100100;
assign LUT_1[52624] = 32'b00000000000000001001010010101101;
assign LUT_1[52625] = 32'b00000000000000000010100100101001;
assign LUT_1[52626] = 32'b00000000000000000101000000111110;
assign LUT_1[52627] = 32'b11111111111111111110010010111010;
assign LUT_1[52628] = 32'b00000000000000010001001100000100;
assign LUT_1[52629] = 32'b00000000000000001010011110000000;
assign LUT_1[52630] = 32'b00000000000000001100111010010101;
assign LUT_1[52631] = 32'b00000000000000000110001100010001;
assign LUT_1[52632] = 32'b00000000000000001000100000100010;
assign LUT_1[52633] = 32'b00000000000000000001110010011110;
assign LUT_1[52634] = 32'b00000000000000000100001110110011;
assign LUT_1[52635] = 32'b11111111111111111101100000101111;
assign LUT_1[52636] = 32'b00000000000000010000011001111001;
assign LUT_1[52637] = 32'b00000000000000001001101011110101;
assign LUT_1[52638] = 32'b00000000000000001100001000001010;
assign LUT_1[52639] = 32'b00000000000000000101011010000110;
assign LUT_1[52640] = 32'b00000000000000001000010010001010;
assign LUT_1[52641] = 32'b00000000000000000001100100000110;
assign LUT_1[52642] = 32'b00000000000000000100000000011011;
assign LUT_1[52643] = 32'b11111111111111111101010010010111;
assign LUT_1[52644] = 32'b00000000000000010000001011100001;
assign LUT_1[52645] = 32'b00000000000000001001011101011101;
assign LUT_1[52646] = 32'b00000000000000001011111001110010;
assign LUT_1[52647] = 32'b00000000000000000101001011101110;
assign LUT_1[52648] = 32'b00000000000000000111011111111111;
assign LUT_1[52649] = 32'b00000000000000000000110001111011;
assign LUT_1[52650] = 32'b00000000000000000011001110010000;
assign LUT_1[52651] = 32'b11111111111111111100100000001100;
assign LUT_1[52652] = 32'b00000000000000001111011001010110;
assign LUT_1[52653] = 32'b00000000000000001000101011010010;
assign LUT_1[52654] = 32'b00000000000000001011000111100111;
assign LUT_1[52655] = 32'b00000000000000000100011001100011;
assign LUT_1[52656] = 32'b00000000000000001010001101101100;
assign LUT_1[52657] = 32'b00000000000000000011011111101000;
assign LUT_1[52658] = 32'b00000000000000000101111011111101;
assign LUT_1[52659] = 32'b11111111111111111111001101111001;
assign LUT_1[52660] = 32'b00000000000000010010000111000011;
assign LUT_1[52661] = 32'b00000000000000001011011000111111;
assign LUT_1[52662] = 32'b00000000000000001101110101010100;
assign LUT_1[52663] = 32'b00000000000000000111000111010000;
assign LUT_1[52664] = 32'b00000000000000001001011011100001;
assign LUT_1[52665] = 32'b00000000000000000010101101011101;
assign LUT_1[52666] = 32'b00000000000000000101001001110010;
assign LUT_1[52667] = 32'b11111111111111111110011011101110;
assign LUT_1[52668] = 32'b00000000000000010001010100111000;
assign LUT_1[52669] = 32'b00000000000000001010100110110100;
assign LUT_1[52670] = 32'b00000000000000001101000011001001;
assign LUT_1[52671] = 32'b00000000000000000110010101000101;
assign LUT_1[52672] = 32'b00000000000000001001010100110011;
assign LUT_1[52673] = 32'b00000000000000000010100110101111;
assign LUT_1[52674] = 32'b00000000000000000101000011000100;
assign LUT_1[52675] = 32'b11111111111111111110010101000000;
assign LUT_1[52676] = 32'b00000000000000010001001110001010;
assign LUT_1[52677] = 32'b00000000000000001010100000000110;
assign LUT_1[52678] = 32'b00000000000000001100111100011011;
assign LUT_1[52679] = 32'b00000000000000000110001110010111;
assign LUT_1[52680] = 32'b00000000000000001000100010101000;
assign LUT_1[52681] = 32'b00000000000000000001110100100100;
assign LUT_1[52682] = 32'b00000000000000000100010000111001;
assign LUT_1[52683] = 32'b11111111111111111101100010110101;
assign LUT_1[52684] = 32'b00000000000000010000011011111111;
assign LUT_1[52685] = 32'b00000000000000001001101101111011;
assign LUT_1[52686] = 32'b00000000000000001100001010010000;
assign LUT_1[52687] = 32'b00000000000000000101011100001100;
assign LUT_1[52688] = 32'b00000000000000001011010000010101;
assign LUT_1[52689] = 32'b00000000000000000100100010010001;
assign LUT_1[52690] = 32'b00000000000000000110111110100110;
assign LUT_1[52691] = 32'b00000000000000000000010000100010;
assign LUT_1[52692] = 32'b00000000000000010011001001101100;
assign LUT_1[52693] = 32'b00000000000000001100011011101000;
assign LUT_1[52694] = 32'b00000000000000001110110111111101;
assign LUT_1[52695] = 32'b00000000000000001000001001111001;
assign LUT_1[52696] = 32'b00000000000000001010011110001010;
assign LUT_1[52697] = 32'b00000000000000000011110000000110;
assign LUT_1[52698] = 32'b00000000000000000110001100011011;
assign LUT_1[52699] = 32'b11111111111111111111011110010111;
assign LUT_1[52700] = 32'b00000000000000010010010111100001;
assign LUT_1[52701] = 32'b00000000000000001011101001011101;
assign LUT_1[52702] = 32'b00000000000000001110000101110010;
assign LUT_1[52703] = 32'b00000000000000000111010111101110;
assign LUT_1[52704] = 32'b00000000000000001010001111110010;
assign LUT_1[52705] = 32'b00000000000000000011100001101110;
assign LUT_1[52706] = 32'b00000000000000000101111110000011;
assign LUT_1[52707] = 32'b11111111111111111111001111111111;
assign LUT_1[52708] = 32'b00000000000000010010001001001001;
assign LUT_1[52709] = 32'b00000000000000001011011011000101;
assign LUT_1[52710] = 32'b00000000000000001101110111011010;
assign LUT_1[52711] = 32'b00000000000000000111001001010110;
assign LUT_1[52712] = 32'b00000000000000001001011101100111;
assign LUT_1[52713] = 32'b00000000000000000010101111100011;
assign LUT_1[52714] = 32'b00000000000000000101001011111000;
assign LUT_1[52715] = 32'b11111111111111111110011101110100;
assign LUT_1[52716] = 32'b00000000000000010001010110111110;
assign LUT_1[52717] = 32'b00000000000000001010101000111010;
assign LUT_1[52718] = 32'b00000000000000001101000101001111;
assign LUT_1[52719] = 32'b00000000000000000110010111001011;
assign LUT_1[52720] = 32'b00000000000000001100001011010100;
assign LUT_1[52721] = 32'b00000000000000000101011101010000;
assign LUT_1[52722] = 32'b00000000000000000111111001100101;
assign LUT_1[52723] = 32'b00000000000000000001001011100001;
assign LUT_1[52724] = 32'b00000000000000010100000100101011;
assign LUT_1[52725] = 32'b00000000000000001101010110100111;
assign LUT_1[52726] = 32'b00000000000000001111110010111100;
assign LUT_1[52727] = 32'b00000000000000001001000100111000;
assign LUT_1[52728] = 32'b00000000000000001011011001001001;
assign LUT_1[52729] = 32'b00000000000000000100101011000101;
assign LUT_1[52730] = 32'b00000000000000000111000111011010;
assign LUT_1[52731] = 32'b00000000000000000000011001010110;
assign LUT_1[52732] = 32'b00000000000000010011010010100000;
assign LUT_1[52733] = 32'b00000000000000001100100100011100;
assign LUT_1[52734] = 32'b00000000000000001111000000110001;
assign LUT_1[52735] = 32'b00000000000000001000010010101101;
assign LUT_1[52736] = 32'b00000000000000000000010001011001;
assign LUT_1[52737] = 32'b11111111111111111001100011010101;
assign LUT_1[52738] = 32'b11111111111111111011111111101010;
assign LUT_1[52739] = 32'b11111111111111110101010001100110;
assign LUT_1[52740] = 32'b00000000000000001000001010110000;
assign LUT_1[52741] = 32'b00000000000000000001011100101100;
assign LUT_1[52742] = 32'b00000000000000000011111001000001;
assign LUT_1[52743] = 32'b11111111111111111101001010111101;
assign LUT_1[52744] = 32'b11111111111111111111011111001110;
assign LUT_1[52745] = 32'b11111111111111111000110001001010;
assign LUT_1[52746] = 32'b11111111111111111011001101011111;
assign LUT_1[52747] = 32'b11111111111111110100011111011011;
assign LUT_1[52748] = 32'b00000000000000000111011000100101;
assign LUT_1[52749] = 32'b00000000000000000000101010100001;
assign LUT_1[52750] = 32'b00000000000000000011000110110110;
assign LUT_1[52751] = 32'b11111111111111111100011000110010;
assign LUT_1[52752] = 32'b00000000000000000010001100111011;
assign LUT_1[52753] = 32'b11111111111111111011011110110111;
assign LUT_1[52754] = 32'b11111111111111111101111011001100;
assign LUT_1[52755] = 32'b11111111111111110111001101001000;
assign LUT_1[52756] = 32'b00000000000000001010000110010010;
assign LUT_1[52757] = 32'b00000000000000000011011000001110;
assign LUT_1[52758] = 32'b00000000000000000101110100100011;
assign LUT_1[52759] = 32'b11111111111111111111000110011111;
assign LUT_1[52760] = 32'b00000000000000000001011010110000;
assign LUT_1[52761] = 32'b11111111111111111010101100101100;
assign LUT_1[52762] = 32'b11111111111111111101001001000001;
assign LUT_1[52763] = 32'b11111111111111110110011010111101;
assign LUT_1[52764] = 32'b00000000000000001001010100000111;
assign LUT_1[52765] = 32'b00000000000000000010100110000011;
assign LUT_1[52766] = 32'b00000000000000000101000010011000;
assign LUT_1[52767] = 32'b11111111111111111110010100010100;
assign LUT_1[52768] = 32'b00000000000000000001001100011000;
assign LUT_1[52769] = 32'b11111111111111111010011110010100;
assign LUT_1[52770] = 32'b11111111111111111100111010101001;
assign LUT_1[52771] = 32'b11111111111111110110001100100101;
assign LUT_1[52772] = 32'b00000000000000001001000101101111;
assign LUT_1[52773] = 32'b00000000000000000010010111101011;
assign LUT_1[52774] = 32'b00000000000000000100110100000000;
assign LUT_1[52775] = 32'b11111111111111111110000101111100;
assign LUT_1[52776] = 32'b00000000000000000000011010001101;
assign LUT_1[52777] = 32'b11111111111111111001101100001001;
assign LUT_1[52778] = 32'b11111111111111111100001000011110;
assign LUT_1[52779] = 32'b11111111111111110101011010011010;
assign LUT_1[52780] = 32'b00000000000000001000010011100100;
assign LUT_1[52781] = 32'b00000000000000000001100101100000;
assign LUT_1[52782] = 32'b00000000000000000100000001110101;
assign LUT_1[52783] = 32'b11111111111111111101010011110001;
assign LUT_1[52784] = 32'b00000000000000000011000111111010;
assign LUT_1[52785] = 32'b11111111111111111100011001110110;
assign LUT_1[52786] = 32'b11111111111111111110110110001011;
assign LUT_1[52787] = 32'b11111111111111111000001000000111;
assign LUT_1[52788] = 32'b00000000000000001011000001010001;
assign LUT_1[52789] = 32'b00000000000000000100010011001101;
assign LUT_1[52790] = 32'b00000000000000000110101111100010;
assign LUT_1[52791] = 32'b00000000000000000000000001011110;
assign LUT_1[52792] = 32'b00000000000000000010010101101111;
assign LUT_1[52793] = 32'b11111111111111111011100111101011;
assign LUT_1[52794] = 32'b11111111111111111110000100000000;
assign LUT_1[52795] = 32'b11111111111111110111010101111100;
assign LUT_1[52796] = 32'b00000000000000001010001111000110;
assign LUT_1[52797] = 32'b00000000000000000011100001000010;
assign LUT_1[52798] = 32'b00000000000000000101111101010111;
assign LUT_1[52799] = 32'b11111111111111111111001111010011;
assign LUT_1[52800] = 32'b00000000000000000010001111000001;
assign LUT_1[52801] = 32'b11111111111111111011100000111101;
assign LUT_1[52802] = 32'b11111111111111111101111101010010;
assign LUT_1[52803] = 32'b11111111111111110111001111001110;
assign LUT_1[52804] = 32'b00000000000000001010001000011000;
assign LUT_1[52805] = 32'b00000000000000000011011010010100;
assign LUT_1[52806] = 32'b00000000000000000101110110101001;
assign LUT_1[52807] = 32'b11111111111111111111001000100101;
assign LUT_1[52808] = 32'b00000000000000000001011100110110;
assign LUT_1[52809] = 32'b11111111111111111010101110110010;
assign LUT_1[52810] = 32'b11111111111111111101001011000111;
assign LUT_1[52811] = 32'b11111111111111110110011101000011;
assign LUT_1[52812] = 32'b00000000000000001001010110001101;
assign LUT_1[52813] = 32'b00000000000000000010101000001001;
assign LUT_1[52814] = 32'b00000000000000000101000100011110;
assign LUT_1[52815] = 32'b11111111111111111110010110011010;
assign LUT_1[52816] = 32'b00000000000000000100001010100011;
assign LUT_1[52817] = 32'b11111111111111111101011100011111;
assign LUT_1[52818] = 32'b11111111111111111111111000110100;
assign LUT_1[52819] = 32'b11111111111111111001001010110000;
assign LUT_1[52820] = 32'b00000000000000001100000011111010;
assign LUT_1[52821] = 32'b00000000000000000101010101110110;
assign LUT_1[52822] = 32'b00000000000000000111110010001011;
assign LUT_1[52823] = 32'b00000000000000000001000100000111;
assign LUT_1[52824] = 32'b00000000000000000011011000011000;
assign LUT_1[52825] = 32'b11111111111111111100101010010100;
assign LUT_1[52826] = 32'b11111111111111111111000110101001;
assign LUT_1[52827] = 32'b11111111111111111000011000100101;
assign LUT_1[52828] = 32'b00000000000000001011010001101111;
assign LUT_1[52829] = 32'b00000000000000000100100011101011;
assign LUT_1[52830] = 32'b00000000000000000111000000000000;
assign LUT_1[52831] = 32'b00000000000000000000010001111100;
assign LUT_1[52832] = 32'b00000000000000000011001010000000;
assign LUT_1[52833] = 32'b11111111111111111100011011111100;
assign LUT_1[52834] = 32'b11111111111111111110111000010001;
assign LUT_1[52835] = 32'b11111111111111111000001010001101;
assign LUT_1[52836] = 32'b00000000000000001011000011010111;
assign LUT_1[52837] = 32'b00000000000000000100010101010011;
assign LUT_1[52838] = 32'b00000000000000000110110001101000;
assign LUT_1[52839] = 32'b00000000000000000000000011100100;
assign LUT_1[52840] = 32'b00000000000000000010010111110101;
assign LUT_1[52841] = 32'b11111111111111111011101001110001;
assign LUT_1[52842] = 32'b11111111111111111110000110000110;
assign LUT_1[52843] = 32'b11111111111111110111011000000010;
assign LUT_1[52844] = 32'b00000000000000001010010001001100;
assign LUT_1[52845] = 32'b00000000000000000011100011001000;
assign LUT_1[52846] = 32'b00000000000000000101111111011101;
assign LUT_1[52847] = 32'b11111111111111111111010001011001;
assign LUT_1[52848] = 32'b00000000000000000101000101100010;
assign LUT_1[52849] = 32'b11111111111111111110010111011110;
assign LUT_1[52850] = 32'b00000000000000000000110011110011;
assign LUT_1[52851] = 32'b11111111111111111010000101101111;
assign LUT_1[52852] = 32'b00000000000000001100111110111001;
assign LUT_1[52853] = 32'b00000000000000000110010000110101;
assign LUT_1[52854] = 32'b00000000000000001000101101001010;
assign LUT_1[52855] = 32'b00000000000000000001111111000110;
assign LUT_1[52856] = 32'b00000000000000000100010011010111;
assign LUT_1[52857] = 32'b11111111111111111101100101010011;
assign LUT_1[52858] = 32'b00000000000000000000000001101000;
assign LUT_1[52859] = 32'b11111111111111111001010011100100;
assign LUT_1[52860] = 32'b00000000000000001100001100101110;
assign LUT_1[52861] = 32'b00000000000000000101011110101010;
assign LUT_1[52862] = 32'b00000000000000000111111010111111;
assign LUT_1[52863] = 32'b00000000000000000001001100111011;
assign LUT_1[52864] = 32'b00000000000000000011010001011100;
assign LUT_1[52865] = 32'b11111111111111111100100011011000;
assign LUT_1[52866] = 32'b11111111111111111110111111101101;
assign LUT_1[52867] = 32'b11111111111111111000010001101001;
assign LUT_1[52868] = 32'b00000000000000001011001010110011;
assign LUT_1[52869] = 32'b00000000000000000100011100101111;
assign LUT_1[52870] = 32'b00000000000000000110111001000100;
assign LUT_1[52871] = 32'b00000000000000000000001011000000;
assign LUT_1[52872] = 32'b00000000000000000010011111010001;
assign LUT_1[52873] = 32'b11111111111111111011110001001101;
assign LUT_1[52874] = 32'b11111111111111111110001101100010;
assign LUT_1[52875] = 32'b11111111111111110111011111011110;
assign LUT_1[52876] = 32'b00000000000000001010011000101000;
assign LUT_1[52877] = 32'b00000000000000000011101010100100;
assign LUT_1[52878] = 32'b00000000000000000110000110111001;
assign LUT_1[52879] = 32'b11111111111111111111011000110101;
assign LUT_1[52880] = 32'b00000000000000000101001100111110;
assign LUT_1[52881] = 32'b11111111111111111110011110111010;
assign LUT_1[52882] = 32'b00000000000000000000111011001111;
assign LUT_1[52883] = 32'b11111111111111111010001101001011;
assign LUT_1[52884] = 32'b00000000000000001101000110010101;
assign LUT_1[52885] = 32'b00000000000000000110011000010001;
assign LUT_1[52886] = 32'b00000000000000001000110100100110;
assign LUT_1[52887] = 32'b00000000000000000010000110100010;
assign LUT_1[52888] = 32'b00000000000000000100011010110011;
assign LUT_1[52889] = 32'b11111111111111111101101100101111;
assign LUT_1[52890] = 32'b00000000000000000000001001000100;
assign LUT_1[52891] = 32'b11111111111111111001011011000000;
assign LUT_1[52892] = 32'b00000000000000001100010100001010;
assign LUT_1[52893] = 32'b00000000000000000101100110000110;
assign LUT_1[52894] = 32'b00000000000000001000000010011011;
assign LUT_1[52895] = 32'b00000000000000000001010100010111;
assign LUT_1[52896] = 32'b00000000000000000100001100011011;
assign LUT_1[52897] = 32'b11111111111111111101011110010111;
assign LUT_1[52898] = 32'b11111111111111111111111010101100;
assign LUT_1[52899] = 32'b11111111111111111001001100101000;
assign LUT_1[52900] = 32'b00000000000000001100000101110010;
assign LUT_1[52901] = 32'b00000000000000000101010111101110;
assign LUT_1[52902] = 32'b00000000000000000111110100000011;
assign LUT_1[52903] = 32'b00000000000000000001000101111111;
assign LUT_1[52904] = 32'b00000000000000000011011010010000;
assign LUT_1[52905] = 32'b11111111111111111100101100001100;
assign LUT_1[52906] = 32'b11111111111111111111001000100001;
assign LUT_1[52907] = 32'b11111111111111111000011010011101;
assign LUT_1[52908] = 32'b00000000000000001011010011100111;
assign LUT_1[52909] = 32'b00000000000000000100100101100011;
assign LUT_1[52910] = 32'b00000000000000000111000001111000;
assign LUT_1[52911] = 32'b00000000000000000000010011110100;
assign LUT_1[52912] = 32'b00000000000000000110000111111101;
assign LUT_1[52913] = 32'b11111111111111111111011001111001;
assign LUT_1[52914] = 32'b00000000000000000001110110001110;
assign LUT_1[52915] = 32'b11111111111111111011001000001010;
assign LUT_1[52916] = 32'b00000000000000001110000001010100;
assign LUT_1[52917] = 32'b00000000000000000111010011010000;
assign LUT_1[52918] = 32'b00000000000000001001101111100101;
assign LUT_1[52919] = 32'b00000000000000000011000001100001;
assign LUT_1[52920] = 32'b00000000000000000101010101110010;
assign LUT_1[52921] = 32'b11111111111111111110100111101110;
assign LUT_1[52922] = 32'b00000000000000000001000100000011;
assign LUT_1[52923] = 32'b11111111111111111010010101111111;
assign LUT_1[52924] = 32'b00000000000000001101001111001001;
assign LUT_1[52925] = 32'b00000000000000000110100001000101;
assign LUT_1[52926] = 32'b00000000000000001000111101011010;
assign LUT_1[52927] = 32'b00000000000000000010001111010110;
assign LUT_1[52928] = 32'b00000000000000000101001111000100;
assign LUT_1[52929] = 32'b11111111111111111110100001000000;
assign LUT_1[52930] = 32'b00000000000000000000111101010101;
assign LUT_1[52931] = 32'b11111111111111111010001111010001;
assign LUT_1[52932] = 32'b00000000000000001101001000011011;
assign LUT_1[52933] = 32'b00000000000000000110011010010111;
assign LUT_1[52934] = 32'b00000000000000001000110110101100;
assign LUT_1[52935] = 32'b00000000000000000010001000101000;
assign LUT_1[52936] = 32'b00000000000000000100011100111001;
assign LUT_1[52937] = 32'b11111111111111111101101110110101;
assign LUT_1[52938] = 32'b00000000000000000000001011001010;
assign LUT_1[52939] = 32'b11111111111111111001011101000110;
assign LUT_1[52940] = 32'b00000000000000001100010110010000;
assign LUT_1[52941] = 32'b00000000000000000101101000001100;
assign LUT_1[52942] = 32'b00000000000000001000000100100001;
assign LUT_1[52943] = 32'b00000000000000000001010110011101;
assign LUT_1[52944] = 32'b00000000000000000111001010100110;
assign LUT_1[52945] = 32'b00000000000000000000011100100010;
assign LUT_1[52946] = 32'b00000000000000000010111000110111;
assign LUT_1[52947] = 32'b11111111111111111100001010110011;
assign LUT_1[52948] = 32'b00000000000000001111000011111101;
assign LUT_1[52949] = 32'b00000000000000001000010101111001;
assign LUT_1[52950] = 32'b00000000000000001010110010001110;
assign LUT_1[52951] = 32'b00000000000000000100000100001010;
assign LUT_1[52952] = 32'b00000000000000000110011000011011;
assign LUT_1[52953] = 32'b11111111111111111111101010010111;
assign LUT_1[52954] = 32'b00000000000000000010000110101100;
assign LUT_1[52955] = 32'b11111111111111111011011000101000;
assign LUT_1[52956] = 32'b00000000000000001110010001110010;
assign LUT_1[52957] = 32'b00000000000000000111100011101110;
assign LUT_1[52958] = 32'b00000000000000001010000000000011;
assign LUT_1[52959] = 32'b00000000000000000011010001111111;
assign LUT_1[52960] = 32'b00000000000000000110001010000011;
assign LUT_1[52961] = 32'b11111111111111111111011011111111;
assign LUT_1[52962] = 32'b00000000000000000001111000010100;
assign LUT_1[52963] = 32'b11111111111111111011001010010000;
assign LUT_1[52964] = 32'b00000000000000001110000011011010;
assign LUT_1[52965] = 32'b00000000000000000111010101010110;
assign LUT_1[52966] = 32'b00000000000000001001110001101011;
assign LUT_1[52967] = 32'b00000000000000000011000011100111;
assign LUT_1[52968] = 32'b00000000000000000101010111111000;
assign LUT_1[52969] = 32'b11111111111111111110101001110100;
assign LUT_1[52970] = 32'b00000000000000000001000110001001;
assign LUT_1[52971] = 32'b11111111111111111010011000000101;
assign LUT_1[52972] = 32'b00000000000000001101010001001111;
assign LUT_1[52973] = 32'b00000000000000000110100011001011;
assign LUT_1[52974] = 32'b00000000000000001000111111100000;
assign LUT_1[52975] = 32'b00000000000000000010010001011100;
assign LUT_1[52976] = 32'b00000000000000001000000101100101;
assign LUT_1[52977] = 32'b00000000000000000001010111100001;
assign LUT_1[52978] = 32'b00000000000000000011110011110110;
assign LUT_1[52979] = 32'b11111111111111111101000101110010;
assign LUT_1[52980] = 32'b00000000000000001111111110111100;
assign LUT_1[52981] = 32'b00000000000000001001010000111000;
assign LUT_1[52982] = 32'b00000000000000001011101101001101;
assign LUT_1[52983] = 32'b00000000000000000100111111001001;
assign LUT_1[52984] = 32'b00000000000000000111010011011010;
assign LUT_1[52985] = 32'b00000000000000000000100101010110;
assign LUT_1[52986] = 32'b00000000000000000011000001101011;
assign LUT_1[52987] = 32'b11111111111111111100010011100111;
assign LUT_1[52988] = 32'b00000000000000001111001100110001;
assign LUT_1[52989] = 32'b00000000000000001000011110101101;
assign LUT_1[52990] = 32'b00000000000000001010111011000010;
assign LUT_1[52991] = 32'b00000000000000000100001100111110;
assign LUT_1[52992] = 32'b11111111111111111110000101100101;
assign LUT_1[52993] = 32'b11111111111111110111010111100001;
assign LUT_1[52994] = 32'b11111111111111111001110011110110;
assign LUT_1[52995] = 32'b11111111111111110011000101110010;
assign LUT_1[52996] = 32'b00000000000000000101111110111100;
assign LUT_1[52997] = 32'b11111111111111111111010000111000;
assign LUT_1[52998] = 32'b00000000000000000001101101001101;
assign LUT_1[52999] = 32'b11111111111111111010111111001001;
assign LUT_1[53000] = 32'b11111111111111111101010011011010;
assign LUT_1[53001] = 32'b11111111111111110110100101010110;
assign LUT_1[53002] = 32'b11111111111111111001000001101011;
assign LUT_1[53003] = 32'b11111111111111110010010011100111;
assign LUT_1[53004] = 32'b00000000000000000101001100110001;
assign LUT_1[53005] = 32'b11111111111111111110011110101101;
assign LUT_1[53006] = 32'b00000000000000000000111011000010;
assign LUT_1[53007] = 32'b11111111111111111010001100111110;
assign LUT_1[53008] = 32'b00000000000000000000000001000111;
assign LUT_1[53009] = 32'b11111111111111111001010011000011;
assign LUT_1[53010] = 32'b11111111111111111011101111011000;
assign LUT_1[53011] = 32'b11111111111111110101000001010100;
assign LUT_1[53012] = 32'b00000000000000000111111010011110;
assign LUT_1[53013] = 32'b00000000000000000001001100011010;
assign LUT_1[53014] = 32'b00000000000000000011101000101111;
assign LUT_1[53015] = 32'b11111111111111111100111010101011;
assign LUT_1[53016] = 32'b11111111111111111111001110111100;
assign LUT_1[53017] = 32'b11111111111111111000100000111000;
assign LUT_1[53018] = 32'b11111111111111111010111101001101;
assign LUT_1[53019] = 32'b11111111111111110100001111001001;
assign LUT_1[53020] = 32'b00000000000000000111001000010011;
assign LUT_1[53021] = 32'b00000000000000000000011010001111;
assign LUT_1[53022] = 32'b00000000000000000010110110100100;
assign LUT_1[53023] = 32'b11111111111111111100001000100000;
assign LUT_1[53024] = 32'b11111111111111111111000000100100;
assign LUT_1[53025] = 32'b11111111111111111000010010100000;
assign LUT_1[53026] = 32'b11111111111111111010101110110101;
assign LUT_1[53027] = 32'b11111111111111110100000000110001;
assign LUT_1[53028] = 32'b00000000000000000110111001111011;
assign LUT_1[53029] = 32'b00000000000000000000001011110111;
assign LUT_1[53030] = 32'b00000000000000000010101000001100;
assign LUT_1[53031] = 32'b11111111111111111011111010001000;
assign LUT_1[53032] = 32'b11111111111111111110001110011001;
assign LUT_1[53033] = 32'b11111111111111110111100000010101;
assign LUT_1[53034] = 32'b11111111111111111001111100101010;
assign LUT_1[53035] = 32'b11111111111111110011001110100110;
assign LUT_1[53036] = 32'b00000000000000000110000111110000;
assign LUT_1[53037] = 32'b11111111111111111111011001101100;
assign LUT_1[53038] = 32'b00000000000000000001110110000001;
assign LUT_1[53039] = 32'b11111111111111111011000111111101;
assign LUT_1[53040] = 32'b00000000000000000000111100000110;
assign LUT_1[53041] = 32'b11111111111111111010001110000010;
assign LUT_1[53042] = 32'b11111111111111111100101010010111;
assign LUT_1[53043] = 32'b11111111111111110101111100010011;
assign LUT_1[53044] = 32'b00000000000000001000110101011101;
assign LUT_1[53045] = 32'b00000000000000000010000111011001;
assign LUT_1[53046] = 32'b00000000000000000100100011101110;
assign LUT_1[53047] = 32'b11111111111111111101110101101010;
assign LUT_1[53048] = 32'b00000000000000000000001001111011;
assign LUT_1[53049] = 32'b11111111111111111001011011110111;
assign LUT_1[53050] = 32'b11111111111111111011111000001100;
assign LUT_1[53051] = 32'b11111111111111110101001010001000;
assign LUT_1[53052] = 32'b00000000000000001000000011010010;
assign LUT_1[53053] = 32'b00000000000000000001010101001110;
assign LUT_1[53054] = 32'b00000000000000000011110001100011;
assign LUT_1[53055] = 32'b11111111111111111101000011011111;
assign LUT_1[53056] = 32'b00000000000000000000000011001101;
assign LUT_1[53057] = 32'b11111111111111111001010101001001;
assign LUT_1[53058] = 32'b11111111111111111011110001011110;
assign LUT_1[53059] = 32'b11111111111111110101000011011010;
assign LUT_1[53060] = 32'b00000000000000000111111100100100;
assign LUT_1[53061] = 32'b00000000000000000001001110100000;
assign LUT_1[53062] = 32'b00000000000000000011101010110101;
assign LUT_1[53063] = 32'b11111111111111111100111100110001;
assign LUT_1[53064] = 32'b11111111111111111111010001000010;
assign LUT_1[53065] = 32'b11111111111111111000100010111110;
assign LUT_1[53066] = 32'b11111111111111111010111111010011;
assign LUT_1[53067] = 32'b11111111111111110100010001001111;
assign LUT_1[53068] = 32'b00000000000000000111001010011001;
assign LUT_1[53069] = 32'b00000000000000000000011100010101;
assign LUT_1[53070] = 32'b00000000000000000010111000101010;
assign LUT_1[53071] = 32'b11111111111111111100001010100110;
assign LUT_1[53072] = 32'b00000000000000000001111110101111;
assign LUT_1[53073] = 32'b11111111111111111011010000101011;
assign LUT_1[53074] = 32'b11111111111111111101101101000000;
assign LUT_1[53075] = 32'b11111111111111110110111110111100;
assign LUT_1[53076] = 32'b00000000000000001001111000000110;
assign LUT_1[53077] = 32'b00000000000000000011001010000010;
assign LUT_1[53078] = 32'b00000000000000000101100110010111;
assign LUT_1[53079] = 32'b11111111111111111110111000010011;
assign LUT_1[53080] = 32'b00000000000000000001001100100100;
assign LUT_1[53081] = 32'b11111111111111111010011110100000;
assign LUT_1[53082] = 32'b11111111111111111100111010110101;
assign LUT_1[53083] = 32'b11111111111111110110001100110001;
assign LUT_1[53084] = 32'b00000000000000001001000101111011;
assign LUT_1[53085] = 32'b00000000000000000010010111110111;
assign LUT_1[53086] = 32'b00000000000000000100110100001100;
assign LUT_1[53087] = 32'b11111111111111111110000110001000;
assign LUT_1[53088] = 32'b00000000000000000000111110001100;
assign LUT_1[53089] = 32'b11111111111111111010010000001000;
assign LUT_1[53090] = 32'b11111111111111111100101100011101;
assign LUT_1[53091] = 32'b11111111111111110101111110011001;
assign LUT_1[53092] = 32'b00000000000000001000110111100011;
assign LUT_1[53093] = 32'b00000000000000000010001001011111;
assign LUT_1[53094] = 32'b00000000000000000100100101110100;
assign LUT_1[53095] = 32'b11111111111111111101110111110000;
assign LUT_1[53096] = 32'b00000000000000000000001100000001;
assign LUT_1[53097] = 32'b11111111111111111001011101111101;
assign LUT_1[53098] = 32'b11111111111111111011111010010010;
assign LUT_1[53099] = 32'b11111111111111110101001100001110;
assign LUT_1[53100] = 32'b00000000000000001000000101011000;
assign LUT_1[53101] = 32'b00000000000000000001010111010100;
assign LUT_1[53102] = 32'b00000000000000000011110011101001;
assign LUT_1[53103] = 32'b11111111111111111101000101100101;
assign LUT_1[53104] = 32'b00000000000000000010111001101110;
assign LUT_1[53105] = 32'b11111111111111111100001011101010;
assign LUT_1[53106] = 32'b11111111111111111110100111111111;
assign LUT_1[53107] = 32'b11111111111111110111111001111011;
assign LUT_1[53108] = 32'b00000000000000001010110011000101;
assign LUT_1[53109] = 32'b00000000000000000100000101000001;
assign LUT_1[53110] = 32'b00000000000000000110100001010110;
assign LUT_1[53111] = 32'b11111111111111111111110011010010;
assign LUT_1[53112] = 32'b00000000000000000010000111100011;
assign LUT_1[53113] = 32'b11111111111111111011011001011111;
assign LUT_1[53114] = 32'b11111111111111111101110101110100;
assign LUT_1[53115] = 32'b11111111111111110111000111110000;
assign LUT_1[53116] = 32'b00000000000000001010000000111010;
assign LUT_1[53117] = 32'b00000000000000000011010010110110;
assign LUT_1[53118] = 32'b00000000000000000101101111001011;
assign LUT_1[53119] = 32'b11111111111111111111000001000111;
assign LUT_1[53120] = 32'b00000000000000000001000101101000;
assign LUT_1[53121] = 32'b11111111111111111010010111100100;
assign LUT_1[53122] = 32'b11111111111111111100110011111001;
assign LUT_1[53123] = 32'b11111111111111110110000101110101;
assign LUT_1[53124] = 32'b00000000000000001000111110111111;
assign LUT_1[53125] = 32'b00000000000000000010010000111011;
assign LUT_1[53126] = 32'b00000000000000000100101101010000;
assign LUT_1[53127] = 32'b11111111111111111101111111001100;
assign LUT_1[53128] = 32'b00000000000000000000010011011101;
assign LUT_1[53129] = 32'b11111111111111111001100101011001;
assign LUT_1[53130] = 32'b11111111111111111100000001101110;
assign LUT_1[53131] = 32'b11111111111111110101010011101010;
assign LUT_1[53132] = 32'b00000000000000001000001100110100;
assign LUT_1[53133] = 32'b00000000000000000001011110110000;
assign LUT_1[53134] = 32'b00000000000000000011111011000101;
assign LUT_1[53135] = 32'b11111111111111111101001101000001;
assign LUT_1[53136] = 32'b00000000000000000011000001001010;
assign LUT_1[53137] = 32'b11111111111111111100010011000110;
assign LUT_1[53138] = 32'b11111111111111111110101111011011;
assign LUT_1[53139] = 32'b11111111111111111000000001010111;
assign LUT_1[53140] = 32'b00000000000000001010111010100001;
assign LUT_1[53141] = 32'b00000000000000000100001100011101;
assign LUT_1[53142] = 32'b00000000000000000110101000110010;
assign LUT_1[53143] = 32'b11111111111111111111111010101110;
assign LUT_1[53144] = 32'b00000000000000000010001110111111;
assign LUT_1[53145] = 32'b11111111111111111011100000111011;
assign LUT_1[53146] = 32'b11111111111111111101111101010000;
assign LUT_1[53147] = 32'b11111111111111110111001111001100;
assign LUT_1[53148] = 32'b00000000000000001010001000010110;
assign LUT_1[53149] = 32'b00000000000000000011011010010010;
assign LUT_1[53150] = 32'b00000000000000000101110110100111;
assign LUT_1[53151] = 32'b11111111111111111111001000100011;
assign LUT_1[53152] = 32'b00000000000000000010000000100111;
assign LUT_1[53153] = 32'b11111111111111111011010010100011;
assign LUT_1[53154] = 32'b11111111111111111101101110111000;
assign LUT_1[53155] = 32'b11111111111111110111000000110100;
assign LUT_1[53156] = 32'b00000000000000001001111001111110;
assign LUT_1[53157] = 32'b00000000000000000011001011111010;
assign LUT_1[53158] = 32'b00000000000000000101101000001111;
assign LUT_1[53159] = 32'b11111111111111111110111010001011;
assign LUT_1[53160] = 32'b00000000000000000001001110011100;
assign LUT_1[53161] = 32'b11111111111111111010100000011000;
assign LUT_1[53162] = 32'b11111111111111111100111100101101;
assign LUT_1[53163] = 32'b11111111111111110110001110101001;
assign LUT_1[53164] = 32'b00000000000000001001000111110011;
assign LUT_1[53165] = 32'b00000000000000000010011001101111;
assign LUT_1[53166] = 32'b00000000000000000100110110000100;
assign LUT_1[53167] = 32'b11111111111111111110001000000000;
assign LUT_1[53168] = 32'b00000000000000000011111100001001;
assign LUT_1[53169] = 32'b11111111111111111101001110000101;
assign LUT_1[53170] = 32'b11111111111111111111101010011010;
assign LUT_1[53171] = 32'b11111111111111111000111100010110;
assign LUT_1[53172] = 32'b00000000000000001011110101100000;
assign LUT_1[53173] = 32'b00000000000000000101000111011100;
assign LUT_1[53174] = 32'b00000000000000000111100011110001;
assign LUT_1[53175] = 32'b00000000000000000000110101101101;
assign LUT_1[53176] = 32'b00000000000000000011001001111110;
assign LUT_1[53177] = 32'b11111111111111111100011011111010;
assign LUT_1[53178] = 32'b11111111111111111110111000001111;
assign LUT_1[53179] = 32'b11111111111111111000001010001011;
assign LUT_1[53180] = 32'b00000000000000001011000011010101;
assign LUT_1[53181] = 32'b00000000000000000100010101010001;
assign LUT_1[53182] = 32'b00000000000000000110110001100110;
assign LUT_1[53183] = 32'b00000000000000000000000011100010;
assign LUT_1[53184] = 32'b00000000000000000011000011010000;
assign LUT_1[53185] = 32'b11111111111111111100010101001100;
assign LUT_1[53186] = 32'b11111111111111111110110001100001;
assign LUT_1[53187] = 32'b11111111111111111000000011011101;
assign LUT_1[53188] = 32'b00000000000000001010111100100111;
assign LUT_1[53189] = 32'b00000000000000000100001110100011;
assign LUT_1[53190] = 32'b00000000000000000110101010111000;
assign LUT_1[53191] = 32'b11111111111111111111111100110100;
assign LUT_1[53192] = 32'b00000000000000000010010001000101;
assign LUT_1[53193] = 32'b11111111111111111011100011000001;
assign LUT_1[53194] = 32'b11111111111111111101111111010110;
assign LUT_1[53195] = 32'b11111111111111110111010001010010;
assign LUT_1[53196] = 32'b00000000000000001010001010011100;
assign LUT_1[53197] = 32'b00000000000000000011011100011000;
assign LUT_1[53198] = 32'b00000000000000000101111000101101;
assign LUT_1[53199] = 32'b11111111111111111111001010101001;
assign LUT_1[53200] = 32'b00000000000000000100111110110010;
assign LUT_1[53201] = 32'b11111111111111111110010000101110;
assign LUT_1[53202] = 32'b00000000000000000000101101000011;
assign LUT_1[53203] = 32'b11111111111111111001111110111111;
assign LUT_1[53204] = 32'b00000000000000001100111000001001;
assign LUT_1[53205] = 32'b00000000000000000110001010000101;
assign LUT_1[53206] = 32'b00000000000000001000100110011010;
assign LUT_1[53207] = 32'b00000000000000000001111000010110;
assign LUT_1[53208] = 32'b00000000000000000100001100100111;
assign LUT_1[53209] = 32'b11111111111111111101011110100011;
assign LUT_1[53210] = 32'b11111111111111111111111010111000;
assign LUT_1[53211] = 32'b11111111111111111001001100110100;
assign LUT_1[53212] = 32'b00000000000000001100000101111110;
assign LUT_1[53213] = 32'b00000000000000000101010111111010;
assign LUT_1[53214] = 32'b00000000000000000111110100001111;
assign LUT_1[53215] = 32'b00000000000000000001000110001011;
assign LUT_1[53216] = 32'b00000000000000000011111110001111;
assign LUT_1[53217] = 32'b11111111111111111101010000001011;
assign LUT_1[53218] = 32'b11111111111111111111101100100000;
assign LUT_1[53219] = 32'b11111111111111111000111110011100;
assign LUT_1[53220] = 32'b00000000000000001011110111100110;
assign LUT_1[53221] = 32'b00000000000000000101001001100010;
assign LUT_1[53222] = 32'b00000000000000000111100101110111;
assign LUT_1[53223] = 32'b00000000000000000000110111110011;
assign LUT_1[53224] = 32'b00000000000000000011001100000100;
assign LUT_1[53225] = 32'b11111111111111111100011110000000;
assign LUT_1[53226] = 32'b11111111111111111110111010010101;
assign LUT_1[53227] = 32'b11111111111111111000001100010001;
assign LUT_1[53228] = 32'b00000000000000001011000101011011;
assign LUT_1[53229] = 32'b00000000000000000100010111010111;
assign LUT_1[53230] = 32'b00000000000000000110110011101100;
assign LUT_1[53231] = 32'b00000000000000000000000101101000;
assign LUT_1[53232] = 32'b00000000000000000101111001110001;
assign LUT_1[53233] = 32'b11111111111111111111001011101101;
assign LUT_1[53234] = 32'b00000000000000000001101000000010;
assign LUT_1[53235] = 32'b11111111111111111010111001111110;
assign LUT_1[53236] = 32'b00000000000000001101110011001000;
assign LUT_1[53237] = 32'b00000000000000000111000101000100;
assign LUT_1[53238] = 32'b00000000000000001001100001011001;
assign LUT_1[53239] = 32'b00000000000000000010110011010101;
assign LUT_1[53240] = 32'b00000000000000000101000111100110;
assign LUT_1[53241] = 32'b11111111111111111110011001100010;
assign LUT_1[53242] = 32'b00000000000000000000110101110111;
assign LUT_1[53243] = 32'b11111111111111111010000111110011;
assign LUT_1[53244] = 32'b00000000000000001101000000111101;
assign LUT_1[53245] = 32'b00000000000000000110010010111001;
assign LUT_1[53246] = 32'b00000000000000001000101111001110;
assign LUT_1[53247] = 32'b00000000000000000010000001001010;
assign LUT_1[53248] = 32'b11111111111111111110111111010111;
assign LUT_1[53249] = 32'b11111111111111111000010001010011;
assign LUT_1[53250] = 32'b11111111111111111010101101101000;
assign LUT_1[53251] = 32'b11111111111111110011111111100100;
assign LUT_1[53252] = 32'b00000000000000000110111000101110;
assign LUT_1[53253] = 32'b00000000000000000000001010101010;
assign LUT_1[53254] = 32'b00000000000000000010100110111111;
assign LUT_1[53255] = 32'b11111111111111111011111000111011;
assign LUT_1[53256] = 32'b11111111111111111110001101001100;
assign LUT_1[53257] = 32'b11111111111111110111011111001000;
assign LUT_1[53258] = 32'b11111111111111111001111011011101;
assign LUT_1[53259] = 32'b11111111111111110011001101011001;
assign LUT_1[53260] = 32'b00000000000000000110000110100011;
assign LUT_1[53261] = 32'b11111111111111111111011000011111;
assign LUT_1[53262] = 32'b00000000000000000001110100110100;
assign LUT_1[53263] = 32'b11111111111111111011000110110000;
assign LUT_1[53264] = 32'b00000000000000000000111010111001;
assign LUT_1[53265] = 32'b11111111111111111010001100110101;
assign LUT_1[53266] = 32'b11111111111111111100101001001010;
assign LUT_1[53267] = 32'b11111111111111110101111011000110;
assign LUT_1[53268] = 32'b00000000000000001000110100010000;
assign LUT_1[53269] = 32'b00000000000000000010000110001100;
assign LUT_1[53270] = 32'b00000000000000000100100010100001;
assign LUT_1[53271] = 32'b11111111111111111101110100011101;
assign LUT_1[53272] = 32'b00000000000000000000001000101110;
assign LUT_1[53273] = 32'b11111111111111111001011010101010;
assign LUT_1[53274] = 32'b11111111111111111011110110111111;
assign LUT_1[53275] = 32'b11111111111111110101001000111011;
assign LUT_1[53276] = 32'b00000000000000001000000010000101;
assign LUT_1[53277] = 32'b00000000000000000001010100000001;
assign LUT_1[53278] = 32'b00000000000000000011110000010110;
assign LUT_1[53279] = 32'b11111111111111111101000010010010;
assign LUT_1[53280] = 32'b11111111111111111111111010010110;
assign LUT_1[53281] = 32'b11111111111111111001001100010010;
assign LUT_1[53282] = 32'b11111111111111111011101000100111;
assign LUT_1[53283] = 32'b11111111111111110100111010100011;
assign LUT_1[53284] = 32'b00000000000000000111110011101101;
assign LUT_1[53285] = 32'b00000000000000000001000101101001;
assign LUT_1[53286] = 32'b00000000000000000011100001111110;
assign LUT_1[53287] = 32'b11111111111111111100110011111010;
assign LUT_1[53288] = 32'b11111111111111111111001000001011;
assign LUT_1[53289] = 32'b11111111111111111000011010000111;
assign LUT_1[53290] = 32'b11111111111111111010110110011100;
assign LUT_1[53291] = 32'b11111111111111110100001000011000;
assign LUT_1[53292] = 32'b00000000000000000111000001100010;
assign LUT_1[53293] = 32'b00000000000000000000010011011110;
assign LUT_1[53294] = 32'b00000000000000000010101111110011;
assign LUT_1[53295] = 32'b11111111111111111100000001101111;
assign LUT_1[53296] = 32'b00000000000000000001110101111000;
assign LUT_1[53297] = 32'b11111111111111111011000111110100;
assign LUT_1[53298] = 32'b11111111111111111101100100001001;
assign LUT_1[53299] = 32'b11111111111111110110110110000101;
assign LUT_1[53300] = 32'b00000000000000001001101111001111;
assign LUT_1[53301] = 32'b00000000000000000011000001001011;
assign LUT_1[53302] = 32'b00000000000000000101011101100000;
assign LUT_1[53303] = 32'b11111111111111111110101111011100;
assign LUT_1[53304] = 32'b00000000000000000001000011101101;
assign LUT_1[53305] = 32'b11111111111111111010010101101001;
assign LUT_1[53306] = 32'b11111111111111111100110001111110;
assign LUT_1[53307] = 32'b11111111111111110110000011111010;
assign LUT_1[53308] = 32'b00000000000000001000111101000100;
assign LUT_1[53309] = 32'b00000000000000000010001111000000;
assign LUT_1[53310] = 32'b00000000000000000100101011010101;
assign LUT_1[53311] = 32'b11111111111111111101111101010001;
assign LUT_1[53312] = 32'b00000000000000000000111100111111;
assign LUT_1[53313] = 32'b11111111111111111010001110111011;
assign LUT_1[53314] = 32'b11111111111111111100101011010000;
assign LUT_1[53315] = 32'b11111111111111110101111101001100;
assign LUT_1[53316] = 32'b00000000000000001000110110010110;
assign LUT_1[53317] = 32'b00000000000000000010001000010010;
assign LUT_1[53318] = 32'b00000000000000000100100100100111;
assign LUT_1[53319] = 32'b11111111111111111101110110100011;
assign LUT_1[53320] = 32'b00000000000000000000001010110100;
assign LUT_1[53321] = 32'b11111111111111111001011100110000;
assign LUT_1[53322] = 32'b11111111111111111011111001000101;
assign LUT_1[53323] = 32'b11111111111111110101001011000001;
assign LUT_1[53324] = 32'b00000000000000001000000100001011;
assign LUT_1[53325] = 32'b00000000000000000001010110000111;
assign LUT_1[53326] = 32'b00000000000000000011110010011100;
assign LUT_1[53327] = 32'b11111111111111111101000100011000;
assign LUT_1[53328] = 32'b00000000000000000010111000100001;
assign LUT_1[53329] = 32'b11111111111111111100001010011101;
assign LUT_1[53330] = 32'b11111111111111111110100110110010;
assign LUT_1[53331] = 32'b11111111111111110111111000101110;
assign LUT_1[53332] = 32'b00000000000000001010110001111000;
assign LUT_1[53333] = 32'b00000000000000000100000011110100;
assign LUT_1[53334] = 32'b00000000000000000110100000001001;
assign LUT_1[53335] = 32'b11111111111111111111110010000101;
assign LUT_1[53336] = 32'b00000000000000000010000110010110;
assign LUT_1[53337] = 32'b11111111111111111011011000010010;
assign LUT_1[53338] = 32'b11111111111111111101110100100111;
assign LUT_1[53339] = 32'b11111111111111110111000110100011;
assign LUT_1[53340] = 32'b00000000000000001001111111101101;
assign LUT_1[53341] = 32'b00000000000000000011010001101001;
assign LUT_1[53342] = 32'b00000000000000000101101101111110;
assign LUT_1[53343] = 32'b11111111111111111110111111111010;
assign LUT_1[53344] = 32'b00000000000000000001110111111110;
assign LUT_1[53345] = 32'b11111111111111111011001001111010;
assign LUT_1[53346] = 32'b11111111111111111101100110001111;
assign LUT_1[53347] = 32'b11111111111111110110111000001011;
assign LUT_1[53348] = 32'b00000000000000001001110001010101;
assign LUT_1[53349] = 32'b00000000000000000011000011010001;
assign LUT_1[53350] = 32'b00000000000000000101011111100110;
assign LUT_1[53351] = 32'b11111111111111111110110001100010;
assign LUT_1[53352] = 32'b00000000000000000001000101110011;
assign LUT_1[53353] = 32'b11111111111111111010010111101111;
assign LUT_1[53354] = 32'b11111111111111111100110100000100;
assign LUT_1[53355] = 32'b11111111111111110110000110000000;
assign LUT_1[53356] = 32'b00000000000000001000111111001010;
assign LUT_1[53357] = 32'b00000000000000000010010001000110;
assign LUT_1[53358] = 32'b00000000000000000100101101011011;
assign LUT_1[53359] = 32'b11111111111111111101111111010111;
assign LUT_1[53360] = 32'b00000000000000000011110011100000;
assign LUT_1[53361] = 32'b11111111111111111101000101011100;
assign LUT_1[53362] = 32'b11111111111111111111100001110001;
assign LUT_1[53363] = 32'b11111111111111111000110011101101;
assign LUT_1[53364] = 32'b00000000000000001011101100110111;
assign LUT_1[53365] = 32'b00000000000000000100111110110011;
assign LUT_1[53366] = 32'b00000000000000000111011011001000;
assign LUT_1[53367] = 32'b00000000000000000000101101000100;
assign LUT_1[53368] = 32'b00000000000000000011000001010101;
assign LUT_1[53369] = 32'b11111111111111111100010011010001;
assign LUT_1[53370] = 32'b11111111111111111110101111100110;
assign LUT_1[53371] = 32'b11111111111111111000000001100010;
assign LUT_1[53372] = 32'b00000000000000001010111010101100;
assign LUT_1[53373] = 32'b00000000000000000100001100101000;
assign LUT_1[53374] = 32'b00000000000000000110101000111101;
assign LUT_1[53375] = 32'b11111111111111111111111010111001;
assign LUT_1[53376] = 32'b00000000000000000001111111011010;
assign LUT_1[53377] = 32'b11111111111111111011010001010110;
assign LUT_1[53378] = 32'b11111111111111111101101101101011;
assign LUT_1[53379] = 32'b11111111111111110110111111100111;
assign LUT_1[53380] = 32'b00000000000000001001111000110001;
assign LUT_1[53381] = 32'b00000000000000000011001010101101;
assign LUT_1[53382] = 32'b00000000000000000101100111000010;
assign LUT_1[53383] = 32'b11111111111111111110111000111110;
assign LUT_1[53384] = 32'b00000000000000000001001101001111;
assign LUT_1[53385] = 32'b11111111111111111010011111001011;
assign LUT_1[53386] = 32'b11111111111111111100111011100000;
assign LUT_1[53387] = 32'b11111111111111110110001101011100;
assign LUT_1[53388] = 32'b00000000000000001001000110100110;
assign LUT_1[53389] = 32'b00000000000000000010011000100010;
assign LUT_1[53390] = 32'b00000000000000000100110100110111;
assign LUT_1[53391] = 32'b11111111111111111110000110110011;
assign LUT_1[53392] = 32'b00000000000000000011111010111100;
assign LUT_1[53393] = 32'b11111111111111111101001100111000;
assign LUT_1[53394] = 32'b11111111111111111111101001001101;
assign LUT_1[53395] = 32'b11111111111111111000111011001001;
assign LUT_1[53396] = 32'b00000000000000001011110100010011;
assign LUT_1[53397] = 32'b00000000000000000101000110001111;
assign LUT_1[53398] = 32'b00000000000000000111100010100100;
assign LUT_1[53399] = 32'b00000000000000000000110100100000;
assign LUT_1[53400] = 32'b00000000000000000011001000110001;
assign LUT_1[53401] = 32'b11111111111111111100011010101101;
assign LUT_1[53402] = 32'b11111111111111111110110111000010;
assign LUT_1[53403] = 32'b11111111111111111000001000111110;
assign LUT_1[53404] = 32'b00000000000000001011000010001000;
assign LUT_1[53405] = 32'b00000000000000000100010100000100;
assign LUT_1[53406] = 32'b00000000000000000110110000011001;
assign LUT_1[53407] = 32'b00000000000000000000000010010101;
assign LUT_1[53408] = 32'b00000000000000000010111010011001;
assign LUT_1[53409] = 32'b11111111111111111100001100010101;
assign LUT_1[53410] = 32'b11111111111111111110101000101010;
assign LUT_1[53411] = 32'b11111111111111110111111010100110;
assign LUT_1[53412] = 32'b00000000000000001010110011110000;
assign LUT_1[53413] = 32'b00000000000000000100000101101100;
assign LUT_1[53414] = 32'b00000000000000000110100010000001;
assign LUT_1[53415] = 32'b11111111111111111111110011111101;
assign LUT_1[53416] = 32'b00000000000000000010001000001110;
assign LUT_1[53417] = 32'b11111111111111111011011010001010;
assign LUT_1[53418] = 32'b11111111111111111101110110011111;
assign LUT_1[53419] = 32'b11111111111111110111001000011011;
assign LUT_1[53420] = 32'b00000000000000001010000001100101;
assign LUT_1[53421] = 32'b00000000000000000011010011100001;
assign LUT_1[53422] = 32'b00000000000000000101101111110110;
assign LUT_1[53423] = 32'b11111111111111111111000001110010;
assign LUT_1[53424] = 32'b00000000000000000100110101111011;
assign LUT_1[53425] = 32'b11111111111111111110000111110111;
assign LUT_1[53426] = 32'b00000000000000000000100100001100;
assign LUT_1[53427] = 32'b11111111111111111001110110001000;
assign LUT_1[53428] = 32'b00000000000000001100101111010010;
assign LUT_1[53429] = 32'b00000000000000000110000001001110;
assign LUT_1[53430] = 32'b00000000000000001000011101100011;
assign LUT_1[53431] = 32'b00000000000000000001101111011111;
assign LUT_1[53432] = 32'b00000000000000000100000011110000;
assign LUT_1[53433] = 32'b11111111111111111101010101101100;
assign LUT_1[53434] = 32'b11111111111111111111110010000001;
assign LUT_1[53435] = 32'b11111111111111111001000011111101;
assign LUT_1[53436] = 32'b00000000000000001011111101000111;
assign LUT_1[53437] = 32'b00000000000000000101001111000011;
assign LUT_1[53438] = 32'b00000000000000000111101011011000;
assign LUT_1[53439] = 32'b00000000000000000000111101010100;
assign LUT_1[53440] = 32'b00000000000000000011111101000010;
assign LUT_1[53441] = 32'b11111111111111111101001110111110;
assign LUT_1[53442] = 32'b11111111111111111111101011010011;
assign LUT_1[53443] = 32'b11111111111111111000111101001111;
assign LUT_1[53444] = 32'b00000000000000001011110110011001;
assign LUT_1[53445] = 32'b00000000000000000101001000010101;
assign LUT_1[53446] = 32'b00000000000000000111100100101010;
assign LUT_1[53447] = 32'b00000000000000000000110110100110;
assign LUT_1[53448] = 32'b00000000000000000011001010110111;
assign LUT_1[53449] = 32'b11111111111111111100011100110011;
assign LUT_1[53450] = 32'b11111111111111111110111001001000;
assign LUT_1[53451] = 32'b11111111111111111000001011000100;
assign LUT_1[53452] = 32'b00000000000000001011000100001110;
assign LUT_1[53453] = 32'b00000000000000000100010110001010;
assign LUT_1[53454] = 32'b00000000000000000110110010011111;
assign LUT_1[53455] = 32'b00000000000000000000000100011011;
assign LUT_1[53456] = 32'b00000000000000000101111000100100;
assign LUT_1[53457] = 32'b11111111111111111111001010100000;
assign LUT_1[53458] = 32'b00000000000000000001100110110101;
assign LUT_1[53459] = 32'b11111111111111111010111000110001;
assign LUT_1[53460] = 32'b00000000000000001101110001111011;
assign LUT_1[53461] = 32'b00000000000000000111000011110111;
assign LUT_1[53462] = 32'b00000000000000001001100000001100;
assign LUT_1[53463] = 32'b00000000000000000010110010001000;
assign LUT_1[53464] = 32'b00000000000000000101000110011001;
assign LUT_1[53465] = 32'b11111111111111111110011000010101;
assign LUT_1[53466] = 32'b00000000000000000000110100101010;
assign LUT_1[53467] = 32'b11111111111111111010000110100110;
assign LUT_1[53468] = 32'b00000000000000001100111111110000;
assign LUT_1[53469] = 32'b00000000000000000110010001101100;
assign LUT_1[53470] = 32'b00000000000000001000101110000001;
assign LUT_1[53471] = 32'b00000000000000000001111111111101;
assign LUT_1[53472] = 32'b00000000000000000100111000000001;
assign LUT_1[53473] = 32'b11111111111111111110001001111101;
assign LUT_1[53474] = 32'b00000000000000000000100110010010;
assign LUT_1[53475] = 32'b11111111111111111001111000001110;
assign LUT_1[53476] = 32'b00000000000000001100110001011000;
assign LUT_1[53477] = 32'b00000000000000000110000011010100;
assign LUT_1[53478] = 32'b00000000000000001000011111101001;
assign LUT_1[53479] = 32'b00000000000000000001110001100101;
assign LUT_1[53480] = 32'b00000000000000000100000101110110;
assign LUT_1[53481] = 32'b11111111111111111101010111110010;
assign LUT_1[53482] = 32'b11111111111111111111110100000111;
assign LUT_1[53483] = 32'b11111111111111111001000110000011;
assign LUT_1[53484] = 32'b00000000000000001011111111001101;
assign LUT_1[53485] = 32'b00000000000000000101010001001001;
assign LUT_1[53486] = 32'b00000000000000000111101101011110;
assign LUT_1[53487] = 32'b00000000000000000000111111011010;
assign LUT_1[53488] = 32'b00000000000000000110110011100011;
assign LUT_1[53489] = 32'b00000000000000000000000101011111;
assign LUT_1[53490] = 32'b00000000000000000010100001110100;
assign LUT_1[53491] = 32'b11111111111111111011110011110000;
assign LUT_1[53492] = 32'b00000000000000001110101100111010;
assign LUT_1[53493] = 32'b00000000000000000111111110110110;
assign LUT_1[53494] = 32'b00000000000000001010011011001011;
assign LUT_1[53495] = 32'b00000000000000000011101101000111;
assign LUT_1[53496] = 32'b00000000000000000110000001011000;
assign LUT_1[53497] = 32'b11111111111111111111010011010100;
assign LUT_1[53498] = 32'b00000000000000000001101111101001;
assign LUT_1[53499] = 32'b11111111111111111011000001100101;
assign LUT_1[53500] = 32'b00000000000000001101111010101111;
assign LUT_1[53501] = 32'b00000000000000000111001100101011;
assign LUT_1[53502] = 32'b00000000000000001001101001000000;
assign LUT_1[53503] = 32'b00000000000000000010111010111100;
assign LUT_1[53504] = 32'b11111111111111111100110011100011;
assign LUT_1[53505] = 32'b11111111111111110110000101011111;
assign LUT_1[53506] = 32'b11111111111111111000100001110100;
assign LUT_1[53507] = 32'b11111111111111110001110011110000;
assign LUT_1[53508] = 32'b00000000000000000100101100111010;
assign LUT_1[53509] = 32'b11111111111111111101111110110110;
assign LUT_1[53510] = 32'b00000000000000000000011011001011;
assign LUT_1[53511] = 32'b11111111111111111001101101000111;
assign LUT_1[53512] = 32'b11111111111111111100000001011000;
assign LUT_1[53513] = 32'b11111111111111110101010011010100;
assign LUT_1[53514] = 32'b11111111111111110111101111101001;
assign LUT_1[53515] = 32'b11111111111111110001000001100101;
assign LUT_1[53516] = 32'b00000000000000000011111010101111;
assign LUT_1[53517] = 32'b11111111111111111101001100101011;
assign LUT_1[53518] = 32'b11111111111111111111101001000000;
assign LUT_1[53519] = 32'b11111111111111111000111010111100;
assign LUT_1[53520] = 32'b11111111111111111110101111000101;
assign LUT_1[53521] = 32'b11111111111111111000000001000001;
assign LUT_1[53522] = 32'b11111111111111111010011101010110;
assign LUT_1[53523] = 32'b11111111111111110011101111010010;
assign LUT_1[53524] = 32'b00000000000000000110101000011100;
assign LUT_1[53525] = 32'b11111111111111111111111010011000;
assign LUT_1[53526] = 32'b00000000000000000010010110101101;
assign LUT_1[53527] = 32'b11111111111111111011101000101001;
assign LUT_1[53528] = 32'b11111111111111111101111100111010;
assign LUT_1[53529] = 32'b11111111111111110111001110110110;
assign LUT_1[53530] = 32'b11111111111111111001101011001011;
assign LUT_1[53531] = 32'b11111111111111110010111101000111;
assign LUT_1[53532] = 32'b00000000000000000101110110010001;
assign LUT_1[53533] = 32'b11111111111111111111001000001101;
assign LUT_1[53534] = 32'b00000000000000000001100100100010;
assign LUT_1[53535] = 32'b11111111111111111010110110011110;
assign LUT_1[53536] = 32'b11111111111111111101101110100010;
assign LUT_1[53537] = 32'b11111111111111110111000000011110;
assign LUT_1[53538] = 32'b11111111111111111001011100110011;
assign LUT_1[53539] = 32'b11111111111111110010101110101111;
assign LUT_1[53540] = 32'b00000000000000000101100111111001;
assign LUT_1[53541] = 32'b11111111111111111110111001110101;
assign LUT_1[53542] = 32'b00000000000000000001010110001010;
assign LUT_1[53543] = 32'b11111111111111111010101000000110;
assign LUT_1[53544] = 32'b11111111111111111100111100010111;
assign LUT_1[53545] = 32'b11111111111111110110001110010011;
assign LUT_1[53546] = 32'b11111111111111111000101010101000;
assign LUT_1[53547] = 32'b11111111111111110001111100100100;
assign LUT_1[53548] = 32'b00000000000000000100110101101110;
assign LUT_1[53549] = 32'b11111111111111111110000111101010;
assign LUT_1[53550] = 32'b00000000000000000000100011111111;
assign LUT_1[53551] = 32'b11111111111111111001110101111011;
assign LUT_1[53552] = 32'b11111111111111111111101010000100;
assign LUT_1[53553] = 32'b11111111111111111000111100000000;
assign LUT_1[53554] = 32'b11111111111111111011011000010101;
assign LUT_1[53555] = 32'b11111111111111110100101010010001;
assign LUT_1[53556] = 32'b00000000000000000111100011011011;
assign LUT_1[53557] = 32'b00000000000000000000110101010111;
assign LUT_1[53558] = 32'b00000000000000000011010001101100;
assign LUT_1[53559] = 32'b11111111111111111100100011101000;
assign LUT_1[53560] = 32'b11111111111111111110110111111001;
assign LUT_1[53561] = 32'b11111111111111111000001001110101;
assign LUT_1[53562] = 32'b11111111111111111010100110001010;
assign LUT_1[53563] = 32'b11111111111111110011111000000110;
assign LUT_1[53564] = 32'b00000000000000000110110001010000;
assign LUT_1[53565] = 32'b00000000000000000000000011001100;
assign LUT_1[53566] = 32'b00000000000000000010011111100001;
assign LUT_1[53567] = 32'b11111111111111111011110001011101;
assign LUT_1[53568] = 32'b11111111111111111110110001001011;
assign LUT_1[53569] = 32'b11111111111111111000000011000111;
assign LUT_1[53570] = 32'b11111111111111111010011111011100;
assign LUT_1[53571] = 32'b11111111111111110011110001011000;
assign LUT_1[53572] = 32'b00000000000000000110101010100010;
assign LUT_1[53573] = 32'b11111111111111111111111100011110;
assign LUT_1[53574] = 32'b00000000000000000010011000110011;
assign LUT_1[53575] = 32'b11111111111111111011101010101111;
assign LUT_1[53576] = 32'b11111111111111111101111111000000;
assign LUT_1[53577] = 32'b11111111111111110111010000111100;
assign LUT_1[53578] = 32'b11111111111111111001101101010001;
assign LUT_1[53579] = 32'b11111111111111110010111111001101;
assign LUT_1[53580] = 32'b00000000000000000101111000010111;
assign LUT_1[53581] = 32'b11111111111111111111001010010011;
assign LUT_1[53582] = 32'b00000000000000000001100110101000;
assign LUT_1[53583] = 32'b11111111111111111010111000100100;
assign LUT_1[53584] = 32'b00000000000000000000101100101101;
assign LUT_1[53585] = 32'b11111111111111111001111110101001;
assign LUT_1[53586] = 32'b11111111111111111100011010111110;
assign LUT_1[53587] = 32'b11111111111111110101101100111010;
assign LUT_1[53588] = 32'b00000000000000001000100110000100;
assign LUT_1[53589] = 32'b00000000000000000001111000000000;
assign LUT_1[53590] = 32'b00000000000000000100010100010101;
assign LUT_1[53591] = 32'b11111111111111111101100110010001;
assign LUT_1[53592] = 32'b11111111111111111111111010100010;
assign LUT_1[53593] = 32'b11111111111111111001001100011110;
assign LUT_1[53594] = 32'b11111111111111111011101000110011;
assign LUT_1[53595] = 32'b11111111111111110100111010101111;
assign LUT_1[53596] = 32'b00000000000000000111110011111001;
assign LUT_1[53597] = 32'b00000000000000000001000101110101;
assign LUT_1[53598] = 32'b00000000000000000011100010001010;
assign LUT_1[53599] = 32'b11111111111111111100110100000110;
assign LUT_1[53600] = 32'b11111111111111111111101100001010;
assign LUT_1[53601] = 32'b11111111111111111000111110000110;
assign LUT_1[53602] = 32'b11111111111111111011011010011011;
assign LUT_1[53603] = 32'b11111111111111110100101100010111;
assign LUT_1[53604] = 32'b00000000000000000111100101100001;
assign LUT_1[53605] = 32'b00000000000000000000110111011101;
assign LUT_1[53606] = 32'b00000000000000000011010011110010;
assign LUT_1[53607] = 32'b11111111111111111100100101101110;
assign LUT_1[53608] = 32'b11111111111111111110111001111111;
assign LUT_1[53609] = 32'b11111111111111111000001011111011;
assign LUT_1[53610] = 32'b11111111111111111010101000010000;
assign LUT_1[53611] = 32'b11111111111111110011111010001100;
assign LUT_1[53612] = 32'b00000000000000000110110011010110;
assign LUT_1[53613] = 32'b00000000000000000000000101010010;
assign LUT_1[53614] = 32'b00000000000000000010100001100111;
assign LUT_1[53615] = 32'b11111111111111111011110011100011;
assign LUT_1[53616] = 32'b00000000000000000001100111101100;
assign LUT_1[53617] = 32'b11111111111111111010111001101000;
assign LUT_1[53618] = 32'b11111111111111111101010101111101;
assign LUT_1[53619] = 32'b11111111111111110110100111111001;
assign LUT_1[53620] = 32'b00000000000000001001100001000011;
assign LUT_1[53621] = 32'b00000000000000000010110010111111;
assign LUT_1[53622] = 32'b00000000000000000101001111010100;
assign LUT_1[53623] = 32'b11111111111111111110100001010000;
assign LUT_1[53624] = 32'b00000000000000000000110101100001;
assign LUT_1[53625] = 32'b11111111111111111010000111011101;
assign LUT_1[53626] = 32'b11111111111111111100100011110010;
assign LUT_1[53627] = 32'b11111111111111110101110101101110;
assign LUT_1[53628] = 32'b00000000000000001000101110111000;
assign LUT_1[53629] = 32'b00000000000000000010000000110100;
assign LUT_1[53630] = 32'b00000000000000000100011101001001;
assign LUT_1[53631] = 32'b11111111111111111101101111000101;
assign LUT_1[53632] = 32'b11111111111111111111110011100110;
assign LUT_1[53633] = 32'b11111111111111111001000101100010;
assign LUT_1[53634] = 32'b11111111111111111011100001110111;
assign LUT_1[53635] = 32'b11111111111111110100110011110011;
assign LUT_1[53636] = 32'b00000000000000000111101100111101;
assign LUT_1[53637] = 32'b00000000000000000000111110111001;
assign LUT_1[53638] = 32'b00000000000000000011011011001110;
assign LUT_1[53639] = 32'b11111111111111111100101101001010;
assign LUT_1[53640] = 32'b11111111111111111111000001011011;
assign LUT_1[53641] = 32'b11111111111111111000010011010111;
assign LUT_1[53642] = 32'b11111111111111111010101111101100;
assign LUT_1[53643] = 32'b11111111111111110100000001101000;
assign LUT_1[53644] = 32'b00000000000000000110111010110010;
assign LUT_1[53645] = 32'b00000000000000000000001100101110;
assign LUT_1[53646] = 32'b00000000000000000010101001000011;
assign LUT_1[53647] = 32'b11111111111111111011111010111111;
assign LUT_1[53648] = 32'b00000000000000000001101111001000;
assign LUT_1[53649] = 32'b11111111111111111011000001000100;
assign LUT_1[53650] = 32'b11111111111111111101011101011001;
assign LUT_1[53651] = 32'b11111111111111110110101111010101;
assign LUT_1[53652] = 32'b00000000000000001001101000011111;
assign LUT_1[53653] = 32'b00000000000000000010111010011011;
assign LUT_1[53654] = 32'b00000000000000000101010110110000;
assign LUT_1[53655] = 32'b11111111111111111110101000101100;
assign LUT_1[53656] = 32'b00000000000000000000111100111101;
assign LUT_1[53657] = 32'b11111111111111111010001110111001;
assign LUT_1[53658] = 32'b11111111111111111100101011001110;
assign LUT_1[53659] = 32'b11111111111111110101111101001010;
assign LUT_1[53660] = 32'b00000000000000001000110110010100;
assign LUT_1[53661] = 32'b00000000000000000010001000010000;
assign LUT_1[53662] = 32'b00000000000000000100100100100101;
assign LUT_1[53663] = 32'b11111111111111111101110110100001;
assign LUT_1[53664] = 32'b00000000000000000000101110100101;
assign LUT_1[53665] = 32'b11111111111111111010000000100001;
assign LUT_1[53666] = 32'b11111111111111111100011100110110;
assign LUT_1[53667] = 32'b11111111111111110101101110110010;
assign LUT_1[53668] = 32'b00000000000000001000100111111100;
assign LUT_1[53669] = 32'b00000000000000000001111001111000;
assign LUT_1[53670] = 32'b00000000000000000100010110001101;
assign LUT_1[53671] = 32'b11111111111111111101101000001001;
assign LUT_1[53672] = 32'b11111111111111111111111100011010;
assign LUT_1[53673] = 32'b11111111111111111001001110010110;
assign LUT_1[53674] = 32'b11111111111111111011101010101011;
assign LUT_1[53675] = 32'b11111111111111110100111100100111;
assign LUT_1[53676] = 32'b00000000000000000111110101110001;
assign LUT_1[53677] = 32'b00000000000000000001000111101101;
assign LUT_1[53678] = 32'b00000000000000000011100100000010;
assign LUT_1[53679] = 32'b11111111111111111100110101111110;
assign LUT_1[53680] = 32'b00000000000000000010101010000111;
assign LUT_1[53681] = 32'b11111111111111111011111100000011;
assign LUT_1[53682] = 32'b11111111111111111110011000011000;
assign LUT_1[53683] = 32'b11111111111111110111101010010100;
assign LUT_1[53684] = 32'b00000000000000001010100011011110;
assign LUT_1[53685] = 32'b00000000000000000011110101011010;
assign LUT_1[53686] = 32'b00000000000000000110010001101111;
assign LUT_1[53687] = 32'b11111111111111111111100011101011;
assign LUT_1[53688] = 32'b00000000000000000001110111111100;
assign LUT_1[53689] = 32'b11111111111111111011001001111000;
assign LUT_1[53690] = 32'b11111111111111111101100110001101;
assign LUT_1[53691] = 32'b11111111111111110110111000001001;
assign LUT_1[53692] = 32'b00000000000000001001110001010011;
assign LUT_1[53693] = 32'b00000000000000000011000011001111;
assign LUT_1[53694] = 32'b00000000000000000101011111100100;
assign LUT_1[53695] = 32'b11111111111111111110110001100000;
assign LUT_1[53696] = 32'b00000000000000000001110001001110;
assign LUT_1[53697] = 32'b11111111111111111011000011001010;
assign LUT_1[53698] = 32'b11111111111111111101011111011111;
assign LUT_1[53699] = 32'b11111111111111110110110001011011;
assign LUT_1[53700] = 32'b00000000000000001001101010100101;
assign LUT_1[53701] = 32'b00000000000000000010111100100001;
assign LUT_1[53702] = 32'b00000000000000000101011000110110;
assign LUT_1[53703] = 32'b11111111111111111110101010110010;
assign LUT_1[53704] = 32'b00000000000000000000111111000011;
assign LUT_1[53705] = 32'b11111111111111111010010000111111;
assign LUT_1[53706] = 32'b11111111111111111100101101010100;
assign LUT_1[53707] = 32'b11111111111111110101111111010000;
assign LUT_1[53708] = 32'b00000000000000001000111000011010;
assign LUT_1[53709] = 32'b00000000000000000010001010010110;
assign LUT_1[53710] = 32'b00000000000000000100100110101011;
assign LUT_1[53711] = 32'b11111111111111111101111000100111;
assign LUT_1[53712] = 32'b00000000000000000011101100110000;
assign LUT_1[53713] = 32'b11111111111111111100111110101100;
assign LUT_1[53714] = 32'b11111111111111111111011011000001;
assign LUT_1[53715] = 32'b11111111111111111000101100111101;
assign LUT_1[53716] = 32'b00000000000000001011100110000111;
assign LUT_1[53717] = 32'b00000000000000000100111000000011;
assign LUT_1[53718] = 32'b00000000000000000111010100011000;
assign LUT_1[53719] = 32'b00000000000000000000100110010100;
assign LUT_1[53720] = 32'b00000000000000000010111010100101;
assign LUT_1[53721] = 32'b11111111111111111100001100100001;
assign LUT_1[53722] = 32'b11111111111111111110101000110110;
assign LUT_1[53723] = 32'b11111111111111110111111010110010;
assign LUT_1[53724] = 32'b00000000000000001010110011111100;
assign LUT_1[53725] = 32'b00000000000000000100000101111000;
assign LUT_1[53726] = 32'b00000000000000000110100010001101;
assign LUT_1[53727] = 32'b11111111111111111111110100001001;
assign LUT_1[53728] = 32'b00000000000000000010101100001101;
assign LUT_1[53729] = 32'b11111111111111111011111110001001;
assign LUT_1[53730] = 32'b11111111111111111110011010011110;
assign LUT_1[53731] = 32'b11111111111111110111101100011010;
assign LUT_1[53732] = 32'b00000000000000001010100101100100;
assign LUT_1[53733] = 32'b00000000000000000011110111100000;
assign LUT_1[53734] = 32'b00000000000000000110010011110101;
assign LUT_1[53735] = 32'b11111111111111111111100101110001;
assign LUT_1[53736] = 32'b00000000000000000001111010000010;
assign LUT_1[53737] = 32'b11111111111111111011001011111110;
assign LUT_1[53738] = 32'b11111111111111111101101000010011;
assign LUT_1[53739] = 32'b11111111111111110110111010001111;
assign LUT_1[53740] = 32'b00000000000000001001110011011001;
assign LUT_1[53741] = 32'b00000000000000000011000101010101;
assign LUT_1[53742] = 32'b00000000000000000101100001101010;
assign LUT_1[53743] = 32'b11111111111111111110110011100110;
assign LUT_1[53744] = 32'b00000000000000000100100111101111;
assign LUT_1[53745] = 32'b11111111111111111101111001101011;
assign LUT_1[53746] = 32'b00000000000000000000010110000000;
assign LUT_1[53747] = 32'b11111111111111111001100111111100;
assign LUT_1[53748] = 32'b00000000000000001100100001000110;
assign LUT_1[53749] = 32'b00000000000000000101110011000010;
assign LUT_1[53750] = 32'b00000000000000001000001111010111;
assign LUT_1[53751] = 32'b00000000000000000001100001010011;
assign LUT_1[53752] = 32'b00000000000000000011110101100100;
assign LUT_1[53753] = 32'b11111111111111111101000111100000;
assign LUT_1[53754] = 32'b11111111111111111111100011110101;
assign LUT_1[53755] = 32'b11111111111111111000110101110001;
assign LUT_1[53756] = 32'b00000000000000001011101110111011;
assign LUT_1[53757] = 32'b00000000000000000101000000110111;
assign LUT_1[53758] = 32'b00000000000000000111011101001100;
assign LUT_1[53759] = 32'b00000000000000000000101111001000;
assign LUT_1[53760] = 32'b11111111111111111000101101110100;
assign LUT_1[53761] = 32'b11111111111111110001111111110000;
assign LUT_1[53762] = 32'b11111111111111110100011100000101;
assign LUT_1[53763] = 32'b11111111111111101101101110000001;
assign LUT_1[53764] = 32'b00000000000000000000100111001011;
assign LUT_1[53765] = 32'b11111111111111111001111001000111;
assign LUT_1[53766] = 32'b11111111111111111100010101011100;
assign LUT_1[53767] = 32'b11111111111111110101100111011000;
assign LUT_1[53768] = 32'b11111111111111110111111011101001;
assign LUT_1[53769] = 32'b11111111111111110001001101100101;
assign LUT_1[53770] = 32'b11111111111111110011101001111010;
assign LUT_1[53771] = 32'b11111111111111101100111011110110;
assign LUT_1[53772] = 32'b11111111111111111111110101000000;
assign LUT_1[53773] = 32'b11111111111111111001000110111100;
assign LUT_1[53774] = 32'b11111111111111111011100011010001;
assign LUT_1[53775] = 32'b11111111111111110100110101001101;
assign LUT_1[53776] = 32'b11111111111111111010101001010110;
assign LUT_1[53777] = 32'b11111111111111110011111011010010;
assign LUT_1[53778] = 32'b11111111111111110110010111100111;
assign LUT_1[53779] = 32'b11111111111111101111101001100011;
assign LUT_1[53780] = 32'b00000000000000000010100010101101;
assign LUT_1[53781] = 32'b11111111111111111011110100101001;
assign LUT_1[53782] = 32'b11111111111111111110010000111110;
assign LUT_1[53783] = 32'b11111111111111110111100010111010;
assign LUT_1[53784] = 32'b11111111111111111001110111001011;
assign LUT_1[53785] = 32'b11111111111111110011001001000111;
assign LUT_1[53786] = 32'b11111111111111110101100101011100;
assign LUT_1[53787] = 32'b11111111111111101110110111011000;
assign LUT_1[53788] = 32'b00000000000000000001110000100010;
assign LUT_1[53789] = 32'b11111111111111111011000010011110;
assign LUT_1[53790] = 32'b11111111111111111101011110110011;
assign LUT_1[53791] = 32'b11111111111111110110110000101111;
assign LUT_1[53792] = 32'b11111111111111111001101000110011;
assign LUT_1[53793] = 32'b11111111111111110010111010101111;
assign LUT_1[53794] = 32'b11111111111111110101010111000100;
assign LUT_1[53795] = 32'b11111111111111101110101001000000;
assign LUT_1[53796] = 32'b00000000000000000001100010001010;
assign LUT_1[53797] = 32'b11111111111111111010110100000110;
assign LUT_1[53798] = 32'b11111111111111111101010000011011;
assign LUT_1[53799] = 32'b11111111111111110110100010010111;
assign LUT_1[53800] = 32'b11111111111111111000110110101000;
assign LUT_1[53801] = 32'b11111111111111110010001000100100;
assign LUT_1[53802] = 32'b11111111111111110100100100111001;
assign LUT_1[53803] = 32'b11111111111111101101110110110101;
assign LUT_1[53804] = 32'b00000000000000000000101111111111;
assign LUT_1[53805] = 32'b11111111111111111010000001111011;
assign LUT_1[53806] = 32'b11111111111111111100011110010000;
assign LUT_1[53807] = 32'b11111111111111110101110000001100;
assign LUT_1[53808] = 32'b11111111111111111011100100010101;
assign LUT_1[53809] = 32'b11111111111111110100110110010001;
assign LUT_1[53810] = 32'b11111111111111110111010010100110;
assign LUT_1[53811] = 32'b11111111111111110000100100100010;
assign LUT_1[53812] = 32'b00000000000000000011011101101100;
assign LUT_1[53813] = 32'b11111111111111111100101111101000;
assign LUT_1[53814] = 32'b11111111111111111111001011111101;
assign LUT_1[53815] = 32'b11111111111111111000011101111001;
assign LUT_1[53816] = 32'b11111111111111111010110010001010;
assign LUT_1[53817] = 32'b11111111111111110100000100000110;
assign LUT_1[53818] = 32'b11111111111111110110100000011011;
assign LUT_1[53819] = 32'b11111111111111101111110010010111;
assign LUT_1[53820] = 32'b00000000000000000010101011100001;
assign LUT_1[53821] = 32'b11111111111111111011111101011101;
assign LUT_1[53822] = 32'b11111111111111111110011001110010;
assign LUT_1[53823] = 32'b11111111111111110111101011101110;
assign LUT_1[53824] = 32'b11111111111111111010101011011100;
assign LUT_1[53825] = 32'b11111111111111110011111101011000;
assign LUT_1[53826] = 32'b11111111111111110110011001101101;
assign LUT_1[53827] = 32'b11111111111111101111101011101001;
assign LUT_1[53828] = 32'b00000000000000000010100100110011;
assign LUT_1[53829] = 32'b11111111111111111011110110101111;
assign LUT_1[53830] = 32'b11111111111111111110010011000100;
assign LUT_1[53831] = 32'b11111111111111110111100101000000;
assign LUT_1[53832] = 32'b11111111111111111001111001010001;
assign LUT_1[53833] = 32'b11111111111111110011001011001101;
assign LUT_1[53834] = 32'b11111111111111110101100111100010;
assign LUT_1[53835] = 32'b11111111111111101110111001011110;
assign LUT_1[53836] = 32'b00000000000000000001110010101000;
assign LUT_1[53837] = 32'b11111111111111111011000100100100;
assign LUT_1[53838] = 32'b11111111111111111101100000111001;
assign LUT_1[53839] = 32'b11111111111111110110110010110101;
assign LUT_1[53840] = 32'b11111111111111111100100110111110;
assign LUT_1[53841] = 32'b11111111111111110101111000111010;
assign LUT_1[53842] = 32'b11111111111111111000010101001111;
assign LUT_1[53843] = 32'b11111111111111110001100111001011;
assign LUT_1[53844] = 32'b00000000000000000100100000010101;
assign LUT_1[53845] = 32'b11111111111111111101110010010001;
assign LUT_1[53846] = 32'b00000000000000000000001110100110;
assign LUT_1[53847] = 32'b11111111111111111001100000100010;
assign LUT_1[53848] = 32'b11111111111111111011110100110011;
assign LUT_1[53849] = 32'b11111111111111110101000110101111;
assign LUT_1[53850] = 32'b11111111111111110111100011000100;
assign LUT_1[53851] = 32'b11111111111111110000110101000000;
assign LUT_1[53852] = 32'b00000000000000000011101110001010;
assign LUT_1[53853] = 32'b11111111111111111101000000000110;
assign LUT_1[53854] = 32'b11111111111111111111011100011011;
assign LUT_1[53855] = 32'b11111111111111111000101110010111;
assign LUT_1[53856] = 32'b11111111111111111011100110011011;
assign LUT_1[53857] = 32'b11111111111111110100111000010111;
assign LUT_1[53858] = 32'b11111111111111110111010100101100;
assign LUT_1[53859] = 32'b11111111111111110000100110101000;
assign LUT_1[53860] = 32'b00000000000000000011011111110010;
assign LUT_1[53861] = 32'b11111111111111111100110001101110;
assign LUT_1[53862] = 32'b11111111111111111111001110000011;
assign LUT_1[53863] = 32'b11111111111111111000011111111111;
assign LUT_1[53864] = 32'b11111111111111111010110100010000;
assign LUT_1[53865] = 32'b11111111111111110100000110001100;
assign LUT_1[53866] = 32'b11111111111111110110100010100001;
assign LUT_1[53867] = 32'b11111111111111101111110100011101;
assign LUT_1[53868] = 32'b00000000000000000010101101100111;
assign LUT_1[53869] = 32'b11111111111111111011111111100011;
assign LUT_1[53870] = 32'b11111111111111111110011011111000;
assign LUT_1[53871] = 32'b11111111111111110111101101110100;
assign LUT_1[53872] = 32'b11111111111111111101100001111101;
assign LUT_1[53873] = 32'b11111111111111110110110011111001;
assign LUT_1[53874] = 32'b11111111111111111001010000001110;
assign LUT_1[53875] = 32'b11111111111111110010100010001010;
assign LUT_1[53876] = 32'b00000000000000000101011011010100;
assign LUT_1[53877] = 32'b11111111111111111110101101010000;
assign LUT_1[53878] = 32'b00000000000000000001001001100101;
assign LUT_1[53879] = 32'b11111111111111111010011011100001;
assign LUT_1[53880] = 32'b11111111111111111100101111110010;
assign LUT_1[53881] = 32'b11111111111111110110000001101110;
assign LUT_1[53882] = 32'b11111111111111111000011110000011;
assign LUT_1[53883] = 32'b11111111111111110001101111111111;
assign LUT_1[53884] = 32'b00000000000000000100101001001001;
assign LUT_1[53885] = 32'b11111111111111111101111011000101;
assign LUT_1[53886] = 32'b00000000000000000000010111011010;
assign LUT_1[53887] = 32'b11111111111111111001101001010110;
assign LUT_1[53888] = 32'b11111111111111111011101101110111;
assign LUT_1[53889] = 32'b11111111111111110100111111110011;
assign LUT_1[53890] = 32'b11111111111111110111011100001000;
assign LUT_1[53891] = 32'b11111111111111110000101110000100;
assign LUT_1[53892] = 32'b00000000000000000011100111001110;
assign LUT_1[53893] = 32'b11111111111111111100111001001010;
assign LUT_1[53894] = 32'b11111111111111111111010101011111;
assign LUT_1[53895] = 32'b11111111111111111000100111011011;
assign LUT_1[53896] = 32'b11111111111111111010111011101100;
assign LUT_1[53897] = 32'b11111111111111110100001101101000;
assign LUT_1[53898] = 32'b11111111111111110110101001111101;
assign LUT_1[53899] = 32'b11111111111111101111111011111001;
assign LUT_1[53900] = 32'b00000000000000000010110101000011;
assign LUT_1[53901] = 32'b11111111111111111100000110111111;
assign LUT_1[53902] = 32'b11111111111111111110100011010100;
assign LUT_1[53903] = 32'b11111111111111110111110101010000;
assign LUT_1[53904] = 32'b11111111111111111101101001011001;
assign LUT_1[53905] = 32'b11111111111111110110111011010101;
assign LUT_1[53906] = 32'b11111111111111111001010111101010;
assign LUT_1[53907] = 32'b11111111111111110010101001100110;
assign LUT_1[53908] = 32'b00000000000000000101100010110000;
assign LUT_1[53909] = 32'b11111111111111111110110100101100;
assign LUT_1[53910] = 32'b00000000000000000001010001000001;
assign LUT_1[53911] = 32'b11111111111111111010100010111101;
assign LUT_1[53912] = 32'b11111111111111111100110111001110;
assign LUT_1[53913] = 32'b11111111111111110110001001001010;
assign LUT_1[53914] = 32'b11111111111111111000100101011111;
assign LUT_1[53915] = 32'b11111111111111110001110111011011;
assign LUT_1[53916] = 32'b00000000000000000100110000100101;
assign LUT_1[53917] = 32'b11111111111111111110000010100001;
assign LUT_1[53918] = 32'b00000000000000000000011110110110;
assign LUT_1[53919] = 32'b11111111111111111001110000110010;
assign LUT_1[53920] = 32'b11111111111111111100101000110110;
assign LUT_1[53921] = 32'b11111111111111110101111010110010;
assign LUT_1[53922] = 32'b11111111111111111000010111000111;
assign LUT_1[53923] = 32'b11111111111111110001101001000011;
assign LUT_1[53924] = 32'b00000000000000000100100010001101;
assign LUT_1[53925] = 32'b11111111111111111101110100001001;
assign LUT_1[53926] = 32'b00000000000000000000010000011110;
assign LUT_1[53927] = 32'b11111111111111111001100010011010;
assign LUT_1[53928] = 32'b11111111111111111011110110101011;
assign LUT_1[53929] = 32'b11111111111111110101001000100111;
assign LUT_1[53930] = 32'b11111111111111110111100100111100;
assign LUT_1[53931] = 32'b11111111111111110000110110111000;
assign LUT_1[53932] = 32'b00000000000000000011110000000010;
assign LUT_1[53933] = 32'b11111111111111111101000001111110;
assign LUT_1[53934] = 32'b11111111111111111111011110010011;
assign LUT_1[53935] = 32'b11111111111111111000110000001111;
assign LUT_1[53936] = 32'b11111111111111111110100100011000;
assign LUT_1[53937] = 32'b11111111111111110111110110010100;
assign LUT_1[53938] = 32'b11111111111111111010010010101001;
assign LUT_1[53939] = 32'b11111111111111110011100100100101;
assign LUT_1[53940] = 32'b00000000000000000110011101101111;
assign LUT_1[53941] = 32'b11111111111111111111101111101011;
assign LUT_1[53942] = 32'b00000000000000000010001100000000;
assign LUT_1[53943] = 32'b11111111111111111011011101111100;
assign LUT_1[53944] = 32'b11111111111111111101110010001101;
assign LUT_1[53945] = 32'b11111111111111110111000100001001;
assign LUT_1[53946] = 32'b11111111111111111001100000011110;
assign LUT_1[53947] = 32'b11111111111111110010110010011010;
assign LUT_1[53948] = 32'b00000000000000000101101011100100;
assign LUT_1[53949] = 32'b11111111111111111110111101100000;
assign LUT_1[53950] = 32'b00000000000000000001011001110101;
assign LUT_1[53951] = 32'b11111111111111111010101011110001;
assign LUT_1[53952] = 32'b11111111111111111101101011011111;
assign LUT_1[53953] = 32'b11111111111111110110111101011011;
assign LUT_1[53954] = 32'b11111111111111111001011001110000;
assign LUT_1[53955] = 32'b11111111111111110010101011101100;
assign LUT_1[53956] = 32'b00000000000000000101100100110110;
assign LUT_1[53957] = 32'b11111111111111111110110110110010;
assign LUT_1[53958] = 32'b00000000000000000001010011000111;
assign LUT_1[53959] = 32'b11111111111111111010100101000011;
assign LUT_1[53960] = 32'b11111111111111111100111001010100;
assign LUT_1[53961] = 32'b11111111111111110110001011010000;
assign LUT_1[53962] = 32'b11111111111111111000100111100101;
assign LUT_1[53963] = 32'b11111111111111110001111001100001;
assign LUT_1[53964] = 32'b00000000000000000100110010101011;
assign LUT_1[53965] = 32'b11111111111111111110000100100111;
assign LUT_1[53966] = 32'b00000000000000000000100000111100;
assign LUT_1[53967] = 32'b11111111111111111001110010111000;
assign LUT_1[53968] = 32'b11111111111111111111100111000001;
assign LUT_1[53969] = 32'b11111111111111111000111000111101;
assign LUT_1[53970] = 32'b11111111111111111011010101010010;
assign LUT_1[53971] = 32'b11111111111111110100100111001110;
assign LUT_1[53972] = 32'b00000000000000000111100000011000;
assign LUT_1[53973] = 32'b00000000000000000000110010010100;
assign LUT_1[53974] = 32'b00000000000000000011001110101001;
assign LUT_1[53975] = 32'b11111111111111111100100000100101;
assign LUT_1[53976] = 32'b11111111111111111110110100110110;
assign LUT_1[53977] = 32'b11111111111111111000000110110010;
assign LUT_1[53978] = 32'b11111111111111111010100011000111;
assign LUT_1[53979] = 32'b11111111111111110011110101000011;
assign LUT_1[53980] = 32'b00000000000000000110101110001101;
assign LUT_1[53981] = 32'b00000000000000000000000000001001;
assign LUT_1[53982] = 32'b00000000000000000010011100011110;
assign LUT_1[53983] = 32'b11111111111111111011101110011010;
assign LUT_1[53984] = 32'b11111111111111111110100110011110;
assign LUT_1[53985] = 32'b11111111111111110111111000011010;
assign LUT_1[53986] = 32'b11111111111111111010010100101111;
assign LUT_1[53987] = 32'b11111111111111110011100110101011;
assign LUT_1[53988] = 32'b00000000000000000110011111110101;
assign LUT_1[53989] = 32'b11111111111111111111110001110001;
assign LUT_1[53990] = 32'b00000000000000000010001110000110;
assign LUT_1[53991] = 32'b11111111111111111011100000000010;
assign LUT_1[53992] = 32'b11111111111111111101110100010011;
assign LUT_1[53993] = 32'b11111111111111110111000110001111;
assign LUT_1[53994] = 32'b11111111111111111001100010100100;
assign LUT_1[53995] = 32'b11111111111111110010110100100000;
assign LUT_1[53996] = 32'b00000000000000000101101101101010;
assign LUT_1[53997] = 32'b11111111111111111110111111100110;
assign LUT_1[53998] = 32'b00000000000000000001011011111011;
assign LUT_1[53999] = 32'b11111111111111111010101101110111;
assign LUT_1[54000] = 32'b00000000000000000000100010000000;
assign LUT_1[54001] = 32'b11111111111111111001110011111100;
assign LUT_1[54002] = 32'b11111111111111111100010000010001;
assign LUT_1[54003] = 32'b11111111111111110101100010001101;
assign LUT_1[54004] = 32'b00000000000000001000011011010111;
assign LUT_1[54005] = 32'b00000000000000000001101101010011;
assign LUT_1[54006] = 32'b00000000000000000100001001101000;
assign LUT_1[54007] = 32'b11111111111111111101011011100100;
assign LUT_1[54008] = 32'b11111111111111111111101111110101;
assign LUT_1[54009] = 32'b11111111111111111001000001110001;
assign LUT_1[54010] = 32'b11111111111111111011011110000110;
assign LUT_1[54011] = 32'b11111111111111110100110000000010;
assign LUT_1[54012] = 32'b00000000000000000111101001001100;
assign LUT_1[54013] = 32'b00000000000000000000111011001000;
assign LUT_1[54014] = 32'b00000000000000000011010111011101;
assign LUT_1[54015] = 32'b11111111111111111100101001011001;
assign LUT_1[54016] = 32'b11111111111111110110100010000000;
assign LUT_1[54017] = 32'b11111111111111101111110011111100;
assign LUT_1[54018] = 32'b11111111111111110010010000010001;
assign LUT_1[54019] = 32'b11111111111111101011100010001101;
assign LUT_1[54020] = 32'b11111111111111111110011011010111;
assign LUT_1[54021] = 32'b11111111111111110111101101010011;
assign LUT_1[54022] = 32'b11111111111111111010001001101000;
assign LUT_1[54023] = 32'b11111111111111110011011011100100;
assign LUT_1[54024] = 32'b11111111111111110101101111110101;
assign LUT_1[54025] = 32'b11111111111111101111000001110001;
assign LUT_1[54026] = 32'b11111111111111110001011110000110;
assign LUT_1[54027] = 32'b11111111111111101010110000000010;
assign LUT_1[54028] = 32'b11111111111111111101101001001100;
assign LUT_1[54029] = 32'b11111111111111110110111011001000;
assign LUT_1[54030] = 32'b11111111111111111001010111011101;
assign LUT_1[54031] = 32'b11111111111111110010101001011001;
assign LUT_1[54032] = 32'b11111111111111111000011101100010;
assign LUT_1[54033] = 32'b11111111111111110001101111011110;
assign LUT_1[54034] = 32'b11111111111111110100001011110011;
assign LUT_1[54035] = 32'b11111111111111101101011101101111;
assign LUT_1[54036] = 32'b00000000000000000000010110111001;
assign LUT_1[54037] = 32'b11111111111111111001101000110101;
assign LUT_1[54038] = 32'b11111111111111111100000101001010;
assign LUT_1[54039] = 32'b11111111111111110101010111000110;
assign LUT_1[54040] = 32'b11111111111111110111101011010111;
assign LUT_1[54041] = 32'b11111111111111110000111101010011;
assign LUT_1[54042] = 32'b11111111111111110011011001101000;
assign LUT_1[54043] = 32'b11111111111111101100101011100100;
assign LUT_1[54044] = 32'b11111111111111111111100100101110;
assign LUT_1[54045] = 32'b11111111111111111000110110101010;
assign LUT_1[54046] = 32'b11111111111111111011010010111111;
assign LUT_1[54047] = 32'b11111111111111110100100100111011;
assign LUT_1[54048] = 32'b11111111111111110111011100111111;
assign LUT_1[54049] = 32'b11111111111111110000101110111011;
assign LUT_1[54050] = 32'b11111111111111110011001011010000;
assign LUT_1[54051] = 32'b11111111111111101100011101001100;
assign LUT_1[54052] = 32'b11111111111111111111010110010110;
assign LUT_1[54053] = 32'b11111111111111111000101000010010;
assign LUT_1[54054] = 32'b11111111111111111011000100100111;
assign LUT_1[54055] = 32'b11111111111111110100010110100011;
assign LUT_1[54056] = 32'b11111111111111110110101010110100;
assign LUT_1[54057] = 32'b11111111111111101111111100110000;
assign LUT_1[54058] = 32'b11111111111111110010011001000101;
assign LUT_1[54059] = 32'b11111111111111101011101011000001;
assign LUT_1[54060] = 32'b11111111111111111110100100001011;
assign LUT_1[54061] = 32'b11111111111111110111110110000111;
assign LUT_1[54062] = 32'b11111111111111111010010010011100;
assign LUT_1[54063] = 32'b11111111111111110011100100011000;
assign LUT_1[54064] = 32'b11111111111111111001011000100001;
assign LUT_1[54065] = 32'b11111111111111110010101010011101;
assign LUT_1[54066] = 32'b11111111111111110101000110110010;
assign LUT_1[54067] = 32'b11111111111111101110011000101110;
assign LUT_1[54068] = 32'b00000000000000000001010001111000;
assign LUT_1[54069] = 32'b11111111111111111010100011110100;
assign LUT_1[54070] = 32'b11111111111111111101000000001001;
assign LUT_1[54071] = 32'b11111111111111110110010010000101;
assign LUT_1[54072] = 32'b11111111111111111000100110010110;
assign LUT_1[54073] = 32'b11111111111111110001111000010010;
assign LUT_1[54074] = 32'b11111111111111110100010100100111;
assign LUT_1[54075] = 32'b11111111111111101101100110100011;
assign LUT_1[54076] = 32'b00000000000000000000011111101101;
assign LUT_1[54077] = 32'b11111111111111111001110001101001;
assign LUT_1[54078] = 32'b11111111111111111100001101111110;
assign LUT_1[54079] = 32'b11111111111111110101011111111010;
assign LUT_1[54080] = 32'b11111111111111111000011111101000;
assign LUT_1[54081] = 32'b11111111111111110001110001100100;
assign LUT_1[54082] = 32'b11111111111111110100001101111001;
assign LUT_1[54083] = 32'b11111111111111101101011111110101;
assign LUT_1[54084] = 32'b00000000000000000000011000111111;
assign LUT_1[54085] = 32'b11111111111111111001101010111011;
assign LUT_1[54086] = 32'b11111111111111111100000111010000;
assign LUT_1[54087] = 32'b11111111111111110101011001001100;
assign LUT_1[54088] = 32'b11111111111111110111101101011101;
assign LUT_1[54089] = 32'b11111111111111110000111111011001;
assign LUT_1[54090] = 32'b11111111111111110011011011101110;
assign LUT_1[54091] = 32'b11111111111111101100101101101010;
assign LUT_1[54092] = 32'b11111111111111111111100110110100;
assign LUT_1[54093] = 32'b11111111111111111000111000110000;
assign LUT_1[54094] = 32'b11111111111111111011010101000101;
assign LUT_1[54095] = 32'b11111111111111110100100111000001;
assign LUT_1[54096] = 32'b11111111111111111010011011001010;
assign LUT_1[54097] = 32'b11111111111111110011101101000110;
assign LUT_1[54098] = 32'b11111111111111110110001001011011;
assign LUT_1[54099] = 32'b11111111111111101111011011010111;
assign LUT_1[54100] = 32'b00000000000000000010010100100001;
assign LUT_1[54101] = 32'b11111111111111111011100110011101;
assign LUT_1[54102] = 32'b11111111111111111110000010110010;
assign LUT_1[54103] = 32'b11111111111111110111010100101110;
assign LUT_1[54104] = 32'b11111111111111111001101000111111;
assign LUT_1[54105] = 32'b11111111111111110010111010111011;
assign LUT_1[54106] = 32'b11111111111111110101010111010000;
assign LUT_1[54107] = 32'b11111111111111101110101001001100;
assign LUT_1[54108] = 32'b00000000000000000001100010010110;
assign LUT_1[54109] = 32'b11111111111111111010110100010010;
assign LUT_1[54110] = 32'b11111111111111111101010000100111;
assign LUT_1[54111] = 32'b11111111111111110110100010100011;
assign LUT_1[54112] = 32'b11111111111111111001011010100111;
assign LUT_1[54113] = 32'b11111111111111110010101100100011;
assign LUT_1[54114] = 32'b11111111111111110101001000111000;
assign LUT_1[54115] = 32'b11111111111111101110011010110100;
assign LUT_1[54116] = 32'b00000000000000000001010011111110;
assign LUT_1[54117] = 32'b11111111111111111010100101111010;
assign LUT_1[54118] = 32'b11111111111111111101000010001111;
assign LUT_1[54119] = 32'b11111111111111110110010100001011;
assign LUT_1[54120] = 32'b11111111111111111000101000011100;
assign LUT_1[54121] = 32'b11111111111111110001111010011000;
assign LUT_1[54122] = 32'b11111111111111110100010110101101;
assign LUT_1[54123] = 32'b11111111111111101101101000101001;
assign LUT_1[54124] = 32'b00000000000000000000100001110011;
assign LUT_1[54125] = 32'b11111111111111111001110011101111;
assign LUT_1[54126] = 32'b11111111111111111100010000000100;
assign LUT_1[54127] = 32'b11111111111111110101100010000000;
assign LUT_1[54128] = 32'b11111111111111111011010110001001;
assign LUT_1[54129] = 32'b11111111111111110100101000000101;
assign LUT_1[54130] = 32'b11111111111111110111000100011010;
assign LUT_1[54131] = 32'b11111111111111110000010110010110;
assign LUT_1[54132] = 32'b00000000000000000011001111100000;
assign LUT_1[54133] = 32'b11111111111111111100100001011100;
assign LUT_1[54134] = 32'b11111111111111111110111101110001;
assign LUT_1[54135] = 32'b11111111111111111000001111101101;
assign LUT_1[54136] = 32'b11111111111111111010100011111110;
assign LUT_1[54137] = 32'b11111111111111110011110101111010;
assign LUT_1[54138] = 32'b11111111111111110110010010001111;
assign LUT_1[54139] = 32'b11111111111111101111100100001011;
assign LUT_1[54140] = 32'b00000000000000000010011101010101;
assign LUT_1[54141] = 32'b11111111111111111011101111010001;
assign LUT_1[54142] = 32'b11111111111111111110001011100110;
assign LUT_1[54143] = 32'b11111111111111110111011101100010;
assign LUT_1[54144] = 32'b11111111111111111001100010000011;
assign LUT_1[54145] = 32'b11111111111111110010110011111111;
assign LUT_1[54146] = 32'b11111111111111110101010000010100;
assign LUT_1[54147] = 32'b11111111111111101110100010010000;
assign LUT_1[54148] = 32'b00000000000000000001011011011010;
assign LUT_1[54149] = 32'b11111111111111111010101101010110;
assign LUT_1[54150] = 32'b11111111111111111101001001101011;
assign LUT_1[54151] = 32'b11111111111111110110011011100111;
assign LUT_1[54152] = 32'b11111111111111111000101111111000;
assign LUT_1[54153] = 32'b11111111111111110010000001110100;
assign LUT_1[54154] = 32'b11111111111111110100011110001001;
assign LUT_1[54155] = 32'b11111111111111101101110000000101;
assign LUT_1[54156] = 32'b00000000000000000000101001001111;
assign LUT_1[54157] = 32'b11111111111111111001111011001011;
assign LUT_1[54158] = 32'b11111111111111111100010111100000;
assign LUT_1[54159] = 32'b11111111111111110101101001011100;
assign LUT_1[54160] = 32'b11111111111111111011011101100101;
assign LUT_1[54161] = 32'b11111111111111110100101111100001;
assign LUT_1[54162] = 32'b11111111111111110111001011110110;
assign LUT_1[54163] = 32'b11111111111111110000011101110010;
assign LUT_1[54164] = 32'b00000000000000000011010110111100;
assign LUT_1[54165] = 32'b11111111111111111100101000111000;
assign LUT_1[54166] = 32'b11111111111111111111000101001101;
assign LUT_1[54167] = 32'b11111111111111111000010111001001;
assign LUT_1[54168] = 32'b11111111111111111010101011011010;
assign LUT_1[54169] = 32'b11111111111111110011111101010110;
assign LUT_1[54170] = 32'b11111111111111110110011001101011;
assign LUT_1[54171] = 32'b11111111111111101111101011100111;
assign LUT_1[54172] = 32'b00000000000000000010100100110001;
assign LUT_1[54173] = 32'b11111111111111111011110110101101;
assign LUT_1[54174] = 32'b11111111111111111110010011000010;
assign LUT_1[54175] = 32'b11111111111111110111100100111110;
assign LUT_1[54176] = 32'b11111111111111111010011101000010;
assign LUT_1[54177] = 32'b11111111111111110011101110111110;
assign LUT_1[54178] = 32'b11111111111111110110001011010011;
assign LUT_1[54179] = 32'b11111111111111101111011101001111;
assign LUT_1[54180] = 32'b00000000000000000010010110011001;
assign LUT_1[54181] = 32'b11111111111111111011101000010101;
assign LUT_1[54182] = 32'b11111111111111111110000100101010;
assign LUT_1[54183] = 32'b11111111111111110111010110100110;
assign LUT_1[54184] = 32'b11111111111111111001101010110111;
assign LUT_1[54185] = 32'b11111111111111110010111100110011;
assign LUT_1[54186] = 32'b11111111111111110101011001001000;
assign LUT_1[54187] = 32'b11111111111111101110101011000100;
assign LUT_1[54188] = 32'b00000000000000000001100100001110;
assign LUT_1[54189] = 32'b11111111111111111010110110001010;
assign LUT_1[54190] = 32'b11111111111111111101010010011111;
assign LUT_1[54191] = 32'b11111111111111110110100100011011;
assign LUT_1[54192] = 32'b11111111111111111100011000100100;
assign LUT_1[54193] = 32'b11111111111111110101101010100000;
assign LUT_1[54194] = 32'b11111111111111111000000110110101;
assign LUT_1[54195] = 32'b11111111111111110001011000110001;
assign LUT_1[54196] = 32'b00000000000000000100010001111011;
assign LUT_1[54197] = 32'b11111111111111111101100011110111;
assign LUT_1[54198] = 32'b00000000000000000000000000001100;
assign LUT_1[54199] = 32'b11111111111111111001010010001000;
assign LUT_1[54200] = 32'b11111111111111111011100110011001;
assign LUT_1[54201] = 32'b11111111111111110100111000010101;
assign LUT_1[54202] = 32'b11111111111111110111010100101010;
assign LUT_1[54203] = 32'b11111111111111110000100110100110;
assign LUT_1[54204] = 32'b00000000000000000011011111110000;
assign LUT_1[54205] = 32'b11111111111111111100110001101100;
assign LUT_1[54206] = 32'b11111111111111111111001110000001;
assign LUT_1[54207] = 32'b11111111111111111000011111111101;
assign LUT_1[54208] = 32'b11111111111111111011011111101011;
assign LUT_1[54209] = 32'b11111111111111110100110001100111;
assign LUT_1[54210] = 32'b11111111111111110111001101111100;
assign LUT_1[54211] = 32'b11111111111111110000011111111000;
assign LUT_1[54212] = 32'b00000000000000000011011001000010;
assign LUT_1[54213] = 32'b11111111111111111100101010111110;
assign LUT_1[54214] = 32'b11111111111111111111000111010011;
assign LUT_1[54215] = 32'b11111111111111111000011001001111;
assign LUT_1[54216] = 32'b11111111111111111010101101100000;
assign LUT_1[54217] = 32'b11111111111111110011111111011100;
assign LUT_1[54218] = 32'b11111111111111110110011011110001;
assign LUT_1[54219] = 32'b11111111111111101111101101101101;
assign LUT_1[54220] = 32'b00000000000000000010100110110111;
assign LUT_1[54221] = 32'b11111111111111111011111000110011;
assign LUT_1[54222] = 32'b11111111111111111110010101001000;
assign LUT_1[54223] = 32'b11111111111111110111100111000100;
assign LUT_1[54224] = 32'b11111111111111111101011011001101;
assign LUT_1[54225] = 32'b11111111111111110110101101001001;
assign LUT_1[54226] = 32'b11111111111111111001001001011110;
assign LUT_1[54227] = 32'b11111111111111110010011011011010;
assign LUT_1[54228] = 32'b00000000000000000101010100100100;
assign LUT_1[54229] = 32'b11111111111111111110100110100000;
assign LUT_1[54230] = 32'b00000000000000000001000010110101;
assign LUT_1[54231] = 32'b11111111111111111010010100110001;
assign LUT_1[54232] = 32'b11111111111111111100101001000010;
assign LUT_1[54233] = 32'b11111111111111110101111010111110;
assign LUT_1[54234] = 32'b11111111111111111000010111010011;
assign LUT_1[54235] = 32'b11111111111111110001101001001111;
assign LUT_1[54236] = 32'b00000000000000000100100010011001;
assign LUT_1[54237] = 32'b11111111111111111101110100010101;
assign LUT_1[54238] = 32'b00000000000000000000010000101010;
assign LUT_1[54239] = 32'b11111111111111111001100010100110;
assign LUT_1[54240] = 32'b11111111111111111100011010101010;
assign LUT_1[54241] = 32'b11111111111111110101101100100110;
assign LUT_1[54242] = 32'b11111111111111111000001000111011;
assign LUT_1[54243] = 32'b11111111111111110001011010110111;
assign LUT_1[54244] = 32'b00000000000000000100010100000001;
assign LUT_1[54245] = 32'b11111111111111111101100101111101;
assign LUT_1[54246] = 32'b00000000000000000000000010010010;
assign LUT_1[54247] = 32'b11111111111111111001010100001110;
assign LUT_1[54248] = 32'b11111111111111111011101000011111;
assign LUT_1[54249] = 32'b11111111111111110100111010011011;
assign LUT_1[54250] = 32'b11111111111111110111010110110000;
assign LUT_1[54251] = 32'b11111111111111110000101000101100;
assign LUT_1[54252] = 32'b00000000000000000011100001110110;
assign LUT_1[54253] = 32'b11111111111111111100110011110010;
assign LUT_1[54254] = 32'b11111111111111111111010000000111;
assign LUT_1[54255] = 32'b11111111111111111000100010000011;
assign LUT_1[54256] = 32'b11111111111111111110010110001100;
assign LUT_1[54257] = 32'b11111111111111110111101000001000;
assign LUT_1[54258] = 32'b11111111111111111010000100011101;
assign LUT_1[54259] = 32'b11111111111111110011010110011001;
assign LUT_1[54260] = 32'b00000000000000000110001111100011;
assign LUT_1[54261] = 32'b11111111111111111111100001011111;
assign LUT_1[54262] = 32'b00000000000000000001111101110100;
assign LUT_1[54263] = 32'b11111111111111111011001111110000;
assign LUT_1[54264] = 32'b11111111111111111101100100000001;
assign LUT_1[54265] = 32'b11111111111111110110110101111101;
assign LUT_1[54266] = 32'b11111111111111111001010010010010;
assign LUT_1[54267] = 32'b11111111111111110010100100001110;
assign LUT_1[54268] = 32'b00000000000000000101011101011000;
assign LUT_1[54269] = 32'b11111111111111111110101111010100;
assign LUT_1[54270] = 32'b00000000000000000001001011101001;
assign LUT_1[54271] = 32'b11111111111111111010011101100101;
assign LUT_1[54272] = 32'b00000000000000000101010110000111;
assign LUT_1[54273] = 32'b11111111111111111110101000000011;
assign LUT_1[54274] = 32'b00000000000000000001000100011000;
assign LUT_1[54275] = 32'b11111111111111111010010110010100;
assign LUT_1[54276] = 32'b00000000000000001101001111011110;
assign LUT_1[54277] = 32'b00000000000000000110100001011010;
assign LUT_1[54278] = 32'b00000000000000001000111101101111;
assign LUT_1[54279] = 32'b00000000000000000010001111101011;
assign LUT_1[54280] = 32'b00000000000000000100100011111100;
assign LUT_1[54281] = 32'b11111111111111111101110101111000;
assign LUT_1[54282] = 32'b00000000000000000000010010001101;
assign LUT_1[54283] = 32'b11111111111111111001100100001001;
assign LUT_1[54284] = 32'b00000000000000001100011101010011;
assign LUT_1[54285] = 32'b00000000000000000101101111001111;
assign LUT_1[54286] = 32'b00000000000000001000001011100100;
assign LUT_1[54287] = 32'b00000000000000000001011101100000;
assign LUT_1[54288] = 32'b00000000000000000111010001101001;
assign LUT_1[54289] = 32'b00000000000000000000100011100101;
assign LUT_1[54290] = 32'b00000000000000000010111111111010;
assign LUT_1[54291] = 32'b11111111111111111100010001110110;
assign LUT_1[54292] = 32'b00000000000000001111001011000000;
assign LUT_1[54293] = 32'b00000000000000001000011100111100;
assign LUT_1[54294] = 32'b00000000000000001010111001010001;
assign LUT_1[54295] = 32'b00000000000000000100001011001101;
assign LUT_1[54296] = 32'b00000000000000000110011111011110;
assign LUT_1[54297] = 32'b11111111111111111111110001011010;
assign LUT_1[54298] = 32'b00000000000000000010001101101111;
assign LUT_1[54299] = 32'b11111111111111111011011111101011;
assign LUT_1[54300] = 32'b00000000000000001110011000110101;
assign LUT_1[54301] = 32'b00000000000000000111101010110001;
assign LUT_1[54302] = 32'b00000000000000001010000111000110;
assign LUT_1[54303] = 32'b00000000000000000011011001000010;
assign LUT_1[54304] = 32'b00000000000000000110010001000110;
assign LUT_1[54305] = 32'b11111111111111111111100011000010;
assign LUT_1[54306] = 32'b00000000000000000001111111010111;
assign LUT_1[54307] = 32'b11111111111111111011010001010011;
assign LUT_1[54308] = 32'b00000000000000001110001010011101;
assign LUT_1[54309] = 32'b00000000000000000111011100011001;
assign LUT_1[54310] = 32'b00000000000000001001111000101110;
assign LUT_1[54311] = 32'b00000000000000000011001010101010;
assign LUT_1[54312] = 32'b00000000000000000101011110111011;
assign LUT_1[54313] = 32'b11111111111111111110110000110111;
assign LUT_1[54314] = 32'b00000000000000000001001101001100;
assign LUT_1[54315] = 32'b11111111111111111010011111001000;
assign LUT_1[54316] = 32'b00000000000000001101011000010010;
assign LUT_1[54317] = 32'b00000000000000000110101010001110;
assign LUT_1[54318] = 32'b00000000000000001001000110100011;
assign LUT_1[54319] = 32'b00000000000000000010011000011111;
assign LUT_1[54320] = 32'b00000000000000001000001100101000;
assign LUT_1[54321] = 32'b00000000000000000001011110100100;
assign LUT_1[54322] = 32'b00000000000000000011111010111001;
assign LUT_1[54323] = 32'b11111111111111111101001100110101;
assign LUT_1[54324] = 32'b00000000000000010000000101111111;
assign LUT_1[54325] = 32'b00000000000000001001010111111011;
assign LUT_1[54326] = 32'b00000000000000001011110100010000;
assign LUT_1[54327] = 32'b00000000000000000101000110001100;
assign LUT_1[54328] = 32'b00000000000000000111011010011101;
assign LUT_1[54329] = 32'b00000000000000000000101100011001;
assign LUT_1[54330] = 32'b00000000000000000011001000101110;
assign LUT_1[54331] = 32'b11111111111111111100011010101010;
assign LUT_1[54332] = 32'b00000000000000001111010011110100;
assign LUT_1[54333] = 32'b00000000000000001000100101110000;
assign LUT_1[54334] = 32'b00000000000000001011000010000101;
assign LUT_1[54335] = 32'b00000000000000000100010100000001;
assign LUT_1[54336] = 32'b00000000000000000111010011101111;
assign LUT_1[54337] = 32'b00000000000000000000100101101011;
assign LUT_1[54338] = 32'b00000000000000000011000010000000;
assign LUT_1[54339] = 32'b11111111111111111100010011111100;
assign LUT_1[54340] = 32'b00000000000000001111001101000110;
assign LUT_1[54341] = 32'b00000000000000001000011111000010;
assign LUT_1[54342] = 32'b00000000000000001010111011010111;
assign LUT_1[54343] = 32'b00000000000000000100001101010011;
assign LUT_1[54344] = 32'b00000000000000000110100001100100;
assign LUT_1[54345] = 32'b11111111111111111111110011100000;
assign LUT_1[54346] = 32'b00000000000000000010001111110101;
assign LUT_1[54347] = 32'b11111111111111111011100001110001;
assign LUT_1[54348] = 32'b00000000000000001110011010111011;
assign LUT_1[54349] = 32'b00000000000000000111101100110111;
assign LUT_1[54350] = 32'b00000000000000001010001001001100;
assign LUT_1[54351] = 32'b00000000000000000011011011001000;
assign LUT_1[54352] = 32'b00000000000000001001001111010001;
assign LUT_1[54353] = 32'b00000000000000000010100001001101;
assign LUT_1[54354] = 32'b00000000000000000100111101100010;
assign LUT_1[54355] = 32'b11111111111111111110001111011110;
assign LUT_1[54356] = 32'b00000000000000010001001000101000;
assign LUT_1[54357] = 32'b00000000000000001010011010100100;
assign LUT_1[54358] = 32'b00000000000000001100110110111001;
assign LUT_1[54359] = 32'b00000000000000000110001000110101;
assign LUT_1[54360] = 32'b00000000000000001000011101000110;
assign LUT_1[54361] = 32'b00000000000000000001101111000010;
assign LUT_1[54362] = 32'b00000000000000000100001011010111;
assign LUT_1[54363] = 32'b11111111111111111101011101010011;
assign LUT_1[54364] = 32'b00000000000000010000010110011101;
assign LUT_1[54365] = 32'b00000000000000001001101000011001;
assign LUT_1[54366] = 32'b00000000000000001100000100101110;
assign LUT_1[54367] = 32'b00000000000000000101010110101010;
assign LUT_1[54368] = 32'b00000000000000001000001110101110;
assign LUT_1[54369] = 32'b00000000000000000001100000101010;
assign LUT_1[54370] = 32'b00000000000000000011111100111111;
assign LUT_1[54371] = 32'b11111111111111111101001110111011;
assign LUT_1[54372] = 32'b00000000000000010000001000000101;
assign LUT_1[54373] = 32'b00000000000000001001011010000001;
assign LUT_1[54374] = 32'b00000000000000001011110110010110;
assign LUT_1[54375] = 32'b00000000000000000101001000010010;
assign LUT_1[54376] = 32'b00000000000000000111011100100011;
assign LUT_1[54377] = 32'b00000000000000000000101110011111;
assign LUT_1[54378] = 32'b00000000000000000011001010110100;
assign LUT_1[54379] = 32'b11111111111111111100011100110000;
assign LUT_1[54380] = 32'b00000000000000001111010101111010;
assign LUT_1[54381] = 32'b00000000000000001000100111110110;
assign LUT_1[54382] = 32'b00000000000000001011000100001011;
assign LUT_1[54383] = 32'b00000000000000000100010110000111;
assign LUT_1[54384] = 32'b00000000000000001010001010010000;
assign LUT_1[54385] = 32'b00000000000000000011011100001100;
assign LUT_1[54386] = 32'b00000000000000000101111000100001;
assign LUT_1[54387] = 32'b11111111111111111111001010011101;
assign LUT_1[54388] = 32'b00000000000000010010000011100111;
assign LUT_1[54389] = 32'b00000000000000001011010101100011;
assign LUT_1[54390] = 32'b00000000000000001101110001111000;
assign LUT_1[54391] = 32'b00000000000000000111000011110100;
assign LUT_1[54392] = 32'b00000000000000001001011000000101;
assign LUT_1[54393] = 32'b00000000000000000010101010000001;
assign LUT_1[54394] = 32'b00000000000000000101000110010110;
assign LUT_1[54395] = 32'b11111111111111111110011000010010;
assign LUT_1[54396] = 32'b00000000000000010001010001011100;
assign LUT_1[54397] = 32'b00000000000000001010100011011000;
assign LUT_1[54398] = 32'b00000000000000001100111111101101;
assign LUT_1[54399] = 32'b00000000000000000110010001101001;
assign LUT_1[54400] = 32'b00000000000000001000010110001010;
assign LUT_1[54401] = 32'b00000000000000000001101000000110;
assign LUT_1[54402] = 32'b00000000000000000100000100011011;
assign LUT_1[54403] = 32'b11111111111111111101010110010111;
assign LUT_1[54404] = 32'b00000000000000010000001111100001;
assign LUT_1[54405] = 32'b00000000000000001001100001011101;
assign LUT_1[54406] = 32'b00000000000000001011111101110010;
assign LUT_1[54407] = 32'b00000000000000000101001111101110;
assign LUT_1[54408] = 32'b00000000000000000111100011111111;
assign LUT_1[54409] = 32'b00000000000000000000110101111011;
assign LUT_1[54410] = 32'b00000000000000000011010010010000;
assign LUT_1[54411] = 32'b11111111111111111100100100001100;
assign LUT_1[54412] = 32'b00000000000000001111011101010110;
assign LUT_1[54413] = 32'b00000000000000001000101111010010;
assign LUT_1[54414] = 32'b00000000000000001011001011100111;
assign LUT_1[54415] = 32'b00000000000000000100011101100011;
assign LUT_1[54416] = 32'b00000000000000001010010001101100;
assign LUT_1[54417] = 32'b00000000000000000011100011101000;
assign LUT_1[54418] = 32'b00000000000000000101111111111101;
assign LUT_1[54419] = 32'b11111111111111111111010001111001;
assign LUT_1[54420] = 32'b00000000000000010010001011000011;
assign LUT_1[54421] = 32'b00000000000000001011011100111111;
assign LUT_1[54422] = 32'b00000000000000001101111001010100;
assign LUT_1[54423] = 32'b00000000000000000111001011010000;
assign LUT_1[54424] = 32'b00000000000000001001011111100001;
assign LUT_1[54425] = 32'b00000000000000000010110001011101;
assign LUT_1[54426] = 32'b00000000000000000101001101110010;
assign LUT_1[54427] = 32'b11111111111111111110011111101110;
assign LUT_1[54428] = 32'b00000000000000010001011000111000;
assign LUT_1[54429] = 32'b00000000000000001010101010110100;
assign LUT_1[54430] = 32'b00000000000000001101000111001001;
assign LUT_1[54431] = 32'b00000000000000000110011001000101;
assign LUT_1[54432] = 32'b00000000000000001001010001001001;
assign LUT_1[54433] = 32'b00000000000000000010100011000101;
assign LUT_1[54434] = 32'b00000000000000000100111111011010;
assign LUT_1[54435] = 32'b11111111111111111110010001010110;
assign LUT_1[54436] = 32'b00000000000000010001001010100000;
assign LUT_1[54437] = 32'b00000000000000001010011100011100;
assign LUT_1[54438] = 32'b00000000000000001100111000110001;
assign LUT_1[54439] = 32'b00000000000000000110001010101101;
assign LUT_1[54440] = 32'b00000000000000001000011110111110;
assign LUT_1[54441] = 32'b00000000000000000001110000111010;
assign LUT_1[54442] = 32'b00000000000000000100001101001111;
assign LUT_1[54443] = 32'b11111111111111111101011111001011;
assign LUT_1[54444] = 32'b00000000000000010000011000010101;
assign LUT_1[54445] = 32'b00000000000000001001101010010001;
assign LUT_1[54446] = 32'b00000000000000001100000110100110;
assign LUT_1[54447] = 32'b00000000000000000101011000100010;
assign LUT_1[54448] = 32'b00000000000000001011001100101011;
assign LUT_1[54449] = 32'b00000000000000000100011110100111;
assign LUT_1[54450] = 32'b00000000000000000110111010111100;
assign LUT_1[54451] = 32'b00000000000000000000001100111000;
assign LUT_1[54452] = 32'b00000000000000010011000110000010;
assign LUT_1[54453] = 32'b00000000000000001100010111111110;
assign LUT_1[54454] = 32'b00000000000000001110110100010011;
assign LUT_1[54455] = 32'b00000000000000001000000110001111;
assign LUT_1[54456] = 32'b00000000000000001010011010100000;
assign LUT_1[54457] = 32'b00000000000000000011101100011100;
assign LUT_1[54458] = 32'b00000000000000000110001000110001;
assign LUT_1[54459] = 32'b11111111111111111111011010101101;
assign LUT_1[54460] = 32'b00000000000000010010010011110111;
assign LUT_1[54461] = 32'b00000000000000001011100101110011;
assign LUT_1[54462] = 32'b00000000000000001110000010001000;
assign LUT_1[54463] = 32'b00000000000000000111010100000100;
assign LUT_1[54464] = 32'b00000000000000001010010011110010;
assign LUT_1[54465] = 32'b00000000000000000011100101101110;
assign LUT_1[54466] = 32'b00000000000000000110000010000011;
assign LUT_1[54467] = 32'b11111111111111111111010011111111;
assign LUT_1[54468] = 32'b00000000000000010010001101001001;
assign LUT_1[54469] = 32'b00000000000000001011011111000101;
assign LUT_1[54470] = 32'b00000000000000001101111011011010;
assign LUT_1[54471] = 32'b00000000000000000111001101010110;
assign LUT_1[54472] = 32'b00000000000000001001100001100111;
assign LUT_1[54473] = 32'b00000000000000000010110011100011;
assign LUT_1[54474] = 32'b00000000000000000101001111111000;
assign LUT_1[54475] = 32'b11111111111111111110100001110100;
assign LUT_1[54476] = 32'b00000000000000010001011010111110;
assign LUT_1[54477] = 32'b00000000000000001010101100111010;
assign LUT_1[54478] = 32'b00000000000000001101001001001111;
assign LUT_1[54479] = 32'b00000000000000000110011011001011;
assign LUT_1[54480] = 32'b00000000000000001100001111010100;
assign LUT_1[54481] = 32'b00000000000000000101100001010000;
assign LUT_1[54482] = 32'b00000000000000000111111101100101;
assign LUT_1[54483] = 32'b00000000000000000001001111100001;
assign LUT_1[54484] = 32'b00000000000000010100001000101011;
assign LUT_1[54485] = 32'b00000000000000001101011010100111;
assign LUT_1[54486] = 32'b00000000000000001111110110111100;
assign LUT_1[54487] = 32'b00000000000000001001001000111000;
assign LUT_1[54488] = 32'b00000000000000001011011101001001;
assign LUT_1[54489] = 32'b00000000000000000100101111000101;
assign LUT_1[54490] = 32'b00000000000000000111001011011010;
assign LUT_1[54491] = 32'b00000000000000000000011101010110;
assign LUT_1[54492] = 32'b00000000000000010011010110100000;
assign LUT_1[54493] = 32'b00000000000000001100101000011100;
assign LUT_1[54494] = 32'b00000000000000001111000100110001;
assign LUT_1[54495] = 32'b00000000000000001000010110101101;
assign LUT_1[54496] = 32'b00000000000000001011001110110001;
assign LUT_1[54497] = 32'b00000000000000000100100000101101;
assign LUT_1[54498] = 32'b00000000000000000110111101000010;
assign LUT_1[54499] = 32'b00000000000000000000001110111110;
assign LUT_1[54500] = 32'b00000000000000010011001000001000;
assign LUT_1[54501] = 32'b00000000000000001100011010000100;
assign LUT_1[54502] = 32'b00000000000000001110110110011001;
assign LUT_1[54503] = 32'b00000000000000001000001000010101;
assign LUT_1[54504] = 32'b00000000000000001010011100100110;
assign LUT_1[54505] = 32'b00000000000000000011101110100010;
assign LUT_1[54506] = 32'b00000000000000000110001010110111;
assign LUT_1[54507] = 32'b11111111111111111111011100110011;
assign LUT_1[54508] = 32'b00000000000000010010010101111101;
assign LUT_1[54509] = 32'b00000000000000001011100111111001;
assign LUT_1[54510] = 32'b00000000000000001110000100001110;
assign LUT_1[54511] = 32'b00000000000000000111010110001010;
assign LUT_1[54512] = 32'b00000000000000001101001010010011;
assign LUT_1[54513] = 32'b00000000000000000110011100001111;
assign LUT_1[54514] = 32'b00000000000000001000111000100100;
assign LUT_1[54515] = 32'b00000000000000000010001010100000;
assign LUT_1[54516] = 32'b00000000000000010101000011101010;
assign LUT_1[54517] = 32'b00000000000000001110010101100110;
assign LUT_1[54518] = 32'b00000000000000010000110001111011;
assign LUT_1[54519] = 32'b00000000000000001010000011110111;
assign LUT_1[54520] = 32'b00000000000000001100011000001000;
assign LUT_1[54521] = 32'b00000000000000000101101010000100;
assign LUT_1[54522] = 32'b00000000000000001000000110011001;
assign LUT_1[54523] = 32'b00000000000000000001011000010101;
assign LUT_1[54524] = 32'b00000000000000010100010001011111;
assign LUT_1[54525] = 32'b00000000000000001101100011011011;
assign LUT_1[54526] = 32'b00000000000000001111111111110000;
assign LUT_1[54527] = 32'b00000000000000001001010001101100;
assign LUT_1[54528] = 32'b00000000000000000011001010010011;
assign LUT_1[54529] = 32'b11111111111111111100011100001111;
assign LUT_1[54530] = 32'b11111111111111111110111000100100;
assign LUT_1[54531] = 32'b11111111111111111000001010100000;
assign LUT_1[54532] = 32'b00000000000000001011000011101010;
assign LUT_1[54533] = 32'b00000000000000000100010101100110;
assign LUT_1[54534] = 32'b00000000000000000110110001111011;
assign LUT_1[54535] = 32'b00000000000000000000000011110111;
assign LUT_1[54536] = 32'b00000000000000000010011000001000;
assign LUT_1[54537] = 32'b11111111111111111011101010000100;
assign LUT_1[54538] = 32'b11111111111111111110000110011001;
assign LUT_1[54539] = 32'b11111111111111110111011000010101;
assign LUT_1[54540] = 32'b00000000000000001010010001011111;
assign LUT_1[54541] = 32'b00000000000000000011100011011011;
assign LUT_1[54542] = 32'b00000000000000000101111111110000;
assign LUT_1[54543] = 32'b11111111111111111111010001101100;
assign LUT_1[54544] = 32'b00000000000000000101000101110101;
assign LUT_1[54545] = 32'b11111111111111111110010111110001;
assign LUT_1[54546] = 32'b00000000000000000000110100000110;
assign LUT_1[54547] = 32'b11111111111111111010000110000010;
assign LUT_1[54548] = 32'b00000000000000001100111111001100;
assign LUT_1[54549] = 32'b00000000000000000110010001001000;
assign LUT_1[54550] = 32'b00000000000000001000101101011101;
assign LUT_1[54551] = 32'b00000000000000000001111111011001;
assign LUT_1[54552] = 32'b00000000000000000100010011101010;
assign LUT_1[54553] = 32'b11111111111111111101100101100110;
assign LUT_1[54554] = 32'b00000000000000000000000001111011;
assign LUT_1[54555] = 32'b11111111111111111001010011110111;
assign LUT_1[54556] = 32'b00000000000000001100001101000001;
assign LUT_1[54557] = 32'b00000000000000000101011110111101;
assign LUT_1[54558] = 32'b00000000000000000111111011010010;
assign LUT_1[54559] = 32'b00000000000000000001001101001110;
assign LUT_1[54560] = 32'b00000000000000000100000101010010;
assign LUT_1[54561] = 32'b11111111111111111101010111001110;
assign LUT_1[54562] = 32'b11111111111111111111110011100011;
assign LUT_1[54563] = 32'b11111111111111111001000101011111;
assign LUT_1[54564] = 32'b00000000000000001011111110101001;
assign LUT_1[54565] = 32'b00000000000000000101010000100101;
assign LUT_1[54566] = 32'b00000000000000000111101100111010;
assign LUT_1[54567] = 32'b00000000000000000000111110110110;
assign LUT_1[54568] = 32'b00000000000000000011010011000111;
assign LUT_1[54569] = 32'b11111111111111111100100101000011;
assign LUT_1[54570] = 32'b11111111111111111111000001011000;
assign LUT_1[54571] = 32'b11111111111111111000010011010100;
assign LUT_1[54572] = 32'b00000000000000001011001100011110;
assign LUT_1[54573] = 32'b00000000000000000100011110011010;
assign LUT_1[54574] = 32'b00000000000000000110111010101111;
assign LUT_1[54575] = 32'b00000000000000000000001100101011;
assign LUT_1[54576] = 32'b00000000000000000110000000110100;
assign LUT_1[54577] = 32'b11111111111111111111010010110000;
assign LUT_1[54578] = 32'b00000000000000000001101111000101;
assign LUT_1[54579] = 32'b11111111111111111011000001000001;
assign LUT_1[54580] = 32'b00000000000000001101111010001011;
assign LUT_1[54581] = 32'b00000000000000000111001100000111;
assign LUT_1[54582] = 32'b00000000000000001001101000011100;
assign LUT_1[54583] = 32'b00000000000000000010111010011000;
assign LUT_1[54584] = 32'b00000000000000000101001110101001;
assign LUT_1[54585] = 32'b11111111111111111110100000100101;
assign LUT_1[54586] = 32'b00000000000000000000111100111010;
assign LUT_1[54587] = 32'b11111111111111111010001110110110;
assign LUT_1[54588] = 32'b00000000000000001101001000000000;
assign LUT_1[54589] = 32'b00000000000000000110011001111100;
assign LUT_1[54590] = 32'b00000000000000001000110110010001;
assign LUT_1[54591] = 32'b00000000000000000010001000001101;
assign LUT_1[54592] = 32'b00000000000000000101000111111011;
assign LUT_1[54593] = 32'b11111111111111111110011001110111;
assign LUT_1[54594] = 32'b00000000000000000000110110001100;
assign LUT_1[54595] = 32'b11111111111111111010001000001000;
assign LUT_1[54596] = 32'b00000000000000001101000001010010;
assign LUT_1[54597] = 32'b00000000000000000110010011001110;
assign LUT_1[54598] = 32'b00000000000000001000101111100011;
assign LUT_1[54599] = 32'b00000000000000000010000001011111;
assign LUT_1[54600] = 32'b00000000000000000100010101110000;
assign LUT_1[54601] = 32'b11111111111111111101100111101100;
assign LUT_1[54602] = 32'b00000000000000000000000100000001;
assign LUT_1[54603] = 32'b11111111111111111001010101111101;
assign LUT_1[54604] = 32'b00000000000000001100001111000111;
assign LUT_1[54605] = 32'b00000000000000000101100001000011;
assign LUT_1[54606] = 32'b00000000000000000111111101011000;
assign LUT_1[54607] = 32'b00000000000000000001001111010100;
assign LUT_1[54608] = 32'b00000000000000000111000011011101;
assign LUT_1[54609] = 32'b00000000000000000000010101011001;
assign LUT_1[54610] = 32'b00000000000000000010110001101110;
assign LUT_1[54611] = 32'b11111111111111111100000011101010;
assign LUT_1[54612] = 32'b00000000000000001110111100110100;
assign LUT_1[54613] = 32'b00000000000000001000001110110000;
assign LUT_1[54614] = 32'b00000000000000001010101011000101;
assign LUT_1[54615] = 32'b00000000000000000011111101000001;
assign LUT_1[54616] = 32'b00000000000000000110010001010010;
assign LUT_1[54617] = 32'b11111111111111111111100011001110;
assign LUT_1[54618] = 32'b00000000000000000001111111100011;
assign LUT_1[54619] = 32'b11111111111111111011010001011111;
assign LUT_1[54620] = 32'b00000000000000001110001010101001;
assign LUT_1[54621] = 32'b00000000000000000111011100100101;
assign LUT_1[54622] = 32'b00000000000000001001111000111010;
assign LUT_1[54623] = 32'b00000000000000000011001010110110;
assign LUT_1[54624] = 32'b00000000000000000110000010111010;
assign LUT_1[54625] = 32'b11111111111111111111010100110110;
assign LUT_1[54626] = 32'b00000000000000000001110001001011;
assign LUT_1[54627] = 32'b11111111111111111011000011000111;
assign LUT_1[54628] = 32'b00000000000000001101111100010001;
assign LUT_1[54629] = 32'b00000000000000000111001110001101;
assign LUT_1[54630] = 32'b00000000000000001001101010100010;
assign LUT_1[54631] = 32'b00000000000000000010111100011110;
assign LUT_1[54632] = 32'b00000000000000000101010000101111;
assign LUT_1[54633] = 32'b11111111111111111110100010101011;
assign LUT_1[54634] = 32'b00000000000000000000111111000000;
assign LUT_1[54635] = 32'b11111111111111111010010000111100;
assign LUT_1[54636] = 32'b00000000000000001101001010000110;
assign LUT_1[54637] = 32'b00000000000000000110011100000010;
assign LUT_1[54638] = 32'b00000000000000001000111000010111;
assign LUT_1[54639] = 32'b00000000000000000010001010010011;
assign LUT_1[54640] = 32'b00000000000000000111111110011100;
assign LUT_1[54641] = 32'b00000000000000000001010000011000;
assign LUT_1[54642] = 32'b00000000000000000011101100101101;
assign LUT_1[54643] = 32'b11111111111111111100111110101001;
assign LUT_1[54644] = 32'b00000000000000001111110111110011;
assign LUT_1[54645] = 32'b00000000000000001001001001101111;
assign LUT_1[54646] = 32'b00000000000000001011100110000100;
assign LUT_1[54647] = 32'b00000000000000000100111000000000;
assign LUT_1[54648] = 32'b00000000000000000111001100010001;
assign LUT_1[54649] = 32'b00000000000000000000011110001101;
assign LUT_1[54650] = 32'b00000000000000000010111010100010;
assign LUT_1[54651] = 32'b11111111111111111100001100011110;
assign LUT_1[54652] = 32'b00000000000000001111000101101000;
assign LUT_1[54653] = 32'b00000000000000001000010111100100;
assign LUT_1[54654] = 32'b00000000000000001010110011111001;
assign LUT_1[54655] = 32'b00000000000000000100000101110101;
assign LUT_1[54656] = 32'b00000000000000000110001010010110;
assign LUT_1[54657] = 32'b11111111111111111111011100010010;
assign LUT_1[54658] = 32'b00000000000000000001111000100111;
assign LUT_1[54659] = 32'b11111111111111111011001010100011;
assign LUT_1[54660] = 32'b00000000000000001110000011101101;
assign LUT_1[54661] = 32'b00000000000000000111010101101001;
assign LUT_1[54662] = 32'b00000000000000001001110001111110;
assign LUT_1[54663] = 32'b00000000000000000011000011111010;
assign LUT_1[54664] = 32'b00000000000000000101011000001011;
assign LUT_1[54665] = 32'b11111111111111111110101010000111;
assign LUT_1[54666] = 32'b00000000000000000001000110011100;
assign LUT_1[54667] = 32'b11111111111111111010011000011000;
assign LUT_1[54668] = 32'b00000000000000001101010001100010;
assign LUT_1[54669] = 32'b00000000000000000110100011011110;
assign LUT_1[54670] = 32'b00000000000000001000111111110011;
assign LUT_1[54671] = 32'b00000000000000000010010001101111;
assign LUT_1[54672] = 32'b00000000000000001000000101111000;
assign LUT_1[54673] = 32'b00000000000000000001010111110100;
assign LUT_1[54674] = 32'b00000000000000000011110100001001;
assign LUT_1[54675] = 32'b11111111111111111101000110000101;
assign LUT_1[54676] = 32'b00000000000000001111111111001111;
assign LUT_1[54677] = 32'b00000000000000001001010001001011;
assign LUT_1[54678] = 32'b00000000000000001011101101100000;
assign LUT_1[54679] = 32'b00000000000000000100111111011100;
assign LUT_1[54680] = 32'b00000000000000000111010011101101;
assign LUT_1[54681] = 32'b00000000000000000000100101101001;
assign LUT_1[54682] = 32'b00000000000000000011000001111110;
assign LUT_1[54683] = 32'b11111111111111111100010011111010;
assign LUT_1[54684] = 32'b00000000000000001111001101000100;
assign LUT_1[54685] = 32'b00000000000000001000011111000000;
assign LUT_1[54686] = 32'b00000000000000001010111011010101;
assign LUT_1[54687] = 32'b00000000000000000100001101010001;
assign LUT_1[54688] = 32'b00000000000000000111000101010101;
assign LUT_1[54689] = 32'b00000000000000000000010111010001;
assign LUT_1[54690] = 32'b00000000000000000010110011100110;
assign LUT_1[54691] = 32'b11111111111111111100000101100010;
assign LUT_1[54692] = 32'b00000000000000001110111110101100;
assign LUT_1[54693] = 32'b00000000000000001000010000101000;
assign LUT_1[54694] = 32'b00000000000000001010101100111101;
assign LUT_1[54695] = 32'b00000000000000000011111110111001;
assign LUT_1[54696] = 32'b00000000000000000110010011001010;
assign LUT_1[54697] = 32'b11111111111111111111100101000110;
assign LUT_1[54698] = 32'b00000000000000000010000001011011;
assign LUT_1[54699] = 32'b11111111111111111011010011010111;
assign LUT_1[54700] = 32'b00000000000000001110001100100001;
assign LUT_1[54701] = 32'b00000000000000000111011110011101;
assign LUT_1[54702] = 32'b00000000000000001001111010110010;
assign LUT_1[54703] = 32'b00000000000000000011001100101110;
assign LUT_1[54704] = 32'b00000000000000001001000000110111;
assign LUT_1[54705] = 32'b00000000000000000010010010110011;
assign LUT_1[54706] = 32'b00000000000000000100101111001000;
assign LUT_1[54707] = 32'b11111111111111111110000001000100;
assign LUT_1[54708] = 32'b00000000000000010000111010001110;
assign LUT_1[54709] = 32'b00000000000000001010001100001010;
assign LUT_1[54710] = 32'b00000000000000001100101000011111;
assign LUT_1[54711] = 32'b00000000000000000101111010011011;
assign LUT_1[54712] = 32'b00000000000000001000001110101100;
assign LUT_1[54713] = 32'b00000000000000000001100000101000;
assign LUT_1[54714] = 32'b00000000000000000011111100111101;
assign LUT_1[54715] = 32'b11111111111111111101001110111001;
assign LUT_1[54716] = 32'b00000000000000010000001000000011;
assign LUT_1[54717] = 32'b00000000000000001001011001111111;
assign LUT_1[54718] = 32'b00000000000000001011110110010100;
assign LUT_1[54719] = 32'b00000000000000000101001000010000;
assign LUT_1[54720] = 32'b00000000000000001000000111111110;
assign LUT_1[54721] = 32'b00000000000000000001011001111010;
assign LUT_1[54722] = 32'b00000000000000000011110110001111;
assign LUT_1[54723] = 32'b11111111111111111101001000001011;
assign LUT_1[54724] = 32'b00000000000000010000000001010101;
assign LUT_1[54725] = 32'b00000000000000001001010011010001;
assign LUT_1[54726] = 32'b00000000000000001011101111100110;
assign LUT_1[54727] = 32'b00000000000000000101000001100010;
assign LUT_1[54728] = 32'b00000000000000000111010101110011;
assign LUT_1[54729] = 32'b00000000000000000000100111101111;
assign LUT_1[54730] = 32'b00000000000000000011000100000100;
assign LUT_1[54731] = 32'b11111111111111111100010110000000;
assign LUT_1[54732] = 32'b00000000000000001111001111001010;
assign LUT_1[54733] = 32'b00000000000000001000100001000110;
assign LUT_1[54734] = 32'b00000000000000001010111101011011;
assign LUT_1[54735] = 32'b00000000000000000100001111010111;
assign LUT_1[54736] = 32'b00000000000000001010000011100000;
assign LUT_1[54737] = 32'b00000000000000000011010101011100;
assign LUT_1[54738] = 32'b00000000000000000101110001110001;
assign LUT_1[54739] = 32'b11111111111111111111000011101101;
assign LUT_1[54740] = 32'b00000000000000010001111100110111;
assign LUT_1[54741] = 32'b00000000000000001011001110110011;
assign LUT_1[54742] = 32'b00000000000000001101101011001000;
assign LUT_1[54743] = 32'b00000000000000000110111101000100;
assign LUT_1[54744] = 32'b00000000000000001001010001010101;
assign LUT_1[54745] = 32'b00000000000000000010100011010001;
assign LUT_1[54746] = 32'b00000000000000000100111111100110;
assign LUT_1[54747] = 32'b11111111111111111110010001100010;
assign LUT_1[54748] = 32'b00000000000000010001001010101100;
assign LUT_1[54749] = 32'b00000000000000001010011100101000;
assign LUT_1[54750] = 32'b00000000000000001100111000111101;
assign LUT_1[54751] = 32'b00000000000000000110001010111001;
assign LUT_1[54752] = 32'b00000000000000001001000010111101;
assign LUT_1[54753] = 32'b00000000000000000010010100111001;
assign LUT_1[54754] = 32'b00000000000000000100110001001110;
assign LUT_1[54755] = 32'b11111111111111111110000011001010;
assign LUT_1[54756] = 32'b00000000000000010000111100010100;
assign LUT_1[54757] = 32'b00000000000000001010001110010000;
assign LUT_1[54758] = 32'b00000000000000001100101010100101;
assign LUT_1[54759] = 32'b00000000000000000101111100100001;
assign LUT_1[54760] = 32'b00000000000000001000010000110010;
assign LUT_1[54761] = 32'b00000000000000000001100010101110;
assign LUT_1[54762] = 32'b00000000000000000011111111000011;
assign LUT_1[54763] = 32'b11111111111111111101010000111111;
assign LUT_1[54764] = 32'b00000000000000010000001010001001;
assign LUT_1[54765] = 32'b00000000000000001001011100000101;
assign LUT_1[54766] = 32'b00000000000000001011111000011010;
assign LUT_1[54767] = 32'b00000000000000000101001010010110;
assign LUT_1[54768] = 32'b00000000000000001010111110011111;
assign LUT_1[54769] = 32'b00000000000000000100010000011011;
assign LUT_1[54770] = 32'b00000000000000000110101100110000;
assign LUT_1[54771] = 32'b11111111111111111111111110101100;
assign LUT_1[54772] = 32'b00000000000000010010110111110110;
assign LUT_1[54773] = 32'b00000000000000001100001001110010;
assign LUT_1[54774] = 32'b00000000000000001110100110000111;
assign LUT_1[54775] = 32'b00000000000000000111111000000011;
assign LUT_1[54776] = 32'b00000000000000001010001100010100;
assign LUT_1[54777] = 32'b00000000000000000011011110010000;
assign LUT_1[54778] = 32'b00000000000000000101111010100101;
assign LUT_1[54779] = 32'b11111111111111111111001100100001;
assign LUT_1[54780] = 32'b00000000000000010010000101101011;
assign LUT_1[54781] = 32'b00000000000000001011010111100111;
assign LUT_1[54782] = 32'b00000000000000001101110011111100;
assign LUT_1[54783] = 32'b00000000000000000111000101111000;
assign LUT_1[54784] = 32'b11111111111111111111000100100100;
assign LUT_1[54785] = 32'b11111111111111111000010110100000;
assign LUT_1[54786] = 32'b11111111111111111010110010110101;
assign LUT_1[54787] = 32'b11111111111111110100000100110001;
assign LUT_1[54788] = 32'b00000000000000000110111101111011;
assign LUT_1[54789] = 32'b00000000000000000000001111110111;
assign LUT_1[54790] = 32'b00000000000000000010101100001100;
assign LUT_1[54791] = 32'b11111111111111111011111110001000;
assign LUT_1[54792] = 32'b11111111111111111110010010011001;
assign LUT_1[54793] = 32'b11111111111111110111100100010101;
assign LUT_1[54794] = 32'b11111111111111111010000000101010;
assign LUT_1[54795] = 32'b11111111111111110011010010100110;
assign LUT_1[54796] = 32'b00000000000000000110001011110000;
assign LUT_1[54797] = 32'b11111111111111111111011101101100;
assign LUT_1[54798] = 32'b00000000000000000001111010000001;
assign LUT_1[54799] = 32'b11111111111111111011001011111101;
assign LUT_1[54800] = 32'b00000000000000000001000000000110;
assign LUT_1[54801] = 32'b11111111111111111010010010000010;
assign LUT_1[54802] = 32'b11111111111111111100101110010111;
assign LUT_1[54803] = 32'b11111111111111110110000000010011;
assign LUT_1[54804] = 32'b00000000000000001000111001011101;
assign LUT_1[54805] = 32'b00000000000000000010001011011001;
assign LUT_1[54806] = 32'b00000000000000000100100111101110;
assign LUT_1[54807] = 32'b11111111111111111101111001101010;
assign LUT_1[54808] = 32'b00000000000000000000001101111011;
assign LUT_1[54809] = 32'b11111111111111111001011111110111;
assign LUT_1[54810] = 32'b11111111111111111011111100001100;
assign LUT_1[54811] = 32'b11111111111111110101001110001000;
assign LUT_1[54812] = 32'b00000000000000001000000111010010;
assign LUT_1[54813] = 32'b00000000000000000001011001001110;
assign LUT_1[54814] = 32'b00000000000000000011110101100011;
assign LUT_1[54815] = 32'b11111111111111111101000111011111;
assign LUT_1[54816] = 32'b11111111111111111111111111100011;
assign LUT_1[54817] = 32'b11111111111111111001010001011111;
assign LUT_1[54818] = 32'b11111111111111111011101101110100;
assign LUT_1[54819] = 32'b11111111111111110100111111110000;
assign LUT_1[54820] = 32'b00000000000000000111111000111010;
assign LUT_1[54821] = 32'b00000000000000000001001010110110;
assign LUT_1[54822] = 32'b00000000000000000011100111001011;
assign LUT_1[54823] = 32'b11111111111111111100111001000111;
assign LUT_1[54824] = 32'b11111111111111111111001101011000;
assign LUT_1[54825] = 32'b11111111111111111000011111010100;
assign LUT_1[54826] = 32'b11111111111111111010111011101001;
assign LUT_1[54827] = 32'b11111111111111110100001101100101;
assign LUT_1[54828] = 32'b00000000000000000111000110101111;
assign LUT_1[54829] = 32'b00000000000000000000011000101011;
assign LUT_1[54830] = 32'b00000000000000000010110101000000;
assign LUT_1[54831] = 32'b11111111111111111100000110111100;
assign LUT_1[54832] = 32'b00000000000000000001111011000101;
assign LUT_1[54833] = 32'b11111111111111111011001101000001;
assign LUT_1[54834] = 32'b11111111111111111101101001010110;
assign LUT_1[54835] = 32'b11111111111111110110111011010010;
assign LUT_1[54836] = 32'b00000000000000001001110100011100;
assign LUT_1[54837] = 32'b00000000000000000011000110011000;
assign LUT_1[54838] = 32'b00000000000000000101100010101101;
assign LUT_1[54839] = 32'b11111111111111111110110100101001;
assign LUT_1[54840] = 32'b00000000000000000001001000111010;
assign LUT_1[54841] = 32'b11111111111111111010011010110110;
assign LUT_1[54842] = 32'b11111111111111111100110111001011;
assign LUT_1[54843] = 32'b11111111111111110110001001000111;
assign LUT_1[54844] = 32'b00000000000000001001000010010001;
assign LUT_1[54845] = 32'b00000000000000000010010100001101;
assign LUT_1[54846] = 32'b00000000000000000100110000100010;
assign LUT_1[54847] = 32'b11111111111111111110000010011110;
assign LUT_1[54848] = 32'b00000000000000000001000010001100;
assign LUT_1[54849] = 32'b11111111111111111010010100001000;
assign LUT_1[54850] = 32'b11111111111111111100110000011101;
assign LUT_1[54851] = 32'b11111111111111110110000010011001;
assign LUT_1[54852] = 32'b00000000000000001000111011100011;
assign LUT_1[54853] = 32'b00000000000000000010001101011111;
assign LUT_1[54854] = 32'b00000000000000000100101001110100;
assign LUT_1[54855] = 32'b11111111111111111101111011110000;
assign LUT_1[54856] = 32'b00000000000000000000010000000001;
assign LUT_1[54857] = 32'b11111111111111111001100001111101;
assign LUT_1[54858] = 32'b11111111111111111011111110010010;
assign LUT_1[54859] = 32'b11111111111111110101010000001110;
assign LUT_1[54860] = 32'b00000000000000001000001001011000;
assign LUT_1[54861] = 32'b00000000000000000001011011010100;
assign LUT_1[54862] = 32'b00000000000000000011110111101001;
assign LUT_1[54863] = 32'b11111111111111111101001001100101;
assign LUT_1[54864] = 32'b00000000000000000010111101101110;
assign LUT_1[54865] = 32'b11111111111111111100001111101010;
assign LUT_1[54866] = 32'b11111111111111111110101011111111;
assign LUT_1[54867] = 32'b11111111111111110111111101111011;
assign LUT_1[54868] = 32'b00000000000000001010110111000101;
assign LUT_1[54869] = 32'b00000000000000000100001001000001;
assign LUT_1[54870] = 32'b00000000000000000110100101010110;
assign LUT_1[54871] = 32'b11111111111111111111110111010010;
assign LUT_1[54872] = 32'b00000000000000000010001011100011;
assign LUT_1[54873] = 32'b11111111111111111011011101011111;
assign LUT_1[54874] = 32'b11111111111111111101111001110100;
assign LUT_1[54875] = 32'b11111111111111110111001011110000;
assign LUT_1[54876] = 32'b00000000000000001010000100111010;
assign LUT_1[54877] = 32'b00000000000000000011010110110110;
assign LUT_1[54878] = 32'b00000000000000000101110011001011;
assign LUT_1[54879] = 32'b11111111111111111111000101000111;
assign LUT_1[54880] = 32'b00000000000000000001111101001011;
assign LUT_1[54881] = 32'b11111111111111111011001111000111;
assign LUT_1[54882] = 32'b11111111111111111101101011011100;
assign LUT_1[54883] = 32'b11111111111111110110111101011000;
assign LUT_1[54884] = 32'b00000000000000001001110110100010;
assign LUT_1[54885] = 32'b00000000000000000011001000011110;
assign LUT_1[54886] = 32'b00000000000000000101100100110011;
assign LUT_1[54887] = 32'b11111111111111111110110110101111;
assign LUT_1[54888] = 32'b00000000000000000001001011000000;
assign LUT_1[54889] = 32'b11111111111111111010011100111100;
assign LUT_1[54890] = 32'b11111111111111111100111001010001;
assign LUT_1[54891] = 32'b11111111111111110110001011001101;
assign LUT_1[54892] = 32'b00000000000000001001000100010111;
assign LUT_1[54893] = 32'b00000000000000000010010110010011;
assign LUT_1[54894] = 32'b00000000000000000100110010101000;
assign LUT_1[54895] = 32'b11111111111111111110000100100100;
assign LUT_1[54896] = 32'b00000000000000000011111000101101;
assign LUT_1[54897] = 32'b11111111111111111101001010101001;
assign LUT_1[54898] = 32'b11111111111111111111100110111110;
assign LUT_1[54899] = 32'b11111111111111111000111000111010;
assign LUT_1[54900] = 32'b00000000000000001011110010000100;
assign LUT_1[54901] = 32'b00000000000000000101000100000000;
assign LUT_1[54902] = 32'b00000000000000000111100000010101;
assign LUT_1[54903] = 32'b00000000000000000000110010010001;
assign LUT_1[54904] = 32'b00000000000000000011000110100010;
assign LUT_1[54905] = 32'b11111111111111111100011000011110;
assign LUT_1[54906] = 32'b11111111111111111110110100110011;
assign LUT_1[54907] = 32'b11111111111111111000000110101111;
assign LUT_1[54908] = 32'b00000000000000001010111111111001;
assign LUT_1[54909] = 32'b00000000000000000100010001110101;
assign LUT_1[54910] = 32'b00000000000000000110101110001010;
assign LUT_1[54911] = 32'b00000000000000000000000000000110;
assign LUT_1[54912] = 32'b00000000000000000010000100100111;
assign LUT_1[54913] = 32'b11111111111111111011010110100011;
assign LUT_1[54914] = 32'b11111111111111111101110010111000;
assign LUT_1[54915] = 32'b11111111111111110111000100110100;
assign LUT_1[54916] = 32'b00000000000000001001111101111110;
assign LUT_1[54917] = 32'b00000000000000000011001111111010;
assign LUT_1[54918] = 32'b00000000000000000101101100001111;
assign LUT_1[54919] = 32'b11111111111111111110111110001011;
assign LUT_1[54920] = 32'b00000000000000000001010010011100;
assign LUT_1[54921] = 32'b11111111111111111010100100011000;
assign LUT_1[54922] = 32'b11111111111111111101000000101101;
assign LUT_1[54923] = 32'b11111111111111110110010010101001;
assign LUT_1[54924] = 32'b00000000000000001001001011110011;
assign LUT_1[54925] = 32'b00000000000000000010011101101111;
assign LUT_1[54926] = 32'b00000000000000000100111010000100;
assign LUT_1[54927] = 32'b11111111111111111110001100000000;
assign LUT_1[54928] = 32'b00000000000000000100000000001001;
assign LUT_1[54929] = 32'b11111111111111111101010010000101;
assign LUT_1[54930] = 32'b11111111111111111111101110011010;
assign LUT_1[54931] = 32'b11111111111111111001000000010110;
assign LUT_1[54932] = 32'b00000000000000001011111001100000;
assign LUT_1[54933] = 32'b00000000000000000101001011011100;
assign LUT_1[54934] = 32'b00000000000000000111100111110001;
assign LUT_1[54935] = 32'b00000000000000000000111001101101;
assign LUT_1[54936] = 32'b00000000000000000011001101111110;
assign LUT_1[54937] = 32'b11111111111111111100011111111010;
assign LUT_1[54938] = 32'b11111111111111111110111100001111;
assign LUT_1[54939] = 32'b11111111111111111000001110001011;
assign LUT_1[54940] = 32'b00000000000000001011000111010101;
assign LUT_1[54941] = 32'b00000000000000000100011001010001;
assign LUT_1[54942] = 32'b00000000000000000110110101100110;
assign LUT_1[54943] = 32'b00000000000000000000000111100010;
assign LUT_1[54944] = 32'b00000000000000000010111111100110;
assign LUT_1[54945] = 32'b11111111111111111100010001100010;
assign LUT_1[54946] = 32'b11111111111111111110101101110111;
assign LUT_1[54947] = 32'b11111111111111110111111111110011;
assign LUT_1[54948] = 32'b00000000000000001010111000111101;
assign LUT_1[54949] = 32'b00000000000000000100001010111001;
assign LUT_1[54950] = 32'b00000000000000000110100111001110;
assign LUT_1[54951] = 32'b11111111111111111111111001001010;
assign LUT_1[54952] = 32'b00000000000000000010001101011011;
assign LUT_1[54953] = 32'b11111111111111111011011111010111;
assign LUT_1[54954] = 32'b11111111111111111101111011101100;
assign LUT_1[54955] = 32'b11111111111111110111001101101000;
assign LUT_1[54956] = 32'b00000000000000001010000110110010;
assign LUT_1[54957] = 32'b00000000000000000011011000101110;
assign LUT_1[54958] = 32'b00000000000000000101110101000011;
assign LUT_1[54959] = 32'b11111111111111111111000110111111;
assign LUT_1[54960] = 32'b00000000000000000100111011001000;
assign LUT_1[54961] = 32'b11111111111111111110001101000100;
assign LUT_1[54962] = 32'b00000000000000000000101001011001;
assign LUT_1[54963] = 32'b11111111111111111001111011010101;
assign LUT_1[54964] = 32'b00000000000000001100110100011111;
assign LUT_1[54965] = 32'b00000000000000000110000110011011;
assign LUT_1[54966] = 32'b00000000000000001000100010110000;
assign LUT_1[54967] = 32'b00000000000000000001110100101100;
assign LUT_1[54968] = 32'b00000000000000000100001000111101;
assign LUT_1[54969] = 32'b11111111111111111101011010111001;
assign LUT_1[54970] = 32'b11111111111111111111110111001110;
assign LUT_1[54971] = 32'b11111111111111111001001001001010;
assign LUT_1[54972] = 32'b00000000000000001100000010010100;
assign LUT_1[54973] = 32'b00000000000000000101010100010000;
assign LUT_1[54974] = 32'b00000000000000000111110000100101;
assign LUT_1[54975] = 32'b00000000000000000001000010100001;
assign LUT_1[54976] = 32'b00000000000000000100000010001111;
assign LUT_1[54977] = 32'b11111111111111111101010100001011;
assign LUT_1[54978] = 32'b11111111111111111111110000100000;
assign LUT_1[54979] = 32'b11111111111111111001000010011100;
assign LUT_1[54980] = 32'b00000000000000001011111011100110;
assign LUT_1[54981] = 32'b00000000000000000101001101100010;
assign LUT_1[54982] = 32'b00000000000000000111101001110111;
assign LUT_1[54983] = 32'b00000000000000000000111011110011;
assign LUT_1[54984] = 32'b00000000000000000011010000000100;
assign LUT_1[54985] = 32'b11111111111111111100100010000000;
assign LUT_1[54986] = 32'b11111111111111111110111110010101;
assign LUT_1[54987] = 32'b11111111111111111000010000010001;
assign LUT_1[54988] = 32'b00000000000000001011001001011011;
assign LUT_1[54989] = 32'b00000000000000000100011011010111;
assign LUT_1[54990] = 32'b00000000000000000110110111101100;
assign LUT_1[54991] = 32'b00000000000000000000001001101000;
assign LUT_1[54992] = 32'b00000000000000000101111101110001;
assign LUT_1[54993] = 32'b11111111111111111111001111101101;
assign LUT_1[54994] = 32'b00000000000000000001101100000010;
assign LUT_1[54995] = 32'b11111111111111111010111101111110;
assign LUT_1[54996] = 32'b00000000000000001101110111001000;
assign LUT_1[54997] = 32'b00000000000000000111001001000100;
assign LUT_1[54998] = 32'b00000000000000001001100101011001;
assign LUT_1[54999] = 32'b00000000000000000010110111010101;
assign LUT_1[55000] = 32'b00000000000000000101001011100110;
assign LUT_1[55001] = 32'b11111111111111111110011101100010;
assign LUT_1[55002] = 32'b00000000000000000000111001110111;
assign LUT_1[55003] = 32'b11111111111111111010001011110011;
assign LUT_1[55004] = 32'b00000000000000001101000100111101;
assign LUT_1[55005] = 32'b00000000000000000110010110111001;
assign LUT_1[55006] = 32'b00000000000000001000110011001110;
assign LUT_1[55007] = 32'b00000000000000000010000101001010;
assign LUT_1[55008] = 32'b00000000000000000100111101001110;
assign LUT_1[55009] = 32'b11111111111111111110001111001010;
assign LUT_1[55010] = 32'b00000000000000000000101011011111;
assign LUT_1[55011] = 32'b11111111111111111001111101011011;
assign LUT_1[55012] = 32'b00000000000000001100110110100101;
assign LUT_1[55013] = 32'b00000000000000000110001000100001;
assign LUT_1[55014] = 32'b00000000000000001000100100110110;
assign LUT_1[55015] = 32'b00000000000000000001110110110010;
assign LUT_1[55016] = 32'b00000000000000000100001011000011;
assign LUT_1[55017] = 32'b11111111111111111101011100111111;
assign LUT_1[55018] = 32'b11111111111111111111111001010100;
assign LUT_1[55019] = 32'b11111111111111111001001011010000;
assign LUT_1[55020] = 32'b00000000000000001100000100011010;
assign LUT_1[55021] = 32'b00000000000000000101010110010110;
assign LUT_1[55022] = 32'b00000000000000000111110010101011;
assign LUT_1[55023] = 32'b00000000000000000001000100100111;
assign LUT_1[55024] = 32'b00000000000000000110111000110000;
assign LUT_1[55025] = 32'b00000000000000000000001010101100;
assign LUT_1[55026] = 32'b00000000000000000010100111000001;
assign LUT_1[55027] = 32'b11111111111111111011111000111101;
assign LUT_1[55028] = 32'b00000000000000001110110010000111;
assign LUT_1[55029] = 32'b00000000000000001000000100000011;
assign LUT_1[55030] = 32'b00000000000000001010100000011000;
assign LUT_1[55031] = 32'b00000000000000000011110010010100;
assign LUT_1[55032] = 32'b00000000000000000110000110100101;
assign LUT_1[55033] = 32'b11111111111111111111011000100001;
assign LUT_1[55034] = 32'b00000000000000000001110100110110;
assign LUT_1[55035] = 32'b11111111111111111011000110110010;
assign LUT_1[55036] = 32'b00000000000000001101111111111100;
assign LUT_1[55037] = 32'b00000000000000000111010001111000;
assign LUT_1[55038] = 32'b00000000000000001001101110001101;
assign LUT_1[55039] = 32'b00000000000000000011000000001001;
assign LUT_1[55040] = 32'b11111111111111111100111000110000;
assign LUT_1[55041] = 32'b11111111111111110110001010101100;
assign LUT_1[55042] = 32'b11111111111111111000100111000001;
assign LUT_1[55043] = 32'b11111111111111110001111000111101;
assign LUT_1[55044] = 32'b00000000000000000100110010000111;
assign LUT_1[55045] = 32'b11111111111111111110000100000011;
assign LUT_1[55046] = 32'b00000000000000000000100000011000;
assign LUT_1[55047] = 32'b11111111111111111001110010010100;
assign LUT_1[55048] = 32'b11111111111111111100000110100101;
assign LUT_1[55049] = 32'b11111111111111110101011000100001;
assign LUT_1[55050] = 32'b11111111111111110111110100110110;
assign LUT_1[55051] = 32'b11111111111111110001000110110010;
assign LUT_1[55052] = 32'b00000000000000000011111111111100;
assign LUT_1[55053] = 32'b11111111111111111101010001111000;
assign LUT_1[55054] = 32'b11111111111111111111101110001101;
assign LUT_1[55055] = 32'b11111111111111111001000000001001;
assign LUT_1[55056] = 32'b11111111111111111110110100010010;
assign LUT_1[55057] = 32'b11111111111111111000000110001110;
assign LUT_1[55058] = 32'b11111111111111111010100010100011;
assign LUT_1[55059] = 32'b11111111111111110011110100011111;
assign LUT_1[55060] = 32'b00000000000000000110101101101001;
assign LUT_1[55061] = 32'b11111111111111111111111111100101;
assign LUT_1[55062] = 32'b00000000000000000010011011111010;
assign LUT_1[55063] = 32'b11111111111111111011101101110110;
assign LUT_1[55064] = 32'b11111111111111111110000010000111;
assign LUT_1[55065] = 32'b11111111111111110111010100000011;
assign LUT_1[55066] = 32'b11111111111111111001110000011000;
assign LUT_1[55067] = 32'b11111111111111110011000010010100;
assign LUT_1[55068] = 32'b00000000000000000101111011011110;
assign LUT_1[55069] = 32'b11111111111111111111001101011010;
assign LUT_1[55070] = 32'b00000000000000000001101001101111;
assign LUT_1[55071] = 32'b11111111111111111010111011101011;
assign LUT_1[55072] = 32'b11111111111111111101110011101111;
assign LUT_1[55073] = 32'b11111111111111110111000101101011;
assign LUT_1[55074] = 32'b11111111111111111001100010000000;
assign LUT_1[55075] = 32'b11111111111111110010110011111100;
assign LUT_1[55076] = 32'b00000000000000000101101101000110;
assign LUT_1[55077] = 32'b11111111111111111110111111000010;
assign LUT_1[55078] = 32'b00000000000000000001011011010111;
assign LUT_1[55079] = 32'b11111111111111111010101101010011;
assign LUT_1[55080] = 32'b11111111111111111101000001100100;
assign LUT_1[55081] = 32'b11111111111111110110010011100000;
assign LUT_1[55082] = 32'b11111111111111111000101111110101;
assign LUT_1[55083] = 32'b11111111111111110010000001110001;
assign LUT_1[55084] = 32'b00000000000000000100111010111011;
assign LUT_1[55085] = 32'b11111111111111111110001100110111;
assign LUT_1[55086] = 32'b00000000000000000000101001001100;
assign LUT_1[55087] = 32'b11111111111111111001111011001000;
assign LUT_1[55088] = 32'b11111111111111111111101111010001;
assign LUT_1[55089] = 32'b11111111111111111001000001001101;
assign LUT_1[55090] = 32'b11111111111111111011011101100010;
assign LUT_1[55091] = 32'b11111111111111110100101111011110;
assign LUT_1[55092] = 32'b00000000000000000111101000101000;
assign LUT_1[55093] = 32'b00000000000000000000111010100100;
assign LUT_1[55094] = 32'b00000000000000000011010110111001;
assign LUT_1[55095] = 32'b11111111111111111100101000110101;
assign LUT_1[55096] = 32'b11111111111111111110111101000110;
assign LUT_1[55097] = 32'b11111111111111111000001111000010;
assign LUT_1[55098] = 32'b11111111111111111010101011010111;
assign LUT_1[55099] = 32'b11111111111111110011111101010011;
assign LUT_1[55100] = 32'b00000000000000000110110110011101;
assign LUT_1[55101] = 32'b00000000000000000000001000011001;
assign LUT_1[55102] = 32'b00000000000000000010100100101110;
assign LUT_1[55103] = 32'b11111111111111111011110110101010;
assign LUT_1[55104] = 32'b11111111111111111110110110011000;
assign LUT_1[55105] = 32'b11111111111111111000001000010100;
assign LUT_1[55106] = 32'b11111111111111111010100100101001;
assign LUT_1[55107] = 32'b11111111111111110011110110100101;
assign LUT_1[55108] = 32'b00000000000000000110101111101111;
assign LUT_1[55109] = 32'b00000000000000000000000001101011;
assign LUT_1[55110] = 32'b00000000000000000010011110000000;
assign LUT_1[55111] = 32'b11111111111111111011101111111100;
assign LUT_1[55112] = 32'b11111111111111111110000100001101;
assign LUT_1[55113] = 32'b11111111111111110111010110001001;
assign LUT_1[55114] = 32'b11111111111111111001110010011110;
assign LUT_1[55115] = 32'b11111111111111110011000100011010;
assign LUT_1[55116] = 32'b00000000000000000101111101100100;
assign LUT_1[55117] = 32'b11111111111111111111001111100000;
assign LUT_1[55118] = 32'b00000000000000000001101011110101;
assign LUT_1[55119] = 32'b11111111111111111010111101110001;
assign LUT_1[55120] = 32'b00000000000000000000110001111010;
assign LUT_1[55121] = 32'b11111111111111111010000011110110;
assign LUT_1[55122] = 32'b11111111111111111100100000001011;
assign LUT_1[55123] = 32'b11111111111111110101110010000111;
assign LUT_1[55124] = 32'b00000000000000001000101011010001;
assign LUT_1[55125] = 32'b00000000000000000001111101001101;
assign LUT_1[55126] = 32'b00000000000000000100011001100010;
assign LUT_1[55127] = 32'b11111111111111111101101011011110;
assign LUT_1[55128] = 32'b11111111111111111111111111101111;
assign LUT_1[55129] = 32'b11111111111111111001010001101011;
assign LUT_1[55130] = 32'b11111111111111111011101110000000;
assign LUT_1[55131] = 32'b11111111111111110100111111111100;
assign LUT_1[55132] = 32'b00000000000000000111111001000110;
assign LUT_1[55133] = 32'b00000000000000000001001011000010;
assign LUT_1[55134] = 32'b00000000000000000011100111010111;
assign LUT_1[55135] = 32'b11111111111111111100111001010011;
assign LUT_1[55136] = 32'b11111111111111111111110001010111;
assign LUT_1[55137] = 32'b11111111111111111001000011010011;
assign LUT_1[55138] = 32'b11111111111111111011011111101000;
assign LUT_1[55139] = 32'b11111111111111110100110001100100;
assign LUT_1[55140] = 32'b00000000000000000111101010101110;
assign LUT_1[55141] = 32'b00000000000000000000111100101010;
assign LUT_1[55142] = 32'b00000000000000000011011000111111;
assign LUT_1[55143] = 32'b11111111111111111100101010111011;
assign LUT_1[55144] = 32'b11111111111111111110111111001100;
assign LUT_1[55145] = 32'b11111111111111111000010001001000;
assign LUT_1[55146] = 32'b11111111111111111010101101011101;
assign LUT_1[55147] = 32'b11111111111111110011111111011001;
assign LUT_1[55148] = 32'b00000000000000000110111000100011;
assign LUT_1[55149] = 32'b00000000000000000000001010011111;
assign LUT_1[55150] = 32'b00000000000000000010100110110100;
assign LUT_1[55151] = 32'b11111111111111111011111000110000;
assign LUT_1[55152] = 32'b00000000000000000001101100111001;
assign LUT_1[55153] = 32'b11111111111111111010111110110101;
assign LUT_1[55154] = 32'b11111111111111111101011011001010;
assign LUT_1[55155] = 32'b11111111111111110110101101000110;
assign LUT_1[55156] = 32'b00000000000000001001100110010000;
assign LUT_1[55157] = 32'b00000000000000000010111000001100;
assign LUT_1[55158] = 32'b00000000000000000101010100100001;
assign LUT_1[55159] = 32'b11111111111111111110100110011101;
assign LUT_1[55160] = 32'b00000000000000000000111010101110;
assign LUT_1[55161] = 32'b11111111111111111010001100101010;
assign LUT_1[55162] = 32'b11111111111111111100101000111111;
assign LUT_1[55163] = 32'b11111111111111110101111010111011;
assign LUT_1[55164] = 32'b00000000000000001000110100000101;
assign LUT_1[55165] = 32'b00000000000000000010000110000001;
assign LUT_1[55166] = 32'b00000000000000000100100010010110;
assign LUT_1[55167] = 32'b11111111111111111101110100010010;
assign LUT_1[55168] = 32'b11111111111111111111111000110011;
assign LUT_1[55169] = 32'b11111111111111111001001010101111;
assign LUT_1[55170] = 32'b11111111111111111011100111000100;
assign LUT_1[55171] = 32'b11111111111111110100111001000000;
assign LUT_1[55172] = 32'b00000000000000000111110010001010;
assign LUT_1[55173] = 32'b00000000000000000001000100000110;
assign LUT_1[55174] = 32'b00000000000000000011100000011011;
assign LUT_1[55175] = 32'b11111111111111111100110010010111;
assign LUT_1[55176] = 32'b11111111111111111111000110101000;
assign LUT_1[55177] = 32'b11111111111111111000011000100100;
assign LUT_1[55178] = 32'b11111111111111111010110100111001;
assign LUT_1[55179] = 32'b11111111111111110100000110110101;
assign LUT_1[55180] = 32'b00000000000000000110111111111111;
assign LUT_1[55181] = 32'b00000000000000000000010001111011;
assign LUT_1[55182] = 32'b00000000000000000010101110010000;
assign LUT_1[55183] = 32'b11111111111111111100000000001100;
assign LUT_1[55184] = 32'b00000000000000000001110100010101;
assign LUT_1[55185] = 32'b11111111111111111011000110010001;
assign LUT_1[55186] = 32'b11111111111111111101100010100110;
assign LUT_1[55187] = 32'b11111111111111110110110100100010;
assign LUT_1[55188] = 32'b00000000000000001001101101101100;
assign LUT_1[55189] = 32'b00000000000000000010111111101000;
assign LUT_1[55190] = 32'b00000000000000000101011011111101;
assign LUT_1[55191] = 32'b11111111111111111110101101111001;
assign LUT_1[55192] = 32'b00000000000000000001000010001010;
assign LUT_1[55193] = 32'b11111111111111111010010100000110;
assign LUT_1[55194] = 32'b11111111111111111100110000011011;
assign LUT_1[55195] = 32'b11111111111111110110000010010111;
assign LUT_1[55196] = 32'b00000000000000001000111011100001;
assign LUT_1[55197] = 32'b00000000000000000010001101011101;
assign LUT_1[55198] = 32'b00000000000000000100101001110010;
assign LUT_1[55199] = 32'b11111111111111111101111011101110;
assign LUT_1[55200] = 32'b00000000000000000000110011110010;
assign LUT_1[55201] = 32'b11111111111111111010000101101110;
assign LUT_1[55202] = 32'b11111111111111111100100010000011;
assign LUT_1[55203] = 32'b11111111111111110101110011111111;
assign LUT_1[55204] = 32'b00000000000000001000101101001001;
assign LUT_1[55205] = 32'b00000000000000000001111111000101;
assign LUT_1[55206] = 32'b00000000000000000100011011011010;
assign LUT_1[55207] = 32'b11111111111111111101101101010110;
assign LUT_1[55208] = 32'b00000000000000000000000001100111;
assign LUT_1[55209] = 32'b11111111111111111001010011100011;
assign LUT_1[55210] = 32'b11111111111111111011101111111000;
assign LUT_1[55211] = 32'b11111111111111110101000001110100;
assign LUT_1[55212] = 32'b00000000000000000111111010111110;
assign LUT_1[55213] = 32'b00000000000000000001001100111010;
assign LUT_1[55214] = 32'b00000000000000000011101001001111;
assign LUT_1[55215] = 32'b11111111111111111100111011001011;
assign LUT_1[55216] = 32'b00000000000000000010101111010100;
assign LUT_1[55217] = 32'b11111111111111111100000001010000;
assign LUT_1[55218] = 32'b11111111111111111110011101100101;
assign LUT_1[55219] = 32'b11111111111111110111101111100001;
assign LUT_1[55220] = 32'b00000000000000001010101000101011;
assign LUT_1[55221] = 32'b00000000000000000011111010100111;
assign LUT_1[55222] = 32'b00000000000000000110010110111100;
assign LUT_1[55223] = 32'b11111111111111111111101000111000;
assign LUT_1[55224] = 32'b00000000000000000001111101001001;
assign LUT_1[55225] = 32'b11111111111111111011001111000101;
assign LUT_1[55226] = 32'b11111111111111111101101011011010;
assign LUT_1[55227] = 32'b11111111111111110110111101010110;
assign LUT_1[55228] = 32'b00000000000000001001110110100000;
assign LUT_1[55229] = 32'b00000000000000000011001000011100;
assign LUT_1[55230] = 32'b00000000000000000101100100110001;
assign LUT_1[55231] = 32'b11111111111111111110110110101101;
assign LUT_1[55232] = 32'b00000000000000000001110110011011;
assign LUT_1[55233] = 32'b11111111111111111011001000010111;
assign LUT_1[55234] = 32'b11111111111111111101100100101100;
assign LUT_1[55235] = 32'b11111111111111110110110110101000;
assign LUT_1[55236] = 32'b00000000000000001001101111110010;
assign LUT_1[55237] = 32'b00000000000000000011000001101110;
assign LUT_1[55238] = 32'b00000000000000000101011110000011;
assign LUT_1[55239] = 32'b11111111111111111110101111111111;
assign LUT_1[55240] = 32'b00000000000000000001000100010000;
assign LUT_1[55241] = 32'b11111111111111111010010110001100;
assign LUT_1[55242] = 32'b11111111111111111100110010100001;
assign LUT_1[55243] = 32'b11111111111111110110000100011101;
assign LUT_1[55244] = 32'b00000000000000001000111101100111;
assign LUT_1[55245] = 32'b00000000000000000010001111100011;
assign LUT_1[55246] = 32'b00000000000000000100101011111000;
assign LUT_1[55247] = 32'b11111111111111111101111101110100;
assign LUT_1[55248] = 32'b00000000000000000011110001111101;
assign LUT_1[55249] = 32'b11111111111111111101000011111001;
assign LUT_1[55250] = 32'b11111111111111111111100000001110;
assign LUT_1[55251] = 32'b11111111111111111000110010001010;
assign LUT_1[55252] = 32'b00000000000000001011101011010100;
assign LUT_1[55253] = 32'b00000000000000000100111101010000;
assign LUT_1[55254] = 32'b00000000000000000111011001100101;
assign LUT_1[55255] = 32'b00000000000000000000101011100001;
assign LUT_1[55256] = 32'b00000000000000000010111111110010;
assign LUT_1[55257] = 32'b11111111111111111100010001101110;
assign LUT_1[55258] = 32'b11111111111111111110101110000011;
assign LUT_1[55259] = 32'b11111111111111110111111111111111;
assign LUT_1[55260] = 32'b00000000000000001010111001001001;
assign LUT_1[55261] = 32'b00000000000000000100001011000101;
assign LUT_1[55262] = 32'b00000000000000000110100111011010;
assign LUT_1[55263] = 32'b11111111111111111111111001010110;
assign LUT_1[55264] = 32'b00000000000000000010110001011010;
assign LUT_1[55265] = 32'b11111111111111111100000011010110;
assign LUT_1[55266] = 32'b11111111111111111110011111101011;
assign LUT_1[55267] = 32'b11111111111111110111110001100111;
assign LUT_1[55268] = 32'b00000000000000001010101010110001;
assign LUT_1[55269] = 32'b00000000000000000011111100101101;
assign LUT_1[55270] = 32'b00000000000000000110011001000010;
assign LUT_1[55271] = 32'b11111111111111111111101010111110;
assign LUT_1[55272] = 32'b00000000000000000001111111001111;
assign LUT_1[55273] = 32'b11111111111111111011010001001011;
assign LUT_1[55274] = 32'b11111111111111111101101101100000;
assign LUT_1[55275] = 32'b11111111111111110110111111011100;
assign LUT_1[55276] = 32'b00000000000000001001111000100110;
assign LUT_1[55277] = 32'b00000000000000000011001010100010;
assign LUT_1[55278] = 32'b00000000000000000101100110110111;
assign LUT_1[55279] = 32'b11111111111111111110111000110011;
assign LUT_1[55280] = 32'b00000000000000000100101100111100;
assign LUT_1[55281] = 32'b11111111111111111101111110111000;
assign LUT_1[55282] = 32'b00000000000000000000011011001101;
assign LUT_1[55283] = 32'b11111111111111111001101101001001;
assign LUT_1[55284] = 32'b00000000000000001100100110010011;
assign LUT_1[55285] = 32'b00000000000000000101111000001111;
assign LUT_1[55286] = 32'b00000000000000001000010100100100;
assign LUT_1[55287] = 32'b00000000000000000001100110100000;
assign LUT_1[55288] = 32'b00000000000000000011111010110001;
assign LUT_1[55289] = 32'b11111111111111111101001100101101;
assign LUT_1[55290] = 32'b11111111111111111111101001000010;
assign LUT_1[55291] = 32'b11111111111111111000111010111110;
assign LUT_1[55292] = 32'b00000000000000001011110100001000;
assign LUT_1[55293] = 32'b00000000000000000101000110000100;
assign LUT_1[55294] = 32'b00000000000000000111100010011001;
assign LUT_1[55295] = 32'b00000000000000000000110100010101;
assign LUT_1[55296] = 32'b00000000000000000000000001010010;
assign LUT_1[55297] = 32'b11111111111111111001010011001110;
assign LUT_1[55298] = 32'b11111111111111111011101111100011;
assign LUT_1[55299] = 32'b11111111111111110101000001011111;
assign LUT_1[55300] = 32'b00000000000000000111111010101001;
assign LUT_1[55301] = 32'b00000000000000000001001100100101;
assign LUT_1[55302] = 32'b00000000000000000011101000111010;
assign LUT_1[55303] = 32'b11111111111111111100111010110110;
assign LUT_1[55304] = 32'b11111111111111111111001111000111;
assign LUT_1[55305] = 32'b11111111111111111000100001000011;
assign LUT_1[55306] = 32'b11111111111111111010111101011000;
assign LUT_1[55307] = 32'b11111111111111110100001111010100;
assign LUT_1[55308] = 32'b00000000000000000111001000011110;
assign LUT_1[55309] = 32'b00000000000000000000011010011010;
assign LUT_1[55310] = 32'b00000000000000000010110110101111;
assign LUT_1[55311] = 32'b11111111111111111100001000101011;
assign LUT_1[55312] = 32'b00000000000000000001111100110100;
assign LUT_1[55313] = 32'b11111111111111111011001110110000;
assign LUT_1[55314] = 32'b11111111111111111101101011000101;
assign LUT_1[55315] = 32'b11111111111111110110111101000001;
assign LUT_1[55316] = 32'b00000000000000001001110110001011;
assign LUT_1[55317] = 32'b00000000000000000011001000000111;
assign LUT_1[55318] = 32'b00000000000000000101100100011100;
assign LUT_1[55319] = 32'b11111111111111111110110110011000;
assign LUT_1[55320] = 32'b00000000000000000001001010101001;
assign LUT_1[55321] = 32'b11111111111111111010011100100101;
assign LUT_1[55322] = 32'b11111111111111111100111000111010;
assign LUT_1[55323] = 32'b11111111111111110110001010110110;
assign LUT_1[55324] = 32'b00000000000000001001000100000000;
assign LUT_1[55325] = 32'b00000000000000000010010101111100;
assign LUT_1[55326] = 32'b00000000000000000100110010010001;
assign LUT_1[55327] = 32'b11111111111111111110000100001101;
assign LUT_1[55328] = 32'b00000000000000000000111100010001;
assign LUT_1[55329] = 32'b11111111111111111010001110001101;
assign LUT_1[55330] = 32'b11111111111111111100101010100010;
assign LUT_1[55331] = 32'b11111111111111110101111100011110;
assign LUT_1[55332] = 32'b00000000000000001000110101101000;
assign LUT_1[55333] = 32'b00000000000000000010000111100100;
assign LUT_1[55334] = 32'b00000000000000000100100011111001;
assign LUT_1[55335] = 32'b11111111111111111101110101110101;
assign LUT_1[55336] = 32'b00000000000000000000001010000110;
assign LUT_1[55337] = 32'b11111111111111111001011100000010;
assign LUT_1[55338] = 32'b11111111111111111011111000010111;
assign LUT_1[55339] = 32'b11111111111111110101001010010011;
assign LUT_1[55340] = 32'b00000000000000001000000011011101;
assign LUT_1[55341] = 32'b00000000000000000001010101011001;
assign LUT_1[55342] = 32'b00000000000000000011110001101110;
assign LUT_1[55343] = 32'b11111111111111111101000011101010;
assign LUT_1[55344] = 32'b00000000000000000010110111110011;
assign LUT_1[55345] = 32'b11111111111111111100001001101111;
assign LUT_1[55346] = 32'b11111111111111111110100110000100;
assign LUT_1[55347] = 32'b11111111111111110111111000000000;
assign LUT_1[55348] = 32'b00000000000000001010110001001010;
assign LUT_1[55349] = 32'b00000000000000000100000011000110;
assign LUT_1[55350] = 32'b00000000000000000110011111011011;
assign LUT_1[55351] = 32'b11111111111111111111110001010111;
assign LUT_1[55352] = 32'b00000000000000000010000101101000;
assign LUT_1[55353] = 32'b11111111111111111011010111100100;
assign LUT_1[55354] = 32'b11111111111111111101110011111001;
assign LUT_1[55355] = 32'b11111111111111110111000101110101;
assign LUT_1[55356] = 32'b00000000000000001001111110111111;
assign LUT_1[55357] = 32'b00000000000000000011010000111011;
assign LUT_1[55358] = 32'b00000000000000000101101101010000;
assign LUT_1[55359] = 32'b11111111111111111110111111001100;
assign LUT_1[55360] = 32'b00000000000000000001111110111010;
assign LUT_1[55361] = 32'b11111111111111111011010000110110;
assign LUT_1[55362] = 32'b11111111111111111101101101001011;
assign LUT_1[55363] = 32'b11111111111111110110111111000111;
assign LUT_1[55364] = 32'b00000000000000001001111000010001;
assign LUT_1[55365] = 32'b00000000000000000011001010001101;
assign LUT_1[55366] = 32'b00000000000000000101100110100010;
assign LUT_1[55367] = 32'b11111111111111111110111000011110;
assign LUT_1[55368] = 32'b00000000000000000001001100101111;
assign LUT_1[55369] = 32'b11111111111111111010011110101011;
assign LUT_1[55370] = 32'b11111111111111111100111011000000;
assign LUT_1[55371] = 32'b11111111111111110110001100111100;
assign LUT_1[55372] = 32'b00000000000000001001000110000110;
assign LUT_1[55373] = 32'b00000000000000000010011000000010;
assign LUT_1[55374] = 32'b00000000000000000100110100010111;
assign LUT_1[55375] = 32'b11111111111111111110000110010011;
assign LUT_1[55376] = 32'b00000000000000000011111010011100;
assign LUT_1[55377] = 32'b11111111111111111101001100011000;
assign LUT_1[55378] = 32'b11111111111111111111101000101101;
assign LUT_1[55379] = 32'b11111111111111111000111010101001;
assign LUT_1[55380] = 32'b00000000000000001011110011110011;
assign LUT_1[55381] = 32'b00000000000000000101000101101111;
assign LUT_1[55382] = 32'b00000000000000000111100010000100;
assign LUT_1[55383] = 32'b00000000000000000000110100000000;
assign LUT_1[55384] = 32'b00000000000000000011001000010001;
assign LUT_1[55385] = 32'b11111111111111111100011010001101;
assign LUT_1[55386] = 32'b11111111111111111110110110100010;
assign LUT_1[55387] = 32'b11111111111111111000001000011110;
assign LUT_1[55388] = 32'b00000000000000001011000001101000;
assign LUT_1[55389] = 32'b00000000000000000100010011100100;
assign LUT_1[55390] = 32'b00000000000000000110101111111001;
assign LUT_1[55391] = 32'b00000000000000000000000001110101;
assign LUT_1[55392] = 32'b00000000000000000010111001111001;
assign LUT_1[55393] = 32'b11111111111111111100001011110101;
assign LUT_1[55394] = 32'b11111111111111111110101000001010;
assign LUT_1[55395] = 32'b11111111111111110111111010000110;
assign LUT_1[55396] = 32'b00000000000000001010110011010000;
assign LUT_1[55397] = 32'b00000000000000000100000101001100;
assign LUT_1[55398] = 32'b00000000000000000110100001100001;
assign LUT_1[55399] = 32'b11111111111111111111110011011101;
assign LUT_1[55400] = 32'b00000000000000000010000111101110;
assign LUT_1[55401] = 32'b11111111111111111011011001101010;
assign LUT_1[55402] = 32'b11111111111111111101110101111111;
assign LUT_1[55403] = 32'b11111111111111110111000111111011;
assign LUT_1[55404] = 32'b00000000000000001010000001000101;
assign LUT_1[55405] = 32'b00000000000000000011010011000001;
assign LUT_1[55406] = 32'b00000000000000000101101111010110;
assign LUT_1[55407] = 32'b11111111111111111111000001010010;
assign LUT_1[55408] = 32'b00000000000000000100110101011011;
assign LUT_1[55409] = 32'b11111111111111111110000111010111;
assign LUT_1[55410] = 32'b00000000000000000000100011101100;
assign LUT_1[55411] = 32'b11111111111111111001110101101000;
assign LUT_1[55412] = 32'b00000000000000001100101110110010;
assign LUT_1[55413] = 32'b00000000000000000110000000101110;
assign LUT_1[55414] = 32'b00000000000000001000011101000011;
assign LUT_1[55415] = 32'b00000000000000000001101110111111;
assign LUT_1[55416] = 32'b00000000000000000100000011010000;
assign LUT_1[55417] = 32'b11111111111111111101010101001100;
assign LUT_1[55418] = 32'b11111111111111111111110001100001;
assign LUT_1[55419] = 32'b11111111111111111001000011011101;
assign LUT_1[55420] = 32'b00000000000000001011111100100111;
assign LUT_1[55421] = 32'b00000000000000000101001110100011;
assign LUT_1[55422] = 32'b00000000000000000111101010111000;
assign LUT_1[55423] = 32'b00000000000000000000111100110100;
assign LUT_1[55424] = 32'b00000000000000000011000001010101;
assign LUT_1[55425] = 32'b11111111111111111100010011010001;
assign LUT_1[55426] = 32'b11111111111111111110101111100110;
assign LUT_1[55427] = 32'b11111111111111111000000001100010;
assign LUT_1[55428] = 32'b00000000000000001010111010101100;
assign LUT_1[55429] = 32'b00000000000000000100001100101000;
assign LUT_1[55430] = 32'b00000000000000000110101000111101;
assign LUT_1[55431] = 32'b11111111111111111111111010111001;
assign LUT_1[55432] = 32'b00000000000000000010001111001010;
assign LUT_1[55433] = 32'b11111111111111111011100001000110;
assign LUT_1[55434] = 32'b11111111111111111101111101011011;
assign LUT_1[55435] = 32'b11111111111111110111001111010111;
assign LUT_1[55436] = 32'b00000000000000001010001000100001;
assign LUT_1[55437] = 32'b00000000000000000011011010011101;
assign LUT_1[55438] = 32'b00000000000000000101110110110010;
assign LUT_1[55439] = 32'b11111111111111111111001000101110;
assign LUT_1[55440] = 32'b00000000000000000100111100110111;
assign LUT_1[55441] = 32'b11111111111111111110001110110011;
assign LUT_1[55442] = 32'b00000000000000000000101011001000;
assign LUT_1[55443] = 32'b11111111111111111001111101000100;
assign LUT_1[55444] = 32'b00000000000000001100110110001110;
assign LUT_1[55445] = 32'b00000000000000000110001000001010;
assign LUT_1[55446] = 32'b00000000000000001000100100011111;
assign LUT_1[55447] = 32'b00000000000000000001110110011011;
assign LUT_1[55448] = 32'b00000000000000000100001010101100;
assign LUT_1[55449] = 32'b11111111111111111101011100101000;
assign LUT_1[55450] = 32'b11111111111111111111111000111101;
assign LUT_1[55451] = 32'b11111111111111111001001010111001;
assign LUT_1[55452] = 32'b00000000000000001100000100000011;
assign LUT_1[55453] = 32'b00000000000000000101010101111111;
assign LUT_1[55454] = 32'b00000000000000000111110010010100;
assign LUT_1[55455] = 32'b00000000000000000001000100010000;
assign LUT_1[55456] = 32'b00000000000000000011111100010100;
assign LUT_1[55457] = 32'b11111111111111111101001110010000;
assign LUT_1[55458] = 32'b11111111111111111111101010100101;
assign LUT_1[55459] = 32'b11111111111111111000111100100001;
assign LUT_1[55460] = 32'b00000000000000001011110101101011;
assign LUT_1[55461] = 32'b00000000000000000101000111100111;
assign LUT_1[55462] = 32'b00000000000000000111100011111100;
assign LUT_1[55463] = 32'b00000000000000000000110101111000;
assign LUT_1[55464] = 32'b00000000000000000011001010001001;
assign LUT_1[55465] = 32'b11111111111111111100011100000101;
assign LUT_1[55466] = 32'b11111111111111111110111000011010;
assign LUT_1[55467] = 32'b11111111111111111000001010010110;
assign LUT_1[55468] = 32'b00000000000000001011000011100000;
assign LUT_1[55469] = 32'b00000000000000000100010101011100;
assign LUT_1[55470] = 32'b00000000000000000110110001110001;
assign LUT_1[55471] = 32'b00000000000000000000000011101101;
assign LUT_1[55472] = 32'b00000000000000000101110111110110;
assign LUT_1[55473] = 32'b11111111111111111111001001110010;
assign LUT_1[55474] = 32'b00000000000000000001100110000111;
assign LUT_1[55475] = 32'b11111111111111111010111000000011;
assign LUT_1[55476] = 32'b00000000000000001101110001001101;
assign LUT_1[55477] = 32'b00000000000000000111000011001001;
assign LUT_1[55478] = 32'b00000000000000001001011111011110;
assign LUT_1[55479] = 32'b00000000000000000010110001011010;
assign LUT_1[55480] = 32'b00000000000000000101000101101011;
assign LUT_1[55481] = 32'b11111111111111111110010111100111;
assign LUT_1[55482] = 32'b00000000000000000000110011111100;
assign LUT_1[55483] = 32'b11111111111111111010000101111000;
assign LUT_1[55484] = 32'b00000000000000001100111111000010;
assign LUT_1[55485] = 32'b00000000000000000110010000111110;
assign LUT_1[55486] = 32'b00000000000000001000101101010011;
assign LUT_1[55487] = 32'b00000000000000000001111111001111;
assign LUT_1[55488] = 32'b00000000000000000100111110111101;
assign LUT_1[55489] = 32'b11111111111111111110010000111001;
assign LUT_1[55490] = 32'b00000000000000000000101101001110;
assign LUT_1[55491] = 32'b11111111111111111001111111001010;
assign LUT_1[55492] = 32'b00000000000000001100111000010100;
assign LUT_1[55493] = 32'b00000000000000000110001010010000;
assign LUT_1[55494] = 32'b00000000000000001000100110100101;
assign LUT_1[55495] = 32'b00000000000000000001111000100001;
assign LUT_1[55496] = 32'b00000000000000000100001100110010;
assign LUT_1[55497] = 32'b11111111111111111101011110101110;
assign LUT_1[55498] = 32'b11111111111111111111111011000011;
assign LUT_1[55499] = 32'b11111111111111111001001100111111;
assign LUT_1[55500] = 32'b00000000000000001100000110001001;
assign LUT_1[55501] = 32'b00000000000000000101011000000101;
assign LUT_1[55502] = 32'b00000000000000000111110100011010;
assign LUT_1[55503] = 32'b00000000000000000001000110010110;
assign LUT_1[55504] = 32'b00000000000000000110111010011111;
assign LUT_1[55505] = 32'b00000000000000000000001100011011;
assign LUT_1[55506] = 32'b00000000000000000010101000110000;
assign LUT_1[55507] = 32'b11111111111111111011111010101100;
assign LUT_1[55508] = 32'b00000000000000001110110011110110;
assign LUT_1[55509] = 32'b00000000000000001000000101110010;
assign LUT_1[55510] = 32'b00000000000000001010100010000111;
assign LUT_1[55511] = 32'b00000000000000000011110100000011;
assign LUT_1[55512] = 32'b00000000000000000110001000010100;
assign LUT_1[55513] = 32'b11111111111111111111011010010000;
assign LUT_1[55514] = 32'b00000000000000000001110110100101;
assign LUT_1[55515] = 32'b11111111111111111011001000100001;
assign LUT_1[55516] = 32'b00000000000000001110000001101011;
assign LUT_1[55517] = 32'b00000000000000000111010011100111;
assign LUT_1[55518] = 32'b00000000000000001001101111111100;
assign LUT_1[55519] = 32'b00000000000000000011000001111000;
assign LUT_1[55520] = 32'b00000000000000000101111001111100;
assign LUT_1[55521] = 32'b11111111111111111111001011111000;
assign LUT_1[55522] = 32'b00000000000000000001101000001101;
assign LUT_1[55523] = 32'b11111111111111111010111010001001;
assign LUT_1[55524] = 32'b00000000000000001101110011010011;
assign LUT_1[55525] = 32'b00000000000000000111000101001111;
assign LUT_1[55526] = 32'b00000000000000001001100001100100;
assign LUT_1[55527] = 32'b00000000000000000010110011100000;
assign LUT_1[55528] = 32'b00000000000000000101000111110001;
assign LUT_1[55529] = 32'b11111111111111111110011001101101;
assign LUT_1[55530] = 32'b00000000000000000000110110000010;
assign LUT_1[55531] = 32'b11111111111111111010000111111110;
assign LUT_1[55532] = 32'b00000000000000001101000001001000;
assign LUT_1[55533] = 32'b00000000000000000110010011000100;
assign LUT_1[55534] = 32'b00000000000000001000101111011001;
assign LUT_1[55535] = 32'b00000000000000000010000001010101;
assign LUT_1[55536] = 32'b00000000000000000111110101011110;
assign LUT_1[55537] = 32'b00000000000000000001000111011010;
assign LUT_1[55538] = 32'b00000000000000000011100011101111;
assign LUT_1[55539] = 32'b11111111111111111100110101101011;
assign LUT_1[55540] = 32'b00000000000000001111101110110101;
assign LUT_1[55541] = 32'b00000000000000001001000000110001;
assign LUT_1[55542] = 32'b00000000000000001011011101000110;
assign LUT_1[55543] = 32'b00000000000000000100101111000010;
assign LUT_1[55544] = 32'b00000000000000000111000011010011;
assign LUT_1[55545] = 32'b00000000000000000000010101001111;
assign LUT_1[55546] = 32'b00000000000000000010110001100100;
assign LUT_1[55547] = 32'b11111111111111111100000011100000;
assign LUT_1[55548] = 32'b00000000000000001110111100101010;
assign LUT_1[55549] = 32'b00000000000000001000001110100110;
assign LUT_1[55550] = 32'b00000000000000001010101010111011;
assign LUT_1[55551] = 32'b00000000000000000011111100110111;
assign LUT_1[55552] = 32'b11111111111111111101110101011110;
assign LUT_1[55553] = 32'b11111111111111110111000111011010;
assign LUT_1[55554] = 32'b11111111111111111001100011101111;
assign LUT_1[55555] = 32'b11111111111111110010110101101011;
assign LUT_1[55556] = 32'b00000000000000000101101110110101;
assign LUT_1[55557] = 32'b11111111111111111111000000110001;
assign LUT_1[55558] = 32'b00000000000000000001011101000110;
assign LUT_1[55559] = 32'b11111111111111111010101111000010;
assign LUT_1[55560] = 32'b11111111111111111101000011010011;
assign LUT_1[55561] = 32'b11111111111111110110010101001111;
assign LUT_1[55562] = 32'b11111111111111111000110001100100;
assign LUT_1[55563] = 32'b11111111111111110010000011100000;
assign LUT_1[55564] = 32'b00000000000000000100111100101010;
assign LUT_1[55565] = 32'b11111111111111111110001110100110;
assign LUT_1[55566] = 32'b00000000000000000000101010111011;
assign LUT_1[55567] = 32'b11111111111111111001111100110111;
assign LUT_1[55568] = 32'b11111111111111111111110001000000;
assign LUT_1[55569] = 32'b11111111111111111001000010111100;
assign LUT_1[55570] = 32'b11111111111111111011011111010001;
assign LUT_1[55571] = 32'b11111111111111110100110001001101;
assign LUT_1[55572] = 32'b00000000000000000111101010010111;
assign LUT_1[55573] = 32'b00000000000000000000111100010011;
assign LUT_1[55574] = 32'b00000000000000000011011000101000;
assign LUT_1[55575] = 32'b11111111111111111100101010100100;
assign LUT_1[55576] = 32'b11111111111111111110111110110101;
assign LUT_1[55577] = 32'b11111111111111111000010000110001;
assign LUT_1[55578] = 32'b11111111111111111010101101000110;
assign LUT_1[55579] = 32'b11111111111111110011111111000010;
assign LUT_1[55580] = 32'b00000000000000000110111000001100;
assign LUT_1[55581] = 32'b00000000000000000000001010001000;
assign LUT_1[55582] = 32'b00000000000000000010100110011101;
assign LUT_1[55583] = 32'b11111111111111111011111000011001;
assign LUT_1[55584] = 32'b11111111111111111110110000011101;
assign LUT_1[55585] = 32'b11111111111111111000000010011001;
assign LUT_1[55586] = 32'b11111111111111111010011110101110;
assign LUT_1[55587] = 32'b11111111111111110011110000101010;
assign LUT_1[55588] = 32'b00000000000000000110101001110100;
assign LUT_1[55589] = 32'b11111111111111111111111011110000;
assign LUT_1[55590] = 32'b00000000000000000010011000000101;
assign LUT_1[55591] = 32'b11111111111111111011101010000001;
assign LUT_1[55592] = 32'b11111111111111111101111110010010;
assign LUT_1[55593] = 32'b11111111111111110111010000001110;
assign LUT_1[55594] = 32'b11111111111111111001101100100011;
assign LUT_1[55595] = 32'b11111111111111110010111110011111;
assign LUT_1[55596] = 32'b00000000000000000101110111101001;
assign LUT_1[55597] = 32'b11111111111111111111001001100101;
assign LUT_1[55598] = 32'b00000000000000000001100101111010;
assign LUT_1[55599] = 32'b11111111111111111010110111110110;
assign LUT_1[55600] = 32'b00000000000000000000101011111111;
assign LUT_1[55601] = 32'b11111111111111111001111101111011;
assign LUT_1[55602] = 32'b11111111111111111100011010010000;
assign LUT_1[55603] = 32'b11111111111111110101101100001100;
assign LUT_1[55604] = 32'b00000000000000001000100101010110;
assign LUT_1[55605] = 32'b00000000000000000001110111010010;
assign LUT_1[55606] = 32'b00000000000000000100010011100111;
assign LUT_1[55607] = 32'b11111111111111111101100101100011;
assign LUT_1[55608] = 32'b11111111111111111111111001110100;
assign LUT_1[55609] = 32'b11111111111111111001001011110000;
assign LUT_1[55610] = 32'b11111111111111111011101000000101;
assign LUT_1[55611] = 32'b11111111111111110100111010000001;
assign LUT_1[55612] = 32'b00000000000000000111110011001011;
assign LUT_1[55613] = 32'b00000000000000000001000101000111;
assign LUT_1[55614] = 32'b00000000000000000011100001011100;
assign LUT_1[55615] = 32'b11111111111111111100110011011000;
assign LUT_1[55616] = 32'b11111111111111111111110011000110;
assign LUT_1[55617] = 32'b11111111111111111001000101000010;
assign LUT_1[55618] = 32'b11111111111111111011100001010111;
assign LUT_1[55619] = 32'b11111111111111110100110011010011;
assign LUT_1[55620] = 32'b00000000000000000111101100011101;
assign LUT_1[55621] = 32'b00000000000000000000111110011001;
assign LUT_1[55622] = 32'b00000000000000000011011010101110;
assign LUT_1[55623] = 32'b11111111111111111100101100101010;
assign LUT_1[55624] = 32'b11111111111111111111000000111011;
assign LUT_1[55625] = 32'b11111111111111111000010010110111;
assign LUT_1[55626] = 32'b11111111111111111010101111001100;
assign LUT_1[55627] = 32'b11111111111111110100000001001000;
assign LUT_1[55628] = 32'b00000000000000000110111010010010;
assign LUT_1[55629] = 32'b00000000000000000000001100001110;
assign LUT_1[55630] = 32'b00000000000000000010101000100011;
assign LUT_1[55631] = 32'b11111111111111111011111010011111;
assign LUT_1[55632] = 32'b00000000000000000001101110101000;
assign LUT_1[55633] = 32'b11111111111111111011000000100100;
assign LUT_1[55634] = 32'b11111111111111111101011100111001;
assign LUT_1[55635] = 32'b11111111111111110110101110110101;
assign LUT_1[55636] = 32'b00000000000000001001100111111111;
assign LUT_1[55637] = 32'b00000000000000000010111001111011;
assign LUT_1[55638] = 32'b00000000000000000101010110010000;
assign LUT_1[55639] = 32'b11111111111111111110101000001100;
assign LUT_1[55640] = 32'b00000000000000000000111100011101;
assign LUT_1[55641] = 32'b11111111111111111010001110011001;
assign LUT_1[55642] = 32'b11111111111111111100101010101110;
assign LUT_1[55643] = 32'b11111111111111110101111100101010;
assign LUT_1[55644] = 32'b00000000000000001000110101110100;
assign LUT_1[55645] = 32'b00000000000000000010000111110000;
assign LUT_1[55646] = 32'b00000000000000000100100100000101;
assign LUT_1[55647] = 32'b11111111111111111101110110000001;
assign LUT_1[55648] = 32'b00000000000000000000101110000101;
assign LUT_1[55649] = 32'b11111111111111111010000000000001;
assign LUT_1[55650] = 32'b11111111111111111100011100010110;
assign LUT_1[55651] = 32'b11111111111111110101101110010010;
assign LUT_1[55652] = 32'b00000000000000001000100111011100;
assign LUT_1[55653] = 32'b00000000000000000001111001011000;
assign LUT_1[55654] = 32'b00000000000000000100010101101101;
assign LUT_1[55655] = 32'b11111111111111111101100111101001;
assign LUT_1[55656] = 32'b11111111111111111111111011111010;
assign LUT_1[55657] = 32'b11111111111111111001001101110110;
assign LUT_1[55658] = 32'b11111111111111111011101010001011;
assign LUT_1[55659] = 32'b11111111111111110100111100000111;
assign LUT_1[55660] = 32'b00000000000000000111110101010001;
assign LUT_1[55661] = 32'b00000000000000000001000111001101;
assign LUT_1[55662] = 32'b00000000000000000011100011100010;
assign LUT_1[55663] = 32'b11111111111111111100110101011110;
assign LUT_1[55664] = 32'b00000000000000000010101001100111;
assign LUT_1[55665] = 32'b11111111111111111011111011100011;
assign LUT_1[55666] = 32'b11111111111111111110010111111000;
assign LUT_1[55667] = 32'b11111111111111110111101001110100;
assign LUT_1[55668] = 32'b00000000000000001010100010111110;
assign LUT_1[55669] = 32'b00000000000000000011110100111010;
assign LUT_1[55670] = 32'b00000000000000000110010001001111;
assign LUT_1[55671] = 32'b11111111111111111111100011001011;
assign LUT_1[55672] = 32'b00000000000000000001110111011100;
assign LUT_1[55673] = 32'b11111111111111111011001001011000;
assign LUT_1[55674] = 32'b11111111111111111101100101101101;
assign LUT_1[55675] = 32'b11111111111111110110110111101001;
assign LUT_1[55676] = 32'b00000000000000001001110000110011;
assign LUT_1[55677] = 32'b00000000000000000011000010101111;
assign LUT_1[55678] = 32'b00000000000000000101011111000100;
assign LUT_1[55679] = 32'b11111111111111111110110001000000;
assign LUT_1[55680] = 32'b00000000000000000000110101100001;
assign LUT_1[55681] = 32'b11111111111111111010000111011101;
assign LUT_1[55682] = 32'b11111111111111111100100011110010;
assign LUT_1[55683] = 32'b11111111111111110101110101101110;
assign LUT_1[55684] = 32'b00000000000000001000101110111000;
assign LUT_1[55685] = 32'b00000000000000000010000000110100;
assign LUT_1[55686] = 32'b00000000000000000100011101001001;
assign LUT_1[55687] = 32'b11111111111111111101101111000101;
assign LUT_1[55688] = 32'b00000000000000000000000011010110;
assign LUT_1[55689] = 32'b11111111111111111001010101010010;
assign LUT_1[55690] = 32'b11111111111111111011110001100111;
assign LUT_1[55691] = 32'b11111111111111110101000011100011;
assign LUT_1[55692] = 32'b00000000000000000111111100101101;
assign LUT_1[55693] = 32'b00000000000000000001001110101001;
assign LUT_1[55694] = 32'b00000000000000000011101010111110;
assign LUT_1[55695] = 32'b11111111111111111100111100111010;
assign LUT_1[55696] = 32'b00000000000000000010110001000011;
assign LUT_1[55697] = 32'b11111111111111111100000010111111;
assign LUT_1[55698] = 32'b11111111111111111110011111010100;
assign LUT_1[55699] = 32'b11111111111111110111110001010000;
assign LUT_1[55700] = 32'b00000000000000001010101010011010;
assign LUT_1[55701] = 32'b00000000000000000011111100010110;
assign LUT_1[55702] = 32'b00000000000000000110011000101011;
assign LUT_1[55703] = 32'b11111111111111111111101010100111;
assign LUT_1[55704] = 32'b00000000000000000001111110111000;
assign LUT_1[55705] = 32'b11111111111111111011010000110100;
assign LUT_1[55706] = 32'b11111111111111111101101101001001;
assign LUT_1[55707] = 32'b11111111111111110110111111000101;
assign LUT_1[55708] = 32'b00000000000000001001111000001111;
assign LUT_1[55709] = 32'b00000000000000000011001010001011;
assign LUT_1[55710] = 32'b00000000000000000101100110100000;
assign LUT_1[55711] = 32'b11111111111111111110111000011100;
assign LUT_1[55712] = 32'b00000000000000000001110000100000;
assign LUT_1[55713] = 32'b11111111111111111011000010011100;
assign LUT_1[55714] = 32'b11111111111111111101011110110001;
assign LUT_1[55715] = 32'b11111111111111110110110000101101;
assign LUT_1[55716] = 32'b00000000000000001001101001110111;
assign LUT_1[55717] = 32'b00000000000000000010111011110011;
assign LUT_1[55718] = 32'b00000000000000000101011000001000;
assign LUT_1[55719] = 32'b11111111111111111110101010000100;
assign LUT_1[55720] = 32'b00000000000000000000111110010101;
assign LUT_1[55721] = 32'b11111111111111111010010000010001;
assign LUT_1[55722] = 32'b11111111111111111100101100100110;
assign LUT_1[55723] = 32'b11111111111111110101111110100010;
assign LUT_1[55724] = 32'b00000000000000001000110111101100;
assign LUT_1[55725] = 32'b00000000000000000010001001101000;
assign LUT_1[55726] = 32'b00000000000000000100100101111101;
assign LUT_1[55727] = 32'b11111111111111111101110111111001;
assign LUT_1[55728] = 32'b00000000000000000011101100000010;
assign LUT_1[55729] = 32'b11111111111111111100111101111110;
assign LUT_1[55730] = 32'b11111111111111111111011010010011;
assign LUT_1[55731] = 32'b11111111111111111000101100001111;
assign LUT_1[55732] = 32'b00000000000000001011100101011001;
assign LUT_1[55733] = 32'b00000000000000000100110111010101;
assign LUT_1[55734] = 32'b00000000000000000111010011101010;
assign LUT_1[55735] = 32'b00000000000000000000100101100110;
assign LUT_1[55736] = 32'b00000000000000000010111001110111;
assign LUT_1[55737] = 32'b11111111111111111100001011110011;
assign LUT_1[55738] = 32'b11111111111111111110101000001000;
assign LUT_1[55739] = 32'b11111111111111110111111010000100;
assign LUT_1[55740] = 32'b00000000000000001010110011001110;
assign LUT_1[55741] = 32'b00000000000000000100000101001010;
assign LUT_1[55742] = 32'b00000000000000000110100001011111;
assign LUT_1[55743] = 32'b11111111111111111111110011011011;
assign LUT_1[55744] = 32'b00000000000000000010110011001001;
assign LUT_1[55745] = 32'b11111111111111111100000101000101;
assign LUT_1[55746] = 32'b11111111111111111110100001011010;
assign LUT_1[55747] = 32'b11111111111111110111110011010110;
assign LUT_1[55748] = 32'b00000000000000001010101100100000;
assign LUT_1[55749] = 32'b00000000000000000011111110011100;
assign LUT_1[55750] = 32'b00000000000000000110011010110001;
assign LUT_1[55751] = 32'b11111111111111111111101100101101;
assign LUT_1[55752] = 32'b00000000000000000010000000111110;
assign LUT_1[55753] = 32'b11111111111111111011010010111010;
assign LUT_1[55754] = 32'b11111111111111111101101111001111;
assign LUT_1[55755] = 32'b11111111111111110111000001001011;
assign LUT_1[55756] = 32'b00000000000000001001111010010101;
assign LUT_1[55757] = 32'b00000000000000000011001100010001;
assign LUT_1[55758] = 32'b00000000000000000101101000100110;
assign LUT_1[55759] = 32'b11111111111111111110111010100010;
assign LUT_1[55760] = 32'b00000000000000000100101110101011;
assign LUT_1[55761] = 32'b11111111111111111110000000100111;
assign LUT_1[55762] = 32'b00000000000000000000011100111100;
assign LUT_1[55763] = 32'b11111111111111111001101110111000;
assign LUT_1[55764] = 32'b00000000000000001100101000000010;
assign LUT_1[55765] = 32'b00000000000000000101111001111110;
assign LUT_1[55766] = 32'b00000000000000001000010110010011;
assign LUT_1[55767] = 32'b00000000000000000001101000001111;
assign LUT_1[55768] = 32'b00000000000000000011111100100000;
assign LUT_1[55769] = 32'b11111111111111111101001110011100;
assign LUT_1[55770] = 32'b11111111111111111111101010110001;
assign LUT_1[55771] = 32'b11111111111111111000111100101101;
assign LUT_1[55772] = 32'b00000000000000001011110101110111;
assign LUT_1[55773] = 32'b00000000000000000101000111110011;
assign LUT_1[55774] = 32'b00000000000000000111100100001000;
assign LUT_1[55775] = 32'b00000000000000000000110110000100;
assign LUT_1[55776] = 32'b00000000000000000011101110001000;
assign LUT_1[55777] = 32'b11111111111111111101000000000100;
assign LUT_1[55778] = 32'b11111111111111111111011100011001;
assign LUT_1[55779] = 32'b11111111111111111000101110010101;
assign LUT_1[55780] = 32'b00000000000000001011100111011111;
assign LUT_1[55781] = 32'b00000000000000000100111001011011;
assign LUT_1[55782] = 32'b00000000000000000111010101110000;
assign LUT_1[55783] = 32'b00000000000000000000100111101100;
assign LUT_1[55784] = 32'b00000000000000000010111011111101;
assign LUT_1[55785] = 32'b11111111111111111100001101111001;
assign LUT_1[55786] = 32'b11111111111111111110101010001110;
assign LUT_1[55787] = 32'b11111111111111110111111100001010;
assign LUT_1[55788] = 32'b00000000000000001010110101010100;
assign LUT_1[55789] = 32'b00000000000000000100000111010000;
assign LUT_1[55790] = 32'b00000000000000000110100011100101;
assign LUT_1[55791] = 32'b11111111111111111111110101100001;
assign LUT_1[55792] = 32'b00000000000000000101101001101010;
assign LUT_1[55793] = 32'b11111111111111111110111011100110;
assign LUT_1[55794] = 32'b00000000000000000001010111111011;
assign LUT_1[55795] = 32'b11111111111111111010101001110111;
assign LUT_1[55796] = 32'b00000000000000001101100011000001;
assign LUT_1[55797] = 32'b00000000000000000110110100111101;
assign LUT_1[55798] = 32'b00000000000000001001010001010010;
assign LUT_1[55799] = 32'b00000000000000000010100011001110;
assign LUT_1[55800] = 32'b00000000000000000100110111011111;
assign LUT_1[55801] = 32'b11111111111111111110001001011011;
assign LUT_1[55802] = 32'b00000000000000000000100101110000;
assign LUT_1[55803] = 32'b11111111111111111001110111101100;
assign LUT_1[55804] = 32'b00000000000000001100110000110110;
assign LUT_1[55805] = 32'b00000000000000000110000010110010;
assign LUT_1[55806] = 32'b00000000000000001000011111000111;
assign LUT_1[55807] = 32'b00000000000000000001110001000011;
assign LUT_1[55808] = 32'b11111111111111111001101111101111;
assign LUT_1[55809] = 32'b11111111111111110011000001101011;
assign LUT_1[55810] = 32'b11111111111111110101011110000000;
assign LUT_1[55811] = 32'b11111111111111101110101111111100;
assign LUT_1[55812] = 32'b00000000000000000001101001000110;
assign LUT_1[55813] = 32'b11111111111111111010111011000010;
assign LUT_1[55814] = 32'b11111111111111111101010111010111;
assign LUT_1[55815] = 32'b11111111111111110110101001010011;
assign LUT_1[55816] = 32'b11111111111111111000111101100100;
assign LUT_1[55817] = 32'b11111111111111110010001111100000;
assign LUT_1[55818] = 32'b11111111111111110100101011110101;
assign LUT_1[55819] = 32'b11111111111111101101111101110001;
assign LUT_1[55820] = 32'b00000000000000000000110110111011;
assign LUT_1[55821] = 32'b11111111111111111010001000110111;
assign LUT_1[55822] = 32'b11111111111111111100100101001100;
assign LUT_1[55823] = 32'b11111111111111110101110111001000;
assign LUT_1[55824] = 32'b11111111111111111011101011010001;
assign LUT_1[55825] = 32'b11111111111111110100111101001101;
assign LUT_1[55826] = 32'b11111111111111110111011001100010;
assign LUT_1[55827] = 32'b11111111111111110000101011011110;
assign LUT_1[55828] = 32'b00000000000000000011100100101000;
assign LUT_1[55829] = 32'b11111111111111111100110110100100;
assign LUT_1[55830] = 32'b11111111111111111111010010111001;
assign LUT_1[55831] = 32'b11111111111111111000100100110101;
assign LUT_1[55832] = 32'b11111111111111111010111001000110;
assign LUT_1[55833] = 32'b11111111111111110100001011000010;
assign LUT_1[55834] = 32'b11111111111111110110100111010111;
assign LUT_1[55835] = 32'b11111111111111101111111001010011;
assign LUT_1[55836] = 32'b00000000000000000010110010011101;
assign LUT_1[55837] = 32'b11111111111111111100000100011001;
assign LUT_1[55838] = 32'b11111111111111111110100000101110;
assign LUT_1[55839] = 32'b11111111111111110111110010101010;
assign LUT_1[55840] = 32'b11111111111111111010101010101110;
assign LUT_1[55841] = 32'b11111111111111110011111100101010;
assign LUT_1[55842] = 32'b11111111111111110110011000111111;
assign LUT_1[55843] = 32'b11111111111111101111101010111011;
assign LUT_1[55844] = 32'b00000000000000000010100100000101;
assign LUT_1[55845] = 32'b11111111111111111011110110000001;
assign LUT_1[55846] = 32'b11111111111111111110010010010110;
assign LUT_1[55847] = 32'b11111111111111110111100100010010;
assign LUT_1[55848] = 32'b11111111111111111001111000100011;
assign LUT_1[55849] = 32'b11111111111111110011001010011111;
assign LUT_1[55850] = 32'b11111111111111110101100110110100;
assign LUT_1[55851] = 32'b11111111111111101110111000110000;
assign LUT_1[55852] = 32'b00000000000000000001110001111010;
assign LUT_1[55853] = 32'b11111111111111111011000011110110;
assign LUT_1[55854] = 32'b11111111111111111101100000001011;
assign LUT_1[55855] = 32'b11111111111111110110110010000111;
assign LUT_1[55856] = 32'b11111111111111111100100110010000;
assign LUT_1[55857] = 32'b11111111111111110101111000001100;
assign LUT_1[55858] = 32'b11111111111111111000010100100001;
assign LUT_1[55859] = 32'b11111111111111110001100110011101;
assign LUT_1[55860] = 32'b00000000000000000100011111100111;
assign LUT_1[55861] = 32'b11111111111111111101110001100011;
assign LUT_1[55862] = 32'b00000000000000000000001101111000;
assign LUT_1[55863] = 32'b11111111111111111001011111110100;
assign LUT_1[55864] = 32'b11111111111111111011110100000101;
assign LUT_1[55865] = 32'b11111111111111110101000110000001;
assign LUT_1[55866] = 32'b11111111111111110111100010010110;
assign LUT_1[55867] = 32'b11111111111111110000110100010010;
assign LUT_1[55868] = 32'b00000000000000000011101101011100;
assign LUT_1[55869] = 32'b11111111111111111100111111011000;
assign LUT_1[55870] = 32'b11111111111111111111011011101101;
assign LUT_1[55871] = 32'b11111111111111111000101101101001;
assign LUT_1[55872] = 32'b11111111111111111011101101010111;
assign LUT_1[55873] = 32'b11111111111111110100111111010011;
assign LUT_1[55874] = 32'b11111111111111110111011011101000;
assign LUT_1[55875] = 32'b11111111111111110000101101100100;
assign LUT_1[55876] = 32'b00000000000000000011100110101110;
assign LUT_1[55877] = 32'b11111111111111111100111000101010;
assign LUT_1[55878] = 32'b11111111111111111111010100111111;
assign LUT_1[55879] = 32'b11111111111111111000100110111011;
assign LUT_1[55880] = 32'b11111111111111111010111011001100;
assign LUT_1[55881] = 32'b11111111111111110100001101001000;
assign LUT_1[55882] = 32'b11111111111111110110101001011101;
assign LUT_1[55883] = 32'b11111111111111101111111011011001;
assign LUT_1[55884] = 32'b00000000000000000010110100100011;
assign LUT_1[55885] = 32'b11111111111111111100000110011111;
assign LUT_1[55886] = 32'b11111111111111111110100010110100;
assign LUT_1[55887] = 32'b11111111111111110111110100110000;
assign LUT_1[55888] = 32'b11111111111111111101101000111001;
assign LUT_1[55889] = 32'b11111111111111110110111010110101;
assign LUT_1[55890] = 32'b11111111111111111001010111001010;
assign LUT_1[55891] = 32'b11111111111111110010101001000110;
assign LUT_1[55892] = 32'b00000000000000000101100010010000;
assign LUT_1[55893] = 32'b11111111111111111110110100001100;
assign LUT_1[55894] = 32'b00000000000000000001010000100001;
assign LUT_1[55895] = 32'b11111111111111111010100010011101;
assign LUT_1[55896] = 32'b11111111111111111100110110101110;
assign LUT_1[55897] = 32'b11111111111111110110001000101010;
assign LUT_1[55898] = 32'b11111111111111111000100100111111;
assign LUT_1[55899] = 32'b11111111111111110001110110111011;
assign LUT_1[55900] = 32'b00000000000000000100110000000101;
assign LUT_1[55901] = 32'b11111111111111111110000010000001;
assign LUT_1[55902] = 32'b00000000000000000000011110010110;
assign LUT_1[55903] = 32'b11111111111111111001110000010010;
assign LUT_1[55904] = 32'b11111111111111111100101000010110;
assign LUT_1[55905] = 32'b11111111111111110101111010010010;
assign LUT_1[55906] = 32'b11111111111111111000010110100111;
assign LUT_1[55907] = 32'b11111111111111110001101000100011;
assign LUT_1[55908] = 32'b00000000000000000100100001101101;
assign LUT_1[55909] = 32'b11111111111111111101110011101001;
assign LUT_1[55910] = 32'b00000000000000000000001111111110;
assign LUT_1[55911] = 32'b11111111111111111001100001111010;
assign LUT_1[55912] = 32'b11111111111111111011110110001011;
assign LUT_1[55913] = 32'b11111111111111110101001000000111;
assign LUT_1[55914] = 32'b11111111111111110111100100011100;
assign LUT_1[55915] = 32'b11111111111111110000110110011000;
assign LUT_1[55916] = 32'b00000000000000000011101111100010;
assign LUT_1[55917] = 32'b11111111111111111101000001011110;
assign LUT_1[55918] = 32'b11111111111111111111011101110011;
assign LUT_1[55919] = 32'b11111111111111111000101111101111;
assign LUT_1[55920] = 32'b11111111111111111110100011111000;
assign LUT_1[55921] = 32'b11111111111111110111110101110100;
assign LUT_1[55922] = 32'b11111111111111111010010010001001;
assign LUT_1[55923] = 32'b11111111111111110011100100000101;
assign LUT_1[55924] = 32'b00000000000000000110011101001111;
assign LUT_1[55925] = 32'b11111111111111111111101111001011;
assign LUT_1[55926] = 32'b00000000000000000010001011100000;
assign LUT_1[55927] = 32'b11111111111111111011011101011100;
assign LUT_1[55928] = 32'b11111111111111111101110001101101;
assign LUT_1[55929] = 32'b11111111111111110111000011101001;
assign LUT_1[55930] = 32'b11111111111111111001011111111110;
assign LUT_1[55931] = 32'b11111111111111110010110001111010;
assign LUT_1[55932] = 32'b00000000000000000101101011000100;
assign LUT_1[55933] = 32'b11111111111111111110111101000000;
assign LUT_1[55934] = 32'b00000000000000000001011001010101;
assign LUT_1[55935] = 32'b11111111111111111010101011010001;
assign LUT_1[55936] = 32'b11111111111111111100101111110010;
assign LUT_1[55937] = 32'b11111111111111110110000001101110;
assign LUT_1[55938] = 32'b11111111111111111000011110000011;
assign LUT_1[55939] = 32'b11111111111111110001101111111111;
assign LUT_1[55940] = 32'b00000000000000000100101001001001;
assign LUT_1[55941] = 32'b11111111111111111101111011000101;
assign LUT_1[55942] = 32'b00000000000000000000010111011010;
assign LUT_1[55943] = 32'b11111111111111111001101001010110;
assign LUT_1[55944] = 32'b11111111111111111011111101100111;
assign LUT_1[55945] = 32'b11111111111111110101001111100011;
assign LUT_1[55946] = 32'b11111111111111110111101011111000;
assign LUT_1[55947] = 32'b11111111111111110000111101110100;
assign LUT_1[55948] = 32'b00000000000000000011110110111110;
assign LUT_1[55949] = 32'b11111111111111111101001000111010;
assign LUT_1[55950] = 32'b11111111111111111111100101001111;
assign LUT_1[55951] = 32'b11111111111111111000110111001011;
assign LUT_1[55952] = 32'b11111111111111111110101011010100;
assign LUT_1[55953] = 32'b11111111111111110111111101010000;
assign LUT_1[55954] = 32'b11111111111111111010011001100101;
assign LUT_1[55955] = 32'b11111111111111110011101011100001;
assign LUT_1[55956] = 32'b00000000000000000110100100101011;
assign LUT_1[55957] = 32'b11111111111111111111110110100111;
assign LUT_1[55958] = 32'b00000000000000000010010010111100;
assign LUT_1[55959] = 32'b11111111111111111011100100111000;
assign LUT_1[55960] = 32'b11111111111111111101111001001001;
assign LUT_1[55961] = 32'b11111111111111110111001011000101;
assign LUT_1[55962] = 32'b11111111111111111001100111011010;
assign LUT_1[55963] = 32'b11111111111111110010111001010110;
assign LUT_1[55964] = 32'b00000000000000000101110010100000;
assign LUT_1[55965] = 32'b11111111111111111111000100011100;
assign LUT_1[55966] = 32'b00000000000000000001100000110001;
assign LUT_1[55967] = 32'b11111111111111111010110010101101;
assign LUT_1[55968] = 32'b11111111111111111101101010110001;
assign LUT_1[55969] = 32'b11111111111111110110111100101101;
assign LUT_1[55970] = 32'b11111111111111111001011001000010;
assign LUT_1[55971] = 32'b11111111111111110010101010111110;
assign LUT_1[55972] = 32'b00000000000000000101100100001000;
assign LUT_1[55973] = 32'b11111111111111111110110110000100;
assign LUT_1[55974] = 32'b00000000000000000001010010011001;
assign LUT_1[55975] = 32'b11111111111111111010100100010101;
assign LUT_1[55976] = 32'b11111111111111111100111000100110;
assign LUT_1[55977] = 32'b11111111111111110110001010100010;
assign LUT_1[55978] = 32'b11111111111111111000100110110111;
assign LUT_1[55979] = 32'b11111111111111110001111000110011;
assign LUT_1[55980] = 32'b00000000000000000100110001111101;
assign LUT_1[55981] = 32'b11111111111111111110000011111001;
assign LUT_1[55982] = 32'b00000000000000000000100000001110;
assign LUT_1[55983] = 32'b11111111111111111001110010001010;
assign LUT_1[55984] = 32'b11111111111111111111100110010011;
assign LUT_1[55985] = 32'b11111111111111111000111000001111;
assign LUT_1[55986] = 32'b11111111111111111011010100100100;
assign LUT_1[55987] = 32'b11111111111111110100100110100000;
assign LUT_1[55988] = 32'b00000000000000000111011111101010;
assign LUT_1[55989] = 32'b00000000000000000000110001100110;
assign LUT_1[55990] = 32'b00000000000000000011001101111011;
assign LUT_1[55991] = 32'b11111111111111111100011111110111;
assign LUT_1[55992] = 32'b11111111111111111110110100001000;
assign LUT_1[55993] = 32'b11111111111111111000000110000100;
assign LUT_1[55994] = 32'b11111111111111111010100010011001;
assign LUT_1[55995] = 32'b11111111111111110011110100010101;
assign LUT_1[55996] = 32'b00000000000000000110101101011111;
assign LUT_1[55997] = 32'b11111111111111111111111111011011;
assign LUT_1[55998] = 32'b00000000000000000010011011110000;
assign LUT_1[55999] = 32'b11111111111111111011101101101100;
assign LUT_1[56000] = 32'b11111111111111111110101101011010;
assign LUT_1[56001] = 32'b11111111111111110111111111010110;
assign LUT_1[56002] = 32'b11111111111111111010011011101011;
assign LUT_1[56003] = 32'b11111111111111110011101101100111;
assign LUT_1[56004] = 32'b00000000000000000110100110110001;
assign LUT_1[56005] = 32'b11111111111111111111111000101101;
assign LUT_1[56006] = 32'b00000000000000000010010101000010;
assign LUT_1[56007] = 32'b11111111111111111011100110111110;
assign LUT_1[56008] = 32'b11111111111111111101111011001111;
assign LUT_1[56009] = 32'b11111111111111110111001101001011;
assign LUT_1[56010] = 32'b11111111111111111001101001100000;
assign LUT_1[56011] = 32'b11111111111111110010111011011100;
assign LUT_1[56012] = 32'b00000000000000000101110100100110;
assign LUT_1[56013] = 32'b11111111111111111111000110100010;
assign LUT_1[56014] = 32'b00000000000000000001100010110111;
assign LUT_1[56015] = 32'b11111111111111111010110100110011;
assign LUT_1[56016] = 32'b00000000000000000000101000111100;
assign LUT_1[56017] = 32'b11111111111111111001111010111000;
assign LUT_1[56018] = 32'b11111111111111111100010111001101;
assign LUT_1[56019] = 32'b11111111111111110101101001001001;
assign LUT_1[56020] = 32'b00000000000000001000100010010011;
assign LUT_1[56021] = 32'b00000000000000000001110100001111;
assign LUT_1[56022] = 32'b00000000000000000100010000100100;
assign LUT_1[56023] = 32'b11111111111111111101100010100000;
assign LUT_1[56024] = 32'b11111111111111111111110110110001;
assign LUT_1[56025] = 32'b11111111111111111001001000101101;
assign LUT_1[56026] = 32'b11111111111111111011100101000010;
assign LUT_1[56027] = 32'b11111111111111110100110110111110;
assign LUT_1[56028] = 32'b00000000000000000111110000001000;
assign LUT_1[56029] = 32'b00000000000000000001000010000100;
assign LUT_1[56030] = 32'b00000000000000000011011110011001;
assign LUT_1[56031] = 32'b11111111111111111100110000010101;
assign LUT_1[56032] = 32'b11111111111111111111101000011001;
assign LUT_1[56033] = 32'b11111111111111111000111010010101;
assign LUT_1[56034] = 32'b11111111111111111011010110101010;
assign LUT_1[56035] = 32'b11111111111111110100101000100110;
assign LUT_1[56036] = 32'b00000000000000000111100001110000;
assign LUT_1[56037] = 32'b00000000000000000000110011101100;
assign LUT_1[56038] = 32'b00000000000000000011010000000001;
assign LUT_1[56039] = 32'b11111111111111111100100001111101;
assign LUT_1[56040] = 32'b11111111111111111110110110001110;
assign LUT_1[56041] = 32'b11111111111111111000001000001010;
assign LUT_1[56042] = 32'b11111111111111111010100100011111;
assign LUT_1[56043] = 32'b11111111111111110011110110011011;
assign LUT_1[56044] = 32'b00000000000000000110101111100101;
assign LUT_1[56045] = 32'b00000000000000000000000001100001;
assign LUT_1[56046] = 32'b00000000000000000010011101110110;
assign LUT_1[56047] = 32'b11111111111111111011101111110010;
assign LUT_1[56048] = 32'b00000000000000000001100011111011;
assign LUT_1[56049] = 32'b11111111111111111010110101110111;
assign LUT_1[56050] = 32'b11111111111111111101010010001100;
assign LUT_1[56051] = 32'b11111111111111110110100100001000;
assign LUT_1[56052] = 32'b00000000000000001001011101010010;
assign LUT_1[56053] = 32'b00000000000000000010101111001110;
assign LUT_1[56054] = 32'b00000000000000000101001011100011;
assign LUT_1[56055] = 32'b11111111111111111110011101011111;
assign LUT_1[56056] = 32'b00000000000000000000110001110000;
assign LUT_1[56057] = 32'b11111111111111111010000011101100;
assign LUT_1[56058] = 32'b11111111111111111100100000000001;
assign LUT_1[56059] = 32'b11111111111111110101110001111101;
assign LUT_1[56060] = 32'b00000000000000001000101011000111;
assign LUT_1[56061] = 32'b00000000000000000001111101000011;
assign LUT_1[56062] = 32'b00000000000000000100011001011000;
assign LUT_1[56063] = 32'b11111111111111111101101011010100;
assign LUT_1[56064] = 32'b11111111111111110111100011111011;
assign LUT_1[56065] = 32'b11111111111111110000110101110111;
assign LUT_1[56066] = 32'b11111111111111110011010010001100;
assign LUT_1[56067] = 32'b11111111111111101100100100001000;
assign LUT_1[56068] = 32'b11111111111111111111011101010010;
assign LUT_1[56069] = 32'b11111111111111111000101111001110;
assign LUT_1[56070] = 32'b11111111111111111011001011100011;
assign LUT_1[56071] = 32'b11111111111111110100011101011111;
assign LUT_1[56072] = 32'b11111111111111110110110001110000;
assign LUT_1[56073] = 32'b11111111111111110000000011101100;
assign LUT_1[56074] = 32'b11111111111111110010100000000001;
assign LUT_1[56075] = 32'b11111111111111101011110001111101;
assign LUT_1[56076] = 32'b11111111111111111110101011000111;
assign LUT_1[56077] = 32'b11111111111111110111111101000011;
assign LUT_1[56078] = 32'b11111111111111111010011001011000;
assign LUT_1[56079] = 32'b11111111111111110011101011010100;
assign LUT_1[56080] = 32'b11111111111111111001011111011101;
assign LUT_1[56081] = 32'b11111111111111110010110001011001;
assign LUT_1[56082] = 32'b11111111111111110101001101101110;
assign LUT_1[56083] = 32'b11111111111111101110011111101010;
assign LUT_1[56084] = 32'b00000000000000000001011000110100;
assign LUT_1[56085] = 32'b11111111111111111010101010110000;
assign LUT_1[56086] = 32'b11111111111111111101000111000101;
assign LUT_1[56087] = 32'b11111111111111110110011001000001;
assign LUT_1[56088] = 32'b11111111111111111000101101010010;
assign LUT_1[56089] = 32'b11111111111111110001111111001110;
assign LUT_1[56090] = 32'b11111111111111110100011011100011;
assign LUT_1[56091] = 32'b11111111111111101101101101011111;
assign LUT_1[56092] = 32'b00000000000000000000100110101001;
assign LUT_1[56093] = 32'b11111111111111111001111000100101;
assign LUT_1[56094] = 32'b11111111111111111100010100111010;
assign LUT_1[56095] = 32'b11111111111111110101100110110110;
assign LUT_1[56096] = 32'b11111111111111111000011110111010;
assign LUT_1[56097] = 32'b11111111111111110001110000110110;
assign LUT_1[56098] = 32'b11111111111111110100001101001011;
assign LUT_1[56099] = 32'b11111111111111101101011111000111;
assign LUT_1[56100] = 32'b00000000000000000000011000010001;
assign LUT_1[56101] = 32'b11111111111111111001101010001101;
assign LUT_1[56102] = 32'b11111111111111111100000110100010;
assign LUT_1[56103] = 32'b11111111111111110101011000011110;
assign LUT_1[56104] = 32'b11111111111111110111101100101111;
assign LUT_1[56105] = 32'b11111111111111110000111110101011;
assign LUT_1[56106] = 32'b11111111111111110011011011000000;
assign LUT_1[56107] = 32'b11111111111111101100101100111100;
assign LUT_1[56108] = 32'b11111111111111111111100110000110;
assign LUT_1[56109] = 32'b11111111111111111000111000000010;
assign LUT_1[56110] = 32'b11111111111111111011010100010111;
assign LUT_1[56111] = 32'b11111111111111110100100110010011;
assign LUT_1[56112] = 32'b11111111111111111010011010011100;
assign LUT_1[56113] = 32'b11111111111111110011101100011000;
assign LUT_1[56114] = 32'b11111111111111110110001000101101;
assign LUT_1[56115] = 32'b11111111111111101111011010101001;
assign LUT_1[56116] = 32'b00000000000000000010010011110011;
assign LUT_1[56117] = 32'b11111111111111111011100101101111;
assign LUT_1[56118] = 32'b11111111111111111110000010000100;
assign LUT_1[56119] = 32'b11111111111111110111010100000000;
assign LUT_1[56120] = 32'b11111111111111111001101000010001;
assign LUT_1[56121] = 32'b11111111111111110010111010001101;
assign LUT_1[56122] = 32'b11111111111111110101010110100010;
assign LUT_1[56123] = 32'b11111111111111101110101000011110;
assign LUT_1[56124] = 32'b00000000000000000001100001101000;
assign LUT_1[56125] = 32'b11111111111111111010110011100100;
assign LUT_1[56126] = 32'b11111111111111111101001111111001;
assign LUT_1[56127] = 32'b11111111111111110110100001110101;
assign LUT_1[56128] = 32'b11111111111111111001100001100011;
assign LUT_1[56129] = 32'b11111111111111110010110011011111;
assign LUT_1[56130] = 32'b11111111111111110101001111110100;
assign LUT_1[56131] = 32'b11111111111111101110100001110000;
assign LUT_1[56132] = 32'b00000000000000000001011010111010;
assign LUT_1[56133] = 32'b11111111111111111010101100110110;
assign LUT_1[56134] = 32'b11111111111111111101001001001011;
assign LUT_1[56135] = 32'b11111111111111110110011011000111;
assign LUT_1[56136] = 32'b11111111111111111000101111011000;
assign LUT_1[56137] = 32'b11111111111111110010000001010100;
assign LUT_1[56138] = 32'b11111111111111110100011101101001;
assign LUT_1[56139] = 32'b11111111111111101101101111100101;
assign LUT_1[56140] = 32'b00000000000000000000101000101111;
assign LUT_1[56141] = 32'b11111111111111111001111010101011;
assign LUT_1[56142] = 32'b11111111111111111100010111000000;
assign LUT_1[56143] = 32'b11111111111111110101101000111100;
assign LUT_1[56144] = 32'b11111111111111111011011101000101;
assign LUT_1[56145] = 32'b11111111111111110100101111000001;
assign LUT_1[56146] = 32'b11111111111111110111001011010110;
assign LUT_1[56147] = 32'b11111111111111110000011101010010;
assign LUT_1[56148] = 32'b00000000000000000011010110011100;
assign LUT_1[56149] = 32'b11111111111111111100101000011000;
assign LUT_1[56150] = 32'b11111111111111111111000100101101;
assign LUT_1[56151] = 32'b11111111111111111000010110101001;
assign LUT_1[56152] = 32'b11111111111111111010101010111010;
assign LUT_1[56153] = 32'b11111111111111110011111100110110;
assign LUT_1[56154] = 32'b11111111111111110110011001001011;
assign LUT_1[56155] = 32'b11111111111111101111101011000111;
assign LUT_1[56156] = 32'b00000000000000000010100100010001;
assign LUT_1[56157] = 32'b11111111111111111011110110001101;
assign LUT_1[56158] = 32'b11111111111111111110010010100010;
assign LUT_1[56159] = 32'b11111111111111110111100100011110;
assign LUT_1[56160] = 32'b11111111111111111010011100100010;
assign LUT_1[56161] = 32'b11111111111111110011101110011110;
assign LUT_1[56162] = 32'b11111111111111110110001010110011;
assign LUT_1[56163] = 32'b11111111111111101111011100101111;
assign LUT_1[56164] = 32'b00000000000000000010010101111001;
assign LUT_1[56165] = 32'b11111111111111111011100111110101;
assign LUT_1[56166] = 32'b11111111111111111110000100001010;
assign LUT_1[56167] = 32'b11111111111111110111010110000110;
assign LUT_1[56168] = 32'b11111111111111111001101010010111;
assign LUT_1[56169] = 32'b11111111111111110010111100010011;
assign LUT_1[56170] = 32'b11111111111111110101011000101000;
assign LUT_1[56171] = 32'b11111111111111101110101010100100;
assign LUT_1[56172] = 32'b00000000000000000001100011101110;
assign LUT_1[56173] = 32'b11111111111111111010110101101010;
assign LUT_1[56174] = 32'b11111111111111111101010001111111;
assign LUT_1[56175] = 32'b11111111111111110110100011111011;
assign LUT_1[56176] = 32'b11111111111111111100011000000100;
assign LUT_1[56177] = 32'b11111111111111110101101010000000;
assign LUT_1[56178] = 32'b11111111111111111000000110010101;
assign LUT_1[56179] = 32'b11111111111111110001011000010001;
assign LUT_1[56180] = 32'b00000000000000000100010001011011;
assign LUT_1[56181] = 32'b11111111111111111101100011010111;
assign LUT_1[56182] = 32'b11111111111111111111111111101100;
assign LUT_1[56183] = 32'b11111111111111111001010001101000;
assign LUT_1[56184] = 32'b11111111111111111011100101111001;
assign LUT_1[56185] = 32'b11111111111111110100110111110101;
assign LUT_1[56186] = 32'b11111111111111110111010100001010;
assign LUT_1[56187] = 32'b11111111111111110000100110000110;
assign LUT_1[56188] = 32'b00000000000000000011011111010000;
assign LUT_1[56189] = 32'b11111111111111111100110001001100;
assign LUT_1[56190] = 32'b11111111111111111111001101100001;
assign LUT_1[56191] = 32'b11111111111111111000011111011101;
assign LUT_1[56192] = 32'b11111111111111111010100011111110;
assign LUT_1[56193] = 32'b11111111111111110011110101111010;
assign LUT_1[56194] = 32'b11111111111111110110010010001111;
assign LUT_1[56195] = 32'b11111111111111101111100100001011;
assign LUT_1[56196] = 32'b00000000000000000010011101010101;
assign LUT_1[56197] = 32'b11111111111111111011101111010001;
assign LUT_1[56198] = 32'b11111111111111111110001011100110;
assign LUT_1[56199] = 32'b11111111111111110111011101100010;
assign LUT_1[56200] = 32'b11111111111111111001110001110011;
assign LUT_1[56201] = 32'b11111111111111110011000011101111;
assign LUT_1[56202] = 32'b11111111111111110101100000000100;
assign LUT_1[56203] = 32'b11111111111111101110110010000000;
assign LUT_1[56204] = 32'b00000000000000000001101011001010;
assign LUT_1[56205] = 32'b11111111111111111010111101000110;
assign LUT_1[56206] = 32'b11111111111111111101011001011011;
assign LUT_1[56207] = 32'b11111111111111110110101011010111;
assign LUT_1[56208] = 32'b11111111111111111100011111100000;
assign LUT_1[56209] = 32'b11111111111111110101110001011100;
assign LUT_1[56210] = 32'b11111111111111111000001101110001;
assign LUT_1[56211] = 32'b11111111111111110001011111101101;
assign LUT_1[56212] = 32'b00000000000000000100011000110111;
assign LUT_1[56213] = 32'b11111111111111111101101010110011;
assign LUT_1[56214] = 32'b00000000000000000000000111001000;
assign LUT_1[56215] = 32'b11111111111111111001011001000100;
assign LUT_1[56216] = 32'b11111111111111111011101101010101;
assign LUT_1[56217] = 32'b11111111111111110100111111010001;
assign LUT_1[56218] = 32'b11111111111111110111011011100110;
assign LUT_1[56219] = 32'b11111111111111110000101101100010;
assign LUT_1[56220] = 32'b00000000000000000011100110101100;
assign LUT_1[56221] = 32'b11111111111111111100111000101000;
assign LUT_1[56222] = 32'b11111111111111111111010100111101;
assign LUT_1[56223] = 32'b11111111111111111000100110111001;
assign LUT_1[56224] = 32'b11111111111111111011011110111101;
assign LUT_1[56225] = 32'b11111111111111110100110000111001;
assign LUT_1[56226] = 32'b11111111111111110111001101001110;
assign LUT_1[56227] = 32'b11111111111111110000011111001010;
assign LUT_1[56228] = 32'b00000000000000000011011000010100;
assign LUT_1[56229] = 32'b11111111111111111100101010010000;
assign LUT_1[56230] = 32'b11111111111111111111000110100101;
assign LUT_1[56231] = 32'b11111111111111111000011000100001;
assign LUT_1[56232] = 32'b11111111111111111010101100110010;
assign LUT_1[56233] = 32'b11111111111111110011111110101110;
assign LUT_1[56234] = 32'b11111111111111110110011011000011;
assign LUT_1[56235] = 32'b11111111111111101111101100111111;
assign LUT_1[56236] = 32'b00000000000000000010100110001001;
assign LUT_1[56237] = 32'b11111111111111111011111000000101;
assign LUT_1[56238] = 32'b11111111111111111110010100011010;
assign LUT_1[56239] = 32'b11111111111111110111100110010110;
assign LUT_1[56240] = 32'b11111111111111111101011010011111;
assign LUT_1[56241] = 32'b11111111111111110110101100011011;
assign LUT_1[56242] = 32'b11111111111111111001001000110000;
assign LUT_1[56243] = 32'b11111111111111110010011010101100;
assign LUT_1[56244] = 32'b00000000000000000101010011110110;
assign LUT_1[56245] = 32'b11111111111111111110100101110010;
assign LUT_1[56246] = 32'b00000000000000000001000010000111;
assign LUT_1[56247] = 32'b11111111111111111010010100000011;
assign LUT_1[56248] = 32'b11111111111111111100101000010100;
assign LUT_1[56249] = 32'b11111111111111110101111010010000;
assign LUT_1[56250] = 32'b11111111111111111000010110100101;
assign LUT_1[56251] = 32'b11111111111111110001101000100001;
assign LUT_1[56252] = 32'b00000000000000000100100001101011;
assign LUT_1[56253] = 32'b11111111111111111101110011100111;
assign LUT_1[56254] = 32'b00000000000000000000001111111100;
assign LUT_1[56255] = 32'b11111111111111111001100001111000;
assign LUT_1[56256] = 32'b11111111111111111100100001100110;
assign LUT_1[56257] = 32'b11111111111111110101110011100010;
assign LUT_1[56258] = 32'b11111111111111111000001111110111;
assign LUT_1[56259] = 32'b11111111111111110001100001110011;
assign LUT_1[56260] = 32'b00000000000000000100011010111101;
assign LUT_1[56261] = 32'b11111111111111111101101100111001;
assign LUT_1[56262] = 32'b00000000000000000000001001001110;
assign LUT_1[56263] = 32'b11111111111111111001011011001010;
assign LUT_1[56264] = 32'b11111111111111111011101111011011;
assign LUT_1[56265] = 32'b11111111111111110101000001010111;
assign LUT_1[56266] = 32'b11111111111111110111011101101100;
assign LUT_1[56267] = 32'b11111111111111110000101111101000;
assign LUT_1[56268] = 32'b00000000000000000011101000110010;
assign LUT_1[56269] = 32'b11111111111111111100111010101110;
assign LUT_1[56270] = 32'b11111111111111111111010111000011;
assign LUT_1[56271] = 32'b11111111111111111000101000111111;
assign LUT_1[56272] = 32'b11111111111111111110011101001000;
assign LUT_1[56273] = 32'b11111111111111110111101111000100;
assign LUT_1[56274] = 32'b11111111111111111010001011011001;
assign LUT_1[56275] = 32'b11111111111111110011011101010101;
assign LUT_1[56276] = 32'b00000000000000000110010110011111;
assign LUT_1[56277] = 32'b11111111111111111111101000011011;
assign LUT_1[56278] = 32'b00000000000000000010000100110000;
assign LUT_1[56279] = 32'b11111111111111111011010110101100;
assign LUT_1[56280] = 32'b11111111111111111101101010111101;
assign LUT_1[56281] = 32'b11111111111111110110111100111001;
assign LUT_1[56282] = 32'b11111111111111111001011001001110;
assign LUT_1[56283] = 32'b11111111111111110010101011001010;
assign LUT_1[56284] = 32'b00000000000000000101100100010100;
assign LUT_1[56285] = 32'b11111111111111111110110110010000;
assign LUT_1[56286] = 32'b00000000000000000001010010100101;
assign LUT_1[56287] = 32'b11111111111111111010100100100001;
assign LUT_1[56288] = 32'b11111111111111111101011100100101;
assign LUT_1[56289] = 32'b11111111111111110110101110100001;
assign LUT_1[56290] = 32'b11111111111111111001001010110110;
assign LUT_1[56291] = 32'b11111111111111110010011100110010;
assign LUT_1[56292] = 32'b00000000000000000101010101111100;
assign LUT_1[56293] = 32'b11111111111111111110100111111000;
assign LUT_1[56294] = 32'b00000000000000000001000100001101;
assign LUT_1[56295] = 32'b11111111111111111010010110001001;
assign LUT_1[56296] = 32'b11111111111111111100101010011010;
assign LUT_1[56297] = 32'b11111111111111110101111100010110;
assign LUT_1[56298] = 32'b11111111111111111000011000101011;
assign LUT_1[56299] = 32'b11111111111111110001101010100111;
assign LUT_1[56300] = 32'b00000000000000000100100011110001;
assign LUT_1[56301] = 32'b11111111111111111101110101101101;
assign LUT_1[56302] = 32'b00000000000000000000010010000010;
assign LUT_1[56303] = 32'b11111111111111111001100011111110;
assign LUT_1[56304] = 32'b11111111111111111111011000000111;
assign LUT_1[56305] = 32'b11111111111111111000101010000011;
assign LUT_1[56306] = 32'b11111111111111111011000110011000;
assign LUT_1[56307] = 32'b11111111111111110100011000010100;
assign LUT_1[56308] = 32'b00000000000000000111010001011110;
assign LUT_1[56309] = 32'b00000000000000000000100011011010;
assign LUT_1[56310] = 32'b00000000000000000010111111101111;
assign LUT_1[56311] = 32'b11111111111111111100010001101011;
assign LUT_1[56312] = 32'b11111111111111111110100101111100;
assign LUT_1[56313] = 32'b11111111111111110111110111111000;
assign LUT_1[56314] = 32'b11111111111111111010010100001101;
assign LUT_1[56315] = 32'b11111111111111110011100110001001;
assign LUT_1[56316] = 32'b00000000000000000110011111010011;
assign LUT_1[56317] = 32'b11111111111111111111110001001111;
assign LUT_1[56318] = 32'b00000000000000000010001101100100;
assign LUT_1[56319] = 32'b11111111111111111011011111100000;
assign LUT_1[56320] = 32'b00000000000000000110011000000010;
assign LUT_1[56321] = 32'b11111111111111111111101001111110;
assign LUT_1[56322] = 32'b00000000000000000010000110010011;
assign LUT_1[56323] = 32'b11111111111111111011011000001111;
assign LUT_1[56324] = 32'b00000000000000001110010001011001;
assign LUT_1[56325] = 32'b00000000000000000111100011010101;
assign LUT_1[56326] = 32'b00000000000000001001111111101010;
assign LUT_1[56327] = 32'b00000000000000000011010001100110;
assign LUT_1[56328] = 32'b00000000000000000101100101110111;
assign LUT_1[56329] = 32'b11111111111111111110110111110011;
assign LUT_1[56330] = 32'b00000000000000000001010100001000;
assign LUT_1[56331] = 32'b11111111111111111010100110000100;
assign LUT_1[56332] = 32'b00000000000000001101011111001110;
assign LUT_1[56333] = 32'b00000000000000000110110001001010;
assign LUT_1[56334] = 32'b00000000000000001001001101011111;
assign LUT_1[56335] = 32'b00000000000000000010011111011011;
assign LUT_1[56336] = 32'b00000000000000001000010011100100;
assign LUT_1[56337] = 32'b00000000000000000001100101100000;
assign LUT_1[56338] = 32'b00000000000000000100000001110101;
assign LUT_1[56339] = 32'b11111111111111111101010011110001;
assign LUT_1[56340] = 32'b00000000000000010000001100111011;
assign LUT_1[56341] = 32'b00000000000000001001011110110111;
assign LUT_1[56342] = 32'b00000000000000001011111011001100;
assign LUT_1[56343] = 32'b00000000000000000101001101001000;
assign LUT_1[56344] = 32'b00000000000000000111100001011001;
assign LUT_1[56345] = 32'b00000000000000000000110011010101;
assign LUT_1[56346] = 32'b00000000000000000011001111101010;
assign LUT_1[56347] = 32'b11111111111111111100100001100110;
assign LUT_1[56348] = 32'b00000000000000001111011010110000;
assign LUT_1[56349] = 32'b00000000000000001000101100101100;
assign LUT_1[56350] = 32'b00000000000000001011001001000001;
assign LUT_1[56351] = 32'b00000000000000000100011010111101;
assign LUT_1[56352] = 32'b00000000000000000111010011000001;
assign LUT_1[56353] = 32'b00000000000000000000100100111101;
assign LUT_1[56354] = 32'b00000000000000000011000001010010;
assign LUT_1[56355] = 32'b11111111111111111100010011001110;
assign LUT_1[56356] = 32'b00000000000000001111001100011000;
assign LUT_1[56357] = 32'b00000000000000001000011110010100;
assign LUT_1[56358] = 32'b00000000000000001010111010101001;
assign LUT_1[56359] = 32'b00000000000000000100001100100101;
assign LUT_1[56360] = 32'b00000000000000000110100000110110;
assign LUT_1[56361] = 32'b11111111111111111111110010110010;
assign LUT_1[56362] = 32'b00000000000000000010001111000111;
assign LUT_1[56363] = 32'b11111111111111111011100001000011;
assign LUT_1[56364] = 32'b00000000000000001110011010001101;
assign LUT_1[56365] = 32'b00000000000000000111101100001001;
assign LUT_1[56366] = 32'b00000000000000001010001000011110;
assign LUT_1[56367] = 32'b00000000000000000011011010011010;
assign LUT_1[56368] = 32'b00000000000000001001001110100011;
assign LUT_1[56369] = 32'b00000000000000000010100000011111;
assign LUT_1[56370] = 32'b00000000000000000100111100110100;
assign LUT_1[56371] = 32'b11111111111111111110001110110000;
assign LUT_1[56372] = 32'b00000000000000010001000111111010;
assign LUT_1[56373] = 32'b00000000000000001010011001110110;
assign LUT_1[56374] = 32'b00000000000000001100110110001011;
assign LUT_1[56375] = 32'b00000000000000000110001000000111;
assign LUT_1[56376] = 32'b00000000000000001000011100011000;
assign LUT_1[56377] = 32'b00000000000000000001101110010100;
assign LUT_1[56378] = 32'b00000000000000000100001010101001;
assign LUT_1[56379] = 32'b11111111111111111101011100100101;
assign LUT_1[56380] = 32'b00000000000000010000010101101111;
assign LUT_1[56381] = 32'b00000000000000001001100111101011;
assign LUT_1[56382] = 32'b00000000000000001100000100000000;
assign LUT_1[56383] = 32'b00000000000000000101010101111100;
assign LUT_1[56384] = 32'b00000000000000001000010101101010;
assign LUT_1[56385] = 32'b00000000000000000001100111100110;
assign LUT_1[56386] = 32'b00000000000000000100000011111011;
assign LUT_1[56387] = 32'b11111111111111111101010101110111;
assign LUT_1[56388] = 32'b00000000000000010000001111000001;
assign LUT_1[56389] = 32'b00000000000000001001100000111101;
assign LUT_1[56390] = 32'b00000000000000001011111101010010;
assign LUT_1[56391] = 32'b00000000000000000101001111001110;
assign LUT_1[56392] = 32'b00000000000000000111100011011111;
assign LUT_1[56393] = 32'b00000000000000000000110101011011;
assign LUT_1[56394] = 32'b00000000000000000011010001110000;
assign LUT_1[56395] = 32'b11111111111111111100100011101100;
assign LUT_1[56396] = 32'b00000000000000001111011100110110;
assign LUT_1[56397] = 32'b00000000000000001000101110110010;
assign LUT_1[56398] = 32'b00000000000000001011001011000111;
assign LUT_1[56399] = 32'b00000000000000000100011101000011;
assign LUT_1[56400] = 32'b00000000000000001010010001001100;
assign LUT_1[56401] = 32'b00000000000000000011100011001000;
assign LUT_1[56402] = 32'b00000000000000000101111111011101;
assign LUT_1[56403] = 32'b11111111111111111111010001011001;
assign LUT_1[56404] = 32'b00000000000000010010001010100011;
assign LUT_1[56405] = 32'b00000000000000001011011100011111;
assign LUT_1[56406] = 32'b00000000000000001101111000110100;
assign LUT_1[56407] = 32'b00000000000000000111001010110000;
assign LUT_1[56408] = 32'b00000000000000001001011111000001;
assign LUT_1[56409] = 32'b00000000000000000010110000111101;
assign LUT_1[56410] = 32'b00000000000000000101001101010010;
assign LUT_1[56411] = 32'b11111111111111111110011111001110;
assign LUT_1[56412] = 32'b00000000000000010001011000011000;
assign LUT_1[56413] = 32'b00000000000000001010101010010100;
assign LUT_1[56414] = 32'b00000000000000001101000110101001;
assign LUT_1[56415] = 32'b00000000000000000110011000100101;
assign LUT_1[56416] = 32'b00000000000000001001010000101001;
assign LUT_1[56417] = 32'b00000000000000000010100010100101;
assign LUT_1[56418] = 32'b00000000000000000100111110111010;
assign LUT_1[56419] = 32'b11111111111111111110010000110110;
assign LUT_1[56420] = 32'b00000000000000010001001010000000;
assign LUT_1[56421] = 32'b00000000000000001010011011111100;
assign LUT_1[56422] = 32'b00000000000000001100111000010001;
assign LUT_1[56423] = 32'b00000000000000000110001010001101;
assign LUT_1[56424] = 32'b00000000000000001000011110011110;
assign LUT_1[56425] = 32'b00000000000000000001110000011010;
assign LUT_1[56426] = 32'b00000000000000000100001100101111;
assign LUT_1[56427] = 32'b11111111111111111101011110101011;
assign LUT_1[56428] = 32'b00000000000000010000010111110101;
assign LUT_1[56429] = 32'b00000000000000001001101001110001;
assign LUT_1[56430] = 32'b00000000000000001100000110000110;
assign LUT_1[56431] = 32'b00000000000000000101011000000010;
assign LUT_1[56432] = 32'b00000000000000001011001100001011;
assign LUT_1[56433] = 32'b00000000000000000100011110000111;
assign LUT_1[56434] = 32'b00000000000000000110111010011100;
assign LUT_1[56435] = 32'b00000000000000000000001100011000;
assign LUT_1[56436] = 32'b00000000000000010011000101100010;
assign LUT_1[56437] = 32'b00000000000000001100010111011110;
assign LUT_1[56438] = 32'b00000000000000001110110011110011;
assign LUT_1[56439] = 32'b00000000000000001000000101101111;
assign LUT_1[56440] = 32'b00000000000000001010011010000000;
assign LUT_1[56441] = 32'b00000000000000000011101011111100;
assign LUT_1[56442] = 32'b00000000000000000110001000010001;
assign LUT_1[56443] = 32'b11111111111111111111011010001101;
assign LUT_1[56444] = 32'b00000000000000010010010011010111;
assign LUT_1[56445] = 32'b00000000000000001011100101010011;
assign LUT_1[56446] = 32'b00000000000000001110000001101000;
assign LUT_1[56447] = 32'b00000000000000000111010011100100;
assign LUT_1[56448] = 32'b00000000000000001001011000000101;
assign LUT_1[56449] = 32'b00000000000000000010101010000001;
assign LUT_1[56450] = 32'b00000000000000000101000110010110;
assign LUT_1[56451] = 32'b11111111111111111110011000010010;
assign LUT_1[56452] = 32'b00000000000000010001010001011100;
assign LUT_1[56453] = 32'b00000000000000001010100011011000;
assign LUT_1[56454] = 32'b00000000000000001100111111101101;
assign LUT_1[56455] = 32'b00000000000000000110010001101001;
assign LUT_1[56456] = 32'b00000000000000001000100101111010;
assign LUT_1[56457] = 32'b00000000000000000001110111110110;
assign LUT_1[56458] = 32'b00000000000000000100010100001011;
assign LUT_1[56459] = 32'b11111111111111111101100110000111;
assign LUT_1[56460] = 32'b00000000000000010000011111010001;
assign LUT_1[56461] = 32'b00000000000000001001110001001101;
assign LUT_1[56462] = 32'b00000000000000001100001101100010;
assign LUT_1[56463] = 32'b00000000000000000101011111011110;
assign LUT_1[56464] = 32'b00000000000000001011010011100111;
assign LUT_1[56465] = 32'b00000000000000000100100101100011;
assign LUT_1[56466] = 32'b00000000000000000111000001111000;
assign LUT_1[56467] = 32'b00000000000000000000010011110100;
assign LUT_1[56468] = 32'b00000000000000010011001100111110;
assign LUT_1[56469] = 32'b00000000000000001100011110111010;
assign LUT_1[56470] = 32'b00000000000000001110111011001111;
assign LUT_1[56471] = 32'b00000000000000001000001101001011;
assign LUT_1[56472] = 32'b00000000000000001010100001011100;
assign LUT_1[56473] = 32'b00000000000000000011110011011000;
assign LUT_1[56474] = 32'b00000000000000000110001111101101;
assign LUT_1[56475] = 32'b11111111111111111111100001101001;
assign LUT_1[56476] = 32'b00000000000000010010011010110011;
assign LUT_1[56477] = 32'b00000000000000001011101100101111;
assign LUT_1[56478] = 32'b00000000000000001110001001000100;
assign LUT_1[56479] = 32'b00000000000000000111011011000000;
assign LUT_1[56480] = 32'b00000000000000001010010011000100;
assign LUT_1[56481] = 32'b00000000000000000011100101000000;
assign LUT_1[56482] = 32'b00000000000000000110000001010101;
assign LUT_1[56483] = 32'b11111111111111111111010011010001;
assign LUT_1[56484] = 32'b00000000000000010010001100011011;
assign LUT_1[56485] = 32'b00000000000000001011011110010111;
assign LUT_1[56486] = 32'b00000000000000001101111010101100;
assign LUT_1[56487] = 32'b00000000000000000111001100101000;
assign LUT_1[56488] = 32'b00000000000000001001100000111001;
assign LUT_1[56489] = 32'b00000000000000000010110010110101;
assign LUT_1[56490] = 32'b00000000000000000101001111001010;
assign LUT_1[56491] = 32'b11111111111111111110100001000110;
assign LUT_1[56492] = 32'b00000000000000010001011010010000;
assign LUT_1[56493] = 32'b00000000000000001010101100001100;
assign LUT_1[56494] = 32'b00000000000000001101001000100001;
assign LUT_1[56495] = 32'b00000000000000000110011010011101;
assign LUT_1[56496] = 32'b00000000000000001100001110100110;
assign LUT_1[56497] = 32'b00000000000000000101100000100010;
assign LUT_1[56498] = 32'b00000000000000000111111100110111;
assign LUT_1[56499] = 32'b00000000000000000001001110110011;
assign LUT_1[56500] = 32'b00000000000000010100000111111101;
assign LUT_1[56501] = 32'b00000000000000001101011001111001;
assign LUT_1[56502] = 32'b00000000000000001111110110001110;
assign LUT_1[56503] = 32'b00000000000000001001001000001010;
assign LUT_1[56504] = 32'b00000000000000001011011100011011;
assign LUT_1[56505] = 32'b00000000000000000100101110010111;
assign LUT_1[56506] = 32'b00000000000000000111001010101100;
assign LUT_1[56507] = 32'b00000000000000000000011100101000;
assign LUT_1[56508] = 32'b00000000000000010011010101110010;
assign LUT_1[56509] = 32'b00000000000000001100100111101110;
assign LUT_1[56510] = 32'b00000000000000001111000100000011;
assign LUT_1[56511] = 32'b00000000000000001000010101111111;
assign LUT_1[56512] = 32'b00000000000000001011010101101101;
assign LUT_1[56513] = 32'b00000000000000000100100111101001;
assign LUT_1[56514] = 32'b00000000000000000111000011111110;
assign LUT_1[56515] = 32'b00000000000000000000010101111010;
assign LUT_1[56516] = 32'b00000000000000010011001111000100;
assign LUT_1[56517] = 32'b00000000000000001100100001000000;
assign LUT_1[56518] = 32'b00000000000000001110111101010101;
assign LUT_1[56519] = 32'b00000000000000001000001111010001;
assign LUT_1[56520] = 32'b00000000000000001010100011100010;
assign LUT_1[56521] = 32'b00000000000000000011110101011110;
assign LUT_1[56522] = 32'b00000000000000000110010001110011;
assign LUT_1[56523] = 32'b11111111111111111111100011101111;
assign LUT_1[56524] = 32'b00000000000000010010011100111001;
assign LUT_1[56525] = 32'b00000000000000001011101110110101;
assign LUT_1[56526] = 32'b00000000000000001110001011001010;
assign LUT_1[56527] = 32'b00000000000000000111011101000110;
assign LUT_1[56528] = 32'b00000000000000001101010001001111;
assign LUT_1[56529] = 32'b00000000000000000110100011001011;
assign LUT_1[56530] = 32'b00000000000000001000111111100000;
assign LUT_1[56531] = 32'b00000000000000000010010001011100;
assign LUT_1[56532] = 32'b00000000000000010101001010100110;
assign LUT_1[56533] = 32'b00000000000000001110011100100010;
assign LUT_1[56534] = 32'b00000000000000010000111000110111;
assign LUT_1[56535] = 32'b00000000000000001010001010110011;
assign LUT_1[56536] = 32'b00000000000000001100011111000100;
assign LUT_1[56537] = 32'b00000000000000000101110001000000;
assign LUT_1[56538] = 32'b00000000000000001000001101010101;
assign LUT_1[56539] = 32'b00000000000000000001011111010001;
assign LUT_1[56540] = 32'b00000000000000010100011000011011;
assign LUT_1[56541] = 32'b00000000000000001101101010010111;
assign LUT_1[56542] = 32'b00000000000000010000000110101100;
assign LUT_1[56543] = 32'b00000000000000001001011000101000;
assign LUT_1[56544] = 32'b00000000000000001100010000101100;
assign LUT_1[56545] = 32'b00000000000000000101100010101000;
assign LUT_1[56546] = 32'b00000000000000000111111110111101;
assign LUT_1[56547] = 32'b00000000000000000001010000111001;
assign LUT_1[56548] = 32'b00000000000000010100001010000011;
assign LUT_1[56549] = 32'b00000000000000001101011011111111;
assign LUT_1[56550] = 32'b00000000000000001111111000010100;
assign LUT_1[56551] = 32'b00000000000000001001001010010000;
assign LUT_1[56552] = 32'b00000000000000001011011110100001;
assign LUT_1[56553] = 32'b00000000000000000100110000011101;
assign LUT_1[56554] = 32'b00000000000000000111001100110010;
assign LUT_1[56555] = 32'b00000000000000000000011110101110;
assign LUT_1[56556] = 32'b00000000000000010011010111111000;
assign LUT_1[56557] = 32'b00000000000000001100101001110100;
assign LUT_1[56558] = 32'b00000000000000001111000110001001;
assign LUT_1[56559] = 32'b00000000000000001000011000000101;
assign LUT_1[56560] = 32'b00000000000000001110001100001110;
assign LUT_1[56561] = 32'b00000000000000000111011110001010;
assign LUT_1[56562] = 32'b00000000000000001001111010011111;
assign LUT_1[56563] = 32'b00000000000000000011001100011011;
assign LUT_1[56564] = 32'b00000000000000010110000101100101;
assign LUT_1[56565] = 32'b00000000000000001111010111100001;
assign LUT_1[56566] = 32'b00000000000000010001110011110110;
assign LUT_1[56567] = 32'b00000000000000001011000101110010;
assign LUT_1[56568] = 32'b00000000000000001101011010000011;
assign LUT_1[56569] = 32'b00000000000000000110101011111111;
assign LUT_1[56570] = 32'b00000000000000001001001000010100;
assign LUT_1[56571] = 32'b00000000000000000010011010010000;
assign LUT_1[56572] = 32'b00000000000000010101010011011010;
assign LUT_1[56573] = 32'b00000000000000001110100101010110;
assign LUT_1[56574] = 32'b00000000000000010001000001101011;
assign LUT_1[56575] = 32'b00000000000000001010010011100111;
assign LUT_1[56576] = 32'b00000000000000000100001100001110;
assign LUT_1[56577] = 32'b11111111111111111101011110001010;
assign LUT_1[56578] = 32'b11111111111111111111111010011111;
assign LUT_1[56579] = 32'b11111111111111111001001100011011;
assign LUT_1[56580] = 32'b00000000000000001100000101100101;
assign LUT_1[56581] = 32'b00000000000000000101010111100001;
assign LUT_1[56582] = 32'b00000000000000000111110011110110;
assign LUT_1[56583] = 32'b00000000000000000001000101110010;
assign LUT_1[56584] = 32'b00000000000000000011011010000011;
assign LUT_1[56585] = 32'b11111111111111111100101011111111;
assign LUT_1[56586] = 32'b11111111111111111111001000010100;
assign LUT_1[56587] = 32'b11111111111111111000011010010000;
assign LUT_1[56588] = 32'b00000000000000001011010011011010;
assign LUT_1[56589] = 32'b00000000000000000100100101010110;
assign LUT_1[56590] = 32'b00000000000000000111000001101011;
assign LUT_1[56591] = 32'b00000000000000000000010011100111;
assign LUT_1[56592] = 32'b00000000000000000110000111110000;
assign LUT_1[56593] = 32'b11111111111111111111011001101100;
assign LUT_1[56594] = 32'b00000000000000000001110110000001;
assign LUT_1[56595] = 32'b11111111111111111011000111111101;
assign LUT_1[56596] = 32'b00000000000000001110000001000111;
assign LUT_1[56597] = 32'b00000000000000000111010011000011;
assign LUT_1[56598] = 32'b00000000000000001001101111011000;
assign LUT_1[56599] = 32'b00000000000000000011000001010100;
assign LUT_1[56600] = 32'b00000000000000000101010101100101;
assign LUT_1[56601] = 32'b11111111111111111110100111100001;
assign LUT_1[56602] = 32'b00000000000000000001000011110110;
assign LUT_1[56603] = 32'b11111111111111111010010101110010;
assign LUT_1[56604] = 32'b00000000000000001101001110111100;
assign LUT_1[56605] = 32'b00000000000000000110100000111000;
assign LUT_1[56606] = 32'b00000000000000001000111101001101;
assign LUT_1[56607] = 32'b00000000000000000010001111001001;
assign LUT_1[56608] = 32'b00000000000000000101000111001101;
assign LUT_1[56609] = 32'b11111111111111111110011001001001;
assign LUT_1[56610] = 32'b00000000000000000000110101011110;
assign LUT_1[56611] = 32'b11111111111111111010000111011010;
assign LUT_1[56612] = 32'b00000000000000001101000000100100;
assign LUT_1[56613] = 32'b00000000000000000110010010100000;
assign LUT_1[56614] = 32'b00000000000000001000101110110101;
assign LUT_1[56615] = 32'b00000000000000000010000000110001;
assign LUT_1[56616] = 32'b00000000000000000100010101000010;
assign LUT_1[56617] = 32'b11111111111111111101100110111110;
assign LUT_1[56618] = 32'b00000000000000000000000011010011;
assign LUT_1[56619] = 32'b11111111111111111001010101001111;
assign LUT_1[56620] = 32'b00000000000000001100001110011001;
assign LUT_1[56621] = 32'b00000000000000000101100000010101;
assign LUT_1[56622] = 32'b00000000000000000111111100101010;
assign LUT_1[56623] = 32'b00000000000000000001001110100110;
assign LUT_1[56624] = 32'b00000000000000000111000010101111;
assign LUT_1[56625] = 32'b00000000000000000000010100101011;
assign LUT_1[56626] = 32'b00000000000000000010110001000000;
assign LUT_1[56627] = 32'b11111111111111111100000010111100;
assign LUT_1[56628] = 32'b00000000000000001110111100000110;
assign LUT_1[56629] = 32'b00000000000000001000001110000010;
assign LUT_1[56630] = 32'b00000000000000001010101010010111;
assign LUT_1[56631] = 32'b00000000000000000011111100010011;
assign LUT_1[56632] = 32'b00000000000000000110010000100100;
assign LUT_1[56633] = 32'b11111111111111111111100010100000;
assign LUT_1[56634] = 32'b00000000000000000001111110110101;
assign LUT_1[56635] = 32'b11111111111111111011010000110001;
assign LUT_1[56636] = 32'b00000000000000001110001001111011;
assign LUT_1[56637] = 32'b00000000000000000111011011110111;
assign LUT_1[56638] = 32'b00000000000000001001111000001100;
assign LUT_1[56639] = 32'b00000000000000000011001010001000;
assign LUT_1[56640] = 32'b00000000000000000110001001110110;
assign LUT_1[56641] = 32'b11111111111111111111011011110010;
assign LUT_1[56642] = 32'b00000000000000000001111000000111;
assign LUT_1[56643] = 32'b11111111111111111011001010000011;
assign LUT_1[56644] = 32'b00000000000000001110000011001101;
assign LUT_1[56645] = 32'b00000000000000000111010101001001;
assign LUT_1[56646] = 32'b00000000000000001001110001011110;
assign LUT_1[56647] = 32'b00000000000000000011000011011010;
assign LUT_1[56648] = 32'b00000000000000000101010111101011;
assign LUT_1[56649] = 32'b11111111111111111110101001100111;
assign LUT_1[56650] = 32'b00000000000000000001000101111100;
assign LUT_1[56651] = 32'b11111111111111111010010111111000;
assign LUT_1[56652] = 32'b00000000000000001101010001000010;
assign LUT_1[56653] = 32'b00000000000000000110100010111110;
assign LUT_1[56654] = 32'b00000000000000001000111111010011;
assign LUT_1[56655] = 32'b00000000000000000010010001001111;
assign LUT_1[56656] = 32'b00000000000000001000000101011000;
assign LUT_1[56657] = 32'b00000000000000000001010111010100;
assign LUT_1[56658] = 32'b00000000000000000011110011101001;
assign LUT_1[56659] = 32'b11111111111111111101000101100101;
assign LUT_1[56660] = 32'b00000000000000001111111110101111;
assign LUT_1[56661] = 32'b00000000000000001001010000101011;
assign LUT_1[56662] = 32'b00000000000000001011101101000000;
assign LUT_1[56663] = 32'b00000000000000000100111110111100;
assign LUT_1[56664] = 32'b00000000000000000111010011001101;
assign LUT_1[56665] = 32'b00000000000000000000100101001001;
assign LUT_1[56666] = 32'b00000000000000000011000001011110;
assign LUT_1[56667] = 32'b11111111111111111100010011011010;
assign LUT_1[56668] = 32'b00000000000000001111001100100100;
assign LUT_1[56669] = 32'b00000000000000001000011110100000;
assign LUT_1[56670] = 32'b00000000000000001010111010110101;
assign LUT_1[56671] = 32'b00000000000000000100001100110001;
assign LUT_1[56672] = 32'b00000000000000000111000100110101;
assign LUT_1[56673] = 32'b00000000000000000000010110110001;
assign LUT_1[56674] = 32'b00000000000000000010110011000110;
assign LUT_1[56675] = 32'b11111111111111111100000101000010;
assign LUT_1[56676] = 32'b00000000000000001110111110001100;
assign LUT_1[56677] = 32'b00000000000000001000010000001000;
assign LUT_1[56678] = 32'b00000000000000001010101100011101;
assign LUT_1[56679] = 32'b00000000000000000011111110011001;
assign LUT_1[56680] = 32'b00000000000000000110010010101010;
assign LUT_1[56681] = 32'b11111111111111111111100100100110;
assign LUT_1[56682] = 32'b00000000000000000010000000111011;
assign LUT_1[56683] = 32'b11111111111111111011010010110111;
assign LUT_1[56684] = 32'b00000000000000001110001100000001;
assign LUT_1[56685] = 32'b00000000000000000111011101111101;
assign LUT_1[56686] = 32'b00000000000000001001111010010010;
assign LUT_1[56687] = 32'b00000000000000000011001100001110;
assign LUT_1[56688] = 32'b00000000000000001001000000010111;
assign LUT_1[56689] = 32'b00000000000000000010010010010011;
assign LUT_1[56690] = 32'b00000000000000000100101110101000;
assign LUT_1[56691] = 32'b11111111111111111110000000100100;
assign LUT_1[56692] = 32'b00000000000000010000111001101110;
assign LUT_1[56693] = 32'b00000000000000001010001011101010;
assign LUT_1[56694] = 32'b00000000000000001100100111111111;
assign LUT_1[56695] = 32'b00000000000000000101111001111011;
assign LUT_1[56696] = 32'b00000000000000001000001110001100;
assign LUT_1[56697] = 32'b00000000000000000001100000001000;
assign LUT_1[56698] = 32'b00000000000000000011111100011101;
assign LUT_1[56699] = 32'b11111111111111111101001110011001;
assign LUT_1[56700] = 32'b00000000000000010000000111100011;
assign LUT_1[56701] = 32'b00000000000000001001011001011111;
assign LUT_1[56702] = 32'b00000000000000001011110101110100;
assign LUT_1[56703] = 32'b00000000000000000101000111110000;
assign LUT_1[56704] = 32'b00000000000000000111001100010001;
assign LUT_1[56705] = 32'b00000000000000000000011110001101;
assign LUT_1[56706] = 32'b00000000000000000010111010100010;
assign LUT_1[56707] = 32'b11111111111111111100001100011110;
assign LUT_1[56708] = 32'b00000000000000001111000101101000;
assign LUT_1[56709] = 32'b00000000000000001000010111100100;
assign LUT_1[56710] = 32'b00000000000000001010110011111001;
assign LUT_1[56711] = 32'b00000000000000000100000101110101;
assign LUT_1[56712] = 32'b00000000000000000110011010000110;
assign LUT_1[56713] = 32'b11111111111111111111101100000010;
assign LUT_1[56714] = 32'b00000000000000000010001000010111;
assign LUT_1[56715] = 32'b11111111111111111011011010010011;
assign LUT_1[56716] = 32'b00000000000000001110010011011101;
assign LUT_1[56717] = 32'b00000000000000000111100101011001;
assign LUT_1[56718] = 32'b00000000000000001010000001101110;
assign LUT_1[56719] = 32'b00000000000000000011010011101010;
assign LUT_1[56720] = 32'b00000000000000001001000111110011;
assign LUT_1[56721] = 32'b00000000000000000010011001101111;
assign LUT_1[56722] = 32'b00000000000000000100110110000100;
assign LUT_1[56723] = 32'b11111111111111111110001000000000;
assign LUT_1[56724] = 32'b00000000000000010001000001001010;
assign LUT_1[56725] = 32'b00000000000000001010010011000110;
assign LUT_1[56726] = 32'b00000000000000001100101111011011;
assign LUT_1[56727] = 32'b00000000000000000110000001010111;
assign LUT_1[56728] = 32'b00000000000000001000010101101000;
assign LUT_1[56729] = 32'b00000000000000000001100111100100;
assign LUT_1[56730] = 32'b00000000000000000100000011111001;
assign LUT_1[56731] = 32'b11111111111111111101010101110101;
assign LUT_1[56732] = 32'b00000000000000010000001110111111;
assign LUT_1[56733] = 32'b00000000000000001001100000111011;
assign LUT_1[56734] = 32'b00000000000000001011111101010000;
assign LUT_1[56735] = 32'b00000000000000000101001111001100;
assign LUT_1[56736] = 32'b00000000000000001000000111010000;
assign LUT_1[56737] = 32'b00000000000000000001011001001100;
assign LUT_1[56738] = 32'b00000000000000000011110101100001;
assign LUT_1[56739] = 32'b11111111111111111101000111011101;
assign LUT_1[56740] = 32'b00000000000000010000000000100111;
assign LUT_1[56741] = 32'b00000000000000001001010010100011;
assign LUT_1[56742] = 32'b00000000000000001011101110111000;
assign LUT_1[56743] = 32'b00000000000000000101000000110100;
assign LUT_1[56744] = 32'b00000000000000000111010101000101;
assign LUT_1[56745] = 32'b00000000000000000000100111000001;
assign LUT_1[56746] = 32'b00000000000000000011000011010110;
assign LUT_1[56747] = 32'b11111111111111111100010101010010;
assign LUT_1[56748] = 32'b00000000000000001111001110011100;
assign LUT_1[56749] = 32'b00000000000000001000100000011000;
assign LUT_1[56750] = 32'b00000000000000001010111100101101;
assign LUT_1[56751] = 32'b00000000000000000100001110101001;
assign LUT_1[56752] = 32'b00000000000000001010000010110010;
assign LUT_1[56753] = 32'b00000000000000000011010100101110;
assign LUT_1[56754] = 32'b00000000000000000101110001000011;
assign LUT_1[56755] = 32'b11111111111111111111000010111111;
assign LUT_1[56756] = 32'b00000000000000010001111100001001;
assign LUT_1[56757] = 32'b00000000000000001011001110000101;
assign LUT_1[56758] = 32'b00000000000000001101101010011010;
assign LUT_1[56759] = 32'b00000000000000000110111100010110;
assign LUT_1[56760] = 32'b00000000000000001001010000100111;
assign LUT_1[56761] = 32'b00000000000000000010100010100011;
assign LUT_1[56762] = 32'b00000000000000000100111110111000;
assign LUT_1[56763] = 32'b11111111111111111110010000110100;
assign LUT_1[56764] = 32'b00000000000000010001001001111110;
assign LUT_1[56765] = 32'b00000000000000001010011011111010;
assign LUT_1[56766] = 32'b00000000000000001100111000001111;
assign LUT_1[56767] = 32'b00000000000000000110001010001011;
assign LUT_1[56768] = 32'b00000000000000001001001001111001;
assign LUT_1[56769] = 32'b00000000000000000010011011110101;
assign LUT_1[56770] = 32'b00000000000000000100111000001010;
assign LUT_1[56771] = 32'b11111111111111111110001010000110;
assign LUT_1[56772] = 32'b00000000000000010001000011010000;
assign LUT_1[56773] = 32'b00000000000000001010010101001100;
assign LUT_1[56774] = 32'b00000000000000001100110001100001;
assign LUT_1[56775] = 32'b00000000000000000110000011011101;
assign LUT_1[56776] = 32'b00000000000000001000010111101110;
assign LUT_1[56777] = 32'b00000000000000000001101001101010;
assign LUT_1[56778] = 32'b00000000000000000100000101111111;
assign LUT_1[56779] = 32'b11111111111111111101010111111011;
assign LUT_1[56780] = 32'b00000000000000010000010001000101;
assign LUT_1[56781] = 32'b00000000000000001001100011000001;
assign LUT_1[56782] = 32'b00000000000000001011111111010110;
assign LUT_1[56783] = 32'b00000000000000000101010001010010;
assign LUT_1[56784] = 32'b00000000000000001011000101011011;
assign LUT_1[56785] = 32'b00000000000000000100010111010111;
assign LUT_1[56786] = 32'b00000000000000000110110011101100;
assign LUT_1[56787] = 32'b00000000000000000000000101101000;
assign LUT_1[56788] = 32'b00000000000000010010111110110010;
assign LUT_1[56789] = 32'b00000000000000001100010000101110;
assign LUT_1[56790] = 32'b00000000000000001110101101000011;
assign LUT_1[56791] = 32'b00000000000000000111111110111111;
assign LUT_1[56792] = 32'b00000000000000001010010011010000;
assign LUT_1[56793] = 32'b00000000000000000011100101001100;
assign LUT_1[56794] = 32'b00000000000000000110000001100001;
assign LUT_1[56795] = 32'b11111111111111111111010011011101;
assign LUT_1[56796] = 32'b00000000000000010010001100100111;
assign LUT_1[56797] = 32'b00000000000000001011011110100011;
assign LUT_1[56798] = 32'b00000000000000001101111010111000;
assign LUT_1[56799] = 32'b00000000000000000111001100110100;
assign LUT_1[56800] = 32'b00000000000000001010000100111000;
assign LUT_1[56801] = 32'b00000000000000000011010110110100;
assign LUT_1[56802] = 32'b00000000000000000101110011001001;
assign LUT_1[56803] = 32'b11111111111111111111000101000101;
assign LUT_1[56804] = 32'b00000000000000010001111110001111;
assign LUT_1[56805] = 32'b00000000000000001011010000001011;
assign LUT_1[56806] = 32'b00000000000000001101101100100000;
assign LUT_1[56807] = 32'b00000000000000000110111110011100;
assign LUT_1[56808] = 32'b00000000000000001001010010101101;
assign LUT_1[56809] = 32'b00000000000000000010100100101001;
assign LUT_1[56810] = 32'b00000000000000000101000000111110;
assign LUT_1[56811] = 32'b11111111111111111110010010111010;
assign LUT_1[56812] = 32'b00000000000000010001001100000100;
assign LUT_1[56813] = 32'b00000000000000001010011110000000;
assign LUT_1[56814] = 32'b00000000000000001100111010010101;
assign LUT_1[56815] = 32'b00000000000000000110001100010001;
assign LUT_1[56816] = 32'b00000000000000001100000000011010;
assign LUT_1[56817] = 32'b00000000000000000101010010010110;
assign LUT_1[56818] = 32'b00000000000000000111101110101011;
assign LUT_1[56819] = 32'b00000000000000000001000000100111;
assign LUT_1[56820] = 32'b00000000000000010011111001110001;
assign LUT_1[56821] = 32'b00000000000000001101001011101101;
assign LUT_1[56822] = 32'b00000000000000001111101000000010;
assign LUT_1[56823] = 32'b00000000000000001000111001111110;
assign LUT_1[56824] = 32'b00000000000000001011001110001111;
assign LUT_1[56825] = 32'b00000000000000000100100000001011;
assign LUT_1[56826] = 32'b00000000000000000110111100100000;
assign LUT_1[56827] = 32'b00000000000000000000001110011100;
assign LUT_1[56828] = 32'b00000000000000010011000111100110;
assign LUT_1[56829] = 32'b00000000000000001100011001100010;
assign LUT_1[56830] = 32'b00000000000000001110110101110111;
assign LUT_1[56831] = 32'b00000000000000001000000111110011;
assign LUT_1[56832] = 32'b00000000000000000000000110011111;
assign LUT_1[56833] = 32'b11111111111111111001011000011011;
assign LUT_1[56834] = 32'b11111111111111111011110100110000;
assign LUT_1[56835] = 32'b11111111111111110101000110101100;
assign LUT_1[56836] = 32'b00000000000000000111111111110110;
assign LUT_1[56837] = 32'b00000000000000000001010001110010;
assign LUT_1[56838] = 32'b00000000000000000011101110000111;
assign LUT_1[56839] = 32'b11111111111111111101000000000011;
assign LUT_1[56840] = 32'b11111111111111111111010100010100;
assign LUT_1[56841] = 32'b11111111111111111000100110010000;
assign LUT_1[56842] = 32'b11111111111111111011000010100101;
assign LUT_1[56843] = 32'b11111111111111110100010100100001;
assign LUT_1[56844] = 32'b00000000000000000111001101101011;
assign LUT_1[56845] = 32'b00000000000000000000011111100111;
assign LUT_1[56846] = 32'b00000000000000000010111011111100;
assign LUT_1[56847] = 32'b11111111111111111100001101111000;
assign LUT_1[56848] = 32'b00000000000000000010000010000001;
assign LUT_1[56849] = 32'b11111111111111111011010011111101;
assign LUT_1[56850] = 32'b11111111111111111101110000010010;
assign LUT_1[56851] = 32'b11111111111111110111000010001110;
assign LUT_1[56852] = 32'b00000000000000001001111011011000;
assign LUT_1[56853] = 32'b00000000000000000011001101010100;
assign LUT_1[56854] = 32'b00000000000000000101101001101001;
assign LUT_1[56855] = 32'b11111111111111111110111011100101;
assign LUT_1[56856] = 32'b00000000000000000001001111110110;
assign LUT_1[56857] = 32'b11111111111111111010100001110010;
assign LUT_1[56858] = 32'b11111111111111111100111110000111;
assign LUT_1[56859] = 32'b11111111111111110110010000000011;
assign LUT_1[56860] = 32'b00000000000000001001001001001101;
assign LUT_1[56861] = 32'b00000000000000000010011011001001;
assign LUT_1[56862] = 32'b00000000000000000100110111011110;
assign LUT_1[56863] = 32'b11111111111111111110001001011010;
assign LUT_1[56864] = 32'b00000000000000000001000001011110;
assign LUT_1[56865] = 32'b11111111111111111010010011011010;
assign LUT_1[56866] = 32'b11111111111111111100101111101111;
assign LUT_1[56867] = 32'b11111111111111110110000001101011;
assign LUT_1[56868] = 32'b00000000000000001000111010110101;
assign LUT_1[56869] = 32'b00000000000000000010001100110001;
assign LUT_1[56870] = 32'b00000000000000000100101001000110;
assign LUT_1[56871] = 32'b11111111111111111101111011000010;
assign LUT_1[56872] = 32'b00000000000000000000001111010011;
assign LUT_1[56873] = 32'b11111111111111111001100001001111;
assign LUT_1[56874] = 32'b11111111111111111011111101100100;
assign LUT_1[56875] = 32'b11111111111111110101001111100000;
assign LUT_1[56876] = 32'b00000000000000001000001000101010;
assign LUT_1[56877] = 32'b00000000000000000001011010100110;
assign LUT_1[56878] = 32'b00000000000000000011110110111011;
assign LUT_1[56879] = 32'b11111111111111111101001000110111;
assign LUT_1[56880] = 32'b00000000000000000010111101000000;
assign LUT_1[56881] = 32'b11111111111111111100001110111100;
assign LUT_1[56882] = 32'b11111111111111111110101011010001;
assign LUT_1[56883] = 32'b11111111111111110111111101001101;
assign LUT_1[56884] = 32'b00000000000000001010110110010111;
assign LUT_1[56885] = 32'b00000000000000000100001000010011;
assign LUT_1[56886] = 32'b00000000000000000110100100101000;
assign LUT_1[56887] = 32'b11111111111111111111110110100100;
assign LUT_1[56888] = 32'b00000000000000000010001010110101;
assign LUT_1[56889] = 32'b11111111111111111011011100110001;
assign LUT_1[56890] = 32'b11111111111111111101111001000110;
assign LUT_1[56891] = 32'b11111111111111110111001011000010;
assign LUT_1[56892] = 32'b00000000000000001010000100001100;
assign LUT_1[56893] = 32'b00000000000000000011010110001000;
assign LUT_1[56894] = 32'b00000000000000000101110010011101;
assign LUT_1[56895] = 32'b11111111111111111111000100011001;
assign LUT_1[56896] = 32'b00000000000000000010000100000111;
assign LUT_1[56897] = 32'b11111111111111111011010110000011;
assign LUT_1[56898] = 32'b11111111111111111101110010011000;
assign LUT_1[56899] = 32'b11111111111111110111000100010100;
assign LUT_1[56900] = 32'b00000000000000001001111101011110;
assign LUT_1[56901] = 32'b00000000000000000011001111011010;
assign LUT_1[56902] = 32'b00000000000000000101101011101111;
assign LUT_1[56903] = 32'b11111111111111111110111101101011;
assign LUT_1[56904] = 32'b00000000000000000001010001111100;
assign LUT_1[56905] = 32'b11111111111111111010100011111000;
assign LUT_1[56906] = 32'b11111111111111111101000000001101;
assign LUT_1[56907] = 32'b11111111111111110110010010001001;
assign LUT_1[56908] = 32'b00000000000000001001001011010011;
assign LUT_1[56909] = 32'b00000000000000000010011101001111;
assign LUT_1[56910] = 32'b00000000000000000100111001100100;
assign LUT_1[56911] = 32'b11111111111111111110001011100000;
assign LUT_1[56912] = 32'b00000000000000000011111111101001;
assign LUT_1[56913] = 32'b11111111111111111101010001100101;
assign LUT_1[56914] = 32'b11111111111111111111101101111010;
assign LUT_1[56915] = 32'b11111111111111111000111111110110;
assign LUT_1[56916] = 32'b00000000000000001011111001000000;
assign LUT_1[56917] = 32'b00000000000000000101001010111100;
assign LUT_1[56918] = 32'b00000000000000000111100111010001;
assign LUT_1[56919] = 32'b00000000000000000000111001001101;
assign LUT_1[56920] = 32'b00000000000000000011001101011110;
assign LUT_1[56921] = 32'b11111111111111111100011111011010;
assign LUT_1[56922] = 32'b11111111111111111110111011101111;
assign LUT_1[56923] = 32'b11111111111111111000001101101011;
assign LUT_1[56924] = 32'b00000000000000001011000110110101;
assign LUT_1[56925] = 32'b00000000000000000100011000110001;
assign LUT_1[56926] = 32'b00000000000000000110110101000110;
assign LUT_1[56927] = 32'b00000000000000000000000111000010;
assign LUT_1[56928] = 32'b00000000000000000010111111000110;
assign LUT_1[56929] = 32'b11111111111111111100010001000010;
assign LUT_1[56930] = 32'b11111111111111111110101101010111;
assign LUT_1[56931] = 32'b11111111111111110111111111010011;
assign LUT_1[56932] = 32'b00000000000000001010111000011101;
assign LUT_1[56933] = 32'b00000000000000000100001010011001;
assign LUT_1[56934] = 32'b00000000000000000110100110101110;
assign LUT_1[56935] = 32'b11111111111111111111111000101010;
assign LUT_1[56936] = 32'b00000000000000000010001100111011;
assign LUT_1[56937] = 32'b11111111111111111011011110110111;
assign LUT_1[56938] = 32'b11111111111111111101111011001100;
assign LUT_1[56939] = 32'b11111111111111110111001101001000;
assign LUT_1[56940] = 32'b00000000000000001010000110010010;
assign LUT_1[56941] = 32'b00000000000000000011011000001110;
assign LUT_1[56942] = 32'b00000000000000000101110100100011;
assign LUT_1[56943] = 32'b11111111111111111111000110011111;
assign LUT_1[56944] = 32'b00000000000000000100111010101000;
assign LUT_1[56945] = 32'b11111111111111111110001100100100;
assign LUT_1[56946] = 32'b00000000000000000000101000111001;
assign LUT_1[56947] = 32'b11111111111111111001111010110101;
assign LUT_1[56948] = 32'b00000000000000001100110011111111;
assign LUT_1[56949] = 32'b00000000000000000110000101111011;
assign LUT_1[56950] = 32'b00000000000000001000100010010000;
assign LUT_1[56951] = 32'b00000000000000000001110100001100;
assign LUT_1[56952] = 32'b00000000000000000100001000011101;
assign LUT_1[56953] = 32'b11111111111111111101011010011001;
assign LUT_1[56954] = 32'b11111111111111111111110110101110;
assign LUT_1[56955] = 32'b11111111111111111001001000101010;
assign LUT_1[56956] = 32'b00000000000000001100000001110100;
assign LUT_1[56957] = 32'b00000000000000000101010011110000;
assign LUT_1[56958] = 32'b00000000000000000111110000000101;
assign LUT_1[56959] = 32'b00000000000000000001000010000001;
assign LUT_1[56960] = 32'b00000000000000000011000110100010;
assign LUT_1[56961] = 32'b11111111111111111100011000011110;
assign LUT_1[56962] = 32'b11111111111111111110110100110011;
assign LUT_1[56963] = 32'b11111111111111111000000110101111;
assign LUT_1[56964] = 32'b00000000000000001010111111111001;
assign LUT_1[56965] = 32'b00000000000000000100010001110101;
assign LUT_1[56966] = 32'b00000000000000000110101110001010;
assign LUT_1[56967] = 32'b00000000000000000000000000000110;
assign LUT_1[56968] = 32'b00000000000000000010010100010111;
assign LUT_1[56969] = 32'b11111111111111111011100110010011;
assign LUT_1[56970] = 32'b11111111111111111110000010101000;
assign LUT_1[56971] = 32'b11111111111111110111010100100100;
assign LUT_1[56972] = 32'b00000000000000001010001101101110;
assign LUT_1[56973] = 32'b00000000000000000011011111101010;
assign LUT_1[56974] = 32'b00000000000000000101111011111111;
assign LUT_1[56975] = 32'b11111111111111111111001101111011;
assign LUT_1[56976] = 32'b00000000000000000101000010000100;
assign LUT_1[56977] = 32'b11111111111111111110010100000000;
assign LUT_1[56978] = 32'b00000000000000000000110000010101;
assign LUT_1[56979] = 32'b11111111111111111010000010010001;
assign LUT_1[56980] = 32'b00000000000000001100111011011011;
assign LUT_1[56981] = 32'b00000000000000000110001101010111;
assign LUT_1[56982] = 32'b00000000000000001000101001101100;
assign LUT_1[56983] = 32'b00000000000000000001111011101000;
assign LUT_1[56984] = 32'b00000000000000000100001111111001;
assign LUT_1[56985] = 32'b11111111111111111101100001110101;
assign LUT_1[56986] = 32'b11111111111111111111111110001010;
assign LUT_1[56987] = 32'b11111111111111111001010000000110;
assign LUT_1[56988] = 32'b00000000000000001100001001010000;
assign LUT_1[56989] = 32'b00000000000000000101011011001100;
assign LUT_1[56990] = 32'b00000000000000000111110111100001;
assign LUT_1[56991] = 32'b00000000000000000001001001011101;
assign LUT_1[56992] = 32'b00000000000000000100000001100001;
assign LUT_1[56993] = 32'b11111111111111111101010011011101;
assign LUT_1[56994] = 32'b11111111111111111111101111110010;
assign LUT_1[56995] = 32'b11111111111111111001000001101110;
assign LUT_1[56996] = 32'b00000000000000001011111010111000;
assign LUT_1[56997] = 32'b00000000000000000101001100110100;
assign LUT_1[56998] = 32'b00000000000000000111101001001001;
assign LUT_1[56999] = 32'b00000000000000000000111011000101;
assign LUT_1[57000] = 32'b00000000000000000011001111010110;
assign LUT_1[57001] = 32'b11111111111111111100100001010010;
assign LUT_1[57002] = 32'b11111111111111111110111101100111;
assign LUT_1[57003] = 32'b11111111111111111000001111100011;
assign LUT_1[57004] = 32'b00000000000000001011001000101101;
assign LUT_1[57005] = 32'b00000000000000000100011010101001;
assign LUT_1[57006] = 32'b00000000000000000110110110111110;
assign LUT_1[57007] = 32'b00000000000000000000001000111010;
assign LUT_1[57008] = 32'b00000000000000000101111101000011;
assign LUT_1[57009] = 32'b11111111111111111111001110111111;
assign LUT_1[57010] = 32'b00000000000000000001101011010100;
assign LUT_1[57011] = 32'b11111111111111111010111101010000;
assign LUT_1[57012] = 32'b00000000000000001101110110011010;
assign LUT_1[57013] = 32'b00000000000000000111001000010110;
assign LUT_1[57014] = 32'b00000000000000001001100100101011;
assign LUT_1[57015] = 32'b00000000000000000010110110100111;
assign LUT_1[57016] = 32'b00000000000000000101001010111000;
assign LUT_1[57017] = 32'b11111111111111111110011100110100;
assign LUT_1[57018] = 32'b00000000000000000000111001001001;
assign LUT_1[57019] = 32'b11111111111111111010001011000101;
assign LUT_1[57020] = 32'b00000000000000001101000100001111;
assign LUT_1[57021] = 32'b00000000000000000110010110001011;
assign LUT_1[57022] = 32'b00000000000000001000110010100000;
assign LUT_1[57023] = 32'b00000000000000000010000100011100;
assign LUT_1[57024] = 32'b00000000000000000101000100001010;
assign LUT_1[57025] = 32'b11111111111111111110010110000110;
assign LUT_1[57026] = 32'b00000000000000000000110010011011;
assign LUT_1[57027] = 32'b11111111111111111010000100010111;
assign LUT_1[57028] = 32'b00000000000000001100111101100001;
assign LUT_1[57029] = 32'b00000000000000000110001111011101;
assign LUT_1[57030] = 32'b00000000000000001000101011110010;
assign LUT_1[57031] = 32'b00000000000000000001111101101110;
assign LUT_1[57032] = 32'b00000000000000000100010001111111;
assign LUT_1[57033] = 32'b11111111111111111101100011111011;
assign LUT_1[57034] = 32'b00000000000000000000000000010000;
assign LUT_1[57035] = 32'b11111111111111111001010010001100;
assign LUT_1[57036] = 32'b00000000000000001100001011010110;
assign LUT_1[57037] = 32'b00000000000000000101011101010010;
assign LUT_1[57038] = 32'b00000000000000000111111001100111;
assign LUT_1[57039] = 32'b00000000000000000001001011100011;
assign LUT_1[57040] = 32'b00000000000000000110111111101100;
assign LUT_1[57041] = 32'b00000000000000000000010001101000;
assign LUT_1[57042] = 32'b00000000000000000010101101111101;
assign LUT_1[57043] = 32'b11111111111111111011111111111001;
assign LUT_1[57044] = 32'b00000000000000001110111001000011;
assign LUT_1[57045] = 32'b00000000000000001000001010111111;
assign LUT_1[57046] = 32'b00000000000000001010100111010100;
assign LUT_1[57047] = 32'b00000000000000000011111001010000;
assign LUT_1[57048] = 32'b00000000000000000110001101100001;
assign LUT_1[57049] = 32'b11111111111111111111011111011101;
assign LUT_1[57050] = 32'b00000000000000000001111011110010;
assign LUT_1[57051] = 32'b11111111111111111011001101101110;
assign LUT_1[57052] = 32'b00000000000000001110000110111000;
assign LUT_1[57053] = 32'b00000000000000000111011000110100;
assign LUT_1[57054] = 32'b00000000000000001001110101001001;
assign LUT_1[57055] = 32'b00000000000000000011000111000101;
assign LUT_1[57056] = 32'b00000000000000000101111111001001;
assign LUT_1[57057] = 32'b11111111111111111111010001000101;
assign LUT_1[57058] = 32'b00000000000000000001101101011010;
assign LUT_1[57059] = 32'b11111111111111111010111111010110;
assign LUT_1[57060] = 32'b00000000000000001101111000100000;
assign LUT_1[57061] = 32'b00000000000000000111001010011100;
assign LUT_1[57062] = 32'b00000000000000001001100110110001;
assign LUT_1[57063] = 32'b00000000000000000010111000101101;
assign LUT_1[57064] = 32'b00000000000000000101001100111110;
assign LUT_1[57065] = 32'b11111111111111111110011110111010;
assign LUT_1[57066] = 32'b00000000000000000000111011001111;
assign LUT_1[57067] = 32'b11111111111111111010001101001011;
assign LUT_1[57068] = 32'b00000000000000001101000110010101;
assign LUT_1[57069] = 32'b00000000000000000110011000010001;
assign LUT_1[57070] = 32'b00000000000000001000110100100110;
assign LUT_1[57071] = 32'b00000000000000000010000110100010;
assign LUT_1[57072] = 32'b00000000000000000111111010101011;
assign LUT_1[57073] = 32'b00000000000000000001001100100111;
assign LUT_1[57074] = 32'b00000000000000000011101000111100;
assign LUT_1[57075] = 32'b11111111111111111100111010111000;
assign LUT_1[57076] = 32'b00000000000000001111110100000010;
assign LUT_1[57077] = 32'b00000000000000001001000101111110;
assign LUT_1[57078] = 32'b00000000000000001011100010010011;
assign LUT_1[57079] = 32'b00000000000000000100110100001111;
assign LUT_1[57080] = 32'b00000000000000000111001000100000;
assign LUT_1[57081] = 32'b00000000000000000000011010011100;
assign LUT_1[57082] = 32'b00000000000000000010110110110001;
assign LUT_1[57083] = 32'b11111111111111111100001000101101;
assign LUT_1[57084] = 32'b00000000000000001111000001110111;
assign LUT_1[57085] = 32'b00000000000000001000010011110011;
assign LUT_1[57086] = 32'b00000000000000001010110000001000;
assign LUT_1[57087] = 32'b00000000000000000100000010000100;
assign LUT_1[57088] = 32'b11111111111111111101111010101011;
assign LUT_1[57089] = 32'b11111111111111110111001100100111;
assign LUT_1[57090] = 32'b11111111111111111001101000111100;
assign LUT_1[57091] = 32'b11111111111111110010111010111000;
assign LUT_1[57092] = 32'b00000000000000000101110100000010;
assign LUT_1[57093] = 32'b11111111111111111111000101111110;
assign LUT_1[57094] = 32'b00000000000000000001100010010011;
assign LUT_1[57095] = 32'b11111111111111111010110100001111;
assign LUT_1[57096] = 32'b11111111111111111101001000100000;
assign LUT_1[57097] = 32'b11111111111111110110011010011100;
assign LUT_1[57098] = 32'b11111111111111111000110110110001;
assign LUT_1[57099] = 32'b11111111111111110010001000101101;
assign LUT_1[57100] = 32'b00000000000000000101000001110111;
assign LUT_1[57101] = 32'b11111111111111111110010011110011;
assign LUT_1[57102] = 32'b00000000000000000000110000001000;
assign LUT_1[57103] = 32'b11111111111111111010000010000100;
assign LUT_1[57104] = 32'b11111111111111111111110110001101;
assign LUT_1[57105] = 32'b11111111111111111001001000001001;
assign LUT_1[57106] = 32'b11111111111111111011100100011110;
assign LUT_1[57107] = 32'b11111111111111110100110110011010;
assign LUT_1[57108] = 32'b00000000000000000111101111100100;
assign LUT_1[57109] = 32'b00000000000000000001000001100000;
assign LUT_1[57110] = 32'b00000000000000000011011101110101;
assign LUT_1[57111] = 32'b11111111111111111100101111110001;
assign LUT_1[57112] = 32'b11111111111111111111000100000010;
assign LUT_1[57113] = 32'b11111111111111111000010101111110;
assign LUT_1[57114] = 32'b11111111111111111010110010010011;
assign LUT_1[57115] = 32'b11111111111111110100000100001111;
assign LUT_1[57116] = 32'b00000000000000000110111101011001;
assign LUT_1[57117] = 32'b00000000000000000000001111010101;
assign LUT_1[57118] = 32'b00000000000000000010101011101010;
assign LUT_1[57119] = 32'b11111111111111111011111101100110;
assign LUT_1[57120] = 32'b11111111111111111110110101101010;
assign LUT_1[57121] = 32'b11111111111111111000000111100110;
assign LUT_1[57122] = 32'b11111111111111111010100011111011;
assign LUT_1[57123] = 32'b11111111111111110011110101110111;
assign LUT_1[57124] = 32'b00000000000000000110101111000001;
assign LUT_1[57125] = 32'b00000000000000000000000000111101;
assign LUT_1[57126] = 32'b00000000000000000010011101010010;
assign LUT_1[57127] = 32'b11111111111111111011101111001110;
assign LUT_1[57128] = 32'b11111111111111111110000011011111;
assign LUT_1[57129] = 32'b11111111111111110111010101011011;
assign LUT_1[57130] = 32'b11111111111111111001110001110000;
assign LUT_1[57131] = 32'b11111111111111110011000011101100;
assign LUT_1[57132] = 32'b00000000000000000101111100110110;
assign LUT_1[57133] = 32'b11111111111111111111001110110010;
assign LUT_1[57134] = 32'b00000000000000000001101011000111;
assign LUT_1[57135] = 32'b11111111111111111010111101000011;
assign LUT_1[57136] = 32'b00000000000000000000110001001100;
assign LUT_1[57137] = 32'b11111111111111111010000011001000;
assign LUT_1[57138] = 32'b11111111111111111100011111011101;
assign LUT_1[57139] = 32'b11111111111111110101110001011001;
assign LUT_1[57140] = 32'b00000000000000001000101010100011;
assign LUT_1[57141] = 32'b00000000000000000001111100011111;
assign LUT_1[57142] = 32'b00000000000000000100011000110100;
assign LUT_1[57143] = 32'b11111111111111111101101010110000;
assign LUT_1[57144] = 32'b11111111111111111111111111000001;
assign LUT_1[57145] = 32'b11111111111111111001010000111101;
assign LUT_1[57146] = 32'b11111111111111111011101101010010;
assign LUT_1[57147] = 32'b11111111111111110100111111001110;
assign LUT_1[57148] = 32'b00000000000000000111111000011000;
assign LUT_1[57149] = 32'b00000000000000000001001010010100;
assign LUT_1[57150] = 32'b00000000000000000011100110101001;
assign LUT_1[57151] = 32'b11111111111111111100111000100101;
assign LUT_1[57152] = 32'b11111111111111111111111000010011;
assign LUT_1[57153] = 32'b11111111111111111001001010001111;
assign LUT_1[57154] = 32'b11111111111111111011100110100100;
assign LUT_1[57155] = 32'b11111111111111110100111000100000;
assign LUT_1[57156] = 32'b00000000000000000111110001101010;
assign LUT_1[57157] = 32'b00000000000000000001000011100110;
assign LUT_1[57158] = 32'b00000000000000000011011111111011;
assign LUT_1[57159] = 32'b11111111111111111100110001110111;
assign LUT_1[57160] = 32'b11111111111111111111000110001000;
assign LUT_1[57161] = 32'b11111111111111111000011000000100;
assign LUT_1[57162] = 32'b11111111111111111010110100011001;
assign LUT_1[57163] = 32'b11111111111111110100000110010101;
assign LUT_1[57164] = 32'b00000000000000000110111111011111;
assign LUT_1[57165] = 32'b00000000000000000000010001011011;
assign LUT_1[57166] = 32'b00000000000000000010101101110000;
assign LUT_1[57167] = 32'b11111111111111111011111111101100;
assign LUT_1[57168] = 32'b00000000000000000001110011110101;
assign LUT_1[57169] = 32'b11111111111111111011000101110001;
assign LUT_1[57170] = 32'b11111111111111111101100010000110;
assign LUT_1[57171] = 32'b11111111111111110110110100000010;
assign LUT_1[57172] = 32'b00000000000000001001101101001100;
assign LUT_1[57173] = 32'b00000000000000000010111111001000;
assign LUT_1[57174] = 32'b00000000000000000101011011011101;
assign LUT_1[57175] = 32'b11111111111111111110101101011001;
assign LUT_1[57176] = 32'b00000000000000000001000001101010;
assign LUT_1[57177] = 32'b11111111111111111010010011100110;
assign LUT_1[57178] = 32'b11111111111111111100101111111011;
assign LUT_1[57179] = 32'b11111111111111110110000001110111;
assign LUT_1[57180] = 32'b00000000000000001000111011000001;
assign LUT_1[57181] = 32'b00000000000000000010001100111101;
assign LUT_1[57182] = 32'b00000000000000000100101001010010;
assign LUT_1[57183] = 32'b11111111111111111101111011001110;
assign LUT_1[57184] = 32'b00000000000000000000110011010010;
assign LUT_1[57185] = 32'b11111111111111111010000101001110;
assign LUT_1[57186] = 32'b11111111111111111100100001100011;
assign LUT_1[57187] = 32'b11111111111111110101110011011111;
assign LUT_1[57188] = 32'b00000000000000001000101100101001;
assign LUT_1[57189] = 32'b00000000000000000001111110100101;
assign LUT_1[57190] = 32'b00000000000000000100011010111010;
assign LUT_1[57191] = 32'b11111111111111111101101100110110;
assign LUT_1[57192] = 32'b00000000000000000000000001000111;
assign LUT_1[57193] = 32'b11111111111111111001010011000011;
assign LUT_1[57194] = 32'b11111111111111111011101111011000;
assign LUT_1[57195] = 32'b11111111111111110101000001010100;
assign LUT_1[57196] = 32'b00000000000000000111111010011110;
assign LUT_1[57197] = 32'b00000000000000000001001100011010;
assign LUT_1[57198] = 32'b00000000000000000011101000101111;
assign LUT_1[57199] = 32'b11111111111111111100111010101011;
assign LUT_1[57200] = 32'b00000000000000000010101110110100;
assign LUT_1[57201] = 32'b11111111111111111100000000110000;
assign LUT_1[57202] = 32'b11111111111111111110011101000101;
assign LUT_1[57203] = 32'b11111111111111110111101111000001;
assign LUT_1[57204] = 32'b00000000000000001010101000001011;
assign LUT_1[57205] = 32'b00000000000000000011111010000111;
assign LUT_1[57206] = 32'b00000000000000000110010110011100;
assign LUT_1[57207] = 32'b11111111111111111111101000011000;
assign LUT_1[57208] = 32'b00000000000000000001111100101001;
assign LUT_1[57209] = 32'b11111111111111111011001110100101;
assign LUT_1[57210] = 32'b11111111111111111101101010111010;
assign LUT_1[57211] = 32'b11111111111111110110111100110110;
assign LUT_1[57212] = 32'b00000000000000001001110110000000;
assign LUT_1[57213] = 32'b00000000000000000011000111111100;
assign LUT_1[57214] = 32'b00000000000000000101100100010001;
assign LUT_1[57215] = 32'b11111111111111111110110110001101;
assign LUT_1[57216] = 32'b00000000000000000000111010101110;
assign LUT_1[57217] = 32'b11111111111111111010001100101010;
assign LUT_1[57218] = 32'b11111111111111111100101000111111;
assign LUT_1[57219] = 32'b11111111111111110101111010111011;
assign LUT_1[57220] = 32'b00000000000000001000110100000101;
assign LUT_1[57221] = 32'b00000000000000000010000110000001;
assign LUT_1[57222] = 32'b00000000000000000100100010010110;
assign LUT_1[57223] = 32'b11111111111111111101110100010010;
assign LUT_1[57224] = 32'b00000000000000000000001000100011;
assign LUT_1[57225] = 32'b11111111111111111001011010011111;
assign LUT_1[57226] = 32'b11111111111111111011110110110100;
assign LUT_1[57227] = 32'b11111111111111110101001000110000;
assign LUT_1[57228] = 32'b00000000000000001000000001111010;
assign LUT_1[57229] = 32'b00000000000000000001010011110110;
assign LUT_1[57230] = 32'b00000000000000000011110000001011;
assign LUT_1[57231] = 32'b11111111111111111101000010000111;
assign LUT_1[57232] = 32'b00000000000000000010110110010000;
assign LUT_1[57233] = 32'b11111111111111111100001000001100;
assign LUT_1[57234] = 32'b11111111111111111110100100100001;
assign LUT_1[57235] = 32'b11111111111111110111110110011101;
assign LUT_1[57236] = 32'b00000000000000001010101111100111;
assign LUT_1[57237] = 32'b00000000000000000100000001100011;
assign LUT_1[57238] = 32'b00000000000000000110011101111000;
assign LUT_1[57239] = 32'b11111111111111111111101111110100;
assign LUT_1[57240] = 32'b00000000000000000010000100000101;
assign LUT_1[57241] = 32'b11111111111111111011010110000001;
assign LUT_1[57242] = 32'b11111111111111111101110010010110;
assign LUT_1[57243] = 32'b11111111111111110111000100010010;
assign LUT_1[57244] = 32'b00000000000000001001111101011100;
assign LUT_1[57245] = 32'b00000000000000000011001111011000;
assign LUT_1[57246] = 32'b00000000000000000101101011101101;
assign LUT_1[57247] = 32'b11111111111111111110111101101001;
assign LUT_1[57248] = 32'b00000000000000000001110101101101;
assign LUT_1[57249] = 32'b11111111111111111011000111101001;
assign LUT_1[57250] = 32'b11111111111111111101100011111110;
assign LUT_1[57251] = 32'b11111111111111110110110101111010;
assign LUT_1[57252] = 32'b00000000000000001001101111000100;
assign LUT_1[57253] = 32'b00000000000000000011000001000000;
assign LUT_1[57254] = 32'b00000000000000000101011101010101;
assign LUT_1[57255] = 32'b11111111111111111110101111010001;
assign LUT_1[57256] = 32'b00000000000000000001000011100010;
assign LUT_1[57257] = 32'b11111111111111111010010101011110;
assign LUT_1[57258] = 32'b11111111111111111100110001110011;
assign LUT_1[57259] = 32'b11111111111111110110000011101111;
assign LUT_1[57260] = 32'b00000000000000001000111100111001;
assign LUT_1[57261] = 32'b00000000000000000010001110110101;
assign LUT_1[57262] = 32'b00000000000000000100101011001010;
assign LUT_1[57263] = 32'b11111111111111111101111101000110;
assign LUT_1[57264] = 32'b00000000000000000011110001001111;
assign LUT_1[57265] = 32'b11111111111111111101000011001011;
assign LUT_1[57266] = 32'b11111111111111111111011111100000;
assign LUT_1[57267] = 32'b11111111111111111000110001011100;
assign LUT_1[57268] = 32'b00000000000000001011101010100110;
assign LUT_1[57269] = 32'b00000000000000000100111100100010;
assign LUT_1[57270] = 32'b00000000000000000111011000110111;
assign LUT_1[57271] = 32'b00000000000000000000101010110011;
assign LUT_1[57272] = 32'b00000000000000000010111111000100;
assign LUT_1[57273] = 32'b11111111111111111100010001000000;
assign LUT_1[57274] = 32'b11111111111111111110101101010101;
assign LUT_1[57275] = 32'b11111111111111110111111111010001;
assign LUT_1[57276] = 32'b00000000000000001010111000011011;
assign LUT_1[57277] = 32'b00000000000000000100001010010111;
assign LUT_1[57278] = 32'b00000000000000000110100110101100;
assign LUT_1[57279] = 32'b11111111111111111111111000101000;
assign LUT_1[57280] = 32'b00000000000000000010111000010110;
assign LUT_1[57281] = 32'b11111111111111111100001010010010;
assign LUT_1[57282] = 32'b11111111111111111110100110100111;
assign LUT_1[57283] = 32'b11111111111111110111111000100011;
assign LUT_1[57284] = 32'b00000000000000001010110001101101;
assign LUT_1[57285] = 32'b00000000000000000100000011101001;
assign LUT_1[57286] = 32'b00000000000000000110011111111110;
assign LUT_1[57287] = 32'b11111111111111111111110001111010;
assign LUT_1[57288] = 32'b00000000000000000010000110001011;
assign LUT_1[57289] = 32'b11111111111111111011011000000111;
assign LUT_1[57290] = 32'b11111111111111111101110100011100;
assign LUT_1[57291] = 32'b11111111111111110111000110011000;
assign LUT_1[57292] = 32'b00000000000000001001111111100010;
assign LUT_1[57293] = 32'b00000000000000000011010001011110;
assign LUT_1[57294] = 32'b00000000000000000101101101110011;
assign LUT_1[57295] = 32'b11111111111111111110111111101111;
assign LUT_1[57296] = 32'b00000000000000000100110011111000;
assign LUT_1[57297] = 32'b11111111111111111110000101110100;
assign LUT_1[57298] = 32'b00000000000000000000100010001001;
assign LUT_1[57299] = 32'b11111111111111111001110100000101;
assign LUT_1[57300] = 32'b00000000000000001100101101001111;
assign LUT_1[57301] = 32'b00000000000000000101111111001011;
assign LUT_1[57302] = 32'b00000000000000001000011011100000;
assign LUT_1[57303] = 32'b00000000000000000001101101011100;
assign LUT_1[57304] = 32'b00000000000000000100000001101101;
assign LUT_1[57305] = 32'b11111111111111111101010011101001;
assign LUT_1[57306] = 32'b11111111111111111111101111111110;
assign LUT_1[57307] = 32'b11111111111111111001000001111010;
assign LUT_1[57308] = 32'b00000000000000001011111011000100;
assign LUT_1[57309] = 32'b00000000000000000101001101000000;
assign LUT_1[57310] = 32'b00000000000000000111101001010101;
assign LUT_1[57311] = 32'b00000000000000000000111011010001;
assign LUT_1[57312] = 32'b00000000000000000011110011010101;
assign LUT_1[57313] = 32'b11111111111111111101000101010001;
assign LUT_1[57314] = 32'b11111111111111111111100001100110;
assign LUT_1[57315] = 32'b11111111111111111000110011100010;
assign LUT_1[57316] = 32'b00000000000000001011101100101100;
assign LUT_1[57317] = 32'b00000000000000000100111110101000;
assign LUT_1[57318] = 32'b00000000000000000111011010111101;
assign LUT_1[57319] = 32'b00000000000000000000101100111001;
assign LUT_1[57320] = 32'b00000000000000000011000001001010;
assign LUT_1[57321] = 32'b11111111111111111100010011000110;
assign LUT_1[57322] = 32'b11111111111111111110101111011011;
assign LUT_1[57323] = 32'b11111111111111111000000001010111;
assign LUT_1[57324] = 32'b00000000000000001010111010100001;
assign LUT_1[57325] = 32'b00000000000000000100001100011101;
assign LUT_1[57326] = 32'b00000000000000000110101000110010;
assign LUT_1[57327] = 32'b11111111111111111111111010101110;
assign LUT_1[57328] = 32'b00000000000000000101101110110111;
assign LUT_1[57329] = 32'b11111111111111111111000000110011;
assign LUT_1[57330] = 32'b00000000000000000001011101001000;
assign LUT_1[57331] = 32'b11111111111111111010101111000100;
assign LUT_1[57332] = 32'b00000000000000001101101000001110;
assign LUT_1[57333] = 32'b00000000000000000110111010001010;
assign LUT_1[57334] = 32'b00000000000000001001010110011111;
assign LUT_1[57335] = 32'b00000000000000000010101000011011;
assign LUT_1[57336] = 32'b00000000000000000100111100101100;
assign LUT_1[57337] = 32'b11111111111111111110001110101000;
assign LUT_1[57338] = 32'b00000000000000000000101010111101;
assign LUT_1[57339] = 32'b11111111111111111001111100111001;
assign LUT_1[57340] = 32'b00000000000000001100110110000011;
assign LUT_1[57341] = 32'b00000000000000000110000111111111;
assign LUT_1[57342] = 32'b00000000000000001000100100010100;
assign LUT_1[57343] = 32'b00000000000000000001110110010000;
assign LUT_1[57344] = 32'b00000000000000000010010010110100;
assign LUT_1[57345] = 32'b11111111111111111011100100110000;
assign LUT_1[57346] = 32'b11111111111111111110000001000101;
assign LUT_1[57347] = 32'b11111111111111110111010011000001;
assign LUT_1[57348] = 32'b00000000000000001010001100001011;
assign LUT_1[57349] = 32'b00000000000000000011011110000111;
assign LUT_1[57350] = 32'b00000000000000000101111010011100;
assign LUT_1[57351] = 32'b11111111111111111111001100011000;
assign LUT_1[57352] = 32'b00000000000000000001100000101001;
assign LUT_1[57353] = 32'b11111111111111111010110010100101;
assign LUT_1[57354] = 32'b11111111111111111101001110111010;
assign LUT_1[57355] = 32'b11111111111111110110100000110110;
assign LUT_1[57356] = 32'b00000000000000001001011010000000;
assign LUT_1[57357] = 32'b00000000000000000010101011111100;
assign LUT_1[57358] = 32'b00000000000000000101001000010001;
assign LUT_1[57359] = 32'b11111111111111111110011010001101;
assign LUT_1[57360] = 32'b00000000000000000100001110010110;
assign LUT_1[57361] = 32'b11111111111111111101100000010010;
assign LUT_1[57362] = 32'b11111111111111111111111100100111;
assign LUT_1[57363] = 32'b11111111111111111001001110100011;
assign LUT_1[57364] = 32'b00000000000000001100000111101101;
assign LUT_1[57365] = 32'b00000000000000000101011001101001;
assign LUT_1[57366] = 32'b00000000000000000111110101111110;
assign LUT_1[57367] = 32'b00000000000000000001000111111010;
assign LUT_1[57368] = 32'b00000000000000000011011100001011;
assign LUT_1[57369] = 32'b11111111111111111100101110000111;
assign LUT_1[57370] = 32'b11111111111111111111001010011100;
assign LUT_1[57371] = 32'b11111111111111111000011100011000;
assign LUT_1[57372] = 32'b00000000000000001011010101100010;
assign LUT_1[57373] = 32'b00000000000000000100100111011110;
assign LUT_1[57374] = 32'b00000000000000000111000011110011;
assign LUT_1[57375] = 32'b00000000000000000000010101101111;
assign LUT_1[57376] = 32'b00000000000000000011001101110011;
assign LUT_1[57377] = 32'b11111111111111111100011111101111;
assign LUT_1[57378] = 32'b11111111111111111110111100000100;
assign LUT_1[57379] = 32'b11111111111111111000001110000000;
assign LUT_1[57380] = 32'b00000000000000001011000111001010;
assign LUT_1[57381] = 32'b00000000000000000100011001000110;
assign LUT_1[57382] = 32'b00000000000000000110110101011011;
assign LUT_1[57383] = 32'b00000000000000000000000111010111;
assign LUT_1[57384] = 32'b00000000000000000010011011101000;
assign LUT_1[57385] = 32'b11111111111111111011101101100100;
assign LUT_1[57386] = 32'b11111111111111111110001001111001;
assign LUT_1[57387] = 32'b11111111111111110111011011110101;
assign LUT_1[57388] = 32'b00000000000000001010010100111111;
assign LUT_1[57389] = 32'b00000000000000000011100110111011;
assign LUT_1[57390] = 32'b00000000000000000110000011010000;
assign LUT_1[57391] = 32'b11111111111111111111010101001100;
assign LUT_1[57392] = 32'b00000000000000000101001001010101;
assign LUT_1[57393] = 32'b11111111111111111110011011010001;
assign LUT_1[57394] = 32'b00000000000000000000110111100110;
assign LUT_1[57395] = 32'b11111111111111111010001001100010;
assign LUT_1[57396] = 32'b00000000000000001101000010101100;
assign LUT_1[57397] = 32'b00000000000000000110010100101000;
assign LUT_1[57398] = 32'b00000000000000001000110000111101;
assign LUT_1[57399] = 32'b00000000000000000010000010111001;
assign LUT_1[57400] = 32'b00000000000000000100010111001010;
assign LUT_1[57401] = 32'b11111111111111111101101001000110;
assign LUT_1[57402] = 32'b00000000000000000000000101011011;
assign LUT_1[57403] = 32'b11111111111111111001010111010111;
assign LUT_1[57404] = 32'b00000000000000001100010000100001;
assign LUT_1[57405] = 32'b00000000000000000101100010011101;
assign LUT_1[57406] = 32'b00000000000000000111111110110010;
assign LUT_1[57407] = 32'b00000000000000000001010000101110;
assign LUT_1[57408] = 32'b00000000000000000100010000011100;
assign LUT_1[57409] = 32'b11111111111111111101100010011000;
assign LUT_1[57410] = 32'b11111111111111111111111110101101;
assign LUT_1[57411] = 32'b11111111111111111001010000101001;
assign LUT_1[57412] = 32'b00000000000000001100001001110011;
assign LUT_1[57413] = 32'b00000000000000000101011011101111;
assign LUT_1[57414] = 32'b00000000000000000111111000000100;
assign LUT_1[57415] = 32'b00000000000000000001001010000000;
assign LUT_1[57416] = 32'b00000000000000000011011110010001;
assign LUT_1[57417] = 32'b11111111111111111100110000001101;
assign LUT_1[57418] = 32'b11111111111111111111001100100010;
assign LUT_1[57419] = 32'b11111111111111111000011110011110;
assign LUT_1[57420] = 32'b00000000000000001011010111101000;
assign LUT_1[57421] = 32'b00000000000000000100101001100100;
assign LUT_1[57422] = 32'b00000000000000000111000101111001;
assign LUT_1[57423] = 32'b00000000000000000000010111110101;
assign LUT_1[57424] = 32'b00000000000000000110001011111110;
assign LUT_1[57425] = 32'b11111111111111111111011101111010;
assign LUT_1[57426] = 32'b00000000000000000001111010001111;
assign LUT_1[57427] = 32'b11111111111111111011001100001011;
assign LUT_1[57428] = 32'b00000000000000001110000101010101;
assign LUT_1[57429] = 32'b00000000000000000111010111010001;
assign LUT_1[57430] = 32'b00000000000000001001110011100110;
assign LUT_1[57431] = 32'b00000000000000000011000101100010;
assign LUT_1[57432] = 32'b00000000000000000101011001110011;
assign LUT_1[57433] = 32'b11111111111111111110101011101111;
assign LUT_1[57434] = 32'b00000000000000000001001000000100;
assign LUT_1[57435] = 32'b11111111111111111010011010000000;
assign LUT_1[57436] = 32'b00000000000000001101010011001010;
assign LUT_1[57437] = 32'b00000000000000000110100101000110;
assign LUT_1[57438] = 32'b00000000000000001001000001011011;
assign LUT_1[57439] = 32'b00000000000000000010010011010111;
assign LUT_1[57440] = 32'b00000000000000000101001011011011;
assign LUT_1[57441] = 32'b11111111111111111110011101010111;
assign LUT_1[57442] = 32'b00000000000000000000111001101100;
assign LUT_1[57443] = 32'b11111111111111111010001011101000;
assign LUT_1[57444] = 32'b00000000000000001101000100110010;
assign LUT_1[57445] = 32'b00000000000000000110010110101110;
assign LUT_1[57446] = 32'b00000000000000001000110011000011;
assign LUT_1[57447] = 32'b00000000000000000010000100111111;
assign LUT_1[57448] = 32'b00000000000000000100011001010000;
assign LUT_1[57449] = 32'b11111111111111111101101011001100;
assign LUT_1[57450] = 32'b00000000000000000000000111100001;
assign LUT_1[57451] = 32'b11111111111111111001011001011101;
assign LUT_1[57452] = 32'b00000000000000001100010010100111;
assign LUT_1[57453] = 32'b00000000000000000101100100100011;
assign LUT_1[57454] = 32'b00000000000000001000000000111000;
assign LUT_1[57455] = 32'b00000000000000000001010010110100;
assign LUT_1[57456] = 32'b00000000000000000111000110111101;
assign LUT_1[57457] = 32'b00000000000000000000011000111001;
assign LUT_1[57458] = 32'b00000000000000000010110101001110;
assign LUT_1[57459] = 32'b11111111111111111100000111001010;
assign LUT_1[57460] = 32'b00000000000000001111000000010100;
assign LUT_1[57461] = 32'b00000000000000001000010010010000;
assign LUT_1[57462] = 32'b00000000000000001010101110100101;
assign LUT_1[57463] = 32'b00000000000000000100000000100001;
assign LUT_1[57464] = 32'b00000000000000000110010100110010;
assign LUT_1[57465] = 32'b11111111111111111111100110101110;
assign LUT_1[57466] = 32'b00000000000000000010000011000011;
assign LUT_1[57467] = 32'b11111111111111111011010100111111;
assign LUT_1[57468] = 32'b00000000000000001110001110001001;
assign LUT_1[57469] = 32'b00000000000000000111100000000101;
assign LUT_1[57470] = 32'b00000000000000001001111100011010;
assign LUT_1[57471] = 32'b00000000000000000011001110010110;
assign LUT_1[57472] = 32'b00000000000000000101010010110111;
assign LUT_1[57473] = 32'b11111111111111111110100100110011;
assign LUT_1[57474] = 32'b00000000000000000001000001001000;
assign LUT_1[57475] = 32'b11111111111111111010010011000100;
assign LUT_1[57476] = 32'b00000000000000001101001100001110;
assign LUT_1[57477] = 32'b00000000000000000110011110001010;
assign LUT_1[57478] = 32'b00000000000000001000111010011111;
assign LUT_1[57479] = 32'b00000000000000000010001100011011;
assign LUT_1[57480] = 32'b00000000000000000100100000101100;
assign LUT_1[57481] = 32'b11111111111111111101110010101000;
assign LUT_1[57482] = 32'b00000000000000000000001110111101;
assign LUT_1[57483] = 32'b11111111111111111001100000111001;
assign LUT_1[57484] = 32'b00000000000000001100011010000011;
assign LUT_1[57485] = 32'b00000000000000000101101011111111;
assign LUT_1[57486] = 32'b00000000000000001000001000010100;
assign LUT_1[57487] = 32'b00000000000000000001011010010000;
assign LUT_1[57488] = 32'b00000000000000000111001110011001;
assign LUT_1[57489] = 32'b00000000000000000000100000010101;
assign LUT_1[57490] = 32'b00000000000000000010111100101010;
assign LUT_1[57491] = 32'b11111111111111111100001110100110;
assign LUT_1[57492] = 32'b00000000000000001111000111110000;
assign LUT_1[57493] = 32'b00000000000000001000011001101100;
assign LUT_1[57494] = 32'b00000000000000001010110110000001;
assign LUT_1[57495] = 32'b00000000000000000100000111111101;
assign LUT_1[57496] = 32'b00000000000000000110011100001110;
assign LUT_1[57497] = 32'b11111111111111111111101110001010;
assign LUT_1[57498] = 32'b00000000000000000010001010011111;
assign LUT_1[57499] = 32'b11111111111111111011011100011011;
assign LUT_1[57500] = 32'b00000000000000001110010101100101;
assign LUT_1[57501] = 32'b00000000000000000111100111100001;
assign LUT_1[57502] = 32'b00000000000000001010000011110110;
assign LUT_1[57503] = 32'b00000000000000000011010101110010;
assign LUT_1[57504] = 32'b00000000000000000110001101110110;
assign LUT_1[57505] = 32'b11111111111111111111011111110010;
assign LUT_1[57506] = 32'b00000000000000000001111100000111;
assign LUT_1[57507] = 32'b11111111111111111011001110000011;
assign LUT_1[57508] = 32'b00000000000000001110000111001101;
assign LUT_1[57509] = 32'b00000000000000000111011001001001;
assign LUT_1[57510] = 32'b00000000000000001001110101011110;
assign LUT_1[57511] = 32'b00000000000000000011000111011010;
assign LUT_1[57512] = 32'b00000000000000000101011011101011;
assign LUT_1[57513] = 32'b11111111111111111110101101100111;
assign LUT_1[57514] = 32'b00000000000000000001001001111100;
assign LUT_1[57515] = 32'b11111111111111111010011011111000;
assign LUT_1[57516] = 32'b00000000000000001101010101000010;
assign LUT_1[57517] = 32'b00000000000000000110100110111110;
assign LUT_1[57518] = 32'b00000000000000001001000011010011;
assign LUT_1[57519] = 32'b00000000000000000010010101001111;
assign LUT_1[57520] = 32'b00000000000000001000001001011000;
assign LUT_1[57521] = 32'b00000000000000000001011011010100;
assign LUT_1[57522] = 32'b00000000000000000011110111101001;
assign LUT_1[57523] = 32'b11111111111111111101001001100101;
assign LUT_1[57524] = 32'b00000000000000010000000010101111;
assign LUT_1[57525] = 32'b00000000000000001001010100101011;
assign LUT_1[57526] = 32'b00000000000000001011110001000000;
assign LUT_1[57527] = 32'b00000000000000000101000010111100;
assign LUT_1[57528] = 32'b00000000000000000111010111001101;
assign LUT_1[57529] = 32'b00000000000000000000101001001001;
assign LUT_1[57530] = 32'b00000000000000000011000101011110;
assign LUT_1[57531] = 32'b11111111111111111100010111011010;
assign LUT_1[57532] = 32'b00000000000000001111010000100100;
assign LUT_1[57533] = 32'b00000000000000001000100010100000;
assign LUT_1[57534] = 32'b00000000000000001010111110110101;
assign LUT_1[57535] = 32'b00000000000000000100010000110001;
assign LUT_1[57536] = 32'b00000000000000000111010000011111;
assign LUT_1[57537] = 32'b00000000000000000000100010011011;
assign LUT_1[57538] = 32'b00000000000000000010111110110000;
assign LUT_1[57539] = 32'b11111111111111111100010000101100;
assign LUT_1[57540] = 32'b00000000000000001111001001110110;
assign LUT_1[57541] = 32'b00000000000000001000011011110010;
assign LUT_1[57542] = 32'b00000000000000001010111000000111;
assign LUT_1[57543] = 32'b00000000000000000100001010000011;
assign LUT_1[57544] = 32'b00000000000000000110011110010100;
assign LUT_1[57545] = 32'b11111111111111111111110000010000;
assign LUT_1[57546] = 32'b00000000000000000010001100100101;
assign LUT_1[57547] = 32'b11111111111111111011011110100001;
assign LUT_1[57548] = 32'b00000000000000001110010111101011;
assign LUT_1[57549] = 32'b00000000000000000111101001100111;
assign LUT_1[57550] = 32'b00000000000000001010000101111100;
assign LUT_1[57551] = 32'b00000000000000000011010111111000;
assign LUT_1[57552] = 32'b00000000000000001001001100000001;
assign LUT_1[57553] = 32'b00000000000000000010011101111101;
assign LUT_1[57554] = 32'b00000000000000000100111010010010;
assign LUT_1[57555] = 32'b11111111111111111110001100001110;
assign LUT_1[57556] = 32'b00000000000000010001000101011000;
assign LUT_1[57557] = 32'b00000000000000001010010111010100;
assign LUT_1[57558] = 32'b00000000000000001100110011101001;
assign LUT_1[57559] = 32'b00000000000000000110000101100101;
assign LUT_1[57560] = 32'b00000000000000001000011001110110;
assign LUT_1[57561] = 32'b00000000000000000001101011110010;
assign LUT_1[57562] = 32'b00000000000000000100001000000111;
assign LUT_1[57563] = 32'b11111111111111111101011010000011;
assign LUT_1[57564] = 32'b00000000000000010000010011001101;
assign LUT_1[57565] = 32'b00000000000000001001100101001001;
assign LUT_1[57566] = 32'b00000000000000001100000001011110;
assign LUT_1[57567] = 32'b00000000000000000101010011011010;
assign LUT_1[57568] = 32'b00000000000000001000001011011110;
assign LUT_1[57569] = 32'b00000000000000000001011101011010;
assign LUT_1[57570] = 32'b00000000000000000011111001101111;
assign LUT_1[57571] = 32'b11111111111111111101001011101011;
assign LUT_1[57572] = 32'b00000000000000010000000100110101;
assign LUT_1[57573] = 32'b00000000000000001001010110110001;
assign LUT_1[57574] = 32'b00000000000000001011110011000110;
assign LUT_1[57575] = 32'b00000000000000000101000101000010;
assign LUT_1[57576] = 32'b00000000000000000111011001010011;
assign LUT_1[57577] = 32'b00000000000000000000101011001111;
assign LUT_1[57578] = 32'b00000000000000000011000111100100;
assign LUT_1[57579] = 32'b11111111111111111100011001100000;
assign LUT_1[57580] = 32'b00000000000000001111010010101010;
assign LUT_1[57581] = 32'b00000000000000001000100100100110;
assign LUT_1[57582] = 32'b00000000000000001011000000111011;
assign LUT_1[57583] = 32'b00000000000000000100010010110111;
assign LUT_1[57584] = 32'b00000000000000001010000111000000;
assign LUT_1[57585] = 32'b00000000000000000011011000111100;
assign LUT_1[57586] = 32'b00000000000000000101110101010001;
assign LUT_1[57587] = 32'b11111111111111111111000111001101;
assign LUT_1[57588] = 32'b00000000000000010010000000010111;
assign LUT_1[57589] = 32'b00000000000000001011010010010011;
assign LUT_1[57590] = 32'b00000000000000001101101110101000;
assign LUT_1[57591] = 32'b00000000000000000111000000100100;
assign LUT_1[57592] = 32'b00000000000000001001010100110101;
assign LUT_1[57593] = 32'b00000000000000000010100110110001;
assign LUT_1[57594] = 32'b00000000000000000101000011000110;
assign LUT_1[57595] = 32'b11111111111111111110010101000010;
assign LUT_1[57596] = 32'b00000000000000010001001110001100;
assign LUT_1[57597] = 32'b00000000000000001010100000001000;
assign LUT_1[57598] = 32'b00000000000000001100111100011101;
assign LUT_1[57599] = 32'b00000000000000000110001110011001;
assign LUT_1[57600] = 32'b00000000000000000000000111000000;
assign LUT_1[57601] = 32'b11111111111111111001011000111100;
assign LUT_1[57602] = 32'b11111111111111111011110101010001;
assign LUT_1[57603] = 32'b11111111111111110101000111001101;
assign LUT_1[57604] = 32'b00000000000000001000000000010111;
assign LUT_1[57605] = 32'b00000000000000000001010010010011;
assign LUT_1[57606] = 32'b00000000000000000011101110101000;
assign LUT_1[57607] = 32'b11111111111111111101000000100100;
assign LUT_1[57608] = 32'b11111111111111111111010100110101;
assign LUT_1[57609] = 32'b11111111111111111000100110110001;
assign LUT_1[57610] = 32'b11111111111111111011000011000110;
assign LUT_1[57611] = 32'b11111111111111110100010101000010;
assign LUT_1[57612] = 32'b00000000000000000111001110001100;
assign LUT_1[57613] = 32'b00000000000000000000100000001000;
assign LUT_1[57614] = 32'b00000000000000000010111100011101;
assign LUT_1[57615] = 32'b11111111111111111100001110011001;
assign LUT_1[57616] = 32'b00000000000000000010000010100010;
assign LUT_1[57617] = 32'b11111111111111111011010100011110;
assign LUT_1[57618] = 32'b11111111111111111101110000110011;
assign LUT_1[57619] = 32'b11111111111111110111000010101111;
assign LUT_1[57620] = 32'b00000000000000001001111011111001;
assign LUT_1[57621] = 32'b00000000000000000011001101110101;
assign LUT_1[57622] = 32'b00000000000000000101101010001010;
assign LUT_1[57623] = 32'b11111111111111111110111100000110;
assign LUT_1[57624] = 32'b00000000000000000001010000010111;
assign LUT_1[57625] = 32'b11111111111111111010100010010011;
assign LUT_1[57626] = 32'b11111111111111111100111110101000;
assign LUT_1[57627] = 32'b11111111111111110110010000100100;
assign LUT_1[57628] = 32'b00000000000000001001001001101110;
assign LUT_1[57629] = 32'b00000000000000000010011011101010;
assign LUT_1[57630] = 32'b00000000000000000100110111111111;
assign LUT_1[57631] = 32'b11111111111111111110001001111011;
assign LUT_1[57632] = 32'b00000000000000000001000001111111;
assign LUT_1[57633] = 32'b11111111111111111010010011111011;
assign LUT_1[57634] = 32'b11111111111111111100110000010000;
assign LUT_1[57635] = 32'b11111111111111110110000010001100;
assign LUT_1[57636] = 32'b00000000000000001000111011010110;
assign LUT_1[57637] = 32'b00000000000000000010001101010010;
assign LUT_1[57638] = 32'b00000000000000000100101001100111;
assign LUT_1[57639] = 32'b11111111111111111101111011100011;
assign LUT_1[57640] = 32'b00000000000000000000001111110100;
assign LUT_1[57641] = 32'b11111111111111111001100001110000;
assign LUT_1[57642] = 32'b11111111111111111011111110000101;
assign LUT_1[57643] = 32'b11111111111111110101010000000001;
assign LUT_1[57644] = 32'b00000000000000001000001001001011;
assign LUT_1[57645] = 32'b00000000000000000001011011000111;
assign LUT_1[57646] = 32'b00000000000000000011110111011100;
assign LUT_1[57647] = 32'b11111111111111111101001001011000;
assign LUT_1[57648] = 32'b00000000000000000010111101100001;
assign LUT_1[57649] = 32'b11111111111111111100001111011101;
assign LUT_1[57650] = 32'b11111111111111111110101011110010;
assign LUT_1[57651] = 32'b11111111111111110111111101101110;
assign LUT_1[57652] = 32'b00000000000000001010110110111000;
assign LUT_1[57653] = 32'b00000000000000000100001000110100;
assign LUT_1[57654] = 32'b00000000000000000110100101001001;
assign LUT_1[57655] = 32'b11111111111111111111110111000101;
assign LUT_1[57656] = 32'b00000000000000000010001011010110;
assign LUT_1[57657] = 32'b11111111111111111011011101010010;
assign LUT_1[57658] = 32'b11111111111111111101111001100111;
assign LUT_1[57659] = 32'b11111111111111110111001011100011;
assign LUT_1[57660] = 32'b00000000000000001010000100101101;
assign LUT_1[57661] = 32'b00000000000000000011010110101001;
assign LUT_1[57662] = 32'b00000000000000000101110010111110;
assign LUT_1[57663] = 32'b11111111111111111111000100111010;
assign LUT_1[57664] = 32'b00000000000000000010000100101000;
assign LUT_1[57665] = 32'b11111111111111111011010110100100;
assign LUT_1[57666] = 32'b11111111111111111101110010111001;
assign LUT_1[57667] = 32'b11111111111111110111000100110101;
assign LUT_1[57668] = 32'b00000000000000001001111101111111;
assign LUT_1[57669] = 32'b00000000000000000011001111111011;
assign LUT_1[57670] = 32'b00000000000000000101101100010000;
assign LUT_1[57671] = 32'b11111111111111111110111110001100;
assign LUT_1[57672] = 32'b00000000000000000001010010011101;
assign LUT_1[57673] = 32'b11111111111111111010100100011001;
assign LUT_1[57674] = 32'b11111111111111111101000000101110;
assign LUT_1[57675] = 32'b11111111111111110110010010101010;
assign LUT_1[57676] = 32'b00000000000000001001001011110100;
assign LUT_1[57677] = 32'b00000000000000000010011101110000;
assign LUT_1[57678] = 32'b00000000000000000100111010000101;
assign LUT_1[57679] = 32'b11111111111111111110001100000001;
assign LUT_1[57680] = 32'b00000000000000000100000000001010;
assign LUT_1[57681] = 32'b11111111111111111101010010000110;
assign LUT_1[57682] = 32'b11111111111111111111101110011011;
assign LUT_1[57683] = 32'b11111111111111111001000000010111;
assign LUT_1[57684] = 32'b00000000000000001011111001100001;
assign LUT_1[57685] = 32'b00000000000000000101001011011101;
assign LUT_1[57686] = 32'b00000000000000000111100111110010;
assign LUT_1[57687] = 32'b00000000000000000000111001101110;
assign LUT_1[57688] = 32'b00000000000000000011001101111111;
assign LUT_1[57689] = 32'b11111111111111111100011111111011;
assign LUT_1[57690] = 32'b11111111111111111110111100010000;
assign LUT_1[57691] = 32'b11111111111111111000001110001100;
assign LUT_1[57692] = 32'b00000000000000001011000111010110;
assign LUT_1[57693] = 32'b00000000000000000100011001010010;
assign LUT_1[57694] = 32'b00000000000000000110110101100111;
assign LUT_1[57695] = 32'b00000000000000000000000111100011;
assign LUT_1[57696] = 32'b00000000000000000010111111100111;
assign LUT_1[57697] = 32'b11111111111111111100010001100011;
assign LUT_1[57698] = 32'b11111111111111111110101101111000;
assign LUT_1[57699] = 32'b11111111111111110111111111110100;
assign LUT_1[57700] = 32'b00000000000000001010111000111110;
assign LUT_1[57701] = 32'b00000000000000000100001010111010;
assign LUT_1[57702] = 32'b00000000000000000110100111001111;
assign LUT_1[57703] = 32'b11111111111111111111111001001011;
assign LUT_1[57704] = 32'b00000000000000000010001101011100;
assign LUT_1[57705] = 32'b11111111111111111011011111011000;
assign LUT_1[57706] = 32'b11111111111111111101111011101101;
assign LUT_1[57707] = 32'b11111111111111110111001101101001;
assign LUT_1[57708] = 32'b00000000000000001010000110110011;
assign LUT_1[57709] = 32'b00000000000000000011011000101111;
assign LUT_1[57710] = 32'b00000000000000000101110101000100;
assign LUT_1[57711] = 32'b11111111111111111111000111000000;
assign LUT_1[57712] = 32'b00000000000000000100111011001001;
assign LUT_1[57713] = 32'b11111111111111111110001101000101;
assign LUT_1[57714] = 32'b00000000000000000000101001011010;
assign LUT_1[57715] = 32'b11111111111111111001111011010110;
assign LUT_1[57716] = 32'b00000000000000001100110100100000;
assign LUT_1[57717] = 32'b00000000000000000110000110011100;
assign LUT_1[57718] = 32'b00000000000000001000100010110001;
assign LUT_1[57719] = 32'b00000000000000000001110100101101;
assign LUT_1[57720] = 32'b00000000000000000100001000111110;
assign LUT_1[57721] = 32'b11111111111111111101011010111010;
assign LUT_1[57722] = 32'b11111111111111111111110111001111;
assign LUT_1[57723] = 32'b11111111111111111001001001001011;
assign LUT_1[57724] = 32'b00000000000000001100000010010101;
assign LUT_1[57725] = 32'b00000000000000000101010100010001;
assign LUT_1[57726] = 32'b00000000000000000111110000100110;
assign LUT_1[57727] = 32'b00000000000000000001000010100010;
assign LUT_1[57728] = 32'b00000000000000000011000111000011;
assign LUT_1[57729] = 32'b11111111111111111100011000111111;
assign LUT_1[57730] = 32'b11111111111111111110110101010100;
assign LUT_1[57731] = 32'b11111111111111111000000111010000;
assign LUT_1[57732] = 32'b00000000000000001011000000011010;
assign LUT_1[57733] = 32'b00000000000000000100010010010110;
assign LUT_1[57734] = 32'b00000000000000000110101110101011;
assign LUT_1[57735] = 32'b00000000000000000000000000100111;
assign LUT_1[57736] = 32'b00000000000000000010010100111000;
assign LUT_1[57737] = 32'b11111111111111111011100110110100;
assign LUT_1[57738] = 32'b11111111111111111110000011001001;
assign LUT_1[57739] = 32'b11111111111111110111010101000101;
assign LUT_1[57740] = 32'b00000000000000001010001110001111;
assign LUT_1[57741] = 32'b00000000000000000011100000001011;
assign LUT_1[57742] = 32'b00000000000000000101111100100000;
assign LUT_1[57743] = 32'b11111111111111111111001110011100;
assign LUT_1[57744] = 32'b00000000000000000101000010100101;
assign LUT_1[57745] = 32'b11111111111111111110010100100001;
assign LUT_1[57746] = 32'b00000000000000000000110000110110;
assign LUT_1[57747] = 32'b11111111111111111010000010110010;
assign LUT_1[57748] = 32'b00000000000000001100111011111100;
assign LUT_1[57749] = 32'b00000000000000000110001101111000;
assign LUT_1[57750] = 32'b00000000000000001000101010001101;
assign LUT_1[57751] = 32'b00000000000000000001111100001001;
assign LUT_1[57752] = 32'b00000000000000000100010000011010;
assign LUT_1[57753] = 32'b11111111111111111101100010010110;
assign LUT_1[57754] = 32'b11111111111111111111111110101011;
assign LUT_1[57755] = 32'b11111111111111111001010000100111;
assign LUT_1[57756] = 32'b00000000000000001100001001110001;
assign LUT_1[57757] = 32'b00000000000000000101011011101101;
assign LUT_1[57758] = 32'b00000000000000000111111000000010;
assign LUT_1[57759] = 32'b00000000000000000001001001111110;
assign LUT_1[57760] = 32'b00000000000000000100000010000010;
assign LUT_1[57761] = 32'b11111111111111111101010011111110;
assign LUT_1[57762] = 32'b11111111111111111111110000010011;
assign LUT_1[57763] = 32'b11111111111111111001000010001111;
assign LUT_1[57764] = 32'b00000000000000001011111011011001;
assign LUT_1[57765] = 32'b00000000000000000101001101010101;
assign LUT_1[57766] = 32'b00000000000000000111101001101010;
assign LUT_1[57767] = 32'b00000000000000000000111011100110;
assign LUT_1[57768] = 32'b00000000000000000011001111110111;
assign LUT_1[57769] = 32'b11111111111111111100100001110011;
assign LUT_1[57770] = 32'b11111111111111111110111110001000;
assign LUT_1[57771] = 32'b11111111111111111000010000000100;
assign LUT_1[57772] = 32'b00000000000000001011001001001110;
assign LUT_1[57773] = 32'b00000000000000000100011011001010;
assign LUT_1[57774] = 32'b00000000000000000110110111011111;
assign LUT_1[57775] = 32'b00000000000000000000001001011011;
assign LUT_1[57776] = 32'b00000000000000000101111101100100;
assign LUT_1[57777] = 32'b11111111111111111111001111100000;
assign LUT_1[57778] = 32'b00000000000000000001101011110101;
assign LUT_1[57779] = 32'b11111111111111111010111101110001;
assign LUT_1[57780] = 32'b00000000000000001101110110111011;
assign LUT_1[57781] = 32'b00000000000000000111001000110111;
assign LUT_1[57782] = 32'b00000000000000001001100101001100;
assign LUT_1[57783] = 32'b00000000000000000010110111001000;
assign LUT_1[57784] = 32'b00000000000000000101001011011001;
assign LUT_1[57785] = 32'b11111111111111111110011101010101;
assign LUT_1[57786] = 32'b00000000000000000000111001101010;
assign LUT_1[57787] = 32'b11111111111111111010001011100110;
assign LUT_1[57788] = 32'b00000000000000001101000100110000;
assign LUT_1[57789] = 32'b00000000000000000110010110101100;
assign LUT_1[57790] = 32'b00000000000000001000110011000001;
assign LUT_1[57791] = 32'b00000000000000000010000100111101;
assign LUT_1[57792] = 32'b00000000000000000101000100101011;
assign LUT_1[57793] = 32'b11111111111111111110010110100111;
assign LUT_1[57794] = 32'b00000000000000000000110010111100;
assign LUT_1[57795] = 32'b11111111111111111010000100111000;
assign LUT_1[57796] = 32'b00000000000000001100111110000010;
assign LUT_1[57797] = 32'b00000000000000000110001111111110;
assign LUT_1[57798] = 32'b00000000000000001000101100010011;
assign LUT_1[57799] = 32'b00000000000000000001111110001111;
assign LUT_1[57800] = 32'b00000000000000000100010010100000;
assign LUT_1[57801] = 32'b11111111111111111101100100011100;
assign LUT_1[57802] = 32'b00000000000000000000000000110001;
assign LUT_1[57803] = 32'b11111111111111111001010010101101;
assign LUT_1[57804] = 32'b00000000000000001100001011110111;
assign LUT_1[57805] = 32'b00000000000000000101011101110011;
assign LUT_1[57806] = 32'b00000000000000000111111010001000;
assign LUT_1[57807] = 32'b00000000000000000001001100000100;
assign LUT_1[57808] = 32'b00000000000000000111000000001101;
assign LUT_1[57809] = 32'b00000000000000000000010010001001;
assign LUT_1[57810] = 32'b00000000000000000010101110011110;
assign LUT_1[57811] = 32'b11111111111111111100000000011010;
assign LUT_1[57812] = 32'b00000000000000001110111001100100;
assign LUT_1[57813] = 32'b00000000000000001000001011100000;
assign LUT_1[57814] = 32'b00000000000000001010100111110101;
assign LUT_1[57815] = 32'b00000000000000000011111001110001;
assign LUT_1[57816] = 32'b00000000000000000110001110000010;
assign LUT_1[57817] = 32'b11111111111111111111011111111110;
assign LUT_1[57818] = 32'b00000000000000000001111100010011;
assign LUT_1[57819] = 32'b11111111111111111011001110001111;
assign LUT_1[57820] = 32'b00000000000000001110000111011001;
assign LUT_1[57821] = 32'b00000000000000000111011001010101;
assign LUT_1[57822] = 32'b00000000000000001001110101101010;
assign LUT_1[57823] = 32'b00000000000000000011000111100110;
assign LUT_1[57824] = 32'b00000000000000000101111111101010;
assign LUT_1[57825] = 32'b11111111111111111111010001100110;
assign LUT_1[57826] = 32'b00000000000000000001101101111011;
assign LUT_1[57827] = 32'b11111111111111111010111111110111;
assign LUT_1[57828] = 32'b00000000000000001101111001000001;
assign LUT_1[57829] = 32'b00000000000000000111001010111101;
assign LUT_1[57830] = 32'b00000000000000001001100111010010;
assign LUT_1[57831] = 32'b00000000000000000010111001001110;
assign LUT_1[57832] = 32'b00000000000000000101001101011111;
assign LUT_1[57833] = 32'b11111111111111111110011111011011;
assign LUT_1[57834] = 32'b00000000000000000000111011110000;
assign LUT_1[57835] = 32'b11111111111111111010001101101100;
assign LUT_1[57836] = 32'b00000000000000001101000110110110;
assign LUT_1[57837] = 32'b00000000000000000110011000110010;
assign LUT_1[57838] = 32'b00000000000000001000110101000111;
assign LUT_1[57839] = 32'b00000000000000000010000111000011;
assign LUT_1[57840] = 32'b00000000000000000111111011001100;
assign LUT_1[57841] = 32'b00000000000000000001001101001000;
assign LUT_1[57842] = 32'b00000000000000000011101001011101;
assign LUT_1[57843] = 32'b11111111111111111100111011011001;
assign LUT_1[57844] = 32'b00000000000000001111110100100011;
assign LUT_1[57845] = 32'b00000000000000001001000110011111;
assign LUT_1[57846] = 32'b00000000000000001011100010110100;
assign LUT_1[57847] = 32'b00000000000000000100110100110000;
assign LUT_1[57848] = 32'b00000000000000000111001001000001;
assign LUT_1[57849] = 32'b00000000000000000000011010111101;
assign LUT_1[57850] = 32'b00000000000000000010110111010010;
assign LUT_1[57851] = 32'b11111111111111111100001001001110;
assign LUT_1[57852] = 32'b00000000000000001111000010011000;
assign LUT_1[57853] = 32'b00000000000000001000010100010100;
assign LUT_1[57854] = 32'b00000000000000001010110000101001;
assign LUT_1[57855] = 32'b00000000000000000100000010100101;
assign LUT_1[57856] = 32'b11111111111111111100000001010001;
assign LUT_1[57857] = 32'b11111111111111110101010011001101;
assign LUT_1[57858] = 32'b11111111111111110111101111100010;
assign LUT_1[57859] = 32'b11111111111111110001000001011110;
assign LUT_1[57860] = 32'b00000000000000000011111010101000;
assign LUT_1[57861] = 32'b11111111111111111101001100100100;
assign LUT_1[57862] = 32'b11111111111111111111101000111001;
assign LUT_1[57863] = 32'b11111111111111111000111010110101;
assign LUT_1[57864] = 32'b11111111111111111011001111000110;
assign LUT_1[57865] = 32'b11111111111111110100100001000010;
assign LUT_1[57866] = 32'b11111111111111110110111101010111;
assign LUT_1[57867] = 32'b11111111111111110000001111010011;
assign LUT_1[57868] = 32'b00000000000000000011001000011101;
assign LUT_1[57869] = 32'b11111111111111111100011010011001;
assign LUT_1[57870] = 32'b11111111111111111110110110101110;
assign LUT_1[57871] = 32'b11111111111111111000001000101010;
assign LUT_1[57872] = 32'b11111111111111111101111100110011;
assign LUT_1[57873] = 32'b11111111111111110111001110101111;
assign LUT_1[57874] = 32'b11111111111111111001101011000100;
assign LUT_1[57875] = 32'b11111111111111110010111101000000;
assign LUT_1[57876] = 32'b00000000000000000101110110001010;
assign LUT_1[57877] = 32'b11111111111111111111001000000110;
assign LUT_1[57878] = 32'b00000000000000000001100100011011;
assign LUT_1[57879] = 32'b11111111111111111010110110010111;
assign LUT_1[57880] = 32'b11111111111111111101001010101000;
assign LUT_1[57881] = 32'b11111111111111110110011100100100;
assign LUT_1[57882] = 32'b11111111111111111000111000111001;
assign LUT_1[57883] = 32'b11111111111111110010001010110101;
assign LUT_1[57884] = 32'b00000000000000000101000011111111;
assign LUT_1[57885] = 32'b11111111111111111110010101111011;
assign LUT_1[57886] = 32'b00000000000000000000110010010000;
assign LUT_1[57887] = 32'b11111111111111111010000100001100;
assign LUT_1[57888] = 32'b11111111111111111100111100010000;
assign LUT_1[57889] = 32'b11111111111111110110001110001100;
assign LUT_1[57890] = 32'b11111111111111111000101010100001;
assign LUT_1[57891] = 32'b11111111111111110001111100011101;
assign LUT_1[57892] = 32'b00000000000000000100110101100111;
assign LUT_1[57893] = 32'b11111111111111111110000111100011;
assign LUT_1[57894] = 32'b00000000000000000000100011111000;
assign LUT_1[57895] = 32'b11111111111111111001110101110100;
assign LUT_1[57896] = 32'b11111111111111111100001010000101;
assign LUT_1[57897] = 32'b11111111111111110101011100000001;
assign LUT_1[57898] = 32'b11111111111111110111111000010110;
assign LUT_1[57899] = 32'b11111111111111110001001010010010;
assign LUT_1[57900] = 32'b00000000000000000100000011011100;
assign LUT_1[57901] = 32'b11111111111111111101010101011000;
assign LUT_1[57902] = 32'b11111111111111111111110001101101;
assign LUT_1[57903] = 32'b11111111111111111001000011101001;
assign LUT_1[57904] = 32'b11111111111111111110110111110010;
assign LUT_1[57905] = 32'b11111111111111111000001001101110;
assign LUT_1[57906] = 32'b11111111111111111010100110000011;
assign LUT_1[57907] = 32'b11111111111111110011110111111111;
assign LUT_1[57908] = 32'b00000000000000000110110001001001;
assign LUT_1[57909] = 32'b00000000000000000000000011000101;
assign LUT_1[57910] = 32'b00000000000000000010011111011010;
assign LUT_1[57911] = 32'b11111111111111111011110001010110;
assign LUT_1[57912] = 32'b11111111111111111110000101100111;
assign LUT_1[57913] = 32'b11111111111111110111010111100011;
assign LUT_1[57914] = 32'b11111111111111111001110011111000;
assign LUT_1[57915] = 32'b11111111111111110011000101110100;
assign LUT_1[57916] = 32'b00000000000000000101111110111110;
assign LUT_1[57917] = 32'b11111111111111111111010000111010;
assign LUT_1[57918] = 32'b00000000000000000001101101001111;
assign LUT_1[57919] = 32'b11111111111111111010111111001011;
assign LUT_1[57920] = 32'b11111111111111111101111110111001;
assign LUT_1[57921] = 32'b11111111111111110111010000110101;
assign LUT_1[57922] = 32'b11111111111111111001101101001010;
assign LUT_1[57923] = 32'b11111111111111110010111111000110;
assign LUT_1[57924] = 32'b00000000000000000101111000010000;
assign LUT_1[57925] = 32'b11111111111111111111001010001100;
assign LUT_1[57926] = 32'b00000000000000000001100110100001;
assign LUT_1[57927] = 32'b11111111111111111010111000011101;
assign LUT_1[57928] = 32'b11111111111111111101001100101110;
assign LUT_1[57929] = 32'b11111111111111110110011110101010;
assign LUT_1[57930] = 32'b11111111111111111000111010111111;
assign LUT_1[57931] = 32'b11111111111111110010001100111011;
assign LUT_1[57932] = 32'b00000000000000000101000110000101;
assign LUT_1[57933] = 32'b11111111111111111110011000000001;
assign LUT_1[57934] = 32'b00000000000000000000110100010110;
assign LUT_1[57935] = 32'b11111111111111111010000110010010;
assign LUT_1[57936] = 32'b11111111111111111111111010011011;
assign LUT_1[57937] = 32'b11111111111111111001001100010111;
assign LUT_1[57938] = 32'b11111111111111111011101000101100;
assign LUT_1[57939] = 32'b11111111111111110100111010101000;
assign LUT_1[57940] = 32'b00000000000000000111110011110010;
assign LUT_1[57941] = 32'b00000000000000000001000101101110;
assign LUT_1[57942] = 32'b00000000000000000011100010000011;
assign LUT_1[57943] = 32'b11111111111111111100110011111111;
assign LUT_1[57944] = 32'b11111111111111111111001000010000;
assign LUT_1[57945] = 32'b11111111111111111000011010001100;
assign LUT_1[57946] = 32'b11111111111111111010110110100001;
assign LUT_1[57947] = 32'b11111111111111110100001000011101;
assign LUT_1[57948] = 32'b00000000000000000111000001100111;
assign LUT_1[57949] = 32'b00000000000000000000010011100011;
assign LUT_1[57950] = 32'b00000000000000000010101111111000;
assign LUT_1[57951] = 32'b11111111111111111100000001110100;
assign LUT_1[57952] = 32'b11111111111111111110111001111000;
assign LUT_1[57953] = 32'b11111111111111111000001011110100;
assign LUT_1[57954] = 32'b11111111111111111010101000001001;
assign LUT_1[57955] = 32'b11111111111111110011111010000101;
assign LUT_1[57956] = 32'b00000000000000000110110011001111;
assign LUT_1[57957] = 32'b00000000000000000000000101001011;
assign LUT_1[57958] = 32'b00000000000000000010100001100000;
assign LUT_1[57959] = 32'b11111111111111111011110011011100;
assign LUT_1[57960] = 32'b11111111111111111110000111101101;
assign LUT_1[57961] = 32'b11111111111111110111011001101001;
assign LUT_1[57962] = 32'b11111111111111111001110101111110;
assign LUT_1[57963] = 32'b11111111111111110011000111111010;
assign LUT_1[57964] = 32'b00000000000000000110000001000100;
assign LUT_1[57965] = 32'b11111111111111111111010011000000;
assign LUT_1[57966] = 32'b00000000000000000001101111010101;
assign LUT_1[57967] = 32'b11111111111111111011000001010001;
assign LUT_1[57968] = 32'b00000000000000000000110101011010;
assign LUT_1[57969] = 32'b11111111111111111010000111010110;
assign LUT_1[57970] = 32'b11111111111111111100100011101011;
assign LUT_1[57971] = 32'b11111111111111110101110101100111;
assign LUT_1[57972] = 32'b00000000000000001000101110110001;
assign LUT_1[57973] = 32'b00000000000000000010000000101101;
assign LUT_1[57974] = 32'b00000000000000000100011101000010;
assign LUT_1[57975] = 32'b11111111111111111101101110111110;
assign LUT_1[57976] = 32'b00000000000000000000000011001111;
assign LUT_1[57977] = 32'b11111111111111111001010101001011;
assign LUT_1[57978] = 32'b11111111111111111011110001100000;
assign LUT_1[57979] = 32'b11111111111111110101000011011100;
assign LUT_1[57980] = 32'b00000000000000000111111100100110;
assign LUT_1[57981] = 32'b00000000000000000001001110100010;
assign LUT_1[57982] = 32'b00000000000000000011101010110111;
assign LUT_1[57983] = 32'b11111111111111111100111100110011;
assign LUT_1[57984] = 32'b11111111111111111111000001010100;
assign LUT_1[57985] = 32'b11111111111111111000010011010000;
assign LUT_1[57986] = 32'b11111111111111111010101111100101;
assign LUT_1[57987] = 32'b11111111111111110100000001100001;
assign LUT_1[57988] = 32'b00000000000000000110111010101011;
assign LUT_1[57989] = 32'b00000000000000000000001100100111;
assign LUT_1[57990] = 32'b00000000000000000010101000111100;
assign LUT_1[57991] = 32'b11111111111111111011111010111000;
assign LUT_1[57992] = 32'b11111111111111111110001111001001;
assign LUT_1[57993] = 32'b11111111111111110111100001000101;
assign LUT_1[57994] = 32'b11111111111111111001111101011010;
assign LUT_1[57995] = 32'b11111111111111110011001111010110;
assign LUT_1[57996] = 32'b00000000000000000110001000100000;
assign LUT_1[57997] = 32'b11111111111111111111011010011100;
assign LUT_1[57998] = 32'b00000000000000000001110110110001;
assign LUT_1[57999] = 32'b11111111111111111011001000101101;
assign LUT_1[58000] = 32'b00000000000000000000111100110110;
assign LUT_1[58001] = 32'b11111111111111111010001110110010;
assign LUT_1[58002] = 32'b11111111111111111100101011000111;
assign LUT_1[58003] = 32'b11111111111111110101111101000011;
assign LUT_1[58004] = 32'b00000000000000001000110110001101;
assign LUT_1[58005] = 32'b00000000000000000010001000001001;
assign LUT_1[58006] = 32'b00000000000000000100100100011110;
assign LUT_1[58007] = 32'b11111111111111111101110110011010;
assign LUT_1[58008] = 32'b00000000000000000000001010101011;
assign LUT_1[58009] = 32'b11111111111111111001011100100111;
assign LUT_1[58010] = 32'b11111111111111111011111000111100;
assign LUT_1[58011] = 32'b11111111111111110101001010111000;
assign LUT_1[58012] = 32'b00000000000000001000000100000010;
assign LUT_1[58013] = 32'b00000000000000000001010101111110;
assign LUT_1[58014] = 32'b00000000000000000011110010010011;
assign LUT_1[58015] = 32'b11111111111111111101000100001111;
assign LUT_1[58016] = 32'b11111111111111111111111100010011;
assign LUT_1[58017] = 32'b11111111111111111001001110001111;
assign LUT_1[58018] = 32'b11111111111111111011101010100100;
assign LUT_1[58019] = 32'b11111111111111110100111100100000;
assign LUT_1[58020] = 32'b00000000000000000111110101101010;
assign LUT_1[58021] = 32'b00000000000000000001000111100110;
assign LUT_1[58022] = 32'b00000000000000000011100011111011;
assign LUT_1[58023] = 32'b11111111111111111100110101110111;
assign LUT_1[58024] = 32'b11111111111111111111001010001000;
assign LUT_1[58025] = 32'b11111111111111111000011100000100;
assign LUT_1[58026] = 32'b11111111111111111010111000011001;
assign LUT_1[58027] = 32'b11111111111111110100001010010101;
assign LUT_1[58028] = 32'b00000000000000000111000011011111;
assign LUT_1[58029] = 32'b00000000000000000000010101011011;
assign LUT_1[58030] = 32'b00000000000000000010110001110000;
assign LUT_1[58031] = 32'b11111111111111111100000011101100;
assign LUT_1[58032] = 32'b00000000000000000001110111110101;
assign LUT_1[58033] = 32'b11111111111111111011001001110001;
assign LUT_1[58034] = 32'b11111111111111111101100110000110;
assign LUT_1[58035] = 32'b11111111111111110110111000000010;
assign LUT_1[58036] = 32'b00000000000000001001110001001100;
assign LUT_1[58037] = 32'b00000000000000000011000011001000;
assign LUT_1[58038] = 32'b00000000000000000101011111011101;
assign LUT_1[58039] = 32'b11111111111111111110110001011001;
assign LUT_1[58040] = 32'b00000000000000000001000101101010;
assign LUT_1[58041] = 32'b11111111111111111010010111100110;
assign LUT_1[58042] = 32'b11111111111111111100110011111011;
assign LUT_1[58043] = 32'b11111111111111110110000101110111;
assign LUT_1[58044] = 32'b00000000000000001000111111000001;
assign LUT_1[58045] = 32'b00000000000000000010010000111101;
assign LUT_1[58046] = 32'b00000000000000000100101101010010;
assign LUT_1[58047] = 32'b11111111111111111101111111001110;
assign LUT_1[58048] = 32'b00000000000000000000111110111100;
assign LUT_1[58049] = 32'b11111111111111111010010000111000;
assign LUT_1[58050] = 32'b11111111111111111100101101001101;
assign LUT_1[58051] = 32'b11111111111111110101111111001001;
assign LUT_1[58052] = 32'b00000000000000001000111000010011;
assign LUT_1[58053] = 32'b00000000000000000010001010001111;
assign LUT_1[58054] = 32'b00000000000000000100100110100100;
assign LUT_1[58055] = 32'b11111111111111111101111000100000;
assign LUT_1[58056] = 32'b00000000000000000000001100110001;
assign LUT_1[58057] = 32'b11111111111111111001011110101101;
assign LUT_1[58058] = 32'b11111111111111111011111011000010;
assign LUT_1[58059] = 32'b11111111111111110101001100111110;
assign LUT_1[58060] = 32'b00000000000000001000000110001000;
assign LUT_1[58061] = 32'b00000000000000000001011000000100;
assign LUT_1[58062] = 32'b00000000000000000011110100011001;
assign LUT_1[58063] = 32'b11111111111111111101000110010101;
assign LUT_1[58064] = 32'b00000000000000000010111010011110;
assign LUT_1[58065] = 32'b11111111111111111100001100011010;
assign LUT_1[58066] = 32'b11111111111111111110101000101111;
assign LUT_1[58067] = 32'b11111111111111110111111010101011;
assign LUT_1[58068] = 32'b00000000000000001010110011110101;
assign LUT_1[58069] = 32'b00000000000000000100000101110001;
assign LUT_1[58070] = 32'b00000000000000000110100010000110;
assign LUT_1[58071] = 32'b11111111111111111111110100000010;
assign LUT_1[58072] = 32'b00000000000000000010001000010011;
assign LUT_1[58073] = 32'b11111111111111111011011010001111;
assign LUT_1[58074] = 32'b11111111111111111101110110100100;
assign LUT_1[58075] = 32'b11111111111111110111001000100000;
assign LUT_1[58076] = 32'b00000000000000001010000001101010;
assign LUT_1[58077] = 32'b00000000000000000011010011100110;
assign LUT_1[58078] = 32'b00000000000000000101101111111011;
assign LUT_1[58079] = 32'b11111111111111111111000001110111;
assign LUT_1[58080] = 32'b00000000000000000001111001111011;
assign LUT_1[58081] = 32'b11111111111111111011001011110111;
assign LUT_1[58082] = 32'b11111111111111111101101000001100;
assign LUT_1[58083] = 32'b11111111111111110110111010001000;
assign LUT_1[58084] = 32'b00000000000000001001110011010010;
assign LUT_1[58085] = 32'b00000000000000000011000101001110;
assign LUT_1[58086] = 32'b00000000000000000101100001100011;
assign LUT_1[58087] = 32'b11111111111111111110110011011111;
assign LUT_1[58088] = 32'b00000000000000000001000111110000;
assign LUT_1[58089] = 32'b11111111111111111010011001101100;
assign LUT_1[58090] = 32'b11111111111111111100110110000001;
assign LUT_1[58091] = 32'b11111111111111110110000111111101;
assign LUT_1[58092] = 32'b00000000000000001001000001000111;
assign LUT_1[58093] = 32'b00000000000000000010010011000011;
assign LUT_1[58094] = 32'b00000000000000000100101111011000;
assign LUT_1[58095] = 32'b11111111111111111110000001010100;
assign LUT_1[58096] = 32'b00000000000000000011110101011101;
assign LUT_1[58097] = 32'b11111111111111111101000111011001;
assign LUT_1[58098] = 32'b11111111111111111111100011101110;
assign LUT_1[58099] = 32'b11111111111111111000110101101010;
assign LUT_1[58100] = 32'b00000000000000001011101110110100;
assign LUT_1[58101] = 32'b00000000000000000101000000110000;
assign LUT_1[58102] = 32'b00000000000000000111011101000101;
assign LUT_1[58103] = 32'b00000000000000000000101111000001;
assign LUT_1[58104] = 32'b00000000000000000011000011010010;
assign LUT_1[58105] = 32'b11111111111111111100010101001110;
assign LUT_1[58106] = 32'b11111111111111111110110001100011;
assign LUT_1[58107] = 32'b11111111111111111000000011011111;
assign LUT_1[58108] = 32'b00000000000000001010111100101001;
assign LUT_1[58109] = 32'b00000000000000000100001110100101;
assign LUT_1[58110] = 32'b00000000000000000110101010111010;
assign LUT_1[58111] = 32'b11111111111111111111111100110110;
assign LUT_1[58112] = 32'b11111111111111111001110101011101;
assign LUT_1[58113] = 32'b11111111111111110011000111011001;
assign LUT_1[58114] = 32'b11111111111111110101100011101110;
assign LUT_1[58115] = 32'b11111111111111101110110101101010;
assign LUT_1[58116] = 32'b00000000000000000001101110110100;
assign LUT_1[58117] = 32'b11111111111111111011000000110000;
assign LUT_1[58118] = 32'b11111111111111111101011101000101;
assign LUT_1[58119] = 32'b11111111111111110110101111000001;
assign LUT_1[58120] = 32'b11111111111111111001000011010010;
assign LUT_1[58121] = 32'b11111111111111110010010101001110;
assign LUT_1[58122] = 32'b11111111111111110100110001100011;
assign LUT_1[58123] = 32'b11111111111111101110000011011111;
assign LUT_1[58124] = 32'b00000000000000000000111100101001;
assign LUT_1[58125] = 32'b11111111111111111010001110100101;
assign LUT_1[58126] = 32'b11111111111111111100101010111010;
assign LUT_1[58127] = 32'b11111111111111110101111100110110;
assign LUT_1[58128] = 32'b11111111111111111011110000111111;
assign LUT_1[58129] = 32'b11111111111111110101000010111011;
assign LUT_1[58130] = 32'b11111111111111110111011111010000;
assign LUT_1[58131] = 32'b11111111111111110000110001001100;
assign LUT_1[58132] = 32'b00000000000000000011101010010110;
assign LUT_1[58133] = 32'b11111111111111111100111100010010;
assign LUT_1[58134] = 32'b11111111111111111111011000100111;
assign LUT_1[58135] = 32'b11111111111111111000101010100011;
assign LUT_1[58136] = 32'b11111111111111111010111110110100;
assign LUT_1[58137] = 32'b11111111111111110100010000110000;
assign LUT_1[58138] = 32'b11111111111111110110101101000101;
assign LUT_1[58139] = 32'b11111111111111101111111111000001;
assign LUT_1[58140] = 32'b00000000000000000010111000001011;
assign LUT_1[58141] = 32'b11111111111111111100001010000111;
assign LUT_1[58142] = 32'b11111111111111111110100110011100;
assign LUT_1[58143] = 32'b11111111111111110111111000011000;
assign LUT_1[58144] = 32'b11111111111111111010110000011100;
assign LUT_1[58145] = 32'b11111111111111110100000010011000;
assign LUT_1[58146] = 32'b11111111111111110110011110101101;
assign LUT_1[58147] = 32'b11111111111111101111110000101001;
assign LUT_1[58148] = 32'b00000000000000000010101001110011;
assign LUT_1[58149] = 32'b11111111111111111011111011101111;
assign LUT_1[58150] = 32'b11111111111111111110011000000100;
assign LUT_1[58151] = 32'b11111111111111110111101010000000;
assign LUT_1[58152] = 32'b11111111111111111001111110010001;
assign LUT_1[58153] = 32'b11111111111111110011010000001101;
assign LUT_1[58154] = 32'b11111111111111110101101100100010;
assign LUT_1[58155] = 32'b11111111111111101110111110011110;
assign LUT_1[58156] = 32'b00000000000000000001110111101000;
assign LUT_1[58157] = 32'b11111111111111111011001001100100;
assign LUT_1[58158] = 32'b11111111111111111101100101111001;
assign LUT_1[58159] = 32'b11111111111111110110110111110101;
assign LUT_1[58160] = 32'b11111111111111111100101011111110;
assign LUT_1[58161] = 32'b11111111111111110101111101111010;
assign LUT_1[58162] = 32'b11111111111111111000011010001111;
assign LUT_1[58163] = 32'b11111111111111110001101100001011;
assign LUT_1[58164] = 32'b00000000000000000100100101010101;
assign LUT_1[58165] = 32'b11111111111111111101110111010001;
assign LUT_1[58166] = 32'b00000000000000000000010011100110;
assign LUT_1[58167] = 32'b11111111111111111001100101100010;
assign LUT_1[58168] = 32'b11111111111111111011111001110011;
assign LUT_1[58169] = 32'b11111111111111110101001011101111;
assign LUT_1[58170] = 32'b11111111111111110111101000000100;
assign LUT_1[58171] = 32'b11111111111111110000111010000000;
assign LUT_1[58172] = 32'b00000000000000000011110011001010;
assign LUT_1[58173] = 32'b11111111111111111101000101000110;
assign LUT_1[58174] = 32'b11111111111111111111100001011011;
assign LUT_1[58175] = 32'b11111111111111111000110011010111;
assign LUT_1[58176] = 32'b11111111111111111011110011000101;
assign LUT_1[58177] = 32'b11111111111111110101000101000001;
assign LUT_1[58178] = 32'b11111111111111110111100001010110;
assign LUT_1[58179] = 32'b11111111111111110000110011010010;
assign LUT_1[58180] = 32'b00000000000000000011101100011100;
assign LUT_1[58181] = 32'b11111111111111111100111110011000;
assign LUT_1[58182] = 32'b11111111111111111111011010101101;
assign LUT_1[58183] = 32'b11111111111111111000101100101001;
assign LUT_1[58184] = 32'b11111111111111111011000000111010;
assign LUT_1[58185] = 32'b11111111111111110100010010110110;
assign LUT_1[58186] = 32'b11111111111111110110101111001011;
assign LUT_1[58187] = 32'b11111111111111110000000001000111;
assign LUT_1[58188] = 32'b00000000000000000010111010010001;
assign LUT_1[58189] = 32'b11111111111111111100001100001101;
assign LUT_1[58190] = 32'b11111111111111111110101000100010;
assign LUT_1[58191] = 32'b11111111111111110111111010011110;
assign LUT_1[58192] = 32'b11111111111111111101101110100111;
assign LUT_1[58193] = 32'b11111111111111110111000000100011;
assign LUT_1[58194] = 32'b11111111111111111001011100111000;
assign LUT_1[58195] = 32'b11111111111111110010101110110100;
assign LUT_1[58196] = 32'b00000000000000000101100111111110;
assign LUT_1[58197] = 32'b11111111111111111110111001111010;
assign LUT_1[58198] = 32'b00000000000000000001010110001111;
assign LUT_1[58199] = 32'b11111111111111111010101000001011;
assign LUT_1[58200] = 32'b11111111111111111100111100011100;
assign LUT_1[58201] = 32'b11111111111111110110001110011000;
assign LUT_1[58202] = 32'b11111111111111111000101010101101;
assign LUT_1[58203] = 32'b11111111111111110001111100101001;
assign LUT_1[58204] = 32'b00000000000000000100110101110011;
assign LUT_1[58205] = 32'b11111111111111111110000111101111;
assign LUT_1[58206] = 32'b00000000000000000000100100000100;
assign LUT_1[58207] = 32'b11111111111111111001110110000000;
assign LUT_1[58208] = 32'b11111111111111111100101110000100;
assign LUT_1[58209] = 32'b11111111111111110110000000000000;
assign LUT_1[58210] = 32'b11111111111111111000011100010101;
assign LUT_1[58211] = 32'b11111111111111110001101110010001;
assign LUT_1[58212] = 32'b00000000000000000100100111011011;
assign LUT_1[58213] = 32'b11111111111111111101111001010111;
assign LUT_1[58214] = 32'b00000000000000000000010101101100;
assign LUT_1[58215] = 32'b11111111111111111001100111101000;
assign LUT_1[58216] = 32'b11111111111111111011111011111001;
assign LUT_1[58217] = 32'b11111111111111110101001101110101;
assign LUT_1[58218] = 32'b11111111111111110111101010001010;
assign LUT_1[58219] = 32'b11111111111111110000111100000110;
assign LUT_1[58220] = 32'b00000000000000000011110101010000;
assign LUT_1[58221] = 32'b11111111111111111101000111001100;
assign LUT_1[58222] = 32'b11111111111111111111100011100001;
assign LUT_1[58223] = 32'b11111111111111111000110101011101;
assign LUT_1[58224] = 32'b11111111111111111110101001100110;
assign LUT_1[58225] = 32'b11111111111111110111111011100010;
assign LUT_1[58226] = 32'b11111111111111111010010111110111;
assign LUT_1[58227] = 32'b11111111111111110011101001110011;
assign LUT_1[58228] = 32'b00000000000000000110100010111101;
assign LUT_1[58229] = 32'b11111111111111111111110100111001;
assign LUT_1[58230] = 32'b00000000000000000010010001001110;
assign LUT_1[58231] = 32'b11111111111111111011100011001010;
assign LUT_1[58232] = 32'b11111111111111111101110111011011;
assign LUT_1[58233] = 32'b11111111111111110111001001010111;
assign LUT_1[58234] = 32'b11111111111111111001100101101100;
assign LUT_1[58235] = 32'b11111111111111110010110111101000;
assign LUT_1[58236] = 32'b00000000000000000101110000110010;
assign LUT_1[58237] = 32'b11111111111111111111000010101110;
assign LUT_1[58238] = 32'b00000000000000000001011111000011;
assign LUT_1[58239] = 32'b11111111111111111010110000111111;
assign LUT_1[58240] = 32'b11111111111111111100110101100000;
assign LUT_1[58241] = 32'b11111111111111110110000111011100;
assign LUT_1[58242] = 32'b11111111111111111000100011110001;
assign LUT_1[58243] = 32'b11111111111111110001110101101101;
assign LUT_1[58244] = 32'b00000000000000000100101110110111;
assign LUT_1[58245] = 32'b11111111111111111110000000110011;
assign LUT_1[58246] = 32'b00000000000000000000011101001000;
assign LUT_1[58247] = 32'b11111111111111111001101111000100;
assign LUT_1[58248] = 32'b11111111111111111100000011010101;
assign LUT_1[58249] = 32'b11111111111111110101010101010001;
assign LUT_1[58250] = 32'b11111111111111110111110001100110;
assign LUT_1[58251] = 32'b11111111111111110001000011100010;
assign LUT_1[58252] = 32'b00000000000000000011111100101100;
assign LUT_1[58253] = 32'b11111111111111111101001110101000;
assign LUT_1[58254] = 32'b11111111111111111111101010111101;
assign LUT_1[58255] = 32'b11111111111111111000111100111001;
assign LUT_1[58256] = 32'b11111111111111111110110001000010;
assign LUT_1[58257] = 32'b11111111111111111000000010111110;
assign LUT_1[58258] = 32'b11111111111111111010011111010011;
assign LUT_1[58259] = 32'b11111111111111110011110001001111;
assign LUT_1[58260] = 32'b00000000000000000110101010011001;
assign LUT_1[58261] = 32'b11111111111111111111111100010101;
assign LUT_1[58262] = 32'b00000000000000000010011000101010;
assign LUT_1[58263] = 32'b11111111111111111011101010100110;
assign LUT_1[58264] = 32'b11111111111111111101111110110111;
assign LUT_1[58265] = 32'b11111111111111110111010000110011;
assign LUT_1[58266] = 32'b11111111111111111001101101001000;
assign LUT_1[58267] = 32'b11111111111111110010111111000100;
assign LUT_1[58268] = 32'b00000000000000000101111000001110;
assign LUT_1[58269] = 32'b11111111111111111111001010001010;
assign LUT_1[58270] = 32'b00000000000000000001100110011111;
assign LUT_1[58271] = 32'b11111111111111111010111000011011;
assign LUT_1[58272] = 32'b11111111111111111101110000011111;
assign LUT_1[58273] = 32'b11111111111111110111000010011011;
assign LUT_1[58274] = 32'b11111111111111111001011110110000;
assign LUT_1[58275] = 32'b11111111111111110010110000101100;
assign LUT_1[58276] = 32'b00000000000000000101101001110110;
assign LUT_1[58277] = 32'b11111111111111111110111011110010;
assign LUT_1[58278] = 32'b00000000000000000001011000000111;
assign LUT_1[58279] = 32'b11111111111111111010101010000011;
assign LUT_1[58280] = 32'b11111111111111111100111110010100;
assign LUT_1[58281] = 32'b11111111111111110110010000010000;
assign LUT_1[58282] = 32'b11111111111111111000101100100101;
assign LUT_1[58283] = 32'b11111111111111110001111110100001;
assign LUT_1[58284] = 32'b00000000000000000100110111101011;
assign LUT_1[58285] = 32'b11111111111111111110001001100111;
assign LUT_1[58286] = 32'b00000000000000000000100101111100;
assign LUT_1[58287] = 32'b11111111111111111001110111111000;
assign LUT_1[58288] = 32'b11111111111111111111101100000001;
assign LUT_1[58289] = 32'b11111111111111111000111101111101;
assign LUT_1[58290] = 32'b11111111111111111011011010010010;
assign LUT_1[58291] = 32'b11111111111111110100101100001110;
assign LUT_1[58292] = 32'b00000000000000000111100101011000;
assign LUT_1[58293] = 32'b00000000000000000000110111010100;
assign LUT_1[58294] = 32'b00000000000000000011010011101001;
assign LUT_1[58295] = 32'b11111111111111111100100101100101;
assign LUT_1[58296] = 32'b11111111111111111110111001110110;
assign LUT_1[58297] = 32'b11111111111111111000001011110010;
assign LUT_1[58298] = 32'b11111111111111111010101000000111;
assign LUT_1[58299] = 32'b11111111111111110011111010000011;
assign LUT_1[58300] = 32'b00000000000000000110110011001101;
assign LUT_1[58301] = 32'b00000000000000000000000101001001;
assign LUT_1[58302] = 32'b00000000000000000010100001011110;
assign LUT_1[58303] = 32'b11111111111111111011110011011010;
assign LUT_1[58304] = 32'b11111111111111111110110011001000;
assign LUT_1[58305] = 32'b11111111111111111000000101000100;
assign LUT_1[58306] = 32'b11111111111111111010100001011001;
assign LUT_1[58307] = 32'b11111111111111110011110011010101;
assign LUT_1[58308] = 32'b00000000000000000110101100011111;
assign LUT_1[58309] = 32'b11111111111111111111111110011011;
assign LUT_1[58310] = 32'b00000000000000000010011010110000;
assign LUT_1[58311] = 32'b11111111111111111011101100101100;
assign LUT_1[58312] = 32'b11111111111111111110000000111101;
assign LUT_1[58313] = 32'b11111111111111110111010010111001;
assign LUT_1[58314] = 32'b11111111111111111001101111001110;
assign LUT_1[58315] = 32'b11111111111111110011000001001010;
assign LUT_1[58316] = 32'b00000000000000000101111010010100;
assign LUT_1[58317] = 32'b11111111111111111111001100010000;
assign LUT_1[58318] = 32'b00000000000000000001101000100101;
assign LUT_1[58319] = 32'b11111111111111111010111010100001;
assign LUT_1[58320] = 32'b00000000000000000000101110101010;
assign LUT_1[58321] = 32'b11111111111111111010000000100110;
assign LUT_1[58322] = 32'b11111111111111111100011100111011;
assign LUT_1[58323] = 32'b11111111111111110101101110110111;
assign LUT_1[58324] = 32'b00000000000000001000101000000001;
assign LUT_1[58325] = 32'b00000000000000000001111001111101;
assign LUT_1[58326] = 32'b00000000000000000100010110010010;
assign LUT_1[58327] = 32'b11111111111111111101101000001110;
assign LUT_1[58328] = 32'b11111111111111111111111100011111;
assign LUT_1[58329] = 32'b11111111111111111001001110011011;
assign LUT_1[58330] = 32'b11111111111111111011101010110000;
assign LUT_1[58331] = 32'b11111111111111110100111100101100;
assign LUT_1[58332] = 32'b00000000000000000111110101110110;
assign LUT_1[58333] = 32'b00000000000000000001000111110010;
assign LUT_1[58334] = 32'b00000000000000000011100100000111;
assign LUT_1[58335] = 32'b11111111111111111100110110000011;
assign LUT_1[58336] = 32'b11111111111111111111101110000111;
assign LUT_1[58337] = 32'b11111111111111111001000000000011;
assign LUT_1[58338] = 32'b11111111111111111011011100011000;
assign LUT_1[58339] = 32'b11111111111111110100101110010100;
assign LUT_1[58340] = 32'b00000000000000000111100111011110;
assign LUT_1[58341] = 32'b00000000000000000000111001011010;
assign LUT_1[58342] = 32'b00000000000000000011010101101111;
assign LUT_1[58343] = 32'b11111111111111111100100111101011;
assign LUT_1[58344] = 32'b11111111111111111110111011111100;
assign LUT_1[58345] = 32'b11111111111111111000001101111000;
assign LUT_1[58346] = 32'b11111111111111111010101010001101;
assign LUT_1[58347] = 32'b11111111111111110011111100001001;
assign LUT_1[58348] = 32'b00000000000000000110110101010011;
assign LUT_1[58349] = 32'b00000000000000000000000111001111;
assign LUT_1[58350] = 32'b00000000000000000010100011100100;
assign LUT_1[58351] = 32'b11111111111111111011110101100000;
assign LUT_1[58352] = 32'b00000000000000000001101001101001;
assign LUT_1[58353] = 32'b11111111111111111010111011100101;
assign LUT_1[58354] = 32'b11111111111111111101010111111010;
assign LUT_1[58355] = 32'b11111111111111110110101001110110;
assign LUT_1[58356] = 32'b00000000000000001001100011000000;
assign LUT_1[58357] = 32'b00000000000000000010110100111100;
assign LUT_1[58358] = 32'b00000000000000000101010001010001;
assign LUT_1[58359] = 32'b11111111111111111110100011001101;
assign LUT_1[58360] = 32'b00000000000000000000110111011110;
assign LUT_1[58361] = 32'b11111111111111111010001001011010;
assign LUT_1[58362] = 32'b11111111111111111100100101101111;
assign LUT_1[58363] = 32'b11111111111111110101110111101011;
assign LUT_1[58364] = 32'b00000000000000001000110000110101;
assign LUT_1[58365] = 32'b00000000000000000010000010110001;
assign LUT_1[58366] = 32'b00000000000000000100011111000110;
assign LUT_1[58367] = 32'b11111111111111111101110001000010;
assign LUT_1[58368] = 32'b00000000000000001000101001100100;
assign LUT_1[58369] = 32'b00000000000000000001111011100000;
assign LUT_1[58370] = 32'b00000000000000000100010111110101;
assign LUT_1[58371] = 32'b11111111111111111101101001110001;
assign LUT_1[58372] = 32'b00000000000000010000100010111011;
assign LUT_1[58373] = 32'b00000000000000001001110100110111;
assign LUT_1[58374] = 32'b00000000000000001100010001001100;
assign LUT_1[58375] = 32'b00000000000000000101100011001000;
assign LUT_1[58376] = 32'b00000000000000000111110111011001;
assign LUT_1[58377] = 32'b00000000000000000001001001010101;
assign LUT_1[58378] = 32'b00000000000000000011100101101010;
assign LUT_1[58379] = 32'b11111111111111111100110111100110;
assign LUT_1[58380] = 32'b00000000000000001111110000110000;
assign LUT_1[58381] = 32'b00000000000000001001000010101100;
assign LUT_1[58382] = 32'b00000000000000001011011111000001;
assign LUT_1[58383] = 32'b00000000000000000100110000111101;
assign LUT_1[58384] = 32'b00000000000000001010100101000110;
assign LUT_1[58385] = 32'b00000000000000000011110111000010;
assign LUT_1[58386] = 32'b00000000000000000110010011010111;
assign LUT_1[58387] = 32'b11111111111111111111100101010011;
assign LUT_1[58388] = 32'b00000000000000010010011110011101;
assign LUT_1[58389] = 32'b00000000000000001011110000011001;
assign LUT_1[58390] = 32'b00000000000000001110001100101110;
assign LUT_1[58391] = 32'b00000000000000000111011110101010;
assign LUT_1[58392] = 32'b00000000000000001001110010111011;
assign LUT_1[58393] = 32'b00000000000000000011000100110111;
assign LUT_1[58394] = 32'b00000000000000000101100001001100;
assign LUT_1[58395] = 32'b11111111111111111110110011001000;
assign LUT_1[58396] = 32'b00000000000000010001101100010010;
assign LUT_1[58397] = 32'b00000000000000001010111110001110;
assign LUT_1[58398] = 32'b00000000000000001101011010100011;
assign LUT_1[58399] = 32'b00000000000000000110101100011111;
assign LUT_1[58400] = 32'b00000000000000001001100100100011;
assign LUT_1[58401] = 32'b00000000000000000010110110011111;
assign LUT_1[58402] = 32'b00000000000000000101010010110100;
assign LUT_1[58403] = 32'b11111111111111111110100100110000;
assign LUT_1[58404] = 32'b00000000000000010001011101111010;
assign LUT_1[58405] = 32'b00000000000000001010101111110110;
assign LUT_1[58406] = 32'b00000000000000001101001100001011;
assign LUT_1[58407] = 32'b00000000000000000110011110000111;
assign LUT_1[58408] = 32'b00000000000000001000110010011000;
assign LUT_1[58409] = 32'b00000000000000000010000100010100;
assign LUT_1[58410] = 32'b00000000000000000100100000101001;
assign LUT_1[58411] = 32'b11111111111111111101110010100101;
assign LUT_1[58412] = 32'b00000000000000010000101011101111;
assign LUT_1[58413] = 32'b00000000000000001001111101101011;
assign LUT_1[58414] = 32'b00000000000000001100011010000000;
assign LUT_1[58415] = 32'b00000000000000000101101011111100;
assign LUT_1[58416] = 32'b00000000000000001011100000000101;
assign LUT_1[58417] = 32'b00000000000000000100110010000001;
assign LUT_1[58418] = 32'b00000000000000000111001110010110;
assign LUT_1[58419] = 32'b00000000000000000000100000010010;
assign LUT_1[58420] = 32'b00000000000000010011011001011100;
assign LUT_1[58421] = 32'b00000000000000001100101011011000;
assign LUT_1[58422] = 32'b00000000000000001111000111101101;
assign LUT_1[58423] = 32'b00000000000000001000011001101001;
assign LUT_1[58424] = 32'b00000000000000001010101101111010;
assign LUT_1[58425] = 32'b00000000000000000011111111110110;
assign LUT_1[58426] = 32'b00000000000000000110011100001011;
assign LUT_1[58427] = 32'b11111111111111111111101110000111;
assign LUT_1[58428] = 32'b00000000000000010010100111010001;
assign LUT_1[58429] = 32'b00000000000000001011111001001101;
assign LUT_1[58430] = 32'b00000000000000001110010101100010;
assign LUT_1[58431] = 32'b00000000000000000111100111011110;
assign LUT_1[58432] = 32'b00000000000000001010100111001100;
assign LUT_1[58433] = 32'b00000000000000000011111001001000;
assign LUT_1[58434] = 32'b00000000000000000110010101011101;
assign LUT_1[58435] = 32'b11111111111111111111100111011001;
assign LUT_1[58436] = 32'b00000000000000010010100000100011;
assign LUT_1[58437] = 32'b00000000000000001011110010011111;
assign LUT_1[58438] = 32'b00000000000000001110001110110100;
assign LUT_1[58439] = 32'b00000000000000000111100000110000;
assign LUT_1[58440] = 32'b00000000000000001001110101000001;
assign LUT_1[58441] = 32'b00000000000000000011000110111101;
assign LUT_1[58442] = 32'b00000000000000000101100011010010;
assign LUT_1[58443] = 32'b11111111111111111110110101001110;
assign LUT_1[58444] = 32'b00000000000000010001101110011000;
assign LUT_1[58445] = 32'b00000000000000001011000000010100;
assign LUT_1[58446] = 32'b00000000000000001101011100101001;
assign LUT_1[58447] = 32'b00000000000000000110101110100101;
assign LUT_1[58448] = 32'b00000000000000001100100010101110;
assign LUT_1[58449] = 32'b00000000000000000101110100101010;
assign LUT_1[58450] = 32'b00000000000000001000010000111111;
assign LUT_1[58451] = 32'b00000000000000000001100010111011;
assign LUT_1[58452] = 32'b00000000000000010100011100000101;
assign LUT_1[58453] = 32'b00000000000000001101101110000001;
assign LUT_1[58454] = 32'b00000000000000010000001010010110;
assign LUT_1[58455] = 32'b00000000000000001001011100010010;
assign LUT_1[58456] = 32'b00000000000000001011110000100011;
assign LUT_1[58457] = 32'b00000000000000000101000010011111;
assign LUT_1[58458] = 32'b00000000000000000111011110110100;
assign LUT_1[58459] = 32'b00000000000000000000110000110000;
assign LUT_1[58460] = 32'b00000000000000010011101001111010;
assign LUT_1[58461] = 32'b00000000000000001100111011110110;
assign LUT_1[58462] = 32'b00000000000000001111011000001011;
assign LUT_1[58463] = 32'b00000000000000001000101010000111;
assign LUT_1[58464] = 32'b00000000000000001011100010001011;
assign LUT_1[58465] = 32'b00000000000000000100110100000111;
assign LUT_1[58466] = 32'b00000000000000000111010000011100;
assign LUT_1[58467] = 32'b00000000000000000000100010011000;
assign LUT_1[58468] = 32'b00000000000000010011011011100010;
assign LUT_1[58469] = 32'b00000000000000001100101101011110;
assign LUT_1[58470] = 32'b00000000000000001111001001110011;
assign LUT_1[58471] = 32'b00000000000000001000011011101111;
assign LUT_1[58472] = 32'b00000000000000001010110000000000;
assign LUT_1[58473] = 32'b00000000000000000100000001111100;
assign LUT_1[58474] = 32'b00000000000000000110011110010001;
assign LUT_1[58475] = 32'b11111111111111111111110000001101;
assign LUT_1[58476] = 32'b00000000000000010010101001010111;
assign LUT_1[58477] = 32'b00000000000000001011111011010011;
assign LUT_1[58478] = 32'b00000000000000001110010111101000;
assign LUT_1[58479] = 32'b00000000000000000111101001100100;
assign LUT_1[58480] = 32'b00000000000000001101011101101101;
assign LUT_1[58481] = 32'b00000000000000000110101111101001;
assign LUT_1[58482] = 32'b00000000000000001001001011111110;
assign LUT_1[58483] = 32'b00000000000000000010011101111010;
assign LUT_1[58484] = 32'b00000000000000010101010111000100;
assign LUT_1[58485] = 32'b00000000000000001110101001000000;
assign LUT_1[58486] = 32'b00000000000000010001000101010101;
assign LUT_1[58487] = 32'b00000000000000001010010111010001;
assign LUT_1[58488] = 32'b00000000000000001100101011100010;
assign LUT_1[58489] = 32'b00000000000000000101111101011110;
assign LUT_1[58490] = 32'b00000000000000001000011001110011;
assign LUT_1[58491] = 32'b00000000000000000001101011101111;
assign LUT_1[58492] = 32'b00000000000000010100100100111001;
assign LUT_1[58493] = 32'b00000000000000001101110110110101;
assign LUT_1[58494] = 32'b00000000000000010000010011001010;
assign LUT_1[58495] = 32'b00000000000000001001100101000110;
assign LUT_1[58496] = 32'b00000000000000001011101001100111;
assign LUT_1[58497] = 32'b00000000000000000100111011100011;
assign LUT_1[58498] = 32'b00000000000000000111010111111000;
assign LUT_1[58499] = 32'b00000000000000000000101001110100;
assign LUT_1[58500] = 32'b00000000000000010011100010111110;
assign LUT_1[58501] = 32'b00000000000000001100110100111010;
assign LUT_1[58502] = 32'b00000000000000001111010001001111;
assign LUT_1[58503] = 32'b00000000000000001000100011001011;
assign LUT_1[58504] = 32'b00000000000000001010110111011100;
assign LUT_1[58505] = 32'b00000000000000000100001001011000;
assign LUT_1[58506] = 32'b00000000000000000110100101101101;
assign LUT_1[58507] = 32'b11111111111111111111110111101001;
assign LUT_1[58508] = 32'b00000000000000010010110000110011;
assign LUT_1[58509] = 32'b00000000000000001100000010101111;
assign LUT_1[58510] = 32'b00000000000000001110011111000100;
assign LUT_1[58511] = 32'b00000000000000000111110001000000;
assign LUT_1[58512] = 32'b00000000000000001101100101001001;
assign LUT_1[58513] = 32'b00000000000000000110110111000101;
assign LUT_1[58514] = 32'b00000000000000001001010011011010;
assign LUT_1[58515] = 32'b00000000000000000010100101010110;
assign LUT_1[58516] = 32'b00000000000000010101011110100000;
assign LUT_1[58517] = 32'b00000000000000001110110000011100;
assign LUT_1[58518] = 32'b00000000000000010001001100110001;
assign LUT_1[58519] = 32'b00000000000000001010011110101101;
assign LUT_1[58520] = 32'b00000000000000001100110010111110;
assign LUT_1[58521] = 32'b00000000000000000110000100111010;
assign LUT_1[58522] = 32'b00000000000000001000100001001111;
assign LUT_1[58523] = 32'b00000000000000000001110011001011;
assign LUT_1[58524] = 32'b00000000000000010100101100010101;
assign LUT_1[58525] = 32'b00000000000000001101111110010001;
assign LUT_1[58526] = 32'b00000000000000010000011010100110;
assign LUT_1[58527] = 32'b00000000000000001001101100100010;
assign LUT_1[58528] = 32'b00000000000000001100100100100110;
assign LUT_1[58529] = 32'b00000000000000000101110110100010;
assign LUT_1[58530] = 32'b00000000000000001000010010110111;
assign LUT_1[58531] = 32'b00000000000000000001100100110011;
assign LUT_1[58532] = 32'b00000000000000010100011101111101;
assign LUT_1[58533] = 32'b00000000000000001101101111111001;
assign LUT_1[58534] = 32'b00000000000000010000001100001110;
assign LUT_1[58535] = 32'b00000000000000001001011110001010;
assign LUT_1[58536] = 32'b00000000000000001011110010011011;
assign LUT_1[58537] = 32'b00000000000000000101000100010111;
assign LUT_1[58538] = 32'b00000000000000000111100000101100;
assign LUT_1[58539] = 32'b00000000000000000000110010101000;
assign LUT_1[58540] = 32'b00000000000000010011101011110010;
assign LUT_1[58541] = 32'b00000000000000001100111101101110;
assign LUT_1[58542] = 32'b00000000000000001111011010000011;
assign LUT_1[58543] = 32'b00000000000000001000101011111111;
assign LUT_1[58544] = 32'b00000000000000001110100000001000;
assign LUT_1[58545] = 32'b00000000000000000111110010000100;
assign LUT_1[58546] = 32'b00000000000000001010001110011001;
assign LUT_1[58547] = 32'b00000000000000000011100000010101;
assign LUT_1[58548] = 32'b00000000000000010110011001011111;
assign LUT_1[58549] = 32'b00000000000000001111101011011011;
assign LUT_1[58550] = 32'b00000000000000010010000111110000;
assign LUT_1[58551] = 32'b00000000000000001011011001101100;
assign LUT_1[58552] = 32'b00000000000000001101101101111101;
assign LUT_1[58553] = 32'b00000000000000000110111111111001;
assign LUT_1[58554] = 32'b00000000000000001001011100001110;
assign LUT_1[58555] = 32'b00000000000000000010101110001010;
assign LUT_1[58556] = 32'b00000000000000010101100111010100;
assign LUT_1[58557] = 32'b00000000000000001110111001010000;
assign LUT_1[58558] = 32'b00000000000000010001010101100101;
assign LUT_1[58559] = 32'b00000000000000001010100111100001;
assign LUT_1[58560] = 32'b00000000000000001101100111001111;
assign LUT_1[58561] = 32'b00000000000000000110111001001011;
assign LUT_1[58562] = 32'b00000000000000001001010101100000;
assign LUT_1[58563] = 32'b00000000000000000010100111011100;
assign LUT_1[58564] = 32'b00000000000000010101100000100110;
assign LUT_1[58565] = 32'b00000000000000001110110010100010;
assign LUT_1[58566] = 32'b00000000000000010001001110110111;
assign LUT_1[58567] = 32'b00000000000000001010100000110011;
assign LUT_1[58568] = 32'b00000000000000001100110101000100;
assign LUT_1[58569] = 32'b00000000000000000110000111000000;
assign LUT_1[58570] = 32'b00000000000000001000100011010101;
assign LUT_1[58571] = 32'b00000000000000000001110101010001;
assign LUT_1[58572] = 32'b00000000000000010100101110011011;
assign LUT_1[58573] = 32'b00000000000000001110000000010111;
assign LUT_1[58574] = 32'b00000000000000010000011100101100;
assign LUT_1[58575] = 32'b00000000000000001001101110101000;
assign LUT_1[58576] = 32'b00000000000000001111100010110001;
assign LUT_1[58577] = 32'b00000000000000001000110100101101;
assign LUT_1[58578] = 32'b00000000000000001011010001000010;
assign LUT_1[58579] = 32'b00000000000000000100100010111110;
assign LUT_1[58580] = 32'b00000000000000010111011100001000;
assign LUT_1[58581] = 32'b00000000000000010000101110000100;
assign LUT_1[58582] = 32'b00000000000000010011001010011001;
assign LUT_1[58583] = 32'b00000000000000001100011100010101;
assign LUT_1[58584] = 32'b00000000000000001110110000100110;
assign LUT_1[58585] = 32'b00000000000000001000000010100010;
assign LUT_1[58586] = 32'b00000000000000001010011110110111;
assign LUT_1[58587] = 32'b00000000000000000011110000110011;
assign LUT_1[58588] = 32'b00000000000000010110101001111101;
assign LUT_1[58589] = 32'b00000000000000001111111011111001;
assign LUT_1[58590] = 32'b00000000000000010010011000001110;
assign LUT_1[58591] = 32'b00000000000000001011101010001010;
assign LUT_1[58592] = 32'b00000000000000001110100010001110;
assign LUT_1[58593] = 32'b00000000000000000111110100001010;
assign LUT_1[58594] = 32'b00000000000000001010010000011111;
assign LUT_1[58595] = 32'b00000000000000000011100010011011;
assign LUT_1[58596] = 32'b00000000000000010110011011100101;
assign LUT_1[58597] = 32'b00000000000000001111101101100001;
assign LUT_1[58598] = 32'b00000000000000010010001001110110;
assign LUT_1[58599] = 32'b00000000000000001011011011110010;
assign LUT_1[58600] = 32'b00000000000000001101110000000011;
assign LUT_1[58601] = 32'b00000000000000000111000001111111;
assign LUT_1[58602] = 32'b00000000000000001001011110010100;
assign LUT_1[58603] = 32'b00000000000000000010110000010000;
assign LUT_1[58604] = 32'b00000000000000010101101001011010;
assign LUT_1[58605] = 32'b00000000000000001110111011010110;
assign LUT_1[58606] = 32'b00000000000000010001010111101011;
assign LUT_1[58607] = 32'b00000000000000001010101001100111;
assign LUT_1[58608] = 32'b00000000000000010000011101110000;
assign LUT_1[58609] = 32'b00000000000000001001101111101100;
assign LUT_1[58610] = 32'b00000000000000001100001100000001;
assign LUT_1[58611] = 32'b00000000000000000101011101111101;
assign LUT_1[58612] = 32'b00000000000000011000010111000111;
assign LUT_1[58613] = 32'b00000000000000010001101001000011;
assign LUT_1[58614] = 32'b00000000000000010100000101011000;
assign LUT_1[58615] = 32'b00000000000000001101010111010100;
assign LUT_1[58616] = 32'b00000000000000001111101011100101;
assign LUT_1[58617] = 32'b00000000000000001000111101100001;
assign LUT_1[58618] = 32'b00000000000000001011011001110110;
assign LUT_1[58619] = 32'b00000000000000000100101011110010;
assign LUT_1[58620] = 32'b00000000000000010111100100111100;
assign LUT_1[58621] = 32'b00000000000000010000110110111000;
assign LUT_1[58622] = 32'b00000000000000010011010011001101;
assign LUT_1[58623] = 32'b00000000000000001100100101001001;
assign LUT_1[58624] = 32'b00000000000000000110011101110000;
assign LUT_1[58625] = 32'b11111111111111111111101111101100;
assign LUT_1[58626] = 32'b00000000000000000010001100000001;
assign LUT_1[58627] = 32'b11111111111111111011011101111101;
assign LUT_1[58628] = 32'b00000000000000001110010111000111;
assign LUT_1[58629] = 32'b00000000000000000111101001000011;
assign LUT_1[58630] = 32'b00000000000000001010000101011000;
assign LUT_1[58631] = 32'b00000000000000000011010111010100;
assign LUT_1[58632] = 32'b00000000000000000101101011100101;
assign LUT_1[58633] = 32'b11111111111111111110111101100001;
assign LUT_1[58634] = 32'b00000000000000000001011001110110;
assign LUT_1[58635] = 32'b11111111111111111010101011110010;
assign LUT_1[58636] = 32'b00000000000000001101100100111100;
assign LUT_1[58637] = 32'b00000000000000000110110110111000;
assign LUT_1[58638] = 32'b00000000000000001001010011001101;
assign LUT_1[58639] = 32'b00000000000000000010100101001001;
assign LUT_1[58640] = 32'b00000000000000001000011001010010;
assign LUT_1[58641] = 32'b00000000000000000001101011001110;
assign LUT_1[58642] = 32'b00000000000000000100000111100011;
assign LUT_1[58643] = 32'b11111111111111111101011001011111;
assign LUT_1[58644] = 32'b00000000000000010000010010101001;
assign LUT_1[58645] = 32'b00000000000000001001100100100101;
assign LUT_1[58646] = 32'b00000000000000001100000000111010;
assign LUT_1[58647] = 32'b00000000000000000101010010110110;
assign LUT_1[58648] = 32'b00000000000000000111100111000111;
assign LUT_1[58649] = 32'b00000000000000000000111001000011;
assign LUT_1[58650] = 32'b00000000000000000011010101011000;
assign LUT_1[58651] = 32'b11111111111111111100100111010100;
assign LUT_1[58652] = 32'b00000000000000001111100000011110;
assign LUT_1[58653] = 32'b00000000000000001000110010011010;
assign LUT_1[58654] = 32'b00000000000000001011001110101111;
assign LUT_1[58655] = 32'b00000000000000000100100000101011;
assign LUT_1[58656] = 32'b00000000000000000111011000101111;
assign LUT_1[58657] = 32'b00000000000000000000101010101011;
assign LUT_1[58658] = 32'b00000000000000000011000111000000;
assign LUT_1[58659] = 32'b11111111111111111100011000111100;
assign LUT_1[58660] = 32'b00000000000000001111010010000110;
assign LUT_1[58661] = 32'b00000000000000001000100100000010;
assign LUT_1[58662] = 32'b00000000000000001011000000010111;
assign LUT_1[58663] = 32'b00000000000000000100010010010011;
assign LUT_1[58664] = 32'b00000000000000000110100110100100;
assign LUT_1[58665] = 32'b11111111111111111111111000100000;
assign LUT_1[58666] = 32'b00000000000000000010010100110101;
assign LUT_1[58667] = 32'b11111111111111111011100110110001;
assign LUT_1[58668] = 32'b00000000000000001110011111111011;
assign LUT_1[58669] = 32'b00000000000000000111110001110111;
assign LUT_1[58670] = 32'b00000000000000001010001110001100;
assign LUT_1[58671] = 32'b00000000000000000011100000001000;
assign LUT_1[58672] = 32'b00000000000000001001010100010001;
assign LUT_1[58673] = 32'b00000000000000000010100110001101;
assign LUT_1[58674] = 32'b00000000000000000101000010100010;
assign LUT_1[58675] = 32'b11111111111111111110010100011110;
assign LUT_1[58676] = 32'b00000000000000010001001101101000;
assign LUT_1[58677] = 32'b00000000000000001010011111100100;
assign LUT_1[58678] = 32'b00000000000000001100111011111001;
assign LUT_1[58679] = 32'b00000000000000000110001101110101;
assign LUT_1[58680] = 32'b00000000000000001000100010000110;
assign LUT_1[58681] = 32'b00000000000000000001110100000010;
assign LUT_1[58682] = 32'b00000000000000000100010000010111;
assign LUT_1[58683] = 32'b11111111111111111101100010010011;
assign LUT_1[58684] = 32'b00000000000000010000011011011101;
assign LUT_1[58685] = 32'b00000000000000001001101101011001;
assign LUT_1[58686] = 32'b00000000000000001100001001101110;
assign LUT_1[58687] = 32'b00000000000000000101011011101010;
assign LUT_1[58688] = 32'b00000000000000001000011011011000;
assign LUT_1[58689] = 32'b00000000000000000001101101010100;
assign LUT_1[58690] = 32'b00000000000000000100001001101001;
assign LUT_1[58691] = 32'b11111111111111111101011011100101;
assign LUT_1[58692] = 32'b00000000000000010000010100101111;
assign LUT_1[58693] = 32'b00000000000000001001100110101011;
assign LUT_1[58694] = 32'b00000000000000001100000011000000;
assign LUT_1[58695] = 32'b00000000000000000101010100111100;
assign LUT_1[58696] = 32'b00000000000000000111101001001101;
assign LUT_1[58697] = 32'b00000000000000000000111011001001;
assign LUT_1[58698] = 32'b00000000000000000011010111011110;
assign LUT_1[58699] = 32'b11111111111111111100101001011010;
assign LUT_1[58700] = 32'b00000000000000001111100010100100;
assign LUT_1[58701] = 32'b00000000000000001000110100100000;
assign LUT_1[58702] = 32'b00000000000000001011010000110101;
assign LUT_1[58703] = 32'b00000000000000000100100010110001;
assign LUT_1[58704] = 32'b00000000000000001010010110111010;
assign LUT_1[58705] = 32'b00000000000000000011101000110110;
assign LUT_1[58706] = 32'b00000000000000000110000101001011;
assign LUT_1[58707] = 32'b11111111111111111111010111000111;
assign LUT_1[58708] = 32'b00000000000000010010010000010001;
assign LUT_1[58709] = 32'b00000000000000001011100010001101;
assign LUT_1[58710] = 32'b00000000000000001101111110100010;
assign LUT_1[58711] = 32'b00000000000000000111010000011110;
assign LUT_1[58712] = 32'b00000000000000001001100100101111;
assign LUT_1[58713] = 32'b00000000000000000010110110101011;
assign LUT_1[58714] = 32'b00000000000000000101010011000000;
assign LUT_1[58715] = 32'b11111111111111111110100100111100;
assign LUT_1[58716] = 32'b00000000000000010001011110000110;
assign LUT_1[58717] = 32'b00000000000000001010110000000010;
assign LUT_1[58718] = 32'b00000000000000001101001100010111;
assign LUT_1[58719] = 32'b00000000000000000110011110010011;
assign LUT_1[58720] = 32'b00000000000000001001010110010111;
assign LUT_1[58721] = 32'b00000000000000000010101000010011;
assign LUT_1[58722] = 32'b00000000000000000101000100101000;
assign LUT_1[58723] = 32'b11111111111111111110010110100100;
assign LUT_1[58724] = 32'b00000000000000010001001111101110;
assign LUT_1[58725] = 32'b00000000000000001010100001101010;
assign LUT_1[58726] = 32'b00000000000000001100111101111111;
assign LUT_1[58727] = 32'b00000000000000000110001111111011;
assign LUT_1[58728] = 32'b00000000000000001000100100001100;
assign LUT_1[58729] = 32'b00000000000000000001110110001000;
assign LUT_1[58730] = 32'b00000000000000000100010010011101;
assign LUT_1[58731] = 32'b11111111111111111101100100011001;
assign LUT_1[58732] = 32'b00000000000000010000011101100011;
assign LUT_1[58733] = 32'b00000000000000001001101111011111;
assign LUT_1[58734] = 32'b00000000000000001100001011110100;
assign LUT_1[58735] = 32'b00000000000000000101011101110000;
assign LUT_1[58736] = 32'b00000000000000001011010001111001;
assign LUT_1[58737] = 32'b00000000000000000100100011110101;
assign LUT_1[58738] = 32'b00000000000000000111000000001010;
assign LUT_1[58739] = 32'b00000000000000000000010010000110;
assign LUT_1[58740] = 32'b00000000000000010011001011010000;
assign LUT_1[58741] = 32'b00000000000000001100011101001100;
assign LUT_1[58742] = 32'b00000000000000001110111001100001;
assign LUT_1[58743] = 32'b00000000000000001000001011011101;
assign LUT_1[58744] = 32'b00000000000000001010011111101110;
assign LUT_1[58745] = 32'b00000000000000000011110001101010;
assign LUT_1[58746] = 32'b00000000000000000110001101111111;
assign LUT_1[58747] = 32'b11111111111111111111011111111011;
assign LUT_1[58748] = 32'b00000000000000010010011001000101;
assign LUT_1[58749] = 32'b00000000000000001011101011000001;
assign LUT_1[58750] = 32'b00000000000000001110000111010110;
assign LUT_1[58751] = 32'b00000000000000000111011001010010;
assign LUT_1[58752] = 32'b00000000000000001001011101110011;
assign LUT_1[58753] = 32'b00000000000000000010101111101111;
assign LUT_1[58754] = 32'b00000000000000000101001100000100;
assign LUT_1[58755] = 32'b11111111111111111110011110000000;
assign LUT_1[58756] = 32'b00000000000000010001010111001010;
assign LUT_1[58757] = 32'b00000000000000001010101001000110;
assign LUT_1[58758] = 32'b00000000000000001101000101011011;
assign LUT_1[58759] = 32'b00000000000000000110010111010111;
assign LUT_1[58760] = 32'b00000000000000001000101011101000;
assign LUT_1[58761] = 32'b00000000000000000001111101100100;
assign LUT_1[58762] = 32'b00000000000000000100011001111001;
assign LUT_1[58763] = 32'b11111111111111111101101011110101;
assign LUT_1[58764] = 32'b00000000000000010000100100111111;
assign LUT_1[58765] = 32'b00000000000000001001110110111011;
assign LUT_1[58766] = 32'b00000000000000001100010011010000;
assign LUT_1[58767] = 32'b00000000000000000101100101001100;
assign LUT_1[58768] = 32'b00000000000000001011011001010101;
assign LUT_1[58769] = 32'b00000000000000000100101011010001;
assign LUT_1[58770] = 32'b00000000000000000111000111100110;
assign LUT_1[58771] = 32'b00000000000000000000011001100010;
assign LUT_1[58772] = 32'b00000000000000010011010010101100;
assign LUT_1[58773] = 32'b00000000000000001100100100101000;
assign LUT_1[58774] = 32'b00000000000000001111000000111101;
assign LUT_1[58775] = 32'b00000000000000001000010010111001;
assign LUT_1[58776] = 32'b00000000000000001010100111001010;
assign LUT_1[58777] = 32'b00000000000000000011111001000110;
assign LUT_1[58778] = 32'b00000000000000000110010101011011;
assign LUT_1[58779] = 32'b11111111111111111111100111010111;
assign LUT_1[58780] = 32'b00000000000000010010100000100001;
assign LUT_1[58781] = 32'b00000000000000001011110010011101;
assign LUT_1[58782] = 32'b00000000000000001110001110110010;
assign LUT_1[58783] = 32'b00000000000000000111100000101110;
assign LUT_1[58784] = 32'b00000000000000001010011000110010;
assign LUT_1[58785] = 32'b00000000000000000011101010101110;
assign LUT_1[58786] = 32'b00000000000000000110000111000011;
assign LUT_1[58787] = 32'b11111111111111111111011000111111;
assign LUT_1[58788] = 32'b00000000000000010010010010001001;
assign LUT_1[58789] = 32'b00000000000000001011100100000101;
assign LUT_1[58790] = 32'b00000000000000001110000000011010;
assign LUT_1[58791] = 32'b00000000000000000111010010010110;
assign LUT_1[58792] = 32'b00000000000000001001100110100111;
assign LUT_1[58793] = 32'b00000000000000000010111000100011;
assign LUT_1[58794] = 32'b00000000000000000101010100111000;
assign LUT_1[58795] = 32'b11111111111111111110100110110100;
assign LUT_1[58796] = 32'b00000000000000010001011111111110;
assign LUT_1[58797] = 32'b00000000000000001010110001111010;
assign LUT_1[58798] = 32'b00000000000000001101001110001111;
assign LUT_1[58799] = 32'b00000000000000000110100000001011;
assign LUT_1[58800] = 32'b00000000000000001100010100010100;
assign LUT_1[58801] = 32'b00000000000000000101100110010000;
assign LUT_1[58802] = 32'b00000000000000001000000010100101;
assign LUT_1[58803] = 32'b00000000000000000001010100100001;
assign LUT_1[58804] = 32'b00000000000000010100001101101011;
assign LUT_1[58805] = 32'b00000000000000001101011111100111;
assign LUT_1[58806] = 32'b00000000000000001111111011111100;
assign LUT_1[58807] = 32'b00000000000000001001001101111000;
assign LUT_1[58808] = 32'b00000000000000001011100010001001;
assign LUT_1[58809] = 32'b00000000000000000100110100000101;
assign LUT_1[58810] = 32'b00000000000000000111010000011010;
assign LUT_1[58811] = 32'b00000000000000000000100010010110;
assign LUT_1[58812] = 32'b00000000000000010011011011100000;
assign LUT_1[58813] = 32'b00000000000000001100101101011100;
assign LUT_1[58814] = 32'b00000000000000001111001001110001;
assign LUT_1[58815] = 32'b00000000000000001000011011101101;
assign LUT_1[58816] = 32'b00000000000000001011011011011011;
assign LUT_1[58817] = 32'b00000000000000000100101101010111;
assign LUT_1[58818] = 32'b00000000000000000111001001101100;
assign LUT_1[58819] = 32'b00000000000000000000011011101000;
assign LUT_1[58820] = 32'b00000000000000010011010100110010;
assign LUT_1[58821] = 32'b00000000000000001100100110101110;
assign LUT_1[58822] = 32'b00000000000000001111000011000011;
assign LUT_1[58823] = 32'b00000000000000001000010100111111;
assign LUT_1[58824] = 32'b00000000000000001010101001010000;
assign LUT_1[58825] = 32'b00000000000000000011111011001100;
assign LUT_1[58826] = 32'b00000000000000000110010111100001;
assign LUT_1[58827] = 32'b11111111111111111111101001011101;
assign LUT_1[58828] = 32'b00000000000000010010100010100111;
assign LUT_1[58829] = 32'b00000000000000001011110100100011;
assign LUT_1[58830] = 32'b00000000000000001110010000111000;
assign LUT_1[58831] = 32'b00000000000000000111100010110100;
assign LUT_1[58832] = 32'b00000000000000001101010110111101;
assign LUT_1[58833] = 32'b00000000000000000110101000111001;
assign LUT_1[58834] = 32'b00000000000000001001000101001110;
assign LUT_1[58835] = 32'b00000000000000000010010111001010;
assign LUT_1[58836] = 32'b00000000000000010101010000010100;
assign LUT_1[58837] = 32'b00000000000000001110100010010000;
assign LUT_1[58838] = 32'b00000000000000010000111110100101;
assign LUT_1[58839] = 32'b00000000000000001010010000100001;
assign LUT_1[58840] = 32'b00000000000000001100100100110010;
assign LUT_1[58841] = 32'b00000000000000000101110110101110;
assign LUT_1[58842] = 32'b00000000000000001000010011000011;
assign LUT_1[58843] = 32'b00000000000000000001100100111111;
assign LUT_1[58844] = 32'b00000000000000010100011110001001;
assign LUT_1[58845] = 32'b00000000000000001101110000000101;
assign LUT_1[58846] = 32'b00000000000000010000001100011010;
assign LUT_1[58847] = 32'b00000000000000001001011110010110;
assign LUT_1[58848] = 32'b00000000000000001100010110011010;
assign LUT_1[58849] = 32'b00000000000000000101101000010110;
assign LUT_1[58850] = 32'b00000000000000001000000100101011;
assign LUT_1[58851] = 32'b00000000000000000001010110100111;
assign LUT_1[58852] = 32'b00000000000000010100001111110001;
assign LUT_1[58853] = 32'b00000000000000001101100001101101;
assign LUT_1[58854] = 32'b00000000000000001111111110000010;
assign LUT_1[58855] = 32'b00000000000000001001001111111110;
assign LUT_1[58856] = 32'b00000000000000001011100100001111;
assign LUT_1[58857] = 32'b00000000000000000100110110001011;
assign LUT_1[58858] = 32'b00000000000000000111010010100000;
assign LUT_1[58859] = 32'b00000000000000000000100100011100;
assign LUT_1[58860] = 32'b00000000000000010011011101100110;
assign LUT_1[58861] = 32'b00000000000000001100101111100010;
assign LUT_1[58862] = 32'b00000000000000001111001011110111;
assign LUT_1[58863] = 32'b00000000000000001000011101110011;
assign LUT_1[58864] = 32'b00000000000000001110010001111100;
assign LUT_1[58865] = 32'b00000000000000000111100011111000;
assign LUT_1[58866] = 32'b00000000000000001010000000001101;
assign LUT_1[58867] = 32'b00000000000000000011010010001001;
assign LUT_1[58868] = 32'b00000000000000010110001011010011;
assign LUT_1[58869] = 32'b00000000000000001111011101001111;
assign LUT_1[58870] = 32'b00000000000000010001111001100100;
assign LUT_1[58871] = 32'b00000000000000001011001011100000;
assign LUT_1[58872] = 32'b00000000000000001101011111110001;
assign LUT_1[58873] = 32'b00000000000000000110110001101101;
assign LUT_1[58874] = 32'b00000000000000001001001110000010;
assign LUT_1[58875] = 32'b00000000000000000010011111111110;
assign LUT_1[58876] = 32'b00000000000000010101011001001000;
assign LUT_1[58877] = 32'b00000000000000001110101011000100;
assign LUT_1[58878] = 32'b00000000000000010001000111011001;
assign LUT_1[58879] = 32'b00000000000000001010011001010101;
assign LUT_1[58880] = 32'b00000000000000000010011000000001;
assign LUT_1[58881] = 32'b11111111111111111011101001111101;
assign LUT_1[58882] = 32'b11111111111111111110000110010010;
assign LUT_1[58883] = 32'b11111111111111110111011000001110;
assign LUT_1[58884] = 32'b00000000000000001010010001011000;
assign LUT_1[58885] = 32'b00000000000000000011100011010100;
assign LUT_1[58886] = 32'b00000000000000000101111111101001;
assign LUT_1[58887] = 32'b11111111111111111111010001100101;
assign LUT_1[58888] = 32'b00000000000000000001100101110110;
assign LUT_1[58889] = 32'b11111111111111111010110111110010;
assign LUT_1[58890] = 32'b11111111111111111101010100000111;
assign LUT_1[58891] = 32'b11111111111111110110100110000011;
assign LUT_1[58892] = 32'b00000000000000001001011111001101;
assign LUT_1[58893] = 32'b00000000000000000010110001001001;
assign LUT_1[58894] = 32'b00000000000000000101001101011110;
assign LUT_1[58895] = 32'b11111111111111111110011111011010;
assign LUT_1[58896] = 32'b00000000000000000100010011100011;
assign LUT_1[58897] = 32'b11111111111111111101100101011111;
assign LUT_1[58898] = 32'b00000000000000000000000001110100;
assign LUT_1[58899] = 32'b11111111111111111001010011110000;
assign LUT_1[58900] = 32'b00000000000000001100001100111010;
assign LUT_1[58901] = 32'b00000000000000000101011110110110;
assign LUT_1[58902] = 32'b00000000000000000111111011001011;
assign LUT_1[58903] = 32'b00000000000000000001001101000111;
assign LUT_1[58904] = 32'b00000000000000000011100001011000;
assign LUT_1[58905] = 32'b11111111111111111100110011010100;
assign LUT_1[58906] = 32'b11111111111111111111001111101001;
assign LUT_1[58907] = 32'b11111111111111111000100001100101;
assign LUT_1[58908] = 32'b00000000000000001011011010101111;
assign LUT_1[58909] = 32'b00000000000000000100101100101011;
assign LUT_1[58910] = 32'b00000000000000000111001001000000;
assign LUT_1[58911] = 32'b00000000000000000000011010111100;
assign LUT_1[58912] = 32'b00000000000000000011010011000000;
assign LUT_1[58913] = 32'b11111111111111111100100100111100;
assign LUT_1[58914] = 32'b11111111111111111111000001010001;
assign LUT_1[58915] = 32'b11111111111111111000010011001101;
assign LUT_1[58916] = 32'b00000000000000001011001100010111;
assign LUT_1[58917] = 32'b00000000000000000100011110010011;
assign LUT_1[58918] = 32'b00000000000000000110111010101000;
assign LUT_1[58919] = 32'b00000000000000000000001100100100;
assign LUT_1[58920] = 32'b00000000000000000010100000110101;
assign LUT_1[58921] = 32'b11111111111111111011110010110001;
assign LUT_1[58922] = 32'b11111111111111111110001111000110;
assign LUT_1[58923] = 32'b11111111111111110111100001000010;
assign LUT_1[58924] = 32'b00000000000000001010011010001100;
assign LUT_1[58925] = 32'b00000000000000000011101100001000;
assign LUT_1[58926] = 32'b00000000000000000110001000011101;
assign LUT_1[58927] = 32'b11111111111111111111011010011001;
assign LUT_1[58928] = 32'b00000000000000000101001110100010;
assign LUT_1[58929] = 32'b11111111111111111110100000011110;
assign LUT_1[58930] = 32'b00000000000000000000111100110011;
assign LUT_1[58931] = 32'b11111111111111111010001110101111;
assign LUT_1[58932] = 32'b00000000000000001101000111111001;
assign LUT_1[58933] = 32'b00000000000000000110011001110101;
assign LUT_1[58934] = 32'b00000000000000001000110110001010;
assign LUT_1[58935] = 32'b00000000000000000010001000000110;
assign LUT_1[58936] = 32'b00000000000000000100011100010111;
assign LUT_1[58937] = 32'b11111111111111111101101110010011;
assign LUT_1[58938] = 32'b00000000000000000000001010101000;
assign LUT_1[58939] = 32'b11111111111111111001011100100100;
assign LUT_1[58940] = 32'b00000000000000001100010101101110;
assign LUT_1[58941] = 32'b00000000000000000101100111101010;
assign LUT_1[58942] = 32'b00000000000000001000000011111111;
assign LUT_1[58943] = 32'b00000000000000000001010101111011;
assign LUT_1[58944] = 32'b00000000000000000100010101101001;
assign LUT_1[58945] = 32'b11111111111111111101100111100101;
assign LUT_1[58946] = 32'b00000000000000000000000011111010;
assign LUT_1[58947] = 32'b11111111111111111001010101110110;
assign LUT_1[58948] = 32'b00000000000000001100001111000000;
assign LUT_1[58949] = 32'b00000000000000000101100000111100;
assign LUT_1[58950] = 32'b00000000000000000111111101010001;
assign LUT_1[58951] = 32'b00000000000000000001001111001101;
assign LUT_1[58952] = 32'b00000000000000000011100011011110;
assign LUT_1[58953] = 32'b11111111111111111100110101011010;
assign LUT_1[58954] = 32'b11111111111111111111010001101111;
assign LUT_1[58955] = 32'b11111111111111111000100011101011;
assign LUT_1[58956] = 32'b00000000000000001011011100110101;
assign LUT_1[58957] = 32'b00000000000000000100101110110001;
assign LUT_1[58958] = 32'b00000000000000000111001011000110;
assign LUT_1[58959] = 32'b00000000000000000000011101000010;
assign LUT_1[58960] = 32'b00000000000000000110010001001011;
assign LUT_1[58961] = 32'b11111111111111111111100011000111;
assign LUT_1[58962] = 32'b00000000000000000001111111011100;
assign LUT_1[58963] = 32'b11111111111111111011010001011000;
assign LUT_1[58964] = 32'b00000000000000001110001010100010;
assign LUT_1[58965] = 32'b00000000000000000111011100011110;
assign LUT_1[58966] = 32'b00000000000000001001111000110011;
assign LUT_1[58967] = 32'b00000000000000000011001010101111;
assign LUT_1[58968] = 32'b00000000000000000101011111000000;
assign LUT_1[58969] = 32'b11111111111111111110110000111100;
assign LUT_1[58970] = 32'b00000000000000000001001101010001;
assign LUT_1[58971] = 32'b11111111111111111010011111001101;
assign LUT_1[58972] = 32'b00000000000000001101011000010111;
assign LUT_1[58973] = 32'b00000000000000000110101010010011;
assign LUT_1[58974] = 32'b00000000000000001001000110101000;
assign LUT_1[58975] = 32'b00000000000000000010011000100100;
assign LUT_1[58976] = 32'b00000000000000000101010000101000;
assign LUT_1[58977] = 32'b11111111111111111110100010100100;
assign LUT_1[58978] = 32'b00000000000000000000111110111001;
assign LUT_1[58979] = 32'b11111111111111111010010000110101;
assign LUT_1[58980] = 32'b00000000000000001101001001111111;
assign LUT_1[58981] = 32'b00000000000000000110011011111011;
assign LUT_1[58982] = 32'b00000000000000001000111000010000;
assign LUT_1[58983] = 32'b00000000000000000010001010001100;
assign LUT_1[58984] = 32'b00000000000000000100011110011101;
assign LUT_1[58985] = 32'b11111111111111111101110000011001;
assign LUT_1[58986] = 32'b00000000000000000000001100101110;
assign LUT_1[58987] = 32'b11111111111111111001011110101010;
assign LUT_1[58988] = 32'b00000000000000001100010111110100;
assign LUT_1[58989] = 32'b00000000000000000101101001110000;
assign LUT_1[58990] = 32'b00000000000000001000000110000101;
assign LUT_1[58991] = 32'b00000000000000000001011000000001;
assign LUT_1[58992] = 32'b00000000000000000111001100001010;
assign LUT_1[58993] = 32'b00000000000000000000011110000110;
assign LUT_1[58994] = 32'b00000000000000000010111010011011;
assign LUT_1[58995] = 32'b11111111111111111100001100010111;
assign LUT_1[58996] = 32'b00000000000000001111000101100001;
assign LUT_1[58997] = 32'b00000000000000001000010111011101;
assign LUT_1[58998] = 32'b00000000000000001010110011110010;
assign LUT_1[58999] = 32'b00000000000000000100000101101110;
assign LUT_1[59000] = 32'b00000000000000000110011001111111;
assign LUT_1[59001] = 32'b11111111111111111111101011111011;
assign LUT_1[59002] = 32'b00000000000000000010001000010000;
assign LUT_1[59003] = 32'b11111111111111111011011010001100;
assign LUT_1[59004] = 32'b00000000000000001110010011010110;
assign LUT_1[59005] = 32'b00000000000000000111100101010010;
assign LUT_1[59006] = 32'b00000000000000001010000001100111;
assign LUT_1[59007] = 32'b00000000000000000011010011100011;
assign LUT_1[59008] = 32'b00000000000000000101011000000100;
assign LUT_1[59009] = 32'b11111111111111111110101010000000;
assign LUT_1[59010] = 32'b00000000000000000001000110010101;
assign LUT_1[59011] = 32'b11111111111111111010011000010001;
assign LUT_1[59012] = 32'b00000000000000001101010001011011;
assign LUT_1[59013] = 32'b00000000000000000110100011010111;
assign LUT_1[59014] = 32'b00000000000000001000111111101100;
assign LUT_1[59015] = 32'b00000000000000000010010001101000;
assign LUT_1[59016] = 32'b00000000000000000100100101111001;
assign LUT_1[59017] = 32'b11111111111111111101110111110101;
assign LUT_1[59018] = 32'b00000000000000000000010100001010;
assign LUT_1[59019] = 32'b11111111111111111001100110000110;
assign LUT_1[59020] = 32'b00000000000000001100011111010000;
assign LUT_1[59021] = 32'b00000000000000000101110001001100;
assign LUT_1[59022] = 32'b00000000000000001000001101100001;
assign LUT_1[59023] = 32'b00000000000000000001011111011101;
assign LUT_1[59024] = 32'b00000000000000000111010011100110;
assign LUT_1[59025] = 32'b00000000000000000000100101100010;
assign LUT_1[59026] = 32'b00000000000000000011000001110111;
assign LUT_1[59027] = 32'b11111111111111111100010011110011;
assign LUT_1[59028] = 32'b00000000000000001111001100111101;
assign LUT_1[59029] = 32'b00000000000000001000011110111001;
assign LUT_1[59030] = 32'b00000000000000001010111011001110;
assign LUT_1[59031] = 32'b00000000000000000100001101001010;
assign LUT_1[59032] = 32'b00000000000000000110100001011011;
assign LUT_1[59033] = 32'b11111111111111111111110011010111;
assign LUT_1[59034] = 32'b00000000000000000010001111101100;
assign LUT_1[59035] = 32'b11111111111111111011100001101000;
assign LUT_1[59036] = 32'b00000000000000001110011010110010;
assign LUT_1[59037] = 32'b00000000000000000111101100101110;
assign LUT_1[59038] = 32'b00000000000000001010001001000011;
assign LUT_1[59039] = 32'b00000000000000000011011010111111;
assign LUT_1[59040] = 32'b00000000000000000110010011000011;
assign LUT_1[59041] = 32'b11111111111111111111100100111111;
assign LUT_1[59042] = 32'b00000000000000000010000001010100;
assign LUT_1[59043] = 32'b11111111111111111011010011010000;
assign LUT_1[59044] = 32'b00000000000000001110001100011010;
assign LUT_1[59045] = 32'b00000000000000000111011110010110;
assign LUT_1[59046] = 32'b00000000000000001001111010101011;
assign LUT_1[59047] = 32'b00000000000000000011001100100111;
assign LUT_1[59048] = 32'b00000000000000000101100000111000;
assign LUT_1[59049] = 32'b11111111111111111110110010110100;
assign LUT_1[59050] = 32'b00000000000000000001001111001001;
assign LUT_1[59051] = 32'b11111111111111111010100001000101;
assign LUT_1[59052] = 32'b00000000000000001101011010001111;
assign LUT_1[59053] = 32'b00000000000000000110101100001011;
assign LUT_1[59054] = 32'b00000000000000001001001000100000;
assign LUT_1[59055] = 32'b00000000000000000010011010011100;
assign LUT_1[59056] = 32'b00000000000000001000001110100101;
assign LUT_1[59057] = 32'b00000000000000000001100000100001;
assign LUT_1[59058] = 32'b00000000000000000011111100110110;
assign LUT_1[59059] = 32'b11111111111111111101001110110010;
assign LUT_1[59060] = 32'b00000000000000010000000111111100;
assign LUT_1[59061] = 32'b00000000000000001001011001111000;
assign LUT_1[59062] = 32'b00000000000000001011110110001101;
assign LUT_1[59063] = 32'b00000000000000000101001000001001;
assign LUT_1[59064] = 32'b00000000000000000111011100011010;
assign LUT_1[59065] = 32'b00000000000000000000101110010110;
assign LUT_1[59066] = 32'b00000000000000000011001010101011;
assign LUT_1[59067] = 32'b11111111111111111100011100100111;
assign LUT_1[59068] = 32'b00000000000000001111010101110001;
assign LUT_1[59069] = 32'b00000000000000001000100111101101;
assign LUT_1[59070] = 32'b00000000000000001011000100000010;
assign LUT_1[59071] = 32'b00000000000000000100010101111110;
assign LUT_1[59072] = 32'b00000000000000000111010101101100;
assign LUT_1[59073] = 32'b00000000000000000000100111101000;
assign LUT_1[59074] = 32'b00000000000000000011000011111101;
assign LUT_1[59075] = 32'b11111111111111111100010101111001;
assign LUT_1[59076] = 32'b00000000000000001111001111000011;
assign LUT_1[59077] = 32'b00000000000000001000100000111111;
assign LUT_1[59078] = 32'b00000000000000001010111101010100;
assign LUT_1[59079] = 32'b00000000000000000100001111010000;
assign LUT_1[59080] = 32'b00000000000000000110100011100001;
assign LUT_1[59081] = 32'b11111111111111111111110101011101;
assign LUT_1[59082] = 32'b00000000000000000010010001110010;
assign LUT_1[59083] = 32'b11111111111111111011100011101110;
assign LUT_1[59084] = 32'b00000000000000001110011100111000;
assign LUT_1[59085] = 32'b00000000000000000111101110110100;
assign LUT_1[59086] = 32'b00000000000000001010001011001001;
assign LUT_1[59087] = 32'b00000000000000000011011101000101;
assign LUT_1[59088] = 32'b00000000000000001001010001001110;
assign LUT_1[59089] = 32'b00000000000000000010100011001010;
assign LUT_1[59090] = 32'b00000000000000000100111111011111;
assign LUT_1[59091] = 32'b11111111111111111110010001011011;
assign LUT_1[59092] = 32'b00000000000000010001001010100101;
assign LUT_1[59093] = 32'b00000000000000001010011100100001;
assign LUT_1[59094] = 32'b00000000000000001100111000110110;
assign LUT_1[59095] = 32'b00000000000000000110001010110010;
assign LUT_1[59096] = 32'b00000000000000001000011111000011;
assign LUT_1[59097] = 32'b00000000000000000001110000111111;
assign LUT_1[59098] = 32'b00000000000000000100001101010100;
assign LUT_1[59099] = 32'b11111111111111111101011111010000;
assign LUT_1[59100] = 32'b00000000000000010000011000011010;
assign LUT_1[59101] = 32'b00000000000000001001101010010110;
assign LUT_1[59102] = 32'b00000000000000001100000110101011;
assign LUT_1[59103] = 32'b00000000000000000101011000100111;
assign LUT_1[59104] = 32'b00000000000000001000010000101011;
assign LUT_1[59105] = 32'b00000000000000000001100010100111;
assign LUT_1[59106] = 32'b00000000000000000011111110111100;
assign LUT_1[59107] = 32'b11111111111111111101010000111000;
assign LUT_1[59108] = 32'b00000000000000010000001010000010;
assign LUT_1[59109] = 32'b00000000000000001001011011111110;
assign LUT_1[59110] = 32'b00000000000000001011111000010011;
assign LUT_1[59111] = 32'b00000000000000000101001010001111;
assign LUT_1[59112] = 32'b00000000000000000111011110100000;
assign LUT_1[59113] = 32'b00000000000000000000110000011100;
assign LUT_1[59114] = 32'b00000000000000000011001100110001;
assign LUT_1[59115] = 32'b11111111111111111100011110101101;
assign LUT_1[59116] = 32'b00000000000000001111010111110111;
assign LUT_1[59117] = 32'b00000000000000001000101001110011;
assign LUT_1[59118] = 32'b00000000000000001011000110001000;
assign LUT_1[59119] = 32'b00000000000000000100011000000100;
assign LUT_1[59120] = 32'b00000000000000001010001100001101;
assign LUT_1[59121] = 32'b00000000000000000011011110001001;
assign LUT_1[59122] = 32'b00000000000000000101111010011110;
assign LUT_1[59123] = 32'b11111111111111111111001100011010;
assign LUT_1[59124] = 32'b00000000000000010010000101100100;
assign LUT_1[59125] = 32'b00000000000000001011010111100000;
assign LUT_1[59126] = 32'b00000000000000001101110011110101;
assign LUT_1[59127] = 32'b00000000000000000111000101110001;
assign LUT_1[59128] = 32'b00000000000000001001011010000010;
assign LUT_1[59129] = 32'b00000000000000000010101011111110;
assign LUT_1[59130] = 32'b00000000000000000101001000010011;
assign LUT_1[59131] = 32'b11111111111111111110011010001111;
assign LUT_1[59132] = 32'b00000000000000010001010011011001;
assign LUT_1[59133] = 32'b00000000000000001010100101010101;
assign LUT_1[59134] = 32'b00000000000000001101000001101010;
assign LUT_1[59135] = 32'b00000000000000000110010011100110;
assign LUT_1[59136] = 32'b00000000000000000000001100001101;
assign LUT_1[59137] = 32'b11111111111111111001011110001001;
assign LUT_1[59138] = 32'b11111111111111111011111010011110;
assign LUT_1[59139] = 32'b11111111111111110101001100011010;
assign LUT_1[59140] = 32'b00000000000000001000000101100100;
assign LUT_1[59141] = 32'b00000000000000000001010111100000;
assign LUT_1[59142] = 32'b00000000000000000011110011110101;
assign LUT_1[59143] = 32'b11111111111111111101000101110001;
assign LUT_1[59144] = 32'b11111111111111111111011010000010;
assign LUT_1[59145] = 32'b11111111111111111000101011111110;
assign LUT_1[59146] = 32'b11111111111111111011001000010011;
assign LUT_1[59147] = 32'b11111111111111110100011010001111;
assign LUT_1[59148] = 32'b00000000000000000111010011011001;
assign LUT_1[59149] = 32'b00000000000000000000100101010101;
assign LUT_1[59150] = 32'b00000000000000000011000001101010;
assign LUT_1[59151] = 32'b11111111111111111100010011100110;
assign LUT_1[59152] = 32'b00000000000000000010000111101111;
assign LUT_1[59153] = 32'b11111111111111111011011001101011;
assign LUT_1[59154] = 32'b11111111111111111101110110000000;
assign LUT_1[59155] = 32'b11111111111111110111000111111100;
assign LUT_1[59156] = 32'b00000000000000001010000001000110;
assign LUT_1[59157] = 32'b00000000000000000011010011000010;
assign LUT_1[59158] = 32'b00000000000000000101101111010111;
assign LUT_1[59159] = 32'b11111111111111111111000001010011;
assign LUT_1[59160] = 32'b00000000000000000001010101100100;
assign LUT_1[59161] = 32'b11111111111111111010100111100000;
assign LUT_1[59162] = 32'b11111111111111111101000011110101;
assign LUT_1[59163] = 32'b11111111111111110110010101110001;
assign LUT_1[59164] = 32'b00000000000000001001001110111011;
assign LUT_1[59165] = 32'b00000000000000000010100000110111;
assign LUT_1[59166] = 32'b00000000000000000100111101001100;
assign LUT_1[59167] = 32'b11111111111111111110001111001000;
assign LUT_1[59168] = 32'b00000000000000000001000111001100;
assign LUT_1[59169] = 32'b11111111111111111010011001001000;
assign LUT_1[59170] = 32'b11111111111111111100110101011101;
assign LUT_1[59171] = 32'b11111111111111110110000111011001;
assign LUT_1[59172] = 32'b00000000000000001001000000100011;
assign LUT_1[59173] = 32'b00000000000000000010010010011111;
assign LUT_1[59174] = 32'b00000000000000000100101110110100;
assign LUT_1[59175] = 32'b11111111111111111110000000110000;
assign LUT_1[59176] = 32'b00000000000000000000010101000001;
assign LUT_1[59177] = 32'b11111111111111111001100110111101;
assign LUT_1[59178] = 32'b11111111111111111100000011010010;
assign LUT_1[59179] = 32'b11111111111111110101010101001110;
assign LUT_1[59180] = 32'b00000000000000001000001110011000;
assign LUT_1[59181] = 32'b00000000000000000001100000010100;
assign LUT_1[59182] = 32'b00000000000000000011111100101001;
assign LUT_1[59183] = 32'b11111111111111111101001110100101;
assign LUT_1[59184] = 32'b00000000000000000011000010101110;
assign LUT_1[59185] = 32'b11111111111111111100010100101010;
assign LUT_1[59186] = 32'b11111111111111111110110000111111;
assign LUT_1[59187] = 32'b11111111111111111000000010111011;
assign LUT_1[59188] = 32'b00000000000000001010111100000101;
assign LUT_1[59189] = 32'b00000000000000000100001110000001;
assign LUT_1[59190] = 32'b00000000000000000110101010010110;
assign LUT_1[59191] = 32'b11111111111111111111111100010010;
assign LUT_1[59192] = 32'b00000000000000000010010000100011;
assign LUT_1[59193] = 32'b11111111111111111011100010011111;
assign LUT_1[59194] = 32'b11111111111111111101111110110100;
assign LUT_1[59195] = 32'b11111111111111110111010000110000;
assign LUT_1[59196] = 32'b00000000000000001010001001111010;
assign LUT_1[59197] = 32'b00000000000000000011011011110110;
assign LUT_1[59198] = 32'b00000000000000000101111000001011;
assign LUT_1[59199] = 32'b11111111111111111111001010000111;
assign LUT_1[59200] = 32'b00000000000000000010001001110101;
assign LUT_1[59201] = 32'b11111111111111111011011011110001;
assign LUT_1[59202] = 32'b11111111111111111101111000000110;
assign LUT_1[59203] = 32'b11111111111111110111001010000010;
assign LUT_1[59204] = 32'b00000000000000001010000011001100;
assign LUT_1[59205] = 32'b00000000000000000011010101001000;
assign LUT_1[59206] = 32'b00000000000000000101110001011101;
assign LUT_1[59207] = 32'b11111111111111111111000011011001;
assign LUT_1[59208] = 32'b00000000000000000001010111101010;
assign LUT_1[59209] = 32'b11111111111111111010101001100110;
assign LUT_1[59210] = 32'b11111111111111111101000101111011;
assign LUT_1[59211] = 32'b11111111111111110110010111110111;
assign LUT_1[59212] = 32'b00000000000000001001010001000001;
assign LUT_1[59213] = 32'b00000000000000000010100010111101;
assign LUT_1[59214] = 32'b00000000000000000100111111010010;
assign LUT_1[59215] = 32'b11111111111111111110010001001110;
assign LUT_1[59216] = 32'b00000000000000000100000101010111;
assign LUT_1[59217] = 32'b11111111111111111101010111010011;
assign LUT_1[59218] = 32'b11111111111111111111110011101000;
assign LUT_1[59219] = 32'b11111111111111111001000101100100;
assign LUT_1[59220] = 32'b00000000000000001011111110101110;
assign LUT_1[59221] = 32'b00000000000000000101010000101010;
assign LUT_1[59222] = 32'b00000000000000000111101100111111;
assign LUT_1[59223] = 32'b00000000000000000000111110111011;
assign LUT_1[59224] = 32'b00000000000000000011010011001100;
assign LUT_1[59225] = 32'b11111111111111111100100101001000;
assign LUT_1[59226] = 32'b11111111111111111111000001011101;
assign LUT_1[59227] = 32'b11111111111111111000010011011001;
assign LUT_1[59228] = 32'b00000000000000001011001100100011;
assign LUT_1[59229] = 32'b00000000000000000100011110011111;
assign LUT_1[59230] = 32'b00000000000000000110111010110100;
assign LUT_1[59231] = 32'b00000000000000000000001100110000;
assign LUT_1[59232] = 32'b00000000000000000011000100110100;
assign LUT_1[59233] = 32'b11111111111111111100010110110000;
assign LUT_1[59234] = 32'b11111111111111111110110011000101;
assign LUT_1[59235] = 32'b11111111111111111000000101000001;
assign LUT_1[59236] = 32'b00000000000000001010111110001011;
assign LUT_1[59237] = 32'b00000000000000000100010000000111;
assign LUT_1[59238] = 32'b00000000000000000110101100011100;
assign LUT_1[59239] = 32'b11111111111111111111111110011000;
assign LUT_1[59240] = 32'b00000000000000000010010010101001;
assign LUT_1[59241] = 32'b11111111111111111011100100100101;
assign LUT_1[59242] = 32'b11111111111111111110000000111010;
assign LUT_1[59243] = 32'b11111111111111110111010010110110;
assign LUT_1[59244] = 32'b00000000000000001010001100000000;
assign LUT_1[59245] = 32'b00000000000000000011011101111100;
assign LUT_1[59246] = 32'b00000000000000000101111010010001;
assign LUT_1[59247] = 32'b11111111111111111111001100001101;
assign LUT_1[59248] = 32'b00000000000000000101000000010110;
assign LUT_1[59249] = 32'b11111111111111111110010010010010;
assign LUT_1[59250] = 32'b00000000000000000000101110100111;
assign LUT_1[59251] = 32'b11111111111111111010000000100011;
assign LUT_1[59252] = 32'b00000000000000001100111001101101;
assign LUT_1[59253] = 32'b00000000000000000110001011101001;
assign LUT_1[59254] = 32'b00000000000000001000100111111110;
assign LUT_1[59255] = 32'b00000000000000000001111001111010;
assign LUT_1[59256] = 32'b00000000000000000100001110001011;
assign LUT_1[59257] = 32'b11111111111111111101100000000111;
assign LUT_1[59258] = 32'b11111111111111111111111100011100;
assign LUT_1[59259] = 32'b11111111111111111001001110011000;
assign LUT_1[59260] = 32'b00000000000000001100000111100010;
assign LUT_1[59261] = 32'b00000000000000000101011001011110;
assign LUT_1[59262] = 32'b00000000000000000111110101110011;
assign LUT_1[59263] = 32'b00000000000000000001000111101111;
assign LUT_1[59264] = 32'b00000000000000000011001100010000;
assign LUT_1[59265] = 32'b11111111111111111100011110001100;
assign LUT_1[59266] = 32'b11111111111111111110111010100001;
assign LUT_1[59267] = 32'b11111111111111111000001100011101;
assign LUT_1[59268] = 32'b00000000000000001011000101100111;
assign LUT_1[59269] = 32'b00000000000000000100010111100011;
assign LUT_1[59270] = 32'b00000000000000000110110011111000;
assign LUT_1[59271] = 32'b00000000000000000000000101110100;
assign LUT_1[59272] = 32'b00000000000000000010011010000101;
assign LUT_1[59273] = 32'b11111111111111111011101100000001;
assign LUT_1[59274] = 32'b11111111111111111110001000010110;
assign LUT_1[59275] = 32'b11111111111111110111011010010010;
assign LUT_1[59276] = 32'b00000000000000001010010011011100;
assign LUT_1[59277] = 32'b00000000000000000011100101011000;
assign LUT_1[59278] = 32'b00000000000000000110000001101101;
assign LUT_1[59279] = 32'b11111111111111111111010011101001;
assign LUT_1[59280] = 32'b00000000000000000101000111110010;
assign LUT_1[59281] = 32'b11111111111111111110011001101110;
assign LUT_1[59282] = 32'b00000000000000000000110110000011;
assign LUT_1[59283] = 32'b11111111111111111010000111111111;
assign LUT_1[59284] = 32'b00000000000000001101000001001001;
assign LUT_1[59285] = 32'b00000000000000000110010011000101;
assign LUT_1[59286] = 32'b00000000000000001000101111011010;
assign LUT_1[59287] = 32'b00000000000000000010000001010110;
assign LUT_1[59288] = 32'b00000000000000000100010101100111;
assign LUT_1[59289] = 32'b11111111111111111101100111100011;
assign LUT_1[59290] = 32'b00000000000000000000000011111000;
assign LUT_1[59291] = 32'b11111111111111111001010101110100;
assign LUT_1[59292] = 32'b00000000000000001100001110111110;
assign LUT_1[59293] = 32'b00000000000000000101100000111010;
assign LUT_1[59294] = 32'b00000000000000000111111101001111;
assign LUT_1[59295] = 32'b00000000000000000001001111001011;
assign LUT_1[59296] = 32'b00000000000000000100000111001111;
assign LUT_1[59297] = 32'b11111111111111111101011001001011;
assign LUT_1[59298] = 32'b11111111111111111111110101100000;
assign LUT_1[59299] = 32'b11111111111111111001000111011100;
assign LUT_1[59300] = 32'b00000000000000001100000000100110;
assign LUT_1[59301] = 32'b00000000000000000101010010100010;
assign LUT_1[59302] = 32'b00000000000000000111101110110111;
assign LUT_1[59303] = 32'b00000000000000000001000000110011;
assign LUT_1[59304] = 32'b00000000000000000011010101000100;
assign LUT_1[59305] = 32'b11111111111111111100100111000000;
assign LUT_1[59306] = 32'b11111111111111111111000011010101;
assign LUT_1[59307] = 32'b11111111111111111000010101010001;
assign LUT_1[59308] = 32'b00000000000000001011001110011011;
assign LUT_1[59309] = 32'b00000000000000000100100000010111;
assign LUT_1[59310] = 32'b00000000000000000110111100101100;
assign LUT_1[59311] = 32'b00000000000000000000001110101000;
assign LUT_1[59312] = 32'b00000000000000000110000010110001;
assign LUT_1[59313] = 32'b11111111111111111111010100101101;
assign LUT_1[59314] = 32'b00000000000000000001110001000010;
assign LUT_1[59315] = 32'b11111111111111111011000010111110;
assign LUT_1[59316] = 32'b00000000000000001101111100001000;
assign LUT_1[59317] = 32'b00000000000000000111001110000100;
assign LUT_1[59318] = 32'b00000000000000001001101010011001;
assign LUT_1[59319] = 32'b00000000000000000010111100010101;
assign LUT_1[59320] = 32'b00000000000000000101010000100110;
assign LUT_1[59321] = 32'b11111111111111111110100010100010;
assign LUT_1[59322] = 32'b00000000000000000000111110110111;
assign LUT_1[59323] = 32'b11111111111111111010010000110011;
assign LUT_1[59324] = 32'b00000000000000001101001001111101;
assign LUT_1[59325] = 32'b00000000000000000110011011111001;
assign LUT_1[59326] = 32'b00000000000000001000111000001110;
assign LUT_1[59327] = 32'b00000000000000000010001010001010;
assign LUT_1[59328] = 32'b00000000000000000101001001111000;
assign LUT_1[59329] = 32'b11111111111111111110011011110100;
assign LUT_1[59330] = 32'b00000000000000000000111000001001;
assign LUT_1[59331] = 32'b11111111111111111010001010000101;
assign LUT_1[59332] = 32'b00000000000000001101000011001111;
assign LUT_1[59333] = 32'b00000000000000000110010101001011;
assign LUT_1[59334] = 32'b00000000000000001000110001100000;
assign LUT_1[59335] = 32'b00000000000000000010000011011100;
assign LUT_1[59336] = 32'b00000000000000000100010111101101;
assign LUT_1[59337] = 32'b11111111111111111101101001101001;
assign LUT_1[59338] = 32'b00000000000000000000000101111110;
assign LUT_1[59339] = 32'b11111111111111111001010111111010;
assign LUT_1[59340] = 32'b00000000000000001100010001000100;
assign LUT_1[59341] = 32'b00000000000000000101100011000000;
assign LUT_1[59342] = 32'b00000000000000000111111111010101;
assign LUT_1[59343] = 32'b00000000000000000001010001010001;
assign LUT_1[59344] = 32'b00000000000000000111000101011010;
assign LUT_1[59345] = 32'b00000000000000000000010111010110;
assign LUT_1[59346] = 32'b00000000000000000010110011101011;
assign LUT_1[59347] = 32'b11111111111111111100000101100111;
assign LUT_1[59348] = 32'b00000000000000001110111110110001;
assign LUT_1[59349] = 32'b00000000000000001000010000101101;
assign LUT_1[59350] = 32'b00000000000000001010101101000010;
assign LUT_1[59351] = 32'b00000000000000000011111110111110;
assign LUT_1[59352] = 32'b00000000000000000110010011001111;
assign LUT_1[59353] = 32'b11111111111111111111100101001011;
assign LUT_1[59354] = 32'b00000000000000000010000001100000;
assign LUT_1[59355] = 32'b11111111111111111011010011011100;
assign LUT_1[59356] = 32'b00000000000000001110001100100110;
assign LUT_1[59357] = 32'b00000000000000000111011110100010;
assign LUT_1[59358] = 32'b00000000000000001001111010110111;
assign LUT_1[59359] = 32'b00000000000000000011001100110011;
assign LUT_1[59360] = 32'b00000000000000000110000100110111;
assign LUT_1[59361] = 32'b11111111111111111111010110110011;
assign LUT_1[59362] = 32'b00000000000000000001110011001000;
assign LUT_1[59363] = 32'b11111111111111111011000101000100;
assign LUT_1[59364] = 32'b00000000000000001101111110001110;
assign LUT_1[59365] = 32'b00000000000000000111010000001010;
assign LUT_1[59366] = 32'b00000000000000001001101100011111;
assign LUT_1[59367] = 32'b00000000000000000010111110011011;
assign LUT_1[59368] = 32'b00000000000000000101010010101100;
assign LUT_1[59369] = 32'b11111111111111111110100100101000;
assign LUT_1[59370] = 32'b00000000000000000001000000111101;
assign LUT_1[59371] = 32'b11111111111111111010010010111001;
assign LUT_1[59372] = 32'b00000000000000001101001100000011;
assign LUT_1[59373] = 32'b00000000000000000110011101111111;
assign LUT_1[59374] = 32'b00000000000000001000111010010100;
assign LUT_1[59375] = 32'b00000000000000000010001100010000;
assign LUT_1[59376] = 32'b00000000000000001000000000011001;
assign LUT_1[59377] = 32'b00000000000000000001010010010101;
assign LUT_1[59378] = 32'b00000000000000000011101110101010;
assign LUT_1[59379] = 32'b11111111111111111101000000100110;
assign LUT_1[59380] = 32'b00000000000000001111111001110000;
assign LUT_1[59381] = 32'b00000000000000001001001011101100;
assign LUT_1[59382] = 32'b00000000000000001011101000000001;
assign LUT_1[59383] = 32'b00000000000000000100111001111101;
assign LUT_1[59384] = 32'b00000000000000000111001110001110;
assign LUT_1[59385] = 32'b00000000000000000000100000001010;
assign LUT_1[59386] = 32'b00000000000000000010111100011111;
assign LUT_1[59387] = 32'b11111111111111111100001110011011;
assign LUT_1[59388] = 32'b00000000000000001111000111100101;
assign LUT_1[59389] = 32'b00000000000000001000011001100001;
assign LUT_1[59390] = 32'b00000000000000001010110101110110;
assign LUT_1[59391] = 32'b00000000000000000100000111110010;
assign LUT_1[59392] = 32'b00000000000000000011010100101111;
assign LUT_1[59393] = 32'b11111111111111111100100110101011;
assign LUT_1[59394] = 32'b11111111111111111111000011000000;
assign LUT_1[59395] = 32'b11111111111111111000010100111100;
assign LUT_1[59396] = 32'b00000000000000001011001110000110;
assign LUT_1[59397] = 32'b00000000000000000100100000000010;
assign LUT_1[59398] = 32'b00000000000000000110111100010111;
assign LUT_1[59399] = 32'b00000000000000000000001110010011;
assign LUT_1[59400] = 32'b00000000000000000010100010100100;
assign LUT_1[59401] = 32'b11111111111111111011110100100000;
assign LUT_1[59402] = 32'b11111111111111111110010000110101;
assign LUT_1[59403] = 32'b11111111111111110111100010110001;
assign LUT_1[59404] = 32'b00000000000000001010011011111011;
assign LUT_1[59405] = 32'b00000000000000000011101101110111;
assign LUT_1[59406] = 32'b00000000000000000110001010001100;
assign LUT_1[59407] = 32'b11111111111111111111011100001000;
assign LUT_1[59408] = 32'b00000000000000000101010000010001;
assign LUT_1[59409] = 32'b11111111111111111110100010001101;
assign LUT_1[59410] = 32'b00000000000000000000111110100010;
assign LUT_1[59411] = 32'b11111111111111111010010000011110;
assign LUT_1[59412] = 32'b00000000000000001101001001101000;
assign LUT_1[59413] = 32'b00000000000000000110011011100100;
assign LUT_1[59414] = 32'b00000000000000001000110111111001;
assign LUT_1[59415] = 32'b00000000000000000010001001110101;
assign LUT_1[59416] = 32'b00000000000000000100011110000110;
assign LUT_1[59417] = 32'b11111111111111111101110000000010;
assign LUT_1[59418] = 32'b00000000000000000000001100010111;
assign LUT_1[59419] = 32'b11111111111111111001011110010011;
assign LUT_1[59420] = 32'b00000000000000001100010111011101;
assign LUT_1[59421] = 32'b00000000000000000101101001011001;
assign LUT_1[59422] = 32'b00000000000000001000000101101110;
assign LUT_1[59423] = 32'b00000000000000000001010111101010;
assign LUT_1[59424] = 32'b00000000000000000100001111101110;
assign LUT_1[59425] = 32'b11111111111111111101100001101010;
assign LUT_1[59426] = 32'b11111111111111111111111101111111;
assign LUT_1[59427] = 32'b11111111111111111001001111111011;
assign LUT_1[59428] = 32'b00000000000000001100001001000101;
assign LUT_1[59429] = 32'b00000000000000000101011011000001;
assign LUT_1[59430] = 32'b00000000000000000111110111010110;
assign LUT_1[59431] = 32'b00000000000000000001001001010010;
assign LUT_1[59432] = 32'b00000000000000000011011101100011;
assign LUT_1[59433] = 32'b11111111111111111100101111011111;
assign LUT_1[59434] = 32'b11111111111111111111001011110100;
assign LUT_1[59435] = 32'b11111111111111111000011101110000;
assign LUT_1[59436] = 32'b00000000000000001011010110111010;
assign LUT_1[59437] = 32'b00000000000000000100101000110110;
assign LUT_1[59438] = 32'b00000000000000000111000101001011;
assign LUT_1[59439] = 32'b00000000000000000000010111000111;
assign LUT_1[59440] = 32'b00000000000000000110001011010000;
assign LUT_1[59441] = 32'b11111111111111111111011101001100;
assign LUT_1[59442] = 32'b00000000000000000001111001100001;
assign LUT_1[59443] = 32'b11111111111111111011001011011101;
assign LUT_1[59444] = 32'b00000000000000001110000100100111;
assign LUT_1[59445] = 32'b00000000000000000111010110100011;
assign LUT_1[59446] = 32'b00000000000000001001110010111000;
assign LUT_1[59447] = 32'b00000000000000000011000100110100;
assign LUT_1[59448] = 32'b00000000000000000101011001000101;
assign LUT_1[59449] = 32'b11111111111111111110101011000001;
assign LUT_1[59450] = 32'b00000000000000000001000111010110;
assign LUT_1[59451] = 32'b11111111111111111010011001010010;
assign LUT_1[59452] = 32'b00000000000000001101010010011100;
assign LUT_1[59453] = 32'b00000000000000000110100100011000;
assign LUT_1[59454] = 32'b00000000000000001001000000101101;
assign LUT_1[59455] = 32'b00000000000000000010010010101001;
assign LUT_1[59456] = 32'b00000000000000000101010010010111;
assign LUT_1[59457] = 32'b11111111111111111110100100010011;
assign LUT_1[59458] = 32'b00000000000000000001000000101000;
assign LUT_1[59459] = 32'b11111111111111111010010010100100;
assign LUT_1[59460] = 32'b00000000000000001101001011101110;
assign LUT_1[59461] = 32'b00000000000000000110011101101010;
assign LUT_1[59462] = 32'b00000000000000001000111001111111;
assign LUT_1[59463] = 32'b00000000000000000010001011111011;
assign LUT_1[59464] = 32'b00000000000000000100100000001100;
assign LUT_1[59465] = 32'b11111111111111111101110010001000;
assign LUT_1[59466] = 32'b00000000000000000000001110011101;
assign LUT_1[59467] = 32'b11111111111111111001100000011001;
assign LUT_1[59468] = 32'b00000000000000001100011001100011;
assign LUT_1[59469] = 32'b00000000000000000101101011011111;
assign LUT_1[59470] = 32'b00000000000000001000000111110100;
assign LUT_1[59471] = 32'b00000000000000000001011001110000;
assign LUT_1[59472] = 32'b00000000000000000111001101111001;
assign LUT_1[59473] = 32'b00000000000000000000011111110101;
assign LUT_1[59474] = 32'b00000000000000000010111100001010;
assign LUT_1[59475] = 32'b11111111111111111100001110000110;
assign LUT_1[59476] = 32'b00000000000000001111000111010000;
assign LUT_1[59477] = 32'b00000000000000001000011001001100;
assign LUT_1[59478] = 32'b00000000000000001010110101100001;
assign LUT_1[59479] = 32'b00000000000000000100000111011101;
assign LUT_1[59480] = 32'b00000000000000000110011011101110;
assign LUT_1[59481] = 32'b11111111111111111111101101101010;
assign LUT_1[59482] = 32'b00000000000000000010001001111111;
assign LUT_1[59483] = 32'b11111111111111111011011011111011;
assign LUT_1[59484] = 32'b00000000000000001110010101000101;
assign LUT_1[59485] = 32'b00000000000000000111100111000001;
assign LUT_1[59486] = 32'b00000000000000001010000011010110;
assign LUT_1[59487] = 32'b00000000000000000011010101010010;
assign LUT_1[59488] = 32'b00000000000000000110001101010110;
assign LUT_1[59489] = 32'b11111111111111111111011111010010;
assign LUT_1[59490] = 32'b00000000000000000001111011100111;
assign LUT_1[59491] = 32'b11111111111111111011001101100011;
assign LUT_1[59492] = 32'b00000000000000001110000110101101;
assign LUT_1[59493] = 32'b00000000000000000111011000101001;
assign LUT_1[59494] = 32'b00000000000000001001110100111110;
assign LUT_1[59495] = 32'b00000000000000000011000110111010;
assign LUT_1[59496] = 32'b00000000000000000101011011001011;
assign LUT_1[59497] = 32'b11111111111111111110101101000111;
assign LUT_1[59498] = 32'b00000000000000000001001001011100;
assign LUT_1[59499] = 32'b11111111111111111010011011011000;
assign LUT_1[59500] = 32'b00000000000000001101010100100010;
assign LUT_1[59501] = 32'b00000000000000000110100110011110;
assign LUT_1[59502] = 32'b00000000000000001001000010110011;
assign LUT_1[59503] = 32'b00000000000000000010010100101111;
assign LUT_1[59504] = 32'b00000000000000001000001000111000;
assign LUT_1[59505] = 32'b00000000000000000001011010110100;
assign LUT_1[59506] = 32'b00000000000000000011110111001001;
assign LUT_1[59507] = 32'b11111111111111111101001001000101;
assign LUT_1[59508] = 32'b00000000000000010000000010001111;
assign LUT_1[59509] = 32'b00000000000000001001010100001011;
assign LUT_1[59510] = 32'b00000000000000001011110000100000;
assign LUT_1[59511] = 32'b00000000000000000101000010011100;
assign LUT_1[59512] = 32'b00000000000000000111010110101101;
assign LUT_1[59513] = 32'b00000000000000000000101000101001;
assign LUT_1[59514] = 32'b00000000000000000011000100111110;
assign LUT_1[59515] = 32'b11111111111111111100010110111010;
assign LUT_1[59516] = 32'b00000000000000001111010000000100;
assign LUT_1[59517] = 32'b00000000000000001000100010000000;
assign LUT_1[59518] = 32'b00000000000000001010111110010101;
assign LUT_1[59519] = 32'b00000000000000000100010000010001;
assign LUT_1[59520] = 32'b00000000000000000110010100110010;
assign LUT_1[59521] = 32'b11111111111111111111100110101110;
assign LUT_1[59522] = 32'b00000000000000000010000011000011;
assign LUT_1[59523] = 32'b11111111111111111011010100111111;
assign LUT_1[59524] = 32'b00000000000000001110001110001001;
assign LUT_1[59525] = 32'b00000000000000000111100000000101;
assign LUT_1[59526] = 32'b00000000000000001001111100011010;
assign LUT_1[59527] = 32'b00000000000000000011001110010110;
assign LUT_1[59528] = 32'b00000000000000000101100010100111;
assign LUT_1[59529] = 32'b11111111111111111110110100100011;
assign LUT_1[59530] = 32'b00000000000000000001010000111000;
assign LUT_1[59531] = 32'b11111111111111111010100010110100;
assign LUT_1[59532] = 32'b00000000000000001101011011111110;
assign LUT_1[59533] = 32'b00000000000000000110101101111010;
assign LUT_1[59534] = 32'b00000000000000001001001010001111;
assign LUT_1[59535] = 32'b00000000000000000010011100001011;
assign LUT_1[59536] = 32'b00000000000000001000010000010100;
assign LUT_1[59537] = 32'b00000000000000000001100010010000;
assign LUT_1[59538] = 32'b00000000000000000011111110100101;
assign LUT_1[59539] = 32'b11111111111111111101010000100001;
assign LUT_1[59540] = 32'b00000000000000010000001001101011;
assign LUT_1[59541] = 32'b00000000000000001001011011100111;
assign LUT_1[59542] = 32'b00000000000000001011110111111100;
assign LUT_1[59543] = 32'b00000000000000000101001001111000;
assign LUT_1[59544] = 32'b00000000000000000111011110001001;
assign LUT_1[59545] = 32'b00000000000000000000110000000101;
assign LUT_1[59546] = 32'b00000000000000000011001100011010;
assign LUT_1[59547] = 32'b11111111111111111100011110010110;
assign LUT_1[59548] = 32'b00000000000000001111010111100000;
assign LUT_1[59549] = 32'b00000000000000001000101001011100;
assign LUT_1[59550] = 32'b00000000000000001011000101110001;
assign LUT_1[59551] = 32'b00000000000000000100010111101101;
assign LUT_1[59552] = 32'b00000000000000000111001111110001;
assign LUT_1[59553] = 32'b00000000000000000000100001101101;
assign LUT_1[59554] = 32'b00000000000000000010111110000010;
assign LUT_1[59555] = 32'b11111111111111111100001111111110;
assign LUT_1[59556] = 32'b00000000000000001111001001001000;
assign LUT_1[59557] = 32'b00000000000000001000011011000100;
assign LUT_1[59558] = 32'b00000000000000001010110111011001;
assign LUT_1[59559] = 32'b00000000000000000100001001010101;
assign LUT_1[59560] = 32'b00000000000000000110011101100110;
assign LUT_1[59561] = 32'b11111111111111111111101111100010;
assign LUT_1[59562] = 32'b00000000000000000010001011110111;
assign LUT_1[59563] = 32'b11111111111111111011011101110011;
assign LUT_1[59564] = 32'b00000000000000001110010110111101;
assign LUT_1[59565] = 32'b00000000000000000111101000111001;
assign LUT_1[59566] = 32'b00000000000000001010000101001110;
assign LUT_1[59567] = 32'b00000000000000000011010111001010;
assign LUT_1[59568] = 32'b00000000000000001001001011010011;
assign LUT_1[59569] = 32'b00000000000000000010011101001111;
assign LUT_1[59570] = 32'b00000000000000000100111001100100;
assign LUT_1[59571] = 32'b11111111111111111110001011100000;
assign LUT_1[59572] = 32'b00000000000000010001000100101010;
assign LUT_1[59573] = 32'b00000000000000001010010110100110;
assign LUT_1[59574] = 32'b00000000000000001100110010111011;
assign LUT_1[59575] = 32'b00000000000000000110000100110111;
assign LUT_1[59576] = 32'b00000000000000001000011001001000;
assign LUT_1[59577] = 32'b00000000000000000001101011000100;
assign LUT_1[59578] = 32'b00000000000000000100000111011001;
assign LUT_1[59579] = 32'b11111111111111111101011001010101;
assign LUT_1[59580] = 32'b00000000000000010000010010011111;
assign LUT_1[59581] = 32'b00000000000000001001100100011011;
assign LUT_1[59582] = 32'b00000000000000001100000000110000;
assign LUT_1[59583] = 32'b00000000000000000101010010101100;
assign LUT_1[59584] = 32'b00000000000000001000010010011010;
assign LUT_1[59585] = 32'b00000000000000000001100100010110;
assign LUT_1[59586] = 32'b00000000000000000100000000101011;
assign LUT_1[59587] = 32'b11111111111111111101010010100111;
assign LUT_1[59588] = 32'b00000000000000010000001011110001;
assign LUT_1[59589] = 32'b00000000000000001001011101101101;
assign LUT_1[59590] = 32'b00000000000000001011111010000010;
assign LUT_1[59591] = 32'b00000000000000000101001011111110;
assign LUT_1[59592] = 32'b00000000000000000111100000001111;
assign LUT_1[59593] = 32'b00000000000000000000110010001011;
assign LUT_1[59594] = 32'b00000000000000000011001110100000;
assign LUT_1[59595] = 32'b11111111111111111100100000011100;
assign LUT_1[59596] = 32'b00000000000000001111011001100110;
assign LUT_1[59597] = 32'b00000000000000001000101011100010;
assign LUT_1[59598] = 32'b00000000000000001011000111110111;
assign LUT_1[59599] = 32'b00000000000000000100011001110011;
assign LUT_1[59600] = 32'b00000000000000001010001101111100;
assign LUT_1[59601] = 32'b00000000000000000011011111111000;
assign LUT_1[59602] = 32'b00000000000000000101111100001101;
assign LUT_1[59603] = 32'b11111111111111111111001110001001;
assign LUT_1[59604] = 32'b00000000000000010010000111010011;
assign LUT_1[59605] = 32'b00000000000000001011011001001111;
assign LUT_1[59606] = 32'b00000000000000001101110101100100;
assign LUT_1[59607] = 32'b00000000000000000111000111100000;
assign LUT_1[59608] = 32'b00000000000000001001011011110001;
assign LUT_1[59609] = 32'b00000000000000000010101101101101;
assign LUT_1[59610] = 32'b00000000000000000101001010000010;
assign LUT_1[59611] = 32'b11111111111111111110011011111110;
assign LUT_1[59612] = 32'b00000000000000010001010101001000;
assign LUT_1[59613] = 32'b00000000000000001010100111000100;
assign LUT_1[59614] = 32'b00000000000000001101000011011001;
assign LUT_1[59615] = 32'b00000000000000000110010101010101;
assign LUT_1[59616] = 32'b00000000000000001001001101011001;
assign LUT_1[59617] = 32'b00000000000000000010011111010101;
assign LUT_1[59618] = 32'b00000000000000000100111011101010;
assign LUT_1[59619] = 32'b11111111111111111110001101100110;
assign LUT_1[59620] = 32'b00000000000000010001000110110000;
assign LUT_1[59621] = 32'b00000000000000001010011000101100;
assign LUT_1[59622] = 32'b00000000000000001100110101000001;
assign LUT_1[59623] = 32'b00000000000000000110000110111101;
assign LUT_1[59624] = 32'b00000000000000001000011011001110;
assign LUT_1[59625] = 32'b00000000000000000001101101001010;
assign LUT_1[59626] = 32'b00000000000000000100001001011111;
assign LUT_1[59627] = 32'b11111111111111111101011011011011;
assign LUT_1[59628] = 32'b00000000000000010000010100100101;
assign LUT_1[59629] = 32'b00000000000000001001100110100001;
assign LUT_1[59630] = 32'b00000000000000001100000010110110;
assign LUT_1[59631] = 32'b00000000000000000101010100110010;
assign LUT_1[59632] = 32'b00000000000000001011001000111011;
assign LUT_1[59633] = 32'b00000000000000000100011010110111;
assign LUT_1[59634] = 32'b00000000000000000110110111001100;
assign LUT_1[59635] = 32'b00000000000000000000001001001000;
assign LUT_1[59636] = 32'b00000000000000010011000010010010;
assign LUT_1[59637] = 32'b00000000000000001100010100001110;
assign LUT_1[59638] = 32'b00000000000000001110110000100011;
assign LUT_1[59639] = 32'b00000000000000001000000010011111;
assign LUT_1[59640] = 32'b00000000000000001010010110110000;
assign LUT_1[59641] = 32'b00000000000000000011101000101100;
assign LUT_1[59642] = 32'b00000000000000000110000101000001;
assign LUT_1[59643] = 32'b11111111111111111111010110111101;
assign LUT_1[59644] = 32'b00000000000000010010010000000111;
assign LUT_1[59645] = 32'b00000000000000001011100010000011;
assign LUT_1[59646] = 32'b00000000000000001101111110011000;
assign LUT_1[59647] = 32'b00000000000000000111010000010100;
assign LUT_1[59648] = 32'b00000000000000000001001000111011;
assign LUT_1[59649] = 32'b11111111111111111010011010110111;
assign LUT_1[59650] = 32'b11111111111111111100110111001100;
assign LUT_1[59651] = 32'b11111111111111110110001001001000;
assign LUT_1[59652] = 32'b00000000000000001001000010010010;
assign LUT_1[59653] = 32'b00000000000000000010010100001110;
assign LUT_1[59654] = 32'b00000000000000000100110000100011;
assign LUT_1[59655] = 32'b11111111111111111110000010011111;
assign LUT_1[59656] = 32'b00000000000000000000010110110000;
assign LUT_1[59657] = 32'b11111111111111111001101000101100;
assign LUT_1[59658] = 32'b11111111111111111100000101000001;
assign LUT_1[59659] = 32'b11111111111111110101010110111101;
assign LUT_1[59660] = 32'b00000000000000001000010000000111;
assign LUT_1[59661] = 32'b00000000000000000001100010000011;
assign LUT_1[59662] = 32'b00000000000000000011111110011000;
assign LUT_1[59663] = 32'b11111111111111111101010000010100;
assign LUT_1[59664] = 32'b00000000000000000011000100011101;
assign LUT_1[59665] = 32'b11111111111111111100010110011001;
assign LUT_1[59666] = 32'b11111111111111111110110010101110;
assign LUT_1[59667] = 32'b11111111111111111000000100101010;
assign LUT_1[59668] = 32'b00000000000000001010111101110100;
assign LUT_1[59669] = 32'b00000000000000000100001111110000;
assign LUT_1[59670] = 32'b00000000000000000110101100000101;
assign LUT_1[59671] = 32'b11111111111111111111111110000001;
assign LUT_1[59672] = 32'b00000000000000000010010010010010;
assign LUT_1[59673] = 32'b11111111111111111011100100001110;
assign LUT_1[59674] = 32'b11111111111111111110000000100011;
assign LUT_1[59675] = 32'b11111111111111110111010010011111;
assign LUT_1[59676] = 32'b00000000000000001010001011101001;
assign LUT_1[59677] = 32'b00000000000000000011011101100101;
assign LUT_1[59678] = 32'b00000000000000000101111001111010;
assign LUT_1[59679] = 32'b11111111111111111111001011110110;
assign LUT_1[59680] = 32'b00000000000000000010000011111010;
assign LUT_1[59681] = 32'b11111111111111111011010101110110;
assign LUT_1[59682] = 32'b11111111111111111101110010001011;
assign LUT_1[59683] = 32'b11111111111111110111000100000111;
assign LUT_1[59684] = 32'b00000000000000001001111101010001;
assign LUT_1[59685] = 32'b00000000000000000011001111001101;
assign LUT_1[59686] = 32'b00000000000000000101101011100010;
assign LUT_1[59687] = 32'b11111111111111111110111101011110;
assign LUT_1[59688] = 32'b00000000000000000001010001101111;
assign LUT_1[59689] = 32'b11111111111111111010100011101011;
assign LUT_1[59690] = 32'b11111111111111111101000000000000;
assign LUT_1[59691] = 32'b11111111111111110110010001111100;
assign LUT_1[59692] = 32'b00000000000000001001001011000110;
assign LUT_1[59693] = 32'b00000000000000000010011101000010;
assign LUT_1[59694] = 32'b00000000000000000100111001010111;
assign LUT_1[59695] = 32'b11111111111111111110001011010011;
assign LUT_1[59696] = 32'b00000000000000000011111111011100;
assign LUT_1[59697] = 32'b11111111111111111101010001011000;
assign LUT_1[59698] = 32'b11111111111111111111101101101101;
assign LUT_1[59699] = 32'b11111111111111111000111111101001;
assign LUT_1[59700] = 32'b00000000000000001011111000110011;
assign LUT_1[59701] = 32'b00000000000000000101001010101111;
assign LUT_1[59702] = 32'b00000000000000000111100111000100;
assign LUT_1[59703] = 32'b00000000000000000000111001000000;
assign LUT_1[59704] = 32'b00000000000000000011001101010001;
assign LUT_1[59705] = 32'b11111111111111111100011111001101;
assign LUT_1[59706] = 32'b11111111111111111110111011100010;
assign LUT_1[59707] = 32'b11111111111111111000001101011110;
assign LUT_1[59708] = 32'b00000000000000001011000110101000;
assign LUT_1[59709] = 32'b00000000000000000100011000100100;
assign LUT_1[59710] = 32'b00000000000000000110110100111001;
assign LUT_1[59711] = 32'b00000000000000000000000110110101;
assign LUT_1[59712] = 32'b00000000000000000011000110100011;
assign LUT_1[59713] = 32'b11111111111111111100011000011111;
assign LUT_1[59714] = 32'b11111111111111111110110100110100;
assign LUT_1[59715] = 32'b11111111111111111000000110110000;
assign LUT_1[59716] = 32'b00000000000000001010111111111010;
assign LUT_1[59717] = 32'b00000000000000000100010001110110;
assign LUT_1[59718] = 32'b00000000000000000110101110001011;
assign LUT_1[59719] = 32'b00000000000000000000000000000111;
assign LUT_1[59720] = 32'b00000000000000000010010100011000;
assign LUT_1[59721] = 32'b11111111111111111011100110010100;
assign LUT_1[59722] = 32'b11111111111111111110000010101001;
assign LUT_1[59723] = 32'b11111111111111110111010100100101;
assign LUT_1[59724] = 32'b00000000000000001010001101101111;
assign LUT_1[59725] = 32'b00000000000000000011011111101011;
assign LUT_1[59726] = 32'b00000000000000000101111100000000;
assign LUT_1[59727] = 32'b11111111111111111111001101111100;
assign LUT_1[59728] = 32'b00000000000000000101000010000101;
assign LUT_1[59729] = 32'b11111111111111111110010100000001;
assign LUT_1[59730] = 32'b00000000000000000000110000010110;
assign LUT_1[59731] = 32'b11111111111111111010000010010010;
assign LUT_1[59732] = 32'b00000000000000001100111011011100;
assign LUT_1[59733] = 32'b00000000000000000110001101011000;
assign LUT_1[59734] = 32'b00000000000000001000101001101101;
assign LUT_1[59735] = 32'b00000000000000000001111011101001;
assign LUT_1[59736] = 32'b00000000000000000100001111111010;
assign LUT_1[59737] = 32'b11111111111111111101100001110110;
assign LUT_1[59738] = 32'b11111111111111111111111110001011;
assign LUT_1[59739] = 32'b11111111111111111001010000000111;
assign LUT_1[59740] = 32'b00000000000000001100001001010001;
assign LUT_1[59741] = 32'b00000000000000000101011011001101;
assign LUT_1[59742] = 32'b00000000000000000111110111100010;
assign LUT_1[59743] = 32'b00000000000000000001001001011110;
assign LUT_1[59744] = 32'b00000000000000000100000001100010;
assign LUT_1[59745] = 32'b11111111111111111101010011011110;
assign LUT_1[59746] = 32'b11111111111111111111101111110011;
assign LUT_1[59747] = 32'b11111111111111111001000001101111;
assign LUT_1[59748] = 32'b00000000000000001011111010111001;
assign LUT_1[59749] = 32'b00000000000000000101001100110101;
assign LUT_1[59750] = 32'b00000000000000000111101001001010;
assign LUT_1[59751] = 32'b00000000000000000000111011000110;
assign LUT_1[59752] = 32'b00000000000000000011001111010111;
assign LUT_1[59753] = 32'b11111111111111111100100001010011;
assign LUT_1[59754] = 32'b11111111111111111110111101101000;
assign LUT_1[59755] = 32'b11111111111111111000001111100100;
assign LUT_1[59756] = 32'b00000000000000001011001000101110;
assign LUT_1[59757] = 32'b00000000000000000100011010101010;
assign LUT_1[59758] = 32'b00000000000000000110110110111111;
assign LUT_1[59759] = 32'b00000000000000000000001000111011;
assign LUT_1[59760] = 32'b00000000000000000101111101000100;
assign LUT_1[59761] = 32'b11111111111111111111001111000000;
assign LUT_1[59762] = 32'b00000000000000000001101011010101;
assign LUT_1[59763] = 32'b11111111111111111010111101010001;
assign LUT_1[59764] = 32'b00000000000000001101110110011011;
assign LUT_1[59765] = 32'b00000000000000000111001000010111;
assign LUT_1[59766] = 32'b00000000000000001001100100101100;
assign LUT_1[59767] = 32'b00000000000000000010110110101000;
assign LUT_1[59768] = 32'b00000000000000000101001010111001;
assign LUT_1[59769] = 32'b11111111111111111110011100110101;
assign LUT_1[59770] = 32'b00000000000000000000111001001010;
assign LUT_1[59771] = 32'b11111111111111111010001011000110;
assign LUT_1[59772] = 32'b00000000000000001101000100010000;
assign LUT_1[59773] = 32'b00000000000000000110010110001100;
assign LUT_1[59774] = 32'b00000000000000001000110010100001;
assign LUT_1[59775] = 32'b00000000000000000010000100011101;
assign LUT_1[59776] = 32'b00000000000000000100001000111110;
assign LUT_1[59777] = 32'b11111111111111111101011010111010;
assign LUT_1[59778] = 32'b11111111111111111111110111001111;
assign LUT_1[59779] = 32'b11111111111111111001001001001011;
assign LUT_1[59780] = 32'b00000000000000001100000010010101;
assign LUT_1[59781] = 32'b00000000000000000101010100010001;
assign LUT_1[59782] = 32'b00000000000000000111110000100110;
assign LUT_1[59783] = 32'b00000000000000000001000010100010;
assign LUT_1[59784] = 32'b00000000000000000011010110110011;
assign LUT_1[59785] = 32'b11111111111111111100101000101111;
assign LUT_1[59786] = 32'b11111111111111111111000101000100;
assign LUT_1[59787] = 32'b11111111111111111000010111000000;
assign LUT_1[59788] = 32'b00000000000000001011010000001010;
assign LUT_1[59789] = 32'b00000000000000000100100010000110;
assign LUT_1[59790] = 32'b00000000000000000110111110011011;
assign LUT_1[59791] = 32'b00000000000000000000010000010111;
assign LUT_1[59792] = 32'b00000000000000000110000100100000;
assign LUT_1[59793] = 32'b11111111111111111111010110011100;
assign LUT_1[59794] = 32'b00000000000000000001110010110001;
assign LUT_1[59795] = 32'b11111111111111111011000100101101;
assign LUT_1[59796] = 32'b00000000000000001101111101110111;
assign LUT_1[59797] = 32'b00000000000000000111001111110011;
assign LUT_1[59798] = 32'b00000000000000001001101100001000;
assign LUT_1[59799] = 32'b00000000000000000010111110000100;
assign LUT_1[59800] = 32'b00000000000000000101010010010101;
assign LUT_1[59801] = 32'b11111111111111111110100100010001;
assign LUT_1[59802] = 32'b00000000000000000001000000100110;
assign LUT_1[59803] = 32'b11111111111111111010010010100010;
assign LUT_1[59804] = 32'b00000000000000001101001011101100;
assign LUT_1[59805] = 32'b00000000000000000110011101101000;
assign LUT_1[59806] = 32'b00000000000000001000111001111101;
assign LUT_1[59807] = 32'b00000000000000000010001011111001;
assign LUT_1[59808] = 32'b00000000000000000101000011111101;
assign LUT_1[59809] = 32'b11111111111111111110010101111001;
assign LUT_1[59810] = 32'b00000000000000000000110010001110;
assign LUT_1[59811] = 32'b11111111111111111010000100001010;
assign LUT_1[59812] = 32'b00000000000000001100111101010100;
assign LUT_1[59813] = 32'b00000000000000000110001111010000;
assign LUT_1[59814] = 32'b00000000000000001000101011100101;
assign LUT_1[59815] = 32'b00000000000000000001111101100001;
assign LUT_1[59816] = 32'b00000000000000000100010001110010;
assign LUT_1[59817] = 32'b11111111111111111101100011101110;
assign LUT_1[59818] = 32'b00000000000000000000000000000011;
assign LUT_1[59819] = 32'b11111111111111111001010001111111;
assign LUT_1[59820] = 32'b00000000000000001100001011001001;
assign LUT_1[59821] = 32'b00000000000000000101011101000101;
assign LUT_1[59822] = 32'b00000000000000000111111001011010;
assign LUT_1[59823] = 32'b00000000000000000001001011010110;
assign LUT_1[59824] = 32'b00000000000000000110111111011111;
assign LUT_1[59825] = 32'b00000000000000000000010001011011;
assign LUT_1[59826] = 32'b00000000000000000010101101110000;
assign LUT_1[59827] = 32'b11111111111111111011111111101100;
assign LUT_1[59828] = 32'b00000000000000001110111000110110;
assign LUT_1[59829] = 32'b00000000000000001000001010110010;
assign LUT_1[59830] = 32'b00000000000000001010100111000111;
assign LUT_1[59831] = 32'b00000000000000000011111001000011;
assign LUT_1[59832] = 32'b00000000000000000110001101010100;
assign LUT_1[59833] = 32'b11111111111111111111011111010000;
assign LUT_1[59834] = 32'b00000000000000000001111011100101;
assign LUT_1[59835] = 32'b11111111111111111011001101100001;
assign LUT_1[59836] = 32'b00000000000000001110000110101011;
assign LUT_1[59837] = 32'b00000000000000000111011000100111;
assign LUT_1[59838] = 32'b00000000000000001001110100111100;
assign LUT_1[59839] = 32'b00000000000000000011000110111000;
assign LUT_1[59840] = 32'b00000000000000000110000110100110;
assign LUT_1[59841] = 32'b11111111111111111111011000100010;
assign LUT_1[59842] = 32'b00000000000000000001110100110111;
assign LUT_1[59843] = 32'b11111111111111111011000110110011;
assign LUT_1[59844] = 32'b00000000000000001101111111111101;
assign LUT_1[59845] = 32'b00000000000000000111010001111001;
assign LUT_1[59846] = 32'b00000000000000001001101110001110;
assign LUT_1[59847] = 32'b00000000000000000011000000001010;
assign LUT_1[59848] = 32'b00000000000000000101010100011011;
assign LUT_1[59849] = 32'b11111111111111111110100110010111;
assign LUT_1[59850] = 32'b00000000000000000001000010101100;
assign LUT_1[59851] = 32'b11111111111111111010010100101000;
assign LUT_1[59852] = 32'b00000000000000001101001101110010;
assign LUT_1[59853] = 32'b00000000000000000110011111101110;
assign LUT_1[59854] = 32'b00000000000000001000111100000011;
assign LUT_1[59855] = 32'b00000000000000000010001101111111;
assign LUT_1[59856] = 32'b00000000000000001000000010001000;
assign LUT_1[59857] = 32'b00000000000000000001010100000100;
assign LUT_1[59858] = 32'b00000000000000000011110000011001;
assign LUT_1[59859] = 32'b11111111111111111101000010010101;
assign LUT_1[59860] = 32'b00000000000000001111111011011111;
assign LUT_1[59861] = 32'b00000000000000001001001101011011;
assign LUT_1[59862] = 32'b00000000000000001011101001110000;
assign LUT_1[59863] = 32'b00000000000000000100111011101100;
assign LUT_1[59864] = 32'b00000000000000000111001111111101;
assign LUT_1[59865] = 32'b00000000000000000000100001111001;
assign LUT_1[59866] = 32'b00000000000000000010111110001110;
assign LUT_1[59867] = 32'b11111111111111111100010000001010;
assign LUT_1[59868] = 32'b00000000000000001111001001010100;
assign LUT_1[59869] = 32'b00000000000000001000011011010000;
assign LUT_1[59870] = 32'b00000000000000001010110111100101;
assign LUT_1[59871] = 32'b00000000000000000100001001100001;
assign LUT_1[59872] = 32'b00000000000000000111000001100101;
assign LUT_1[59873] = 32'b00000000000000000000010011100001;
assign LUT_1[59874] = 32'b00000000000000000010101111110110;
assign LUT_1[59875] = 32'b11111111111111111100000001110010;
assign LUT_1[59876] = 32'b00000000000000001110111010111100;
assign LUT_1[59877] = 32'b00000000000000001000001100111000;
assign LUT_1[59878] = 32'b00000000000000001010101001001101;
assign LUT_1[59879] = 32'b00000000000000000011111011001001;
assign LUT_1[59880] = 32'b00000000000000000110001111011010;
assign LUT_1[59881] = 32'b11111111111111111111100001010110;
assign LUT_1[59882] = 32'b00000000000000000001111101101011;
assign LUT_1[59883] = 32'b11111111111111111011001111100111;
assign LUT_1[59884] = 32'b00000000000000001110001000110001;
assign LUT_1[59885] = 32'b00000000000000000111011010101101;
assign LUT_1[59886] = 32'b00000000000000001001110111000010;
assign LUT_1[59887] = 32'b00000000000000000011001000111110;
assign LUT_1[59888] = 32'b00000000000000001000111101000111;
assign LUT_1[59889] = 32'b00000000000000000010001111000011;
assign LUT_1[59890] = 32'b00000000000000000100101011011000;
assign LUT_1[59891] = 32'b11111111111111111101111101010100;
assign LUT_1[59892] = 32'b00000000000000010000110110011110;
assign LUT_1[59893] = 32'b00000000000000001010001000011010;
assign LUT_1[59894] = 32'b00000000000000001100100100101111;
assign LUT_1[59895] = 32'b00000000000000000101110110101011;
assign LUT_1[59896] = 32'b00000000000000001000001010111100;
assign LUT_1[59897] = 32'b00000000000000000001011100111000;
assign LUT_1[59898] = 32'b00000000000000000011111001001101;
assign LUT_1[59899] = 32'b11111111111111111101001011001001;
assign LUT_1[59900] = 32'b00000000000000010000000100010011;
assign LUT_1[59901] = 32'b00000000000000001001010110001111;
assign LUT_1[59902] = 32'b00000000000000001011110010100100;
assign LUT_1[59903] = 32'b00000000000000000101000100100000;
assign LUT_1[59904] = 32'b11111111111111111101000011001100;
assign LUT_1[59905] = 32'b11111111111111110110010101001000;
assign LUT_1[59906] = 32'b11111111111111111000110001011101;
assign LUT_1[59907] = 32'b11111111111111110010000011011001;
assign LUT_1[59908] = 32'b00000000000000000100111100100011;
assign LUT_1[59909] = 32'b11111111111111111110001110011111;
assign LUT_1[59910] = 32'b00000000000000000000101010110100;
assign LUT_1[59911] = 32'b11111111111111111001111100110000;
assign LUT_1[59912] = 32'b11111111111111111100010001000001;
assign LUT_1[59913] = 32'b11111111111111110101100010111101;
assign LUT_1[59914] = 32'b11111111111111110111111111010010;
assign LUT_1[59915] = 32'b11111111111111110001010001001110;
assign LUT_1[59916] = 32'b00000000000000000100001010011000;
assign LUT_1[59917] = 32'b11111111111111111101011100010100;
assign LUT_1[59918] = 32'b11111111111111111111111000101001;
assign LUT_1[59919] = 32'b11111111111111111001001010100101;
assign LUT_1[59920] = 32'b11111111111111111110111110101110;
assign LUT_1[59921] = 32'b11111111111111111000010000101010;
assign LUT_1[59922] = 32'b11111111111111111010101100111111;
assign LUT_1[59923] = 32'b11111111111111110011111110111011;
assign LUT_1[59924] = 32'b00000000000000000110111000000101;
assign LUT_1[59925] = 32'b00000000000000000000001010000001;
assign LUT_1[59926] = 32'b00000000000000000010100110010110;
assign LUT_1[59927] = 32'b11111111111111111011111000010010;
assign LUT_1[59928] = 32'b11111111111111111110001100100011;
assign LUT_1[59929] = 32'b11111111111111110111011110011111;
assign LUT_1[59930] = 32'b11111111111111111001111010110100;
assign LUT_1[59931] = 32'b11111111111111110011001100110000;
assign LUT_1[59932] = 32'b00000000000000000110000101111010;
assign LUT_1[59933] = 32'b11111111111111111111010111110110;
assign LUT_1[59934] = 32'b00000000000000000001110100001011;
assign LUT_1[59935] = 32'b11111111111111111011000110000111;
assign LUT_1[59936] = 32'b11111111111111111101111110001011;
assign LUT_1[59937] = 32'b11111111111111110111010000000111;
assign LUT_1[59938] = 32'b11111111111111111001101100011100;
assign LUT_1[59939] = 32'b11111111111111110010111110011000;
assign LUT_1[59940] = 32'b00000000000000000101110111100010;
assign LUT_1[59941] = 32'b11111111111111111111001001011110;
assign LUT_1[59942] = 32'b00000000000000000001100101110011;
assign LUT_1[59943] = 32'b11111111111111111010110111101111;
assign LUT_1[59944] = 32'b11111111111111111101001100000000;
assign LUT_1[59945] = 32'b11111111111111110110011101111100;
assign LUT_1[59946] = 32'b11111111111111111000111010010001;
assign LUT_1[59947] = 32'b11111111111111110010001100001101;
assign LUT_1[59948] = 32'b00000000000000000101000101010111;
assign LUT_1[59949] = 32'b11111111111111111110010111010011;
assign LUT_1[59950] = 32'b00000000000000000000110011101000;
assign LUT_1[59951] = 32'b11111111111111111010000101100100;
assign LUT_1[59952] = 32'b11111111111111111111111001101101;
assign LUT_1[59953] = 32'b11111111111111111001001011101001;
assign LUT_1[59954] = 32'b11111111111111111011100111111110;
assign LUT_1[59955] = 32'b11111111111111110100111001111010;
assign LUT_1[59956] = 32'b00000000000000000111110011000100;
assign LUT_1[59957] = 32'b00000000000000000001000101000000;
assign LUT_1[59958] = 32'b00000000000000000011100001010101;
assign LUT_1[59959] = 32'b11111111111111111100110011010001;
assign LUT_1[59960] = 32'b11111111111111111111000111100010;
assign LUT_1[59961] = 32'b11111111111111111000011001011110;
assign LUT_1[59962] = 32'b11111111111111111010110101110011;
assign LUT_1[59963] = 32'b11111111111111110100000111101111;
assign LUT_1[59964] = 32'b00000000000000000111000000111001;
assign LUT_1[59965] = 32'b00000000000000000000010010110101;
assign LUT_1[59966] = 32'b00000000000000000010101111001010;
assign LUT_1[59967] = 32'b11111111111111111100000001000110;
assign LUT_1[59968] = 32'b11111111111111111111000000110100;
assign LUT_1[59969] = 32'b11111111111111111000010010110000;
assign LUT_1[59970] = 32'b11111111111111111010101111000101;
assign LUT_1[59971] = 32'b11111111111111110100000001000001;
assign LUT_1[59972] = 32'b00000000000000000110111010001011;
assign LUT_1[59973] = 32'b00000000000000000000001100000111;
assign LUT_1[59974] = 32'b00000000000000000010101000011100;
assign LUT_1[59975] = 32'b11111111111111111011111010011000;
assign LUT_1[59976] = 32'b11111111111111111110001110101001;
assign LUT_1[59977] = 32'b11111111111111110111100000100101;
assign LUT_1[59978] = 32'b11111111111111111001111100111010;
assign LUT_1[59979] = 32'b11111111111111110011001110110110;
assign LUT_1[59980] = 32'b00000000000000000110001000000000;
assign LUT_1[59981] = 32'b11111111111111111111011001111100;
assign LUT_1[59982] = 32'b00000000000000000001110110010001;
assign LUT_1[59983] = 32'b11111111111111111011001000001101;
assign LUT_1[59984] = 32'b00000000000000000000111100010110;
assign LUT_1[59985] = 32'b11111111111111111010001110010010;
assign LUT_1[59986] = 32'b11111111111111111100101010100111;
assign LUT_1[59987] = 32'b11111111111111110101111100100011;
assign LUT_1[59988] = 32'b00000000000000001000110101101101;
assign LUT_1[59989] = 32'b00000000000000000010000111101001;
assign LUT_1[59990] = 32'b00000000000000000100100011111110;
assign LUT_1[59991] = 32'b11111111111111111101110101111010;
assign LUT_1[59992] = 32'b00000000000000000000001010001011;
assign LUT_1[59993] = 32'b11111111111111111001011100000111;
assign LUT_1[59994] = 32'b11111111111111111011111000011100;
assign LUT_1[59995] = 32'b11111111111111110101001010011000;
assign LUT_1[59996] = 32'b00000000000000001000000011100010;
assign LUT_1[59997] = 32'b00000000000000000001010101011110;
assign LUT_1[59998] = 32'b00000000000000000011110001110011;
assign LUT_1[59999] = 32'b11111111111111111101000011101111;
assign LUT_1[60000] = 32'b11111111111111111111111011110011;
assign LUT_1[60001] = 32'b11111111111111111001001101101111;
assign LUT_1[60002] = 32'b11111111111111111011101010000100;
assign LUT_1[60003] = 32'b11111111111111110100111100000000;
assign LUT_1[60004] = 32'b00000000000000000111110101001010;
assign LUT_1[60005] = 32'b00000000000000000001000111000110;
assign LUT_1[60006] = 32'b00000000000000000011100011011011;
assign LUT_1[60007] = 32'b11111111111111111100110101010111;
assign LUT_1[60008] = 32'b11111111111111111111001001101000;
assign LUT_1[60009] = 32'b11111111111111111000011011100100;
assign LUT_1[60010] = 32'b11111111111111111010110111111001;
assign LUT_1[60011] = 32'b11111111111111110100001001110101;
assign LUT_1[60012] = 32'b00000000000000000111000010111111;
assign LUT_1[60013] = 32'b00000000000000000000010100111011;
assign LUT_1[60014] = 32'b00000000000000000010110001010000;
assign LUT_1[60015] = 32'b11111111111111111100000011001100;
assign LUT_1[60016] = 32'b00000000000000000001110111010101;
assign LUT_1[60017] = 32'b11111111111111111011001001010001;
assign LUT_1[60018] = 32'b11111111111111111101100101100110;
assign LUT_1[60019] = 32'b11111111111111110110110111100010;
assign LUT_1[60020] = 32'b00000000000000001001110000101100;
assign LUT_1[60021] = 32'b00000000000000000011000010101000;
assign LUT_1[60022] = 32'b00000000000000000101011110111101;
assign LUT_1[60023] = 32'b11111111111111111110110000111001;
assign LUT_1[60024] = 32'b00000000000000000001000101001010;
assign LUT_1[60025] = 32'b11111111111111111010010111000110;
assign LUT_1[60026] = 32'b11111111111111111100110011011011;
assign LUT_1[60027] = 32'b11111111111111110110000101010111;
assign LUT_1[60028] = 32'b00000000000000001000111110100001;
assign LUT_1[60029] = 32'b00000000000000000010010000011101;
assign LUT_1[60030] = 32'b00000000000000000100101100110010;
assign LUT_1[60031] = 32'b11111111111111111101111110101110;
assign LUT_1[60032] = 32'b00000000000000000000000011001111;
assign LUT_1[60033] = 32'b11111111111111111001010101001011;
assign LUT_1[60034] = 32'b11111111111111111011110001100000;
assign LUT_1[60035] = 32'b11111111111111110101000011011100;
assign LUT_1[60036] = 32'b00000000000000000111111100100110;
assign LUT_1[60037] = 32'b00000000000000000001001110100010;
assign LUT_1[60038] = 32'b00000000000000000011101010110111;
assign LUT_1[60039] = 32'b11111111111111111100111100110011;
assign LUT_1[60040] = 32'b11111111111111111111010001000100;
assign LUT_1[60041] = 32'b11111111111111111000100011000000;
assign LUT_1[60042] = 32'b11111111111111111010111111010101;
assign LUT_1[60043] = 32'b11111111111111110100010001010001;
assign LUT_1[60044] = 32'b00000000000000000111001010011011;
assign LUT_1[60045] = 32'b00000000000000000000011100010111;
assign LUT_1[60046] = 32'b00000000000000000010111000101100;
assign LUT_1[60047] = 32'b11111111111111111100001010101000;
assign LUT_1[60048] = 32'b00000000000000000001111110110001;
assign LUT_1[60049] = 32'b11111111111111111011010000101101;
assign LUT_1[60050] = 32'b11111111111111111101101101000010;
assign LUT_1[60051] = 32'b11111111111111110110111110111110;
assign LUT_1[60052] = 32'b00000000000000001001111000001000;
assign LUT_1[60053] = 32'b00000000000000000011001010000100;
assign LUT_1[60054] = 32'b00000000000000000101100110011001;
assign LUT_1[60055] = 32'b11111111111111111110111000010101;
assign LUT_1[60056] = 32'b00000000000000000001001100100110;
assign LUT_1[60057] = 32'b11111111111111111010011110100010;
assign LUT_1[60058] = 32'b11111111111111111100111010110111;
assign LUT_1[60059] = 32'b11111111111111110110001100110011;
assign LUT_1[60060] = 32'b00000000000000001001000101111101;
assign LUT_1[60061] = 32'b00000000000000000010010111111001;
assign LUT_1[60062] = 32'b00000000000000000100110100001110;
assign LUT_1[60063] = 32'b11111111111111111110000110001010;
assign LUT_1[60064] = 32'b00000000000000000000111110001110;
assign LUT_1[60065] = 32'b11111111111111111010010000001010;
assign LUT_1[60066] = 32'b11111111111111111100101100011111;
assign LUT_1[60067] = 32'b11111111111111110101111110011011;
assign LUT_1[60068] = 32'b00000000000000001000110111100101;
assign LUT_1[60069] = 32'b00000000000000000010001001100001;
assign LUT_1[60070] = 32'b00000000000000000100100101110110;
assign LUT_1[60071] = 32'b11111111111111111101110111110010;
assign LUT_1[60072] = 32'b00000000000000000000001100000011;
assign LUT_1[60073] = 32'b11111111111111111001011101111111;
assign LUT_1[60074] = 32'b11111111111111111011111010010100;
assign LUT_1[60075] = 32'b11111111111111110101001100010000;
assign LUT_1[60076] = 32'b00000000000000001000000101011010;
assign LUT_1[60077] = 32'b00000000000000000001010111010110;
assign LUT_1[60078] = 32'b00000000000000000011110011101011;
assign LUT_1[60079] = 32'b11111111111111111101000101100111;
assign LUT_1[60080] = 32'b00000000000000000010111001110000;
assign LUT_1[60081] = 32'b11111111111111111100001011101100;
assign LUT_1[60082] = 32'b11111111111111111110101000000001;
assign LUT_1[60083] = 32'b11111111111111110111111001111101;
assign LUT_1[60084] = 32'b00000000000000001010110011000111;
assign LUT_1[60085] = 32'b00000000000000000100000101000011;
assign LUT_1[60086] = 32'b00000000000000000110100001011000;
assign LUT_1[60087] = 32'b11111111111111111111110011010100;
assign LUT_1[60088] = 32'b00000000000000000010000111100101;
assign LUT_1[60089] = 32'b11111111111111111011011001100001;
assign LUT_1[60090] = 32'b11111111111111111101110101110110;
assign LUT_1[60091] = 32'b11111111111111110111000111110010;
assign LUT_1[60092] = 32'b00000000000000001010000000111100;
assign LUT_1[60093] = 32'b00000000000000000011010010111000;
assign LUT_1[60094] = 32'b00000000000000000101101111001101;
assign LUT_1[60095] = 32'b11111111111111111111000001001001;
assign LUT_1[60096] = 32'b00000000000000000010000000110111;
assign LUT_1[60097] = 32'b11111111111111111011010010110011;
assign LUT_1[60098] = 32'b11111111111111111101101111001000;
assign LUT_1[60099] = 32'b11111111111111110111000001000100;
assign LUT_1[60100] = 32'b00000000000000001001111010001110;
assign LUT_1[60101] = 32'b00000000000000000011001100001010;
assign LUT_1[60102] = 32'b00000000000000000101101000011111;
assign LUT_1[60103] = 32'b11111111111111111110111010011011;
assign LUT_1[60104] = 32'b00000000000000000001001110101100;
assign LUT_1[60105] = 32'b11111111111111111010100000101000;
assign LUT_1[60106] = 32'b11111111111111111100111100111101;
assign LUT_1[60107] = 32'b11111111111111110110001110111001;
assign LUT_1[60108] = 32'b00000000000000001001001000000011;
assign LUT_1[60109] = 32'b00000000000000000010011001111111;
assign LUT_1[60110] = 32'b00000000000000000100110110010100;
assign LUT_1[60111] = 32'b11111111111111111110001000010000;
assign LUT_1[60112] = 32'b00000000000000000011111100011001;
assign LUT_1[60113] = 32'b11111111111111111101001110010101;
assign LUT_1[60114] = 32'b11111111111111111111101010101010;
assign LUT_1[60115] = 32'b11111111111111111000111100100110;
assign LUT_1[60116] = 32'b00000000000000001011110101110000;
assign LUT_1[60117] = 32'b00000000000000000101000111101100;
assign LUT_1[60118] = 32'b00000000000000000111100100000001;
assign LUT_1[60119] = 32'b00000000000000000000110101111101;
assign LUT_1[60120] = 32'b00000000000000000011001010001110;
assign LUT_1[60121] = 32'b11111111111111111100011100001010;
assign LUT_1[60122] = 32'b11111111111111111110111000011111;
assign LUT_1[60123] = 32'b11111111111111111000001010011011;
assign LUT_1[60124] = 32'b00000000000000001011000011100101;
assign LUT_1[60125] = 32'b00000000000000000100010101100001;
assign LUT_1[60126] = 32'b00000000000000000110110001110110;
assign LUT_1[60127] = 32'b00000000000000000000000011110010;
assign LUT_1[60128] = 32'b00000000000000000010111011110110;
assign LUT_1[60129] = 32'b11111111111111111100001101110010;
assign LUT_1[60130] = 32'b11111111111111111110101010000111;
assign LUT_1[60131] = 32'b11111111111111110111111100000011;
assign LUT_1[60132] = 32'b00000000000000001010110101001101;
assign LUT_1[60133] = 32'b00000000000000000100000111001001;
assign LUT_1[60134] = 32'b00000000000000000110100011011110;
assign LUT_1[60135] = 32'b11111111111111111111110101011010;
assign LUT_1[60136] = 32'b00000000000000000010001001101011;
assign LUT_1[60137] = 32'b11111111111111111011011011100111;
assign LUT_1[60138] = 32'b11111111111111111101110111111100;
assign LUT_1[60139] = 32'b11111111111111110111001001111000;
assign LUT_1[60140] = 32'b00000000000000001010000011000010;
assign LUT_1[60141] = 32'b00000000000000000011010100111110;
assign LUT_1[60142] = 32'b00000000000000000101110001010011;
assign LUT_1[60143] = 32'b11111111111111111111000011001111;
assign LUT_1[60144] = 32'b00000000000000000100110111011000;
assign LUT_1[60145] = 32'b11111111111111111110001001010100;
assign LUT_1[60146] = 32'b00000000000000000000100101101001;
assign LUT_1[60147] = 32'b11111111111111111001110111100101;
assign LUT_1[60148] = 32'b00000000000000001100110000101111;
assign LUT_1[60149] = 32'b00000000000000000110000010101011;
assign LUT_1[60150] = 32'b00000000000000001000011111000000;
assign LUT_1[60151] = 32'b00000000000000000001110000111100;
assign LUT_1[60152] = 32'b00000000000000000100000101001101;
assign LUT_1[60153] = 32'b11111111111111111101010111001001;
assign LUT_1[60154] = 32'b11111111111111111111110011011110;
assign LUT_1[60155] = 32'b11111111111111111001000101011010;
assign LUT_1[60156] = 32'b00000000000000001011111110100100;
assign LUT_1[60157] = 32'b00000000000000000101010000100000;
assign LUT_1[60158] = 32'b00000000000000000111101100110101;
assign LUT_1[60159] = 32'b00000000000000000000111110110001;
assign LUT_1[60160] = 32'b11111111111111111010110111011000;
assign LUT_1[60161] = 32'b11111111111111110100001001010100;
assign LUT_1[60162] = 32'b11111111111111110110100101101001;
assign LUT_1[60163] = 32'b11111111111111101111110111100101;
assign LUT_1[60164] = 32'b00000000000000000010110000101111;
assign LUT_1[60165] = 32'b11111111111111111100000010101011;
assign LUT_1[60166] = 32'b11111111111111111110011111000000;
assign LUT_1[60167] = 32'b11111111111111110111110000111100;
assign LUT_1[60168] = 32'b11111111111111111010000101001101;
assign LUT_1[60169] = 32'b11111111111111110011010111001001;
assign LUT_1[60170] = 32'b11111111111111110101110011011110;
assign LUT_1[60171] = 32'b11111111111111101111000101011010;
assign LUT_1[60172] = 32'b00000000000000000001111110100100;
assign LUT_1[60173] = 32'b11111111111111111011010000100000;
assign LUT_1[60174] = 32'b11111111111111111101101100110101;
assign LUT_1[60175] = 32'b11111111111111110110111110110001;
assign LUT_1[60176] = 32'b11111111111111111100110010111010;
assign LUT_1[60177] = 32'b11111111111111110110000100110110;
assign LUT_1[60178] = 32'b11111111111111111000100001001011;
assign LUT_1[60179] = 32'b11111111111111110001110011000111;
assign LUT_1[60180] = 32'b00000000000000000100101100010001;
assign LUT_1[60181] = 32'b11111111111111111101111110001101;
assign LUT_1[60182] = 32'b00000000000000000000011010100010;
assign LUT_1[60183] = 32'b11111111111111111001101100011110;
assign LUT_1[60184] = 32'b11111111111111111100000000101111;
assign LUT_1[60185] = 32'b11111111111111110101010010101011;
assign LUT_1[60186] = 32'b11111111111111110111101111000000;
assign LUT_1[60187] = 32'b11111111111111110001000000111100;
assign LUT_1[60188] = 32'b00000000000000000011111010000110;
assign LUT_1[60189] = 32'b11111111111111111101001100000010;
assign LUT_1[60190] = 32'b11111111111111111111101000010111;
assign LUT_1[60191] = 32'b11111111111111111000111010010011;
assign LUT_1[60192] = 32'b11111111111111111011110010010111;
assign LUT_1[60193] = 32'b11111111111111110101000100010011;
assign LUT_1[60194] = 32'b11111111111111110111100000101000;
assign LUT_1[60195] = 32'b11111111111111110000110010100100;
assign LUT_1[60196] = 32'b00000000000000000011101011101110;
assign LUT_1[60197] = 32'b11111111111111111100111101101010;
assign LUT_1[60198] = 32'b11111111111111111111011001111111;
assign LUT_1[60199] = 32'b11111111111111111000101011111011;
assign LUT_1[60200] = 32'b11111111111111111011000000001100;
assign LUT_1[60201] = 32'b11111111111111110100010010001000;
assign LUT_1[60202] = 32'b11111111111111110110101110011101;
assign LUT_1[60203] = 32'b11111111111111110000000000011001;
assign LUT_1[60204] = 32'b00000000000000000010111001100011;
assign LUT_1[60205] = 32'b11111111111111111100001011011111;
assign LUT_1[60206] = 32'b11111111111111111110100111110100;
assign LUT_1[60207] = 32'b11111111111111110111111001110000;
assign LUT_1[60208] = 32'b11111111111111111101101101111001;
assign LUT_1[60209] = 32'b11111111111111110110111111110101;
assign LUT_1[60210] = 32'b11111111111111111001011100001010;
assign LUT_1[60211] = 32'b11111111111111110010101110000110;
assign LUT_1[60212] = 32'b00000000000000000101100111010000;
assign LUT_1[60213] = 32'b11111111111111111110111001001100;
assign LUT_1[60214] = 32'b00000000000000000001010101100001;
assign LUT_1[60215] = 32'b11111111111111111010100111011101;
assign LUT_1[60216] = 32'b11111111111111111100111011101110;
assign LUT_1[60217] = 32'b11111111111111110110001101101010;
assign LUT_1[60218] = 32'b11111111111111111000101001111111;
assign LUT_1[60219] = 32'b11111111111111110001111011111011;
assign LUT_1[60220] = 32'b00000000000000000100110101000101;
assign LUT_1[60221] = 32'b11111111111111111110000111000001;
assign LUT_1[60222] = 32'b00000000000000000000100011010110;
assign LUT_1[60223] = 32'b11111111111111111001110101010010;
assign LUT_1[60224] = 32'b11111111111111111100110101000000;
assign LUT_1[60225] = 32'b11111111111111110110000110111100;
assign LUT_1[60226] = 32'b11111111111111111000100011010001;
assign LUT_1[60227] = 32'b11111111111111110001110101001101;
assign LUT_1[60228] = 32'b00000000000000000100101110010111;
assign LUT_1[60229] = 32'b11111111111111111110000000010011;
assign LUT_1[60230] = 32'b00000000000000000000011100101000;
assign LUT_1[60231] = 32'b11111111111111111001101110100100;
assign LUT_1[60232] = 32'b11111111111111111100000010110101;
assign LUT_1[60233] = 32'b11111111111111110101010100110001;
assign LUT_1[60234] = 32'b11111111111111110111110001000110;
assign LUT_1[60235] = 32'b11111111111111110001000011000010;
assign LUT_1[60236] = 32'b00000000000000000011111100001100;
assign LUT_1[60237] = 32'b11111111111111111101001110001000;
assign LUT_1[60238] = 32'b11111111111111111111101010011101;
assign LUT_1[60239] = 32'b11111111111111111000111100011001;
assign LUT_1[60240] = 32'b11111111111111111110110000100010;
assign LUT_1[60241] = 32'b11111111111111111000000010011110;
assign LUT_1[60242] = 32'b11111111111111111010011110110011;
assign LUT_1[60243] = 32'b11111111111111110011110000101111;
assign LUT_1[60244] = 32'b00000000000000000110101001111001;
assign LUT_1[60245] = 32'b11111111111111111111111011110101;
assign LUT_1[60246] = 32'b00000000000000000010011000001010;
assign LUT_1[60247] = 32'b11111111111111111011101010000110;
assign LUT_1[60248] = 32'b11111111111111111101111110010111;
assign LUT_1[60249] = 32'b11111111111111110111010000010011;
assign LUT_1[60250] = 32'b11111111111111111001101100101000;
assign LUT_1[60251] = 32'b11111111111111110010111110100100;
assign LUT_1[60252] = 32'b00000000000000000101110111101110;
assign LUT_1[60253] = 32'b11111111111111111111001001101010;
assign LUT_1[60254] = 32'b00000000000000000001100101111111;
assign LUT_1[60255] = 32'b11111111111111111010110111111011;
assign LUT_1[60256] = 32'b11111111111111111101101111111111;
assign LUT_1[60257] = 32'b11111111111111110111000001111011;
assign LUT_1[60258] = 32'b11111111111111111001011110010000;
assign LUT_1[60259] = 32'b11111111111111110010110000001100;
assign LUT_1[60260] = 32'b00000000000000000101101001010110;
assign LUT_1[60261] = 32'b11111111111111111110111011010010;
assign LUT_1[60262] = 32'b00000000000000000001010111100111;
assign LUT_1[60263] = 32'b11111111111111111010101001100011;
assign LUT_1[60264] = 32'b11111111111111111100111101110100;
assign LUT_1[60265] = 32'b11111111111111110110001111110000;
assign LUT_1[60266] = 32'b11111111111111111000101100000101;
assign LUT_1[60267] = 32'b11111111111111110001111110000001;
assign LUT_1[60268] = 32'b00000000000000000100110111001011;
assign LUT_1[60269] = 32'b11111111111111111110001001000111;
assign LUT_1[60270] = 32'b00000000000000000000100101011100;
assign LUT_1[60271] = 32'b11111111111111111001110111011000;
assign LUT_1[60272] = 32'b11111111111111111111101011100001;
assign LUT_1[60273] = 32'b11111111111111111000111101011101;
assign LUT_1[60274] = 32'b11111111111111111011011001110010;
assign LUT_1[60275] = 32'b11111111111111110100101011101110;
assign LUT_1[60276] = 32'b00000000000000000111100100111000;
assign LUT_1[60277] = 32'b00000000000000000000110110110100;
assign LUT_1[60278] = 32'b00000000000000000011010011001001;
assign LUT_1[60279] = 32'b11111111111111111100100101000101;
assign LUT_1[60280] = 32'b11111111111111111110111001010110;
assign LUT_1[60281] = 32'b11111111111111111000001011010010;
assign LUT_1[60282] = 32'b11111111111111111010100111100111;
assign LUT_1[60283] = 32'b11111111111111110011111001100011;
assign LUT_1[60284] = 32'b00000000000000000110110010101101;
assign LUT_1[60285] = 32'b00000000000000000000000100101001;
assign LUT_1[60286] = 32'b00000000000000000010100000111110;
assign LUT_1[60287] = 32'b11111111111111111011110010111010;
assign LUT_1[60288] = 32'b11111111111111111101110111011011;
assign LUT_1[60289] = 32'b11111111111111110111001001010111;
assign LUT_1[60290] = 32'b11111111111111111001100101101100;
assign LUT_1[60291] = 32'b11111111111111110010110111101000;
assign LUT_1[60292] = 32'b00000000000000000101110000110010;
assign LUT_1[60293] = 32'b11111111111111111111000010101110;
assign LUT_1[60294] = 32'b00000000000000000001011111000011;
assign LUT_1[60295] = 32'b11111111111111111010110000111111;
assign LUT_1[60296] = 32'b11111111111111111101000101010000;
assign LUT_1[60297] = 32'b11111111111111110110010111001100;
assign LUT_1[60298] = 32'b11111111111111111000110011100001;
assign LUT_1[60299] = 32'b11111111111111110010000101011101;
assign LUT_1[60300] = 32'b00000000000000000100111110100111;
assign LUT_1[60301] = 32'b11111111111111111110010000100011;
assign LUT_1[60302] = 32'b00000000000000000000101100111000;
assign LUT_1[60303] = 32'b11111111111111111001111110110100;
assign LUT_1[60304] = 32'b11111111111111111111110010111101;
assign LUT_1[60305] = 32'b11111111111111111001000100111001;
assign LUT_1[60306] = 32'b11111111111111111011100001001110;
assign LUT_1[60307] = 32'b11111111111111110100110011001010;
assign LUT_1[60308] = 32'b00000000000000000111101100010100;
assign LUT_1[60309] = 32'b00000000000000000000111110010000;
assign LUT_1[60310] = 32'b00000000000000000011011010100101;
assign LUT_1[60311] = 32'b11111111111111111100101100100001;
assign LUT_1[60312] = 32'b11111111111111111111000000110010;
assign LUT_1[60313] = 32'b11111111111111111000010010101110;
assign LUT_1[60314] = 32'b11111111111111111010101111000011;
assign LUT_1[60315] = 32'b11111111111111110100000000111111;
assign LUT_1[60316] = 32'b00000000000000000110111010001001;
assign LUT_1[60317] = 32'b00000000000000000000001100000101;
assign LUT_1[60318] = 32'b00000000000000000010101000011010;
assign LUT_1[60319] = 32'b11111111111111111011111010010110;
assign LUT_1[60320] = 32'b11111111111111111110110010011010;
assign LUT_1[60321] = 32'b11111111111111111000000100010110;
assign LUT_1[60322] = 32'b11111111111111111010100000101011;
assign LUT_1[60323] = 32'b11111111111111110011110010100111;
assign LUT_1[60324] = 32'b00000000000000000110101011110001;
assign LUT_1[60325] = 32'b11111111111111111111111101101101;
assign LUT_1[60326] = 32'b00000000000000000010011010000010;
assign LUT_1[60327] = 32'b11111111111111111011101011111110;
assign LUT_1[60328] = 32'b11111111111111111110000000001111;
assign LUT_1[60329] = 32'b11111111111111110111010010001011;
assign LUT_1[60330] = 32'b11111111111111111001101110100000;
assign LUT_1[60331] = 32'b11111111111111110011000000011100;
assign LUT_1[60332] = 32'b00000000000000000101111001100110;
assign LUT_1[60333] = 32'b11111111111111111111001011100010;
assign LUT_1[60334] = 32'b00000000000000000001100111110111;
assign LUT_1[60335] = 32'b11111111111111111010111001110011;
assign LUT_1[60336] = 32'b00000000000000000000101101111100;
assign LUT_1[60337] = 32'b11111111111111111001111111111000;
assign LUT_1[60338] = 32'b11111111111111111100011100001101;
assign LUT_1[60339] = 32'b11111111111111110101101110001001;
assign LUT_1[60340] = 32'b00000000000000001000100111010011;
assign LUT_1[60341] = 32'b00000000000000000001111001001111;
assign LUT_1[60342] = 32'b00000000000000000100010101100100;
assign LUT_1[60343] = 32'b11111111111111111101100111100000;
assign LUT_1[60344] = 32'b11111111111111111111111011110001;
assign LUT_1[60345] = 32'b11111111111111111001001101101101;
assign LUT_1[60346] = 32'b11111111111111111011101010000010;
assign LUT_1[60347] = 32'b11111111111111110100111011111110;
assign LUT_1[60348] = 32'b00000000000000000111110101001000;
assign LUT_1[60349] = 32'b00000000000000000001000111000100;
assign LUT_1[60350] = 32'b00000000000000000011100011011001;
assign LUT_1[60351] = 32'b11111111111111111100110101010101;
assign LUT_1[60352] = 32'b11111111111111111111110101000011;
assign LUT_1[60353] = 32'b11111111111111111001000110111111;
assign LUT_1[60354] = 32'b11111111111111111011100011010100;
assign LUT_1[60355] = 32'b11111111111111110100110101010000;
assign LUT_1[60356] = 32'b00000000000000000111101110011010;
assign LUT_1[60357] = 32'b00000000000000000001000000010110;
assign LUT_1[60358] = 32'b00000000000000000011011100101011;
assign LUT_1[60359] = 32'b11111111111111111100101110100111;
assign LUT_1[60360] = 32'b11111111111111111111000010111000;
assign LUT_1[60361] = 32'b11111111111111111000010100110100;
assign LUT_1[60362] = 32'b11111111111111111010110001001001;
assign LUT_1[60363] = 32'b11111111111111110100000011000101;
assign LUT_1[60364] = 32'b00000000000000000110111100001111;
assign LUT_1[60365] = 32'b00000000000000000000001110001011;
assign LUT_1[60366] = 32'b00000000000000000010101010100000;
assign LUT_1[60367] = 32'b11111111111111111011111100011100;
assign LUT_1[60368] = 32'b00000000000000000001110000100101;
assign LUT_1[60369] = 32'b11111111111111111011000010100001;
assign LUT_1[60370] = 32'b11111111111111111101011110110110;
assign LUT_1[60371] = 32'b11111111111111110110110000110010;
assign LUT_1[60372] = 32'b00000000000000001001101001111100;
assign LUT_1[60373] = 32'b00000000000000000010111011111000;
assign LUT_1[60374] = 32'b00000000000000000101011000001101;
assign LUT_1[60375] = 32'b11111111111111111110101010001001;
assign LUT_1[60376] = 32'b00000000000000000000111110011010;
assign LUT_1[60377] = 32'b11111111111111111010010000010110;
assign LUT_1[60378] = 32'b11111111111111111100101100101011;
assign LUT_1[60379] = 32'b11111111111111110101111110100111;
assign LUT_1[60380] = 32'b00000000000000001000110111110001;
assign LUT_1[60381] = 32'b00000000000000000010001001101101;
assign LUT_1[60382] = 32'b00000000000000000100100110000010;
assign LUT_1[60383] = 32'b11111111111111111101110111111110;
assign LUT_1[60384] = 32'b00000000000000000000110000000010;
assign LUT_1[60385] = 32'b11111111111111111010000001111110;
assign LUT_1[60386] = 32'b11111111111111111100011110010011;
assign LUT_1[60387] = 32'b11111111111111110101110000001111;
assign LUT_1[60388] = 32'b00000000000000001000101001011001;
assign LUT_1[60389] = 32'b00000000000000000001111011010101;
assign LUT_1[60390] = 32'b00000000000000000100010111101010;
assign LUT_1[60391] = 32'b11111111111111111101101001100110;
assign LUT_1[60392] = 32'b11111111111111111111111101110111;
assign LUT_1[60393] = 32'b11111111111111111001001111110011;
assign LUT_1[60394] = 32'b11111111111111111011101100001000;
assign LUT_1[60395] = 32'b11111111111111110100111110000100;
assign LUT_1[60396] = 32'b00000000000000000111110111001110;
assign LUT_1[60397] = 32'b00000000000000000001001001001010;
assign LUT_1[60398] = 32'b00000000000000000011100101011111;
assign LUT_1[60399] = 32'b11111111111111111100110111011011;
assign LUT_1[60400] = 32'b00000000000000000010101011100100;
assign LUT_1[60401] = 32'b11111111111111111011111101100000;
assign LUT_1[60402] = 32'b11111111111111111110011001110101;
assign LUT_1[60403] = 32'b11111111111111110111101011110001;
assign LUT_1[60404] = 32'b00000000000000001010100100111011;
assign LUT_1[60405] = 32'b00000000000000000011110110110111;
assign LUT_1[60406] = 32'b00000000000000000110010011001100;
assign LUT_1[60407] = 32'b11111111111111111111100101001000;
assign LUT_1[60408] = 32'b00000000000000000001111001011001;
assign LUT_1[60409] = 32'b11111111111111111011001011010101;
assign LUT_1[60410] = 32'b11111111111111111101100111101010;
assign LUT_1[60411] = 32'b11111111111111110110111001100110;
assign LUT_1[60412] = 32'b00000000000000001001110010110000;
assign LUT_1[60413] = 32'b00000000000000000011000100101100;
assign LUT_1[60414] = 32'b00000000000000000101100001000001;
assign LUT_1[60415] = 32'b11111111111111111110110010111101;
assign LUT_1[60416] = 32'b00000000000000001001101011011111;
assign LUT_1[60417] = 32'b00000000000000000010111101011011;
assign LUT_1[60418] = 32'b00000000000000000101011001110000;
assign LUT_1[60419] = 32'b11111111111111111110101011101100;
assign LUT_1[60420] = 32'b00000000000000010001100100110110;
assign LUT_1[60421] = 32'b00000000000000001010110110110010;
assign LUT_1[60422] = 32'b00000000000000001101010011000111;
assign LUT_1[60423] = 32'b00000000000000000110100101000011;
assign LUT_1[60424] = 32'b00000000000000001000111001010100;
assign LUT_1[60425] = 32'b00000000000000000010001011010000;
assign LUT_1[60426] = 32'b00000000000000000100100111100101;
assign LUT_1[60427] = 32'b11111111111111111101111001100001;
assign LUT_1[60428] = 32'b00000000000000010000110010101011;
assign LUT_1[60429] = 32'b00000000000000001010000100100111;
assign LUT_1[60430] = 32'b00000000000000001100100000111100;
assign LUT_1[60431] = 32'b00000000000000000101110010111000;
assign LUT_1[60432] = 32'b00000000000000001011100111000001;
assign LUT_1[60433] = 32'b00000000000000000100111000111101;
assign LUT_1[60434] = 32'b00000000000000000111010101010010;
assign LUT_1[60435] = 32'b00000000000000000000100111001110;
assign LUT_1[60436] = 32'b00000000000000010011100000011000;
assign LUT_1[60437] = 32'b00000000000000001100110010010100;
assign LUT_1[60438] = 32'b00000000000000001111001110101001;
assign LUT_1[60439] = 32'b00000000000000001000100000100101;
assign LUT_1[60440] = 32'b00000000000000001010110100110110;
assign LUT_1[60441] = 32'b00000000000000000100000110110010;
assign LUT_1[60442] = 32'b00000000000000000110100011000111;
assign LUT_1[60443] = 32'b11111111111111111111110101000011;
assign LUT_1[60444] = 32'b00000000000000010010101110001101;
assign LUT_1[60445] = 32'b00000000000000001100000000001001;
assign LUT_1[60446] = 32'b00000000000000001110011100011110;
assign LUT_1[60447] = 32'b00000000000000000111101110011010;
assign LUT_1[60448] = 32'b00000000000000001010100110011110;
assign LUT_1[60449] = 32'b00000000000000000011111000011010;
assign LUT_1[60450] = 32'b00000000000000000110010100101111;
assign LUT_1[60451] = 32'b11111111111111111111100110101011;
assign LUT_1[60452] = 32'b00000000000000010010011111110101;
assign LUT_1[60453] = 32'b00000000000000001011110001110001;
assign LUT_1[60454] = 32'b00000000000000001110001110000110;
assign LUT_1[60455] = 32'b00000000000000000111100000000010;
assign LUT_1[60456] = 32'b00000000000000001001110100010011;
assign LUT_1[60457] = 32'b00000000000000000011000110001111;
assign LUT_1[60458] = 32'b00000000000000000101100010100100;
assign LUT_1[60459] = 32'b11111111111111111110110100100000;
assign LUT_1[60460] = 32'b00000000000000010001101101101010;
assign LUT_1[60461] = 32'b00000000000000001010111111100110;
assign LUT_1[60462] = 32'b00000000000000001101011011111011;
assign LUT_1[60463] = 32'b00000000000000000110101101110111;
assign LUT_1[60464] = 32'b00000000000000001100100010000000;
assign LUT_1[60465] = 32'b00000000000000000101110011111100;
assign LUT_1[60466] = 32'b00000000000000001000010000010001;
assign LUT_1[60467] = 32'b00000000000000000001100010001101;
assign LUT_1[60468] = 32'b00000000000000010100011011010111;
assign LUT_1[60469] = 32'b00000000000000001101101101010011;
assign LUT_1[60470] = 32'b00000000000000010000001001101000;
assign LUT_1[60471] = 32'b00000000000000001001011011100100;
assign LUT_1[60472] = 32'b00000000000000001011101111110101;
assign LUT_1[60473] = 32'b00000000000000000101000001110001;
assign LUT_1[60474] = 32'b00000000000000000111011110000110;
assign LUT_1[60475] = 32'b00000000000000000000110000000010;
assign LUT_1[60476] = 32'b00000000000000010011101001001100;
assign LUT_1[60477] = 32'b00000000000000001100111011001000;
assign LUT_1[60478] = 32'b00000000000000001111010111011101;
assign LUT_1[60479] = 32'b00000000000000001000101001011001;
assign LUT_1[60480] = 32'b00000000000000001011101001000111;
assign LUT_1[60481] = 32'b00000000000000000100111011000011;
assign LUT_1[60482] = 32'b00000000000000000111010111011000;
assign LUT_1[60483] = 32'b00000000000000000000101001010100;
assign LUT_1[60484] = 32'b00000000000000010011100010011110;
assign LUT_1[60485] = 32'b00000000000000001100110100011010;
assign LUT_1[60486] = 32'b00000000000000001111010000101111;
assign LUT_1[60487] = 32'b00000000000000001000100010101011;
assign LUT_1[60488] = 32'b00000000000000001010110110111100;
assign LUT_1[60489] = 32'b00000000000000000100001000111000;
assign LUT_1[60490] = 32'b00000000000000000110100101001101;
assign LUT_1[60491] = 32'b11111111111111111111110111001001;
assign LUT_1[60492] = 32'b00000000000000010010110000010011;
assign LUT_1[60493] = 32'b00000000000000001100000010001111;
assign LUT_1[60494] = 32'b00000000000000001110011110100100;
assign LUT_1[60495] = 32'b00000000000000000111110000100000;
assign LUT_1[60496] = 32'b00000000000000001101100100101001;
assign LUT_1[60497] = 32'b00000000000000000110110110100101;
assign LUT_1[60498] = 32'b00000000000000001001010010111010;
assign LUT_1[60499] = 32'b00000000000000000010100100110110;
assign LUT_1[60500] = 32'b00000000000000010101011110000000;
assign LUT_1[60501] = 32'b00000000000000001110101111111100;
assign LUT_1[60502] = 32'b00000000000000010001001100010001;
assign LUT_1[60503] = 32'b00000000000000001010011110001101;
assign LUT_1[60504] = 32'b00000000000000001100110010011110;
assign LUT_1[60505] = 32'b00000000000000000110000100011010;
assign LUT_1[60506] = 32'b00000000000000001000100000101111;
assign LUT_1[60507] = 32'b00000000000000000001110010101011;
assign LUT_1[60508] = 32'b00000000000000010100101011110101;
assign LUT_1[60509] = 32'b00000000000000001101111101110001;
assign LUT_1[60510] = 32'b00000000000000010000011010000110;
assign LUT_1[60511] = 32'b00000000000000001001101100000010;
assign LUT_1[60512] = 32'b00000000000000001100100100000110;
assign LUT_1[60513] = 32'b00000000000000000101110110000010;
assign LUT_1[60514] = 32'b00000000000000001000010010010111;
assign LUT_1[60515] = 32'b00000000000000000001100100010011;
assign LUT_1[60516] = 32'b00000000000000010100011101011101;
assign LUT_1[60517] = 32'b00000000000000001101101111011001;
assign LUT_1[60518] = 32'b00000000000000010000001011101110;
assign LUT_1[60519] = 32'b00000000000000001001011101101010;
assign LUT_1[60520] = 32'b00000000000000001011110001111011;
assign LUT_1[60521] = 32'b00000000000000000101000011110111;
assign LUT_1[60522] = 32'b00000000000000000111100000001100;
assign LUT_1[60523] = 32'b00000000000000000000110010001000;
assign LUT_1[60524] = 32'b00000000000000010011101011010010;
assign LUT_1[60525] = 32'b00000000000000001100111101001110;
assign LUT_1[60526] = 32'b00000000000000001111011001100011;
assign LUT_1[60527] = 32'b00000000000000001000101011011111;
assign LUT_1[60528] = 32'b00000000000000001110011111101000;
assign LUT_1[60529] = 32'b00000000000000000111110001100100;
assign LUT_1[60530] = 32'b00000000000000001010001101111001;
assign LUT_1[60531] = 32'b00000000000000000011011111110101;
assign LUT_1[60532] = 32'b00000000000000010110011000111111;
assign LUT_1[60533] = 32'b00000000000000001111101010111011;
assign LUT_1[60534] = 32'b00000000000000010010000111010000;
assign LUT_1[60535] = 32'b00000000000000001011011001001100;
assign LUT_1[60536] = 32'b00000000000000001101101101011101;
assign LUT_1[60537] = 32'b00000000000000000110111111011001;
assign LUT_1[60538] = 32'b00000000000000001001011011101110;
assign LUT_1[60539] = 32'b00000000000000000010101101101010;
assign LUT_1[60540] = 32'b00000000000000010101100110110100;
assign LUT_1[60541] = 32'b00000000000000001110111000110000;
assign LUT_1[60542] = 32'b00000000000000010001010101000101;
assign LUT_1[60543] = 32'b00000000000000001010100111000001;
assign LUT_1[60544] = 32'b00000000000000001100101011100010;
assign LUT_1[60545] = 32'b00000000000000000101111101011110;
assign LUT_1[60546] = 32'b00000000000000001000011001110011;
assign LUT_1[60547] = 32'b00000000000000000001101011101111;
assign LUT_1[60548] = 32'b00000000000000010100100100111001;
assign LUT_1[60549] = 32'b00000000000000001101110110110101;
assign LUT_1[60550] = 32'b00000000000000010000010011001010;
assign LUT_1[60551] = 32'b00000000000000001001100101000110;
assign LUT_1[60552] = 32'b00000000000000001011111001010111;
assign LUT_1[60553] = 32'b00000000000000000101001011010011;
assign LUT_1[60554] = 32'b00000000000000000111100111101000;
assign LUT_1[60555] = 32'b00000000000000000000111001100100;
assign LUT_1[60556] = 32'b00000000000000010011110010101110;
assign LUT_1[60557] = 32'b00000000000000001101000100101010;
assign LUT_1[60558] = 32'b00000000000000001111100000111111;
assign LUT_1[60559] = 32'b00000000000000001000110010111011;
assign LUT_1[60560] = 32'b00000000000000001110100111000100;
assign LUT_1[60561] = 32'b00000000000000000111111001000000;
assign LUT_1[60562] = 32'b00000000000000001010010101010101;
assign LUT_1[60563] = 32'b00000000000000000011100111010001;
assign LUT_1[60564] = 32'b00000000000000010110100000011011;
assign LUT_1[60565] = 32'b00000000000000001111110010010111;
assign LUT_1[60566] = 32'b00000000000000010010001110101100;
assign LUT_1[60567] = 32'b00000000000000001011100000101000;
assign LUT_1[60568] = 32'b00000000000000001101110100111001;
assign LUT_1[60569] = 32'b00000000000000000111000110110101;
assign LUT_1[60570] = 32'b00000000000000001001100011001010;
assign LUT_1[60571] = 32'b00000000000000000010110101000110;
assign LUT_1[60572] = 32'b00000000000000010101101110010000;
assign LUT_1[60573] = 32'b00000000000000001111000000001100;
assign LUT_1[60574] = 32'b00000000000000010001011100100001;
assign LUT_1[60575] = 32'b00000000000000001010101110011101;
assign LUT_1[60576] = 32'b00000000000000001101100110100001;
assign LUT_1[60577] = 32'b00000000000000000110111000011101;
assign LUT_1[60578] = 32'b00000000000000001001010100110010;
assign LUT_1[60579] = 32'b00000000000000000010100110101110;
assign LUT_1[60580] = 32'b00000000000000010101011111111000;
assign LUT_1[60581] = 32'b00000000000000001110110001110100;
assign LUT_1[60582] = 32'b00000000000000010001001110001001;
assign LUT_1[60583] = 32'b00000000000000001010100000000101;
assign LUT_1[60584] = 32'b00000000000000001100110100010110;
assign LUT_1[60585] = 32'b00000000000000000110000110010010;
assign LUT_1[60586] = 32'b00000000000000001000100010100111;
assign LUT_1[60587] = 32'b00000000000000000001110100100011;
assign LUT_1[60588] = 32'b00000000000000010100101101101101;
assign LUT_1[60589] = 32'b00000000000000001101111111101001;
assign LUT_1[60590] = 32'b00000000000000010000011011111110;
assign LUT_1[60591] = 32'b00000000000000001001101101111010;
assign LUT_1[60592] = 32'b00000000000000001111100010000011;
assign LUT_1[60593] = 32'b00000000000000001000110011111111;
assign LUT_1[60594] = 32'b00000000000000001011010000010100;
assign LUT_1[60595] = 32'b00000000000000000100100010010000;
assign LUT_1[60596] = 32'b00000000000000010111011011011010;
assign LUT_1[60597] = 32'b00000000000000010000101101010110;
assign LUT_1[60598] = 32'b00000000000000010011001001101011;
assign LUT_1[60599] = 32'b00000000000000001100011011100111;
assign LUT_1[60600] = 32'b00000000000000001110101111111000;
assign LUT_1[60601] = 32'b00000000000000001000000001110100;
assign LUT_1[60602] = 32'b00000000000000001010011110001001;
assign LUT_1[60603] = 32'b00000000000000000011110000000101;
assign LUT_1[60604] = 32'b00000000000000010110101001001111;
assign LUT_1[60605] = 32'b00000000000000001111111011001011;
assign LUT_1[60606] = 32'b00000000000000010010010111100000;
assign LUT_1[60607] = 32'b00000000000000001011101001011100;
assign LUT_1[60608] = 32'b00000000000000001110101001001010;
assign LUT_1[60609] = 32'b00000000000000000111111011000110;
assign LUT_1[60610] = 32'b00000000000000001010010111011011;
assign LUT_1[60611] = 32'b00000000000000000011101001010111;
assign LUT_1[60612] = 32'b00000000000000010110100010100001;
assign LUT_1[60613] = 32'b00000000000000001111110100011101;
assign LUT_1[60614] = 32'b00000000000000010010010000110010;
assign LUT_1[60615] = 32'b00000000000000001011100010101110;
assign LUT_1[60616] = 32'b00000000000000001101110110111111;
assign LUT_1[60617] = 32'b00000000000000000111001000111011;
assign LUT_1[60618] = 32'b00000000000000001001100101010000;
assign LUT_1[60619] = 32'b00000000000000000010110111001100;
assign LUT_1[60620] = 32'b00000000000000010101110000010110;
assign LUT_1[60621] = 32'b00000000000000001111000010010010;
assign LUT_1[60622] = 32'b00000000000000010001011110100111;
assign LUT_1[60623] = 32'b00000000000000001010110000100011;
assign LUT_1[60624] = 32'b00000000000000010000100100101100;
assign LUT_1[60625] = 32'b00000000000000001001110110101000;
assign LUT_1[60626] = 32'b00000000000000001100010010111101;
assign LUT_1[60627] = 32'b00000000000000000101100100111001;
assign LUT_1[60628] = 32'b00000000000000011000011110000011;
assign LUT_1[60629] = 32'b00000000000000010001101111111111;
assign LUT_1[60630] = 32'b00000000000000010100001100010100;
assign LUT_1[60631] = 32'b00000000000000001101011110010000;
assign LUT_1[60632] = 32'b00000000000000001111110010100001;
assign LUT_1[60633] = 32'b00000000000000001001000100011101;
assign LUT_1[60634] = 32'b00000000000000001011100000110010;
assign LUT_1[60635] = 32'b00000000000000000100110010101110;
assign LUT_1[60636] = 32'b00000000000000010111101011111000;
assign LUT_1[60637] = 32'b00000000000000010000111101110100;
assign LUT_1[60638] = 32'b00000000000000010011011010001001;
assign LUT_1[60639] = 32'b00000000000000001100101100000101;
assign LUT_1[60640] = 32'b00000000000000001111100100001001;
assign LUT_1[60641] = 32'b00000000000000001000110110000101;
assign LUT_1[60642] = 32'b00000000000000001011010010011010;
assign LUT_1[60643] = 32'b00000000000000000100100100010110;
assign LUT_1[60644] = 32'b00000000000000010111011101100000;
assign LUT_1[60645] = 32'b00000000000000010000101111011100;
assign LUT_1[60646] = 32'b00000000000000010011001011110001;
assign LUT_1[60647] = 32'b00000000000000001100011101101101;
assign LUT_1[60648] = 32'b00000000000000001110110001111110;
assign LUT_1[60649] = 32'b00000000000000001000000011111010;
assign LUT_1[60650] = 32'b00000000000000001010100000001111;
assign LUT_1[60651] = 32'b00000000000000000011110010001011;
assign LUT_1[60652] = 32'b00000000000000010110101011010101;
assign LUT_1[60653] = 32'b00000000000000001111111101010001;
assign LUT_1[60654] = 32'b00000000000000010010011001100110;
assign LUT_1[60655] = 32'b00000000000000001011101011100010;
assign LUT_1[60656] = 32'b00000000000000010001011111101011;
assign LUT_1[60657] = 32'b00000000000000001010110001100111;
assign LUT_1[60658] = 32'b00000000000000001101001101111100;
assign LUT_1[60659] = 32'b00000000000000000110011111111000;
assign LUT_1[60660] = 32'b00000000000000011001011001000010;
assign LUT_1[60661] = 32'b00000000000000010010101010111110;
assign LUT_1[60662] = 32'b00000000000000010101000111010011;
assign LUT_1[60663] = 32'b00000000000000001110011001001111;
assign LUT_1[60664] = 32'b00000000000000010000101101100000;
assign LUT_1[60665] = 32'b00000000000000001001111111011100;
assign LUT_1[60666] = 32'b00000000000000001100011011110001;
assign LUT_1[60667] = 32'b00000000000000000101101101101101;
assign LUT_1[60668] = 32'b00000000000000011000100110110111;
assign LUT_1[60669] = 32'b00000000000000010001111000110011;
assign LUT_1[60670] = 32'b00000000000000010100010101001000;
assign LUT_1[60671] = 32'b00000000000000001101100111000100;
assign LUT_1[60672] = 32'b00000000000000000111011111101011;
assign LUT_1[60673] = 32'b00000000000000000000110001100111;
assign LUT_1[60674] = 32'b00000000000000000011001101111100;
assign LUT_1[60675] = 32'b11111111111111111100011111111000;
assign LUT_1[60676] = 32'b00000000000000001111011001000010;
assign LUT_1[60677] = 32'b00000000000000001000101010111110;
assign LUT_1[60678] = 32'b00000000000000001011000111010011;
assign LUT_1[60679] = 32'b00000000000000000100011001001111;
assign LUT_1[60680] = 32'b00000000000000000110101101100000;
assign LUT_1[60681] = 32'b11111111111111111111111111011100;
assign LUT_1[60682] = 32'b00000000000000000010011011110001;
assign LUT_1[60683] = 32'b11111111111111111011101101101101;
assign LUT_1[60684] = 32'b00000000000000001110100110110111;
assign LUT_1[60685] = 32'b00000000000000000111111000110011;
assign LUT_1[60686] = 32'b00000000000000001010010101001000;
assign LUT_1[60687] = 32'b00000000000000000011100111000100;
assign LUT_1[60688] = 32'b00000000000000001001011011001101;
assign LUT_1[60689] = 32'b00000000000000000010101101001001;
assign LUT_1[60690] = 32'b00000000000000000101001001011110;
assign LUT_1[60691] = 32'b11111111111111111110011011011010;
assign LUT_1[60692] = 32'b00000000000000010001010100100100;
assign LUT_1[60693] = 32'b00000000000000001010100110100000;
assign LUT_1[60694] = 32'b00000000000000001101000010110101;
assign LUT_1[60695] = 32'b00000000000000000110010100110001;
assign LUT_1[60696] = 32'b00000000000000001000101001000010;
assign LUT_1[60697] = 32'b00000000000000000001111010111110;
assign LUT_1[60698] = 32'b00000000000000000100010111010011;
assign LUT_1[60699] = 32'b11111111111111111101101001001111;
assign LUT_1[60700] = 32'b00000000000000010000100010011001;
assign LUT_1[60701] = 32'b00000000000000001001110100010101;
assign LUT_1[60702] = 32'b00000000000000001100010000101010;
assign LUT_1[60703] = 32'b00000000000000000101100010100110;
assign LUT_1[60704] = 32'b00000000000000001000011010101010;
assign LUT_1[60705] = 32'b00000000000000000001101100100110;
assign LUT_1[60706] = 32'b00000000000000000100001000111011;
assign LUT_1[60707] = 32'b11111111111111111101011010110111;
assign LUT_1[60708] = 32'b00000000000000010000010100000001;
assign LUT_1[60709] = 32'b00000000000000001001100101111101;
assign LUT_1[60710] = 32'b00000000000000001100000010010010;
assign LUT_1[60711] = 32'b00000000000000000101010100001110;
assign LUT_1[60712] = 32'b00000000000000000111101000011111;
assign LUT_1[60713] = 32'b00000000000000000000111010011011;
assign LUT_1[60714] = 32'b00000000000000000011010110110000;
assign LUT_1[60715] = 32'b11111111111111111100101000101100;
assign LUT_1[60716] = 32'b00000000000000001111100001110110;
assign LUT_1[60717] = 32'b00000000000000001000110011110010;
assign LUT_1[60718] = 32'b00000000000000001011010000000111;
assign LUT_1[60719] = 32'b00000000000000000100100010000011;
assign LUT_1[60720] = 32'b00000000000000001010010110001100;
assign LUT_1[60721] = 32'b00000000000000000011101000001000;
assign LUT_1[60722] = 32'b00000000000000000110000100011101;
assign LUT_1[60723] = 32'b11111111111111111111010110011001;
assign LUT_1[60724] = 32'b00000000000000010010001111100011;
assign LUT_1[60725] = 32'b00000000000000001011100001011111;
assign LUT_1[60726] = 32'b00000000000000001101111101110100;
assign LUT_1[60727] = 32'b00000000000000000111001111110000;
assign LUT_1[60728] = 32'b00000000000000001001100100000001;
assign LUT_1[60729] = 32'b00000000000000000010110101111101;
assign LUT_1[60730] = 32'b00000000000000000101010010010010;
assign LUT_1[60731] = 32'b11111111111111111110100100001110;
assign LUT_1[60732] = 32'b00000000000000010001011101011000;
assign LUT_1[60733] = 32'b00000000000000001010101111010100;
assign LUT_1[60734] = 32'b00000000000000001101001011101001;
assign LUT_1[60735] = 32'b00000000000000000110011101100101;
assign LUT_1[60736] = 32'b00000000000000001001011101010011;
assign LUT_1[60737] = 32'b00000000000000000010101111001111;
assign LUT_1[60738] = 32'b00000000000000000101001011100100;
assign LUT_1[60739] = 32'b11111111111111111110011101100000;
assign LUT_1[60740] = 32'b00000000000000010001010110101010;
assign LUT_1[60741] = 32'b00000000000000001010101000100110;
assign LUT_1[60742] = 32'b00000000000000001101000100111011;
assign LUT_1[60743] = 32'b00000000000000000110010110110111;
assign LUT_1[60744] = 32'b00000000000000001000101011001000;
assign LUT_1[60745] = 32'b00000000000000000001111101000100;
assign LUT_1[60746] = 32'b00000000000000000100011001011001;
assign LUT_1[60747] = 32'b11111111111111111101101011010101;
assign LUT_1[60748] = 32'b00000000000000010000100100011111;
assign LUT_1[60749] = 32'b00000000000000001001110110011011;
assign LUT_1[60750] = 32'b00000000000000001100010010110000;
assign LUT_1[60751] = 32'b00000000000000000101100100101100;
assign LUT_1[60752] = 32'b00000000000000001011011000110101;
assign LUT_1[60753] = 32'b00000000000000000100101010110001;
assign LUT_1[60754] = 32'b00000000000000000111000111000110;
assign LUT_1[60755] = 32'b00000000000000000000011001000010;
assign LUT_1[60756] = 32'b00000000000000010011010010001100;
assign LUT_1[60757] = 32'b00000000000000001100100100001000;
assign LUT_1[60758] = 32'b00000000000000001111000000011101;
assign LUT_1[60759] = 32'b00000000000000001000010010011001;
assign LUT_1[60760] = 32'b00000000000000001010100110101010;
assign LUT_1[60761] = 32'b00000000000000000011111000100110;
assign LUT_1[60762] = 32'b00000000000000000110010100111011;
assign LUT_1[60763] = 32'b11111111111111111111100110110111;
assign LUT_1[60764] = 32'b00000000000000010010100000000001;
assign LUT_1[60765] = 32'b00000000000000001011110001111101;
assign LUT_1[60766] = 32'b00000000000000001110001110010010;
assign LUT_1[60767] = 32'b00000000000000000111100000001110;
assign LUT_1[60768] = 32'b00000000000000001010011000010010;
assign LUT_1[60769] = 32'b00000000000000000011101010001110;
assign LUT_1[60770] = 32'b00000000000000000110000110100011;
assign LUT_1[60771] = 32'b11111111111111111111011000011111;
assign LUT_1[60772] = 32'b00000000000000010010010001101001;
assign LUT_1[60773] = 32'b00000000000000001011100011100101;
assign LUT_1[60774] = 32'b00000000000000001101111111111010;
assign LUT_1[60775] = 32'b00000000000000000111010001110110;
assign LUT_1[60776] = 32'b00000000000000001001100110000111;
assign LUT_1[60777] = 32'b00000000000000000010111000000011;
assign LUT_1[60778] = 32'b00000000000000000101010100011000;
assign LUT_1[60779] = 32'b11111111111111111110100110010100;
assign LUT_1[60780] = 32'b00000000000000010001011111011110;
assign LUT_1[60781] = 32'b00000000000000001010110001011010;
assign LUT_1[60782] = 32'b00000000000000001101001101101111;
assign LUT_1[60783] = 32'b00000000000000000110011111101011;
assign LUT_1[60784] = 32'b00000000000000001100010011110100;
assign LUT_1[60785] = 32'b00000000000000000101100101110000;
assign LUT_1[60786] = 32'b00000000000000001000000010000101;
assign LUT_1[60787] = 32'b00000000000000000001010100000001;
assign LUT_1[60788] = 32'b00000000000000010100001101001011;
assign LUT_1[60789] = 32'b00000000000000001101011111000111;
assign LUT_1[60790] = 32'b00000000000000001111111011011100;
assign LUT_1[60791] = 32'b00000000000000001001001101011000;
assign LUT_1[60792] = 32'b00000000000000001011100001101001;
assign LUT_1[60793] = 32'b00000000000000000100110011100101;
assign LUT_1[60794] = 32'b00000000000000000111001111111010;
assign LUT_1[60795] = 32'b00000000000000000000100001110110;
assign LUT_1[60796] = 32'b00000000000000010011011011000000;
assign LUT_1[60797] = 32'b00000000000000001100101100111100;
assign LUT_1[60798] = 32'b00000000000000001111001001010001;
assign LUT_1[60799] = 32'b00000000000000001000011011001101;
assign LUT_1[60800] = 32'b00000000000000001010011111101110;
assign LUT_1[60801] = 32'b00000000000000000011110001101010;
assign LUT_1[60802] = 32'b00000000000000000110001101111111;
assign LUT_1[60803] = 32'b11111111111111111111011111111011;
assign LUT_1[60804] = 32'b00000000000000010010011001000101;
assign LUT_1[60805] = 32'b00000000000000001011101011000001;
assign LUT_1[60806] = 32'b00000000000000001110000111010110;
assign LUT_1[60807] = 32'b00000000000000000111011001010010;
assign LUT_1[60808] = 32'b00000000000000001001101101100011;
assign LUT_1[60809] = 32'b00000000000000000010111111011111;
assign LUT_1[60810] = 32'b00000000000000000101011011110100;
assign LUT_1[60811] = 32'b11111111111111111110101101110000;
assign LUT_1[60812] = 32'b00000000000000010001100110111010;
assign LUT_1[60813] = 32'b00000000000000001010111000110110;
assign LUT_1[60814] = 32'b00000000000000001101010101001011;
assign LUT_1[60815] = 32'b00000000000000000110100111000111;
assign LUT_1[60816] = 32'b00000000000000001100011011010000;
assign LUT_1[60817] = 32'b00000000000000000101101101001100;
assign LUT_1[60818] = 32'b00000000000000001000001001100001;
assign LUT_1[60819] = 32'b00000000000000000001011011011101;
assign LUT_1[60820] = 32'b00000000000000010100010100100111;
assign LUT_1[60821] = 32'b00000000000000001101100110100011;
assign LUT_1[60822] = 32'b00000000000000010000000010111000;
assign LUT_1[60823] = 32'b00000000000000001001010100110100;
assign LUT_1[60824] = 32'b00000000000000001011101001000101;
assign LUT_1[60825] = 32'b00000000000000000100111011000001;
assign LUT_1[60826] = 32'b00000000000000000111010111010110;
assign LUT_1[60827] = 32'b00000000000000000000101001010010;
assign LUT_1[60828] = 32'b00000000000000010011100010011100;
assign LUT_1[60829] = 32'b00000000000000001100110100011000;
assign LUT_1[60830] = 32'b00000000000000001111010000101101;
assign LUT_1[60831] = 32'b00000000000000001000100010101001;
assign LUT_1[60832] = 32'b00000000000000001011011010101101;
assign LUT_1[60833] = 32'b00000000000000000100101100101001;
assign LUT_1[60834] = 32'b00000000000000000111001000111110;
assign LUT_1[60835] = 32'b00000000000000000000011010111010;
assign LUT_1[60836] = 32'b00000000000000010011010100000100;
assign LUT_1[60837] = 32'b00000000000000001100100110000000;
assign LUT_1[60838] = 32'b00000000000000001111000010010101;
assign LUT_1[60839] = 32'b00000000000000001000010100010001;
assign LUT_1[60840] = 32'b00000000000000001010101000100010;
assign LUT_1[60841] = 32'b00000000000000000011111010011110;
assign LUT_1[60842] = 32'b00000000000000000110010110110011;
assign LUT_1[60843] = 32'b11111111111111111111101000101111;
assign LUT_1[60844] = 32'b00000000000000010010100001111001;
assign LUT_1[60845] = 32'b00000000000000001011110011110101;
assign LUT_1[60846] = 32'b00000000000000001110010000001010;
assign LUT_1[60847] = 32'b00000000000000000111100010000110;
assign LUT_1[60848] = 32'b00000000000000001101010110001111;
assign LUT_1[60849] = 32'b00000000000000000110101000001011;
assign LUT_1[60850] = 32'b00000000000000001001000100100000;
assign LUT_1[60851] = 32'b00000000000000000010010110011100;
assign LUT_1[60852] = 32'b00000000000000010101001111100110;
assign LUT_1[60853] = 32'b00000000000000001110100001100010;
assign LUT_1[60854] = 32'b00000000000000010000111101110111;
assign LUT_1[60855] = 32'b00000000000000001010001111110011;
assign LUT_1[60856] = 32'b00000000000000001100100100000100;
assign LUT_1[60857] = 32'b00000000000000000101110110000000;
assign LUT_1[60858] = 32'b00000000000000001000010010010101;
assign LUT_1[60859] = 32'b00000000000000000001100100010001;
assign LUT_1[60860] = 32'b00000000000000010100011101011011;
assign LUT_1[60861] = 32'b00000000000000001101101111010111;
assign LUT_1[60862] = 32'b00000000000000010000001011101100;
assign LUT_1[60863] = 32'b00000000000000001001011101101000;
assign LUT_1[60864] = 32'b00000000000000001100011101010110;
assign LUT_1[60865] = 32'b00000000000000000101101111010010;
assign LUT_1[60866] = 32'b00000000000000001000001011100111;
assign LUT_1[60867] = 32'b00000000000000000001011101100011;
assign LUT_1[60868] = 32'b00000000000000010100010110101101;
assign LUT_1[60869] = 32'b00000000000000001101101000101001;
assign LUT_1[60870] = 32'b00000000000000010000000100111110;
assign LUT_1[60871] = 32'b00000000000000001001010110111010;
assign LUT_1[60872] = 32'b00000000000000001011101011001011;
assign LUT_1[60873] = 32'b00000000000000000100111101000111;
assign LUT_1[60874] = 32'b00000000000000000111011001011100;
assign LUT_1[60875] = 32'b00000000000000000000101011011000;
assign LUT_1[60876] = 32'b00000000000000010011100100100010;
assign LUT_1[60877] = 32'b00000000000000001100110110011110;
assign LUT_1[60878] = 32'b00000000000000001111010010110011;
assign LUT_1[60879] = 32'b00000000000000001000100100101111;
assign LUT_1[60880] = 32'b00000000000000001110011000111000;
assign LUT_1[60881] = 32'b00000000000000000111101010110100;
assign LUT_1[60882] = 32'b00000000000000001010000111001001;
assign LUT_1[60883] = 32'b00000000000000000011011001000101;
assign LUT_1[60884] = 32'b00000000000000010110010010001111;
assign LUT_1[60885] = 32'b00000000000000001111100100001011;
assign LUT_1[60886] = 32'b00000000000000010010000000100000;
assign LUT_1[60887] = 32'b00000000000000001011010010011100;
assign LUT_1[60888] = 32'b00000000000000001101100110101101;
assign LUT_1[60889] = 32'b00000000000000000110111000101001;
assign LUT_1[60890] = 32'b00000000000000001001010100111110;
assign LUT_1[60891] = 32'b00000000000000000010100110111010;
assign LUT_1[60892] = 32'b00000000000000010101100000000100;
assign LUT_1[60893] = 32'b00000000000000001110110010000000;
assign LUT_1[60894] = 32'b00000000000000010001001110010101;
assign LUT_1[60895] = 32'b00000000000000001010100000010001;
assign LUT_1[60896] = 32'b00000000000000001101011000010101;
assign LUT_1[60897] = 32'b00000000000000000110101010010001;
assign LUT_1[60898] = 32'b00000000000000001001000110100110;
assign LUT_1[60899] = 32'b00000000000000000010011000100010;
assign LUT_1[60900] = 32'b00000000000000010101010001101100;
assign LUT_1[60901] = 32'b00000000000000001110100011101000;
assign LUT_1[60902] = 32'b00000000000000010000111111111101;
assign LUT_1[60903] = 32'b00000000000000001010010001111001;
assign LUT_1[60904] = 32'b00000000000000001100100110001010;
assign LUT_1[60905] = 32'b00000000000000000101111000000110;
assign LUT_1[60906] = 32'b00000000000000001000010100011011;
assign LUT_1[60907] = 32'b00000000000000000001100110010111;
assign LUT_1[60908] = 32'b00000000000000010100011111100001;
assign LUT_1[60909] = 32'b00000000000000001101110001011101;
assign LUT_1[60910] = 32'b00000000000000010000001101110010;
assign LUT_1[60911] = 32'b00000000000000001001011111101110;
assign LUT_1[60912] = 32'b00000000000000001111010011110111;
assign LUT_1[60913] = 32'b00000000000000001000100101110011;
assign LUT_1[60914] = 32'b00000000000000001011000010001000;
assign LUT_1[60915] = 32'b00000000000000000100010100000100;
assign LUT_1[60916] = 32'b00000000000000010111001101001110;
assign LUT_1[60917] = 32'b00000000000000010000011111001010;
assign LUT_1[60918] = 32'b00000000000000010010111011011111;
assign LUT_1[60919] = 32'b00000000000000001100001101011011;
assign LUT_1[60920] = 32'b00000000000000001110100001101100;
assign LUT_1[60921] = 32'b00000000000000000111110011101000;
assign LUT_1[60922] = 32'b00000000000000001010001111111101;
assign LUT_1[60923] = 32'b00000000000000000011100001111001;
assign LUT_1[60924] = 32'b00000000000000010110011011000011;
assign LUT_1[60925] = 32'b00000000000000001111101100111111;
assign LUT_1[60926] = 32'b00000000000000010010001001010100;
assign LUT_1[60927] = 32'b00000000000000001011011011010000;
assign LUT_1[60928] = 32'b00000000000000000011011001111100;
assign LUT_1[60929] = 32'b11111111111111111100101011111000;
assign LUT_1[60930] = 32'b11111111111111111111001000001101;
assign LUT_1[60931] = 32'b11111111111111111000011010001001;
assign LUT_1[60932] = 32'b00000000000000001011010011010011;
assign LUT_1[60933] = 32'b00000000000000000100100101001111;
assign LUT_1[60934] = 32'b00000000000000000111000001100100;
assign LUT_1[60935] = 32'b00000000000000000000010011100000;
assign LUT_1[60936] = 32'b00000000000000000010100111110001;
assign LUT_1[60937] = 32'b11111111111111111011111001101101;
assign LUT_1[60938] = 32'b11111111111111111110010110000010;
assign LUT_1[60939] = 32'b11111111111111110111100111111110;
assign LUT_1[60940] = 32'b00000000000000001010100001001000;
assign LUT_1[60941] = 32'b00000000000000000011110011000100;
assign LUT_1[60942] = 32'b00000000000000000110001111011001;
assign LUT_1[60943] = 32'b11111111111111111111100001010101;
assign LUT_1[60944] = 32'b00000000000000000101010101011110;
assign LUT_1[60945] = 32'b11111111111111111110100111011010;
assign LUT_1[60946] = 32'b00000000000000000001000011101111;
assign LUT_1[60947] = 32'b11111111111111111010010101101011;
assign LUT_1[60948] = 32'b00000000000000001101001110110101;
assign LUT_1[60949] = 32'b00000000000000000110100000110001;
assign LUT_1[60950] = 32'b00000000000000001000111101000110;
assign LUT_1[60951] = 32'b00000000000000000010001111000010;
assign LUT_1[60952] = 32'b00000000000000000100100011010011;
assign LUT_1[60953] = 32'b11111111111111111101110101001111;
assign LUT_1[60954] = 32'b00000000000000000000010001100100;
assign LUT_1[60955] = 32'b11111111111111111001100011100000;
assign LUT_1[60956] = 32'b00000000000000001100011100101010;
assign LUT_1[60957] = 32'b00000000000000000101101110100110;
assign LUT_1[60958] = 32'b00000000000000001000001010111011;
assign LUT_1[60959] = 32'b00000000000000000001011100110111;
assign LUT_1[60960] = 32'b00000000000000000100010100111011;
assign LUT_1[60961] = 32'b11111111111111111101100110110111;
assign LUT_1[60962] = 32'b00000000000000000000000011001100;
assign LUT_1[60963] = 32'b11111111111111111001010101001000;
assign LUT_1[60964] = 32'b00000000000000001100001110010010;
assign LUT_1[60965] = 32'b00000000000000000101100000001110;
assign LUT_1[60966] = 32'b00000000000000000111111100100011;
assign LUT_1[60967] = 32'b00000000000000000001001110011111;
assign LUT_1[60968] = 32'b00000000000000000011100010110000;
assign LUT_1[60969] = 32'b11111111111111111100110100101100;
assign LUT_1[60970] = 32'b11111111111111111111010001000001;
assign LUT_1[60971] = 32'b11111111111111111000100010111101;
assign LUT_1[60972] = 32'b00000000000000001011011100000111;
assign LUT_1[60973] = 32'b00000000000000000100101110000011;
assign LUT_1[60974] = 32'b00000000000000000111001010011000;
assign LUT_1[60975] = 32'b00000000000000000000011100010100;
assign LUT_1[60976] = 32'b00000000000000000110010000011101;
assign LUT_1[60977] = 32'b11111111111111111111100010011001;
assign LUT_1[60978] = 32'b00000000000000000001111110101110;
assign LUT_1[60979] = 32'b11111111111111111011010000101010;
assign LUT_1[60980] = 32'b00000000000000001110001001110100;
assign LUT_1[60981] = 32'b00000000000000000111011011110000;
assign LUT_1[60982] = 32'b00000000000000001001111000000101;
assign LUT_1[60983] = 32'b00000000000000000011001010000001;
assign LUT_1[60984] = 32'b00000000000000000101011110010010;
assign LUT_1[60985] = 32'b11111111111111111110110000001110;
assign LUT_1[60986] = 32'b00000000000000000001001100100011;
assign LUT_1[60987] = 32'b11111111111111111010011110011111;
assign LUT_1[60988] = 32'b00000000000000001101010111101001;
assign LUT_1[60989] = 32'b00000000000000000110101001100101;
assign LUT_1[60990] = 32'b00000000000000001001000101111010;
assign LUT_1[60991] = 32'b00000000000000000010010111110110;
assign LUT_1[60992] = 32'b00000000000000000101010111100100;
assign LUT_1[60993] = 32'b11111111111111111110101001100000;
assign LUT_1[60994] = 32'b00000000000000000001000101110101;
assign LUT_1[60995] = 32'b11111111111111111010010111110001;
assign LUT_1[60996] = 32'b00000000000000001101010000111011;
assign LUT_1[60997] = 32'b00000000000000000110100010110111;
assign LUT_1[60998] = 32'b00000000000000001000111111001100;
assign LUT_1[60999] = 32'b00000000000000000010010001001000;
assign LUT_1[61000] = 32'b00000000000000000100100101011001;
assign LUT_1[61001] = 32'b11111111111111111101110111010101;
assign LUT_1[61002] = 32'b00000000000000000000010011101010;
assign LUT_1[61003] = 32'b11111111111111111001100101100110;
assign LUT_1[61004] = 32'b00000000000000001100011110110000;
assign LUT_1[61005] = 32'b00000000000000000101110000101100;
assign LUT_1[61006] = 32'b00000000000000001000001101000001;
assign LUT_1[61007] = 32'b00000000000000000001011110111101;
assign LUT_1[61008] = 32'b00000000000000000111010011000110;
assign LUT_1[61009] = 32'b00000000000000000000100101000010;
assign LUT_1[61010] = 32'b00000000000000000011000001010111;
assign LUT_1[61011] = 32'b11111111111111111100010011010011;
assign LUT_1[61012] = 32'b00000000000000001111001100011101;
assign LUT_1[61013] = 32'b00000000000000001000011110011001;
assign LUT_1[61014] = 32'b00000000000000001010111010101110;
assign LUT_1[61015] = 32'b00000000000000000100001100101010;
assign LUT_1[61016] = 32'b00000000000000000110100000111011;
assign LUT_1[61017] = 32'b11111111111111111111110010110111;
assign LUT_1[61018] = 32'b00000000000000000010001111001100;
assign LUT_1[61019] = 32'b11111111111111111011100001001000;
assign LUT_1[61020] = 32'b00000000000000001110011010010010;
assign LUT_1[61021] = 32'b00000000000000000111101100001110;
assign LUT_1[61022] = 32'b00000000000000001010001000100011;
assign LUT_1[61023] = 32'b00000000000000000011011010011111;
assign LUT_1[61024] = 32'b00000000000000000110010010100011;
assign LUT_1[61025] = 32'b11111111111111111111100100011111;
assign LUT_1[61026] = 32'b00000000000000000010000000110100;
assign LUT_1[61027] = 32'b11111111111111111011010010110000;
assign LUT_1[61028] = 32'b00000000000000001110001011111010;
assign LUT_1[61029] = 32'b00000000000000000111011101110110;
assign LUT_1[61030] = 32'b00000000000000001001111010001011;
assign LUT_1[61031] = 32'b00000000000000000011001100000111;
assign LUT_1[61032] = 32'b00000000000000000101100000011000;
assign LUT_1[61033] = 32'b11111111111111111110110010010100;
assign LUT_1[61034] = 32'b00000000000000000001001110101001;
assign LUT_1[61035] = 32'b11111111111111111010100000100101;
assign LUT_1[61036] = 32'b00000000000000001101011001101111;
assign LUT_1[61037] = 32'b00000000000000000110101011101011;
assign LUT_1[61038] = 32'b00000000000000001001001000000000;
assign LUT_1[61039] = 32'b00000000000000000010011001111100;
assign LUT_1[61040] = 32'b00000000000000001000001110000101;
assign LUT_1[61041] = 32'b00000000000000000001100000000001;
assign LUT_1[61042] = 32'b00000000000000000011111100010110;
assign LUT_1[61043] = 32'b11111111111111111101001110010010;
assign LUT_1[61044] = 32'b00000000000000010000000111011100;
assign LUT_1[61045] = 32'b00000000000000001001011001011000;
assign LUT_1[61046] = 32'b00000000000000001011110101101101;
assign LUT_1[61047] = 32'b00000000000000000101000111101001;
assign LUT_1[61048] = 32'b00000000000000000111011011111010;
assign LUT_1[61049] = 32'b00000000000000000000101101110110;
assign LUT_1[61050] = 32'b00000000000000000011001010001011;
assign LUT_1[61051] = 32'b11111111111111111100011100000111;
assign LUT_1[61052] = 32'b00000000000000001111010101010001;
assign LUT_1[61053] = 32'b00000000000000001000100111001101;
assign LUT_1[61054] = 32'b00000000000000001011000011100010;
assign LUT_1[61055] = 32'b00000000000000000100010101011110;
assign LUT_1[61056] = 32'b00000000000000000110011001111111;
assign LUT_1[61057] = 32'b11111111111111111111101011111011;
assign LUT_1[61058] = 32'b00000000000000000010001000010000;
assign LUT_1[61059] = 32'b11111111111111111011011010001100;
assign LUT_1[61060] = 32'b00000000000000001110010011010110;
assign LUT_1[61061] = 32'b00000000000000000111100101010010;
assign LUT_1[61062] = 32'b00000000000000001010000001100111;
assign LUT_1[61063] = 32'b00000000000000000011010011100011;
assign LUT_1[61064] = 32'b00000000000000000101100111110100;
assign LUT_1[61065] = 32'b11111111111111111110111001110000;
assign LUT_1[61066] = 32'b00000000000000000001010110000101;
assign LUT_1[61067] = 32'b11111111111111111010101000000001;
assign LUT_1[61068] = 32'b00000000000000001101100001001011;
assign LUT_1[61069] = 32'b00000000000000000110110011000111;
assign LUT_1[61070] = 32'b00000000000000001001001111011100;
assign LUT_1[61071] = 32'b00000000000000000010100001011000;
assign LUT_1[61072] = 32'b00000000000000001000010101100001;
assign LUT_1[61073] = 32'b00000000000000000001100111011101;
assign LUT_1[61074] = 32'b00000000000000000100000011110010;
assign LUT_1[61075] = 32'b11111111111111111101010101101110;
assign LUT_1[61076] = 32'b00000000000000010000001110111000;
assign LUT_1[61077] = 32'b00000000000000001001100000110100;
assign LUT_1[61078] = 32'b00000000000000001011111101001001;
assign LUT_1[61079] = 32'b00000000000000000101001111000101;
assign LUT_1[61080] = 32'b00000000000000000111100011010110;
assign LUT_1[61081] = 32'b00000000000000000000110101010010;
assign LUT_1[61082] = 32'b00000000000000000011010001100111;
assign LUT_1[61083] = 32'b11111111111111111100100011100011;
assign LUT_1[61084] = 32'b00000000000000001111011100101101;
assign LUT_1[61085] = 32'b00000000000000001000101110101001;
assign LUT_1[61086] = 32'b00000000000000001011001010111110;
assign LUT_1[61087] = 32'b00000000000000000100011100111010;
assign LUT_1[61088] = 32'b00000000000000000111010100111110;
assign LUT_1[61089] = 32'b00000000000000000000100110111010;
assign LUT_1[61090] = 32'b00000000000000000011000011001111;
assign LUT_1[61091] = 32'b11111111111111111100010101001011;
assign LUT_1[61092] = 32'b00000000000000001111001110010101;
assign LUT_1[61093] = 32'b00000000000000001000100000010001;
assign LUT_1[61094] = 32'b00000000000000001010111100100110;
assign LUT_1[61095] = 32'b00000000000000000100001110100010;
assign LUT_1[61096] = 32'b00000000000000000110100010110011;
assign LUT_1[61097] = 32'b11111111111111111111110100101111;
assign LUT_1[61098] = 32'b00000000000000000010010001000100;
assign LUT_1[61099] = 32'b11111111111111111011100011000000;
assign LUT_1[61100] = 32'b00000000000000001110011100001010;
assign LUT_1[61101] = 32'b00000000000000000111101110000110;
assign LUT_1[61102] = 32'b00000000000000001010001010011011;
assign LUT_1[61103] = 32'b00000000000000000011011100010111;
assign LUT_1[61104] = 32'b00000000000000001001010000100000;
assign LUT_1[61105] = 32'b00000000000000000010100010011100;
assign LUT_1[61106] = 32'b00000000000000000100111110110001;
assign LUT_1[61107] = 32'b11111111111111111110010000101101;
assign LUT_1[61108] = 32'b00000000000000010001001001110111;
assign LUT_1[61109] = 32'b00000000000000001010011011110011;
assign LUT_1[61110] = 32'b00000000000000001100111000001000;
assign LUT_1[61111] = 32'b00000000000000000110001010000100;
assign LUT_1[61112] = 32'b00000000000000001000011110010101;
assign LUT_1[61113] = 32'b00000000000000000001110000010001;
assign LUT_1[61114] = 32'b00000000000000000100001100100110;
assign LUT_1[61115] = 32'b11111111111111111101011110100010;
assign LUT_1[61116] = 32'b00000000000000010000010111101100;
assign LUT_1[61117] = 32'b00000000000000001001101001101000;
assign LUT_1[61118] = 32'b00000000000000001100000101111101;
assign LUT_1[61119] = 32'b00000000000000000101010111111001;
assign LUT_1[61120] = 32'b00000000000000001000010111100111;
assign LUT_1[61121] = 32'b00000000000000000001101001100011;
assign LUT_1[61122] = 32'b00000000000000000100000101111000;
assign LUT_1[61123] = 32'b11111111111111111101010111110100;
assign LUT_1[61124] = 32'b00000000000000010000010000111110;
assign LUT_1[61125] = 32'b00000000000000001001100010111010;
assign LUT_1[61126] = 32'b00000000000000001011111111001111;
assign LUT_1[61127] = 32'b00000000000000000101010001001011;
assign LUT_1[61128] = 32'b00000000000000000111100101011100;
assign LUT_1[61129] = 32'b00000000000000000000110111011000;
assign LUT_1[61130] = 32'b00000000000000000011010011101101;
assign LUT_1[61131] = 32'b11111111111111111100100101101001;
assign LUT_1[61132] = 32'b00000000000000001111011110110011;
assign LUT_1[61133] = 32'b00000000000000001000110000101111;
assign LUT_1[61134] = 32'b00000000000000001011001101000100;
assign LUT_1[61135] = 32'b00000000000000000100011111000000;
assign LUT_1[61136] = 32'b00000000000000001010010011001001;
assign LUT_1[61137] = 32'b00000000000000000011100101000101;
assign LUT_1[61138] = 32'b00000000000000000110000001011010;
assign LUT_1[61139] = 32'b11111111111111111111010011010110;
assign LUT_1[61140] = 32'b00000000000000010010001100100000;
assign LUT_1[61141] = 32'b00000000000000001011011110011100;
assign LUT_1[61142] = 32'b00000000000000001101111010110001;
assign LUT_1[61143] = 32'b00000000000000000111001100101101;
assign LUT_1[61144] = 32'b00000000000000001001100000111110;
assign LUT_1[61145] = 32'b00000000000000000010110010111010;
assign LUT_1[61146] = 32'b00000000000000000101001111001111;
assign LUT_1[61147] = 32'b11111111111111111110100001001011;
assign LUT_1[61148] = 32'b00000000000000010001011010010101;
assign LUT_1[61149] = 32'b00000000000000001010101100010001;
assign LUT_1[61150] = 32'b00000000000000001101001000100110;
assign LUT_1[61151] = 32'b00000000000000000110011010100010;
assign LUT_1[61152] = 32'b00000000000000001001010010100110;
assign LUT_1[61153] = 32'b00000000000000000010100100100010;
assign LUT_1[61154] = 32'b00000000000000000101000000110111;
assign LUT_1[61155] = 32'b11111111111111111110010010110011;
assign LUT_1[61156] = 32'b00000000000000010001001011111101;
assign LUT_1[61157] = 32'b00000000000000001010011101111001;
assign LUT_1[61158] = 32'b00000000000000001100111010001110;
assign LUT_1[61159] = 32'b00000000000000000110001100001010;
assign LUT_1[61160] = 32'b00000000000000001000100000011011;
assign LUT_1[61161] = 32'b00000000000000000001110010010111;
assign LUT_1[61162] = 32'b00000000000000000100001110101100;
assign LUT_1[61163] = 32'b11111111111111111101100000101000;
assign LUT_1[61164] = 32'b00000000000000010000011001110010;
assign LUT_1[61165] = 32'b00000000000000001001101011101110;
assign LUT_1[61166] = 32'b00000000000000001100001000000011;
assign LUT_1[61167] = 32'b00000000000000000101011001111111;
assign LUT_1[61168] = 32'b00000000000000001011001110001000;
assign LUT_1[61169] = 32'b00000000000000000100100000000100;
assign LUT_1[61170] = 32'b00000000000000000110111100011001;
assign LUT_1[61171] = 32'b00000000000000000000001110010101;
assign LUT_1[61172] = 32'b00000000000000010011000111011111;
assign LUT_1[61173] = 32'b00000000000000001100011001011011;
assign LUT_1[61174] = 32'b00000000000000001110110101110000;
assign LUT_1[61175] = 32'b00000000000000001000000111101100;
assign LUT_1[61176] = 32'b00000000000000001010011011111101;
assign LUT_1[61177] = 32'b00000000000000000011101101111001;
assign LUT_1[61178] = 32'b00000000000000000110001010001110;
assign LUT_1[61179] = 32'b11111111111111111111011100001010;
assign LUT_1[61180] = 32'b00000000000000010010010101010100;
assign LUT_1[61181] = 32'b00000000000000001011100111010000;
assign LUT_1[61182] = 32'b00000000000000001110000011100101;
assign LUT_1[61183] = 32'b00000000000000000111010101100001;
assign LUT_1[61184] = 32'b00000000000000000001001110001000;
assign LUT_1[61185] = 32'b11111111111111111010100000000100;
assign LUT_1[61186] = 32'b11111111111111111100111100011001;
assign LUT_1[61187] = 32'b11111111111111110110001110010101;
assign LUT_1[61188] = 32'b00000000000000001001000111011111;
assign LUT_1[61189] = 32'b00000000000000000010011001011011;
assign LUT_1[61190] = 32'b00000000000000000100110101110000;
assign LUT_1[61191] = 32'b11111111111111111110000111101100;
assign LUT_1[61192] = 32'b00000000000000000000011011111101;
assign LUT_1[61193] = 32'b11111111111111111001101101111001;
assign LUT_1[61194] = 32'b11111111111111111100001010001110;
assign LUT_1[61195] = 32'b11111111111111110101011100001010;
assign LUT_1[61196] = 32'b00000000000000001000010101010100;
assign LUT_1[61197] = 32'b00000000000000000001100111010000;
assign LUT_1[61198] = 32'b00000000000000000100000011100101;
assign LUT_1[61199] = 32'b11111111111111111101010101100001;
assign LUT_1[61200] = 32'b00000000000000000011001001101010;
assign LUT_1[61201] = 32'b11111111111111111100011011100110;
assign LUT_1[61202] = 32'b11111111111111111110110111111011;
assign LUT_1[61203] = 32'b11111111111111111000001001110111;
assign LUT_1[61204] = 32'b00000000000000001011000011000001;
assign LUT_1[61205] = 32'b00000000000000000100010100111101;
assign LUT_1[61206] = 32'b00000000000000000110110001010010;
assign LUT_1[61207] = 32'b00000000000000000000000011001110;
assign LUT_1[61208] = 32'b00000000000000000010010111011111;
assign LUT_1[61209] = 32'b11111111111111111011101001011011;
assign LUT_1[61210] = 32'b11111111111111111110000101110000;
assign LUT_1[61211] = 32'b11111111111111110111010111101100;
assign LUT_1[61212] = 32'b00000000000000001010010000110110;
assign LUT_1[61213] = 32'b00000000000000000011100010110010;
assign LUT_1[61214] = 32'b00000000000000000101111111000111;
assign LUT_1[61215] = 32'b11111111111111111111010001000011;
assign LUT_1[61216] = 32'b00000000000000000010001001000111;
assign LUT_1[61217] = 32'b11111111111111111011011011000011;
assign LUT_1[61218] = 32'b11111111111111111101110111011000;
assign LUT_1[61219] = 32'b11111111111111110111001001010100;
assign LUT_1[61220] = 32'b00000000000000001010000010011110;
assign LUT_1[61221] = 32'b00000000000000000011010100011010;
assign LUT_1[61222] = 32'b00000000000000000101110000101111;
assign LUT_1[61223] = 32'b11111111111111111111000010101011;
assign LUT_1[61224] = 32'b00000000000000000001010110111100;
assign LUT_1[61225] = 32'b11111111111111111010101000111000;
assign LUT_1[61226] = 32'b11111111111111111101000101001101;
assign LUT_1[61227] = 32'b11111111111111110110010111001001;
assign LUT_1[61228] = 32'b00000000000000001001010000010011;
assign LUT_1[61229] = 32'b00000000000000000010100010001111;
assign LUT_1[61230] = 32'b00000000000000000100111110100100;
assign LUT_1[61231] = 32'b11111111111111111110010000100000;
assign LUT_1[61232] = 32'b00000000000000000100000100101001;
assign LUT_1[61233] = 32'b11111111111111111101010110100101;
assign LUT_1[61234] = 32'b11111111111111111111110010111010;
assign LUT_1[61235] = 32'b11111111111111111001000100110110;
assign LUT_1[61236] = 32'b00000000000000001011111110000000;
assign LUT_1[61237] = 32'b00000000000000000101001111111100;
assign LUT_1[61238] = 32'b00000000000000000111101100010001;
assign LUT_1[61239] = 32'b00000000000000000000111110001101;
assign LUT_1[61240] = 32'b00000000000000000011010010011110;
assign LUT_1[61241] = 32'b11111111111111111100100100011010;
assign LUT_1[61242] = 32'b11111111111111111111000000101111;
assign LUT_1[61243] = 32'b11111111111111111000010010101011;
assign LUT_1[61244] = 32'b00000000000000001011001011110101;
assign LUT_1[61245] = 32'b00000000000000000100011101110001;
assign LUT_1[61246] = 32'b00000000000000000110111010000110;
assign LUT_1[61247] = 32'b00000000000000000000001100000010;
assign LUT_1[61248] = 32'b00000000000000000011001011110000;
assign LUT_1[61249] = 32'b11111111111111111100011101101100;
assign LUT_1[61250] = 32'b11111111111111111110111010000001;
assign LUT_1[61251] = 32'b11111111111111111000001011111101;
assign LUT_1[61252] = 32'b00000000000000001011000101000111;
assign LUT_1[61253] = 32'b00000000000000000100010111000011;
assign LUT_1[61254] = 32'b00000000000000000110110011011000;
assign LUT_1[61255] = 32'b00000000000000000000000101010100;
assign LUT_1[61256] = 32'b00000000000000000010011001100101;
assign LUT_1[61257] = 32'b11111111111111111011101011100001;
assign LUT_1[61258] = 32'b11111111111111111110000111110110;
assign LUT_1[61259] = 32'b11111111111111110111011001110010;
assign LUT_1[61260] = 32'b00000000000000001010010010111100;
assign LUT_1[61261] = 32'b00000000000000000011100100111000;
assign LUT_1[61262] = 32'b00000000000000000110000001001101;
assign LUT_1[61263] = 32'b11111111111111111111010011001001;
assign LUT_1[61264] = 32'b00000000000000000101000111010010;
assign LUT_1[61265] = 32'b11111111111111111110011001001110;
assign LUT_1[61266] = 32'b00000000000000000000110101100011;
assign LUT_1[61267] = 32'b11111111111111111010000111011111;
assign LUT_1[61268] = 32'b00000000000000001101000000101001;
assign LUT_1[61269] = 32'b00000000000000000110010010100101;
assign LUT_1[61270] = 32'b00000000000000001000101110111010;
assign LUT_1[61271] = 32'b00000000000000000010000000110110;
assign LUT_1[61272] = 32'b00000000000000000100010101000111;
assign LUT_1[61273] = 32'b11111111111111111101100111000011;
assign LUT_1[61274] = 32'b00000000000000000000000011011000;
assign LUT_1[61275] = 32'b11111111111111111001010101010100;
assign LUT_1[61276] = 32'b00000000000000001100001110011110;
assign LUT_1[61277] = 32'b00000000000000000101100000011010;
assign LUT_1[61278] = 32'b00000000000000000111111100101111;
assign LUT_1[61279] = 32'b00000000000000000001001110101011;
assign LUT_1[61280] = 32'b00000000000000000100000110101111;
assign LUT_1[61281] = 32'b11111111111111111101011000101011;
assign LUT_1[61282] = 32'b11111111111111111111110101000000;
assign LUT_1[61283] = 32'b11111111111111111001000110111100;
assign LUT_1[61284] = 32'b00000000000000001100000000000110;
assign LUT_1[61285] = 32'b00000000000000000101010010000010;
assign LUT_1[61286] = 32'b00000000000000000111101110010111;
assign LUT_1[61287] = 32'b00000000000000000001000000010011;
assign LUT_1[61288] = 32'b00000000000000000011010100100100;
assign LUT_1[61289] = 32'b11111111111111111100100110100000;
assign LUT_1[61290] = 32'b11111111111111111111000010110101;
assign LUT_1[61291] = 32'b11111111111111111000010100110001;
assign LUT_1[61292] = 32'b00000000000000001011001101111011;
assign LUT_1[61293] = 32'b00000000000000000100011111110111;
assign LUT_1[61294] = 32'b00000000000000000110111100001100;
assign LUT_1[61295] = 32'b00000000000000000000001110001000;
assign LUT_1[61296] = 32'b00000000000000000110000010010001;
assign LUT_1[61297] = 32'b11111111111111111111010100001101;
assign LUT_1[61298] = 32'b00000000000000000001110000100010;
assign LUT_1[61299] = 32'b11111111111111111011000010011110;
assign LUT_1[61300] = 32'b00000000000000001101111011101000;
assign LUT_1[61301] = 32'b00000000000000000111001101100100;
assign LUT_1[61302] = 32'b00000000000000001001101001111001;
assign LUT_1[61303] = 32'b00000000000000000010111011110101;
assign LUT_1[61304] = 32'b00000000000000000101010000000110;
assign LUT_1[61305] = 32'b11111111111111111110100010000010;
assign LUT_1[61306] = 32'b00000000000000000000111110010111;
assign LUT_1[61307] = 32'b11111111111111111010010000010011;
assign LUT_1[61308] = 32'b00000000000000001101001001011101;
assign LUT_1[61309] = 32'b00000000000000000110011011011001;
assign LUT_1[61310] = 32'b00000000000000001000110111101110;
assign LUT_1[61311] = 32'b00000000000000000010001001101010;
assign LUT_1[61312] = 32'b00000000000000000100001110001011;
assign LUT_1[61313] = 32'b11111111111111111101100000000111;
assign LUT_1[61314] = 32'b11111111111111111111111100011100;
assign LUT_1[61315] = 32'b11111111111111111001001110011000;
assign LUT_1[61316] = 32'b00000000000000001100000111100010;
assign LUT_1[61317] = 32'b00000000000000000101011001011110;
assign LUT_1[61318] = 32'b00000000000000000111110101110011;
assign LUT_1[61319] = 32'b00000000000000000001000111101111;
assign LUT_1[61320] = 32'b00000000000000000011011100000000;
assign LUT_1[61321] = 32'b11111111111111111100101101111100;
assign LUT_1[61322] = 32'b11111111111111111111001010010001;
assign LUT_1[61323] = 32'b11111111111111111000011100001101;
assign LUT_1[61324] = 32'b00000000000000001011010101010111;
assign LUT_1[61325] = 32'b00000000000000000100100111010011;
assign LUT_1[61326] = 32'b00000000000000000111000011101000;
assign LUT_1[61327] = 32'b00000000000000000000010101100100;
assign LUT_1[61328] = 32'b00000000000000000110001001101101;
assign LUT_1[61329] = 32'b11111111111111111111011011101001;
assign LUT_1[61330] = 32'b00000000000000000001110111111110;
assign LUT_1[61331] = 32'b11111111111111111011001001111010;
assign LUT_1[61332] = 32'b00000000000000001110000011000100;
assign LUT_1[61333] = 32'b00000000000000000111010101000000;
assign LUT_1[61334] = 32'b00000000000000001001110001010101;
assign LUT_1[61335] = 32'b00000000000000000011000011010001;
assign LUT_1[61336] = 32'b00000000000000000101010111100010;
assign LUT_1[61337] = 32'b11111111111111111110101001011110;
assign LUT_1[61338] = 32'b00000000000000000001000101110011;
assign LUT_1[61339] = 32'b11111111111111111010010111101111;
assign LUT_1[61340] = 32'b00000000000000001101010000111001;
assign LUT_1[61341] = 32'b00000000000000000110100010110101;
assign LUT_1[61342] = 32'b00000000000000001000111111001010;
assign LUT_1[61343] = 32'b00000000000000000010010001000110;
assign LUT_1[61344] = 32'b00000000000000000101001001001010;
assign LUT_1[61345] = 32'b11111111111111111110011011000110;
assign LUT_1[61346] = 32'b00000000000000000000110111011011;
assign LUT_1[61347] = 32'b11111111111111111010001001010111;
assign LUT_1[61348] = 32'b00000000000000001101000010100001;
assign LUT_1[61349] = 32'b00000000000000000110010100011101;
assign LUT_1[61350] = 32'b00000000000000001000110000110010;
assign LUT_1[61351] = 32'b00000000000000000010000010101110;
assign LUT_1[61352] = 32'b00000000000000000100010110111111;
assign LUT_1[61353] = 32'b11111111111111111101101000111011;
assign LUT_1[61354] = 32'b00000000000000000000000101010000;
assign LUT_1[61355] = 32'b11111111111111111001010111001100;
assign LUT_1[61356] = 32'b00000000000000001100010000010110;
assign LUT_1[61357] = 32'b00000000000000000101100010010010;
assign LUT_1[61358] = 32'b00000000000000000111111110100111;
assign LUT_1[61359] = 32'b00000000000000000001010000100011;
assign LUT_1[61360] = 32'b00000000000000000111000100101100;
assign LUT_1[61361] = 32'b00000000000000000000010110101000;
assign LUT_1[61362] = 32'b00000000000000000010110010111101;
assign LUT_1[61363] = 32'b11111111111111111100000100111001;
assign LUT_1[61364] = 32'b00000000000000001110111110000011;
assign LUT_1[61365] = 32'b00000000000000001000001111111111;
assign LUT_1[61366] = 32'b00000000000000001010101100010100;
assign LUT_1[61367] = 32'b00000000000000000011111110010000;
assign LUT_1[61368] = 32'b00000000000000000110010010100001;
assign LUT_1[61369] = 32'b11111111111111111111100100011101;
assign LUT_1[61370] = 32'b00000000000000000010000000110010;
assign LUT_1[61371] = 32'b11111111111111111011010010101110;
assign LUT_1[61372] = 32'b00000000000000001110001011111000;
assign LUT_1[61373] = 32'b00000000000000000111011101110100;
assign LUT_1[61374] = 32'b00000000000000001001111010001001;
assign LUT_1[61375] = 32'b00000000000000000011001100000101;
assign LUT_1[61376] = 32'b00000000000000000110001011110011;
assign LUT_1[61377] = 32'b11111111111111111111011101101111;
assign LUT_1[61378] = 32'b00000000000000000001111010000100;
assign LUT_1[61379] = 32'b11111111111111111011001100000000;
assign LUT_1[61380] = 32'b00000000000000001110000101001010;
assign LUT_1[61381] = 32'b00000000000000000111010111000110;
assign LUT_1[61382] = 32'b00000000000000001001110011011011;
assign LUT_1[61383] = 32'b00000000000000000011000101010111;
assign LUT_1[61384] = 32'b00000000000000000101011001101000;
assign LUT_1[61385] = 32'b11111111111111111110101011100100;
assign LUT_1[61386] = 32'b00000000000000000001000111111001;
assign LUT_1[61387] = 32'b11111111111111111010011001110101;
assign LUT_1[61388] = 32'b00000000000000001101010010111111;
assign LUT_1[61389] = 32'b00000000000000000110100100111011;
assign LUT_1[61390] = 32'b00000000000000001001000001010000;
assign LUT_1[61391] = 32'b00000000000000000010010011001100;
assign LUT_1[61392] = 32'b00000000000000001000000111010101;
assign LUT_1[61393] = 32'b00000000000000000001011001010001;
assign LUT_1[61394] = 32'b00000000000000000011110101100110;
assign LUT_1[61395] = 32'b11111111111111111101000111100010;
assign LUT_1[61396] = 32'b00000000000000010000000000101100;
assign LUT_1[61397] = 32'b00000000000000001001010010101000;
assign LUT_1[61398] = 32'b00000000000000001011101110111101;
assign LUT_1[61399] = 32'b00000000000000000101000000111001;
assign LUT_1[61400] = 32'b00000000000000000111010101001010;
assign LUT_1[61401] = 32'b00000000000000000000100111000110;
assign LUT_1[61402] = 32'b00000000000000000011000011011011;
assign LUT_1[61403] = 32'b11111111111111111100010101010111;
assign LUT_1[61404] = 32'b00000000000000001111001110100001;
assign LUT_1[61405] = 32'b00000000000000001000100000011101;
assign LUT_1[61406] = 32'b00000000000000001010111100110010;
assign LUT_1[61407] = 32'b00000000000000000100001110101110;
assign LUT_1[61408] = 32'b00000000000000000111000110110010;
assign LUT_1[61409] = 32'b00000000000000000000011000101110;
assign LUT_1[61410] = 32'b00000000000000000010110101000011;
assign LUT_1[61411] = 32'b11111111111111111100000110111111;
assign LUT_1[61412] = 32'b00000000000000001111000000001001;
assign LUT_1[61413] = 32'b00000000000000001000010010000101;
assign LUT_1[61414] = 32'b00000000000000001010101110011010;
assign LUT_1[61415] = 32'b00000000000000000100000000010110;
assign LUT_1[61416] = 32'b00000000000000000110010100100111;
assign LUT_1[61417] = 32'b11111111111111111111100110100011;
assign LUT_1[61418] = 32'b00000000000000000010000010111000;
assign LUT_1[61419] = 32'b11111111111111111011010100110100;
assign LUT_1[61420] = 32'b00000000000000001110001101111110;
assign LUT_1[61421] = 32'b00000000000000000111011111111010;
assign LUT_1[61422] = 32'b00000000000000001001111100001111;
assign LUT_1[61423] = 32'b00000000000000000011001110001011;
assign LUT_1[61424] = 32'b00000000000000001001000010010100;
assign LUT_1[61425] = 32'b00000000000000000010010100010000;
assign LUT_1[61426] = 32'b00000000000000000100110000100101;
assign LUT_1[61427] = 32'b11111111111111111110000010100001;
assign LUT_1[61428] = 32'b00000000000000010000111011101011;
assign LUT_1[61429] = 32'b00000000000000001010001101100111;
assign LUT_1[61430] = 32'b00000000000000001100101001111100;
assign LUT_1[61431] = 32'b00000000000000000101111011111000;
assign LUT_1[61432] = 32'b00000000000000001000010000001001;
assign LUT_1[61433] = 32'b00000000000000000001100010000101;
assign LUT_1[61434] = 32'b00000000000000000011111110011010;
assign LUT_1[61435] = 32'b11111111111111111101010000010110;
assign LUT_1[61436] = 32'b00000000000000010000001001100000;
assign LUT_1[61437] = 32'b00000000000000001001011011011100;
assign LUT_1[61438] = 32'b00000000000000001011110111110001;
assign LUT_1[61439] = 32'b00000000000000000101001001101101;
assign LUT_1[61440] = 32'b00000000000000000010000111111010;
assign LUT_1[61441] = 32'b11111111111111111011011001110110;
assign LUT_1[61442] = 32'b11111111111111111101110110001011;
assign LUT_1[61443] = 32'b11111111111111110111001000000111;
assign LUT_1[61444] = 32'b00000000000000001010000001010001;
assign LUT_1[61445] = 32'b00000000000000000011010011001101;
assign LUT_1[61446] = 32'b00000000000000000101101111100010;
assign LUT_1[61447] = 32'b11111111111111111111000001011110;
assign LUT_1[61448] = 32'b00000000000000000001010101101111;
assign LUT_1[61449] = 32'b11111111111111111010100111101011;
assign LUT_1[61450] = 32'b11111111111111111101000100000000;
assign LUT_1[61451] = 32'b11111111111111110110010101111100;
assign LUT_1[61452] = 32'b00000000000000001001001111000110;
assign LUT_1[61453] = 32'b00000000000000000010100001000010;
assign LUT_1[61454] = 32'b00000000000000000100111101010111;
assign LUT_1[61455] = 32'b11111111111111111110001111010011;
assign LUT_1[61456] = 32'b00000000000000000100000011011100;
assign LUT_1[61457] = 32'b11111111111111111101010101011000;
assign LUT_1[61458] = 32'b11111111111111111111110001101101;
assign LUT_1[61459] = 32'b11111111111111111001000011101001;
assign LUT_1[61460] = 32'b00000000000000001011111100110011;
assign LUT_1[61461] = 32'b00000000000000000101001110101111;
assign LUT_1[61462] = 32'b00000000000000000111101011000100;
assign LUT_1[61463] = 32'b00000000000000000000111101000000;
assign LUT_1[61464] = 32'b00000000000000000011010001010001;
assign LUT_1[61465] = 32'b11111111111111111100100011001101;
assign LUT_1[61466] = 32'b11111111111111111110111111100010;
assign LUT_1[61467] = 32'b11111111111111111000010001011110;
assign LUT_1[61468] = 32'b00000000000000001011001010101000;
assign LUT_1[61469] = 32'b00000000000000000100011100100100;
assign LUT_1[61470] = 32'b00000000000000000110111000111001;
assign LUT_1[61471] = 32'b00000000000000000000001010110101;
assign LUT_1[61472] = 32'b00000000000000000011000010111001;
assign LUT_1[61473] = 32'b11111111111111111100010100110101;
assign LUT_1[61474] = 32'b11111111111111111110110001001010;
assign LUT_1[61475] = 32'b11111111111111111000000011000110;
assign LUT_1[61476] = 32'b00000000000000001010111100010000;
assign LUT_1[61477] = 32'b00000000000000000100001110001100;
assign LUT_1[61478] = 32'b00000000000000000110101010100001;
assign LUT_1[61479] = 32'b11111111111111111111111100011101;
assign LUT_1[61480] = 32'b00000000000000000010010000101110;
assign LUT_1[61481] = 32'b11111111111111111011100010101010;
assign LUT_1[61482] = 32'b11111111111111111101111110111111;
assign LUT_1[61483] = 32'b11111111111111110111010000111011;
assign LUT_1[61484] = 32'b00000000000000001010001010000101;
assign LUT_1[61485] = 32'b00000000000000000011011100000001;
assign LUT_1[61486] = 32'b00000000000000000101111000010110;
assign LUT_1[61487] = 32'b11111111111111111111001010010010;
assign LUT_1[61488] = 32'b00000000000000000100111110011011;
assign LUT_1[61489] = 32'b11111111111111111110010000010111;
assign LUT_1[61490] = 32'b00000000000000000000101100101100;
assign LUT_1[61491] = 32'b11111111111111111001111110101000;
assign LUT_1[61492] = 32'b00000000000000001100110111110010;
assign LUT_1[61493] = 32'b00000000000000000110001001101110;
assign LUT_1[61494] = 32'b00000000000000001000100110000011;
assign LUT_1[61495] = 32'b00000000000000000001110111111111;
assign LUT_1[61496] = 32'b00000000000000000100001100010000;
assign LUT_1[61497] = 32'b11111111111111111101011110001100;
assign LUT_1[61498] = 32'b11111111111111111111111010100001;
assign LUT_1[61499] = 32'b11111111111111111001001100011101;
assign LUT_1[61500] = 32'b00000000000000001100000101100111;
assign LUT_1[61501] = 32'b00000000000000000101010111100011;
assign LUT_1[61502] = 32'b00000000000000000111110011111000;
assign LUT_1[61503] = 32'b00000000000000000001000101110100;
assign LUT_1[61504] = 32'b00000000000000000100000101100010;
assign LUT_1[61505] = 32'b11111111111111111101010111011110;
assign LUT_1[61506] = 32'b11111111111111111111110011110011;
assign LUT_1[61507] = 32'b11111111111111111001000101101111;
assign LUT_1[61508] = 32'b00000000000000001011111110111001;
assign LUT_1[61509] = 32'b00000000000000000101010000110101;
assign LUT_1[61510] = 32'b00000000000000000111101101001010;
assign LUT_1[61511] = 32'b00000000000000000000111111000110;
assign LUT_1[61512] = 32'b00000000000000000011010011010111;
assign LUT_1[61513] = 32'b11111111111111111100100101010011;
assign LUT_1[61514] = 32'b11111111111111111111000001101000;
assign LUT_1[61515] = 32'b11111111111111111000010011100100;
assign LUT_1[61516] = 32'b00000000000000001011001100101110;
assign LUT_1[61517] = 32'b00000000000000000100011110101010;
assign LUT_1[61518] = 32'b00000000000000000110111010111111;
assign LUT_1[61519] = 32'b00000000000000000000001100111011;
assign LUT_1[61520] = 32'b00000000000000000110000001000100;
assign LUT_1[61521] = 32'b11111111111111111111010011000000;
assign LUT_1[61522] = 32'b00000000000000000001101111010101;
assign LUT_1[61523] = 32'b11111111111111111011000001010001;
assign LUT_1[61524] = 32'b00000000000000001101111010011011;
assign LUT_1[61525] = 32'b00000000000000000111001100010111;
assign LUT_1[61526] = 32'b00000000000000001001101000101100;
assign LUT_1[61527] = 32'b00000000000000000010111010101000;
assign LUT_1[61528] = 32'b00000000000000000101001110111001;
assign LUT_1[61529] = 32'b11111111111111111110100000110101;
assign LUT_1[61530] = 32'b00000000000000000000111101001010;
assign LUT_1[61531] = 32'b11111111111111111010001111000110;
assign LUT_1[61532] = 32'b00000000000000001101001000010000;
assign LUT_1[61533] = 32'b00000000000000000110011010001100;
assign LUT_1[61534] = 32'b00000000000000001000110110100001;
assign LUT_1[61535] = 32'b00000000000000000010001000011101;
assign LUT_1[61536] = 32'b00000000000000000101000000100001;
assign LUT_1[61537] = 32'b11111111111111111110010010011101;
assign LUT_1[61538] = 32'b00000000000000000000101110110010;
assign LUT_1[61539] = 32'b11111111111111111010000000101110;
assign LUT_1[61540] = 32'b00000000000000001100111001111000;
assign LUT_1[61541] = 32'b00000000000000000110001011110100;
assign LUT_1[61542] = 32'b00000000000000001000101000001001;
assign LUT_1[61543] = 32'b00000000000000000001111010000101;
assign LUT_1[61544] = 32'b00000000000000000100001110010110;
assign LUT_1[61545] = 32'b11111111111111111101100000010010;
assign LUT_1[61546] = 32'b11111111111111111111111100100111;
assign LUT_1[61547] = 32'b11111111111111111001001110100011;
assign LUT_1[61548] = 32'b00000000000000001100000111101101;
assign LUT_1[61549] = 32'b00000000000000000101011001101001;
assign LUT_1[61550] = 32'b00000000000000000111110101111110;
assign LUT_1[61551] = 32'b00000000000000000001000111111010;
assign LUT_1[61552] = 32'b00000000000000000110111100000011;
assign LUT_1[61553] = 32'b00000000000000000000001101111111;
assign LUT_1[61554] = 32'b00000000000000000010101010010100;
assign LUT_1[61555] = 32'b11111111111111111011111100010000;
assign LUT_1[61556] = 32'b00000000000000001110110101011010;
assign LUT_1[61557] = 32'b00000000000000001000000111010110;
assign LUT_1[61558] = 32'b00000000000000001010100011101011;
assign LUT_1[61559] = 32'b00000000000000000011110101100111;
assign LUT_1[61560] = 32'b00000000000000000110001001111000;
assign LUT_1[61561] = 32'b11111111111111111111011011110100;
assign LUT_1[61562] = 32'b00000000000000000001111000001001;
assign LUT_1[61563] = 32'b11111111111111111011001010000101;
assign LUT_1[61564] = 32'b00000000000000001110000011001111;
assign LUT_1[61565] = 32'b00000000000000000111010101001011;
assign LUT_1[61566] = 32'b00000000000000001001110001100000;
assign LUT_1[61567] = 32'b00000000000000000011000011011100;
assign LUT_1[61568] = 32'b00000000000000000101000111111101;
assign LUT_1[61569] = 32'b11111111111111111110011001111001;
assign LUT_1[61570] = 32'b00000000000000000000110110001110;
assign LUT_1[61571] = 32'b11111111111111111010001000001010;
assign LUT_1[61572] = 32'b00000000000000001101000001010100;
assign LUT_1[61573] = 32'b00000000000000000110010011010000;
assign LUT_1[61574] = 32'b00000000000000001000101111100101;
assign LUT_1[61575] = 32'b00000000000000000010000001100001;
assign LUT_1[61576] = 32'b00000000000000000100010101110010;
assign LUT_1[61577] = 32'b11111111111111111101100111101110;
assign LUT_1[61578] = 32'b00000000000000000000000100000011;
assign LUT_1[61579] = 32'b11111111111111111001010101111111;
assign LUT_1[61580] = 32'b00000000000000001100001111001001;
assign LUT_1[61581] = 32'b00000000000000000101100001000101;
assign LUT_1[61582] = 32'b00000000000000000111111101011010;
assign LUT_1[61583] = 32'b00000000000000000001001111010110;
assign LUT_1[61584] = 32'b00000000000000000111000011011111;
assign LUT_1[61585] = 32'b00000000000000000000010101011011;
assign LUT_1[61586] = 32'b00000000000000000010110001110000;
assign LUT_1[61587] = 32'b11111111111111111100000011101100;
assign LUT_1[61588] = 32'b00000000000000001110111100110110;
assign LUT_1[61589] = 32'b00000000000000001000001110110010;
assign LUT_1[61590] = 32'b00000000000000001010101011000111;
assign LUT_1[61591] = 32'b00000000000000000011111101000011;
assign LUT_1[61592] = 32'b00000000000000000110010001010100;
assign LUT_1[61593] = 32'b11111111111111111111100011010000;
assign LUT_1[61594] = 32'b00000000000000000001111111100101;
assign LUT_1[61595] = 32'b11111111111111111011010001100001;
assign LUT_1[61596] = 32'b00000000000000001110001010101011;
assign LUT_1[61597] = 32'b00000000000000000111011100100111;
assign LUT_1[61598] = 32'b00000000000000001001111000111100;
assign LUT_1[61599] = 32'b00000000000000000011001010111000;
assign LUT_1[61600] = 32'b00000000000000000110000010111100;
assign LUT_1[61601] = 32'b11111111111111111111010100111000;
assign LUT_1[61602] = 32'b00000000000000000001110001001101;
assign LUT_1[61603] = 32'b11111111111111111011000011001001;
assign LUT_1[61604] = 32'b00000000000000001101111100010011;
assign LUT_1[61605] = 32'b00000000000000000111001110001111;
assign LUT_1[61606] = 32'b00000000000000001001101010100100;
assign LUT_1[61607] = 32'b00000000000000000010111100100000;
assign LUT_1[61608] = 32'b00000000000000000101010000110001;
assign LUT_1[61609] = 32'b11111111111111111110100010101101;
assign LUT_1[61610] = 32'b00000000000000000000111111000010;
assign LUT_1[61611] = 32'b11111111111111111010010000111110;
assign LUT_1[61612] = 32'b00000000000000001101001010001000;
assign LUT_1[61613] = 32'b00000000000000000110011100000100;
assign LUT_1[61614] = 32'b00000000000000001000111000011001;
assign LUT_1[61615] = 32'b00000000000000000010001010010101;
assign LUT_1[61616] = 32'b00000000000000000111111110011110;
assign LUT_1[61617] = 32'b00000000000000000001010000011010;
assign LUT_1[61618] = 32'b00000000000000000011101100101111;
assign LUT_1[61619] = 32'b11111111111111111100111110101011;
assign LUT_1[61620] = 32'b00000000000000001111110111110101;
assign LUT_1[61621] = 32'b00000000000000001001001001110001;
assign LUT_1[61622] = 32'b00000000000000001011100110000110;
assign LUT_1[61623] = 32'b00000000000000000100111000000010;
assign LUT_1[61624] = 32'b00000000000000000111001100010011;
assign LUT_1[61625] = 32'b00000000000000000000011110001111;
assign LUT_1[61626] = 32'b00000000000000000010111010100100;
assign LUT_1[61627] = 32'b11111111111111111100001100100000;
assign LUT_1[61628] = 32'b00000000000000001111000101101010;
assign LUT_1[61629] = 32'b00000000000000001000010111100110;
assign LUT_1[61630] = 32'b00000000000000001010110011111011;
assign LUT_1[61631] = 32'b00000000000000000100000101110111;
assign LUT_1[61632] = 32'b00000000000000000111000101100101;
assign LUT_1[61633] = 32'b00000000000000000000010111100001;
assign LUT_1[61634] = 32'b00000000000000000010110011110110;
assign LUT_1[61635] = 32'b11111111111111111100000101110010;
assign LUT_1[61636] = 32'b00000000000000001110111110111100;
assign LUT_1[61637] = 32'b00000000000000001000010000111000;
assign LUT_1[61638] = 32'b00000000000000001010101101001101;
assign LUT_1[61639] = 32'b00000000000000000011111111001001;
assign LUT_1[61640] = 32'b00000000000000000110010011011010;
assign LUT_1[61641] = 32'b11111111111111111111100101010110;
assign LUT_1[61642] = 32'b00000000000000000010000001101011;
assign LUT_1[61643] = 32'b11111111111111111011010011100111;
assign LUT_1[61644] = 32'b00000000000000001110001100110001;
assign LUT_1[61645] = 32'b00000000000000000111011110101101;
assign LUT_1[61646] = 32'b00000000000000001001111011000010;
assign LUT_1[61647] = 32'b00000000000000000011001100111110;
assign LUT_1[61648] = 32'b00000000000000001001000001000111;
assign LUT_1[61649] = 32'b00000000000000000010010011000011;
assign LUT_1[61650] = 32'b00000000000000000100101111011000;
assign LUT_1[61651] = 32'b11111111111111111110000001010100;
assign LUT_1[61652] = 32'b00000000000000010000111010011110;
assign LUT_1[61653] = 32'b00000000000000001010001100011010;
assign LUT_1[61654] = 32'b00000000000000001100101000101111;
assign LUT_1[61655] = 32'b00000000000000000101111010101011;
assign LUT_1[61656] = 32'b00000000000000001000001110111100;
assign LUT_1[61657] = 32'b00000000000000000001100000111000;
assign LUT_1[61658] = 32'b00000000000000000011111101001101;
assign LUT_1[61659] = 32'b11111111111111111101001111001001;
assign LUT_1[61660] = 32'b00000000000000010000001000010011;
assign LUT_1[61661] = 32'b00000000000000001001011010001111;
assign LUT_1[61662] = 32'b00000000000000001011110110100100;
assign LUT_1[61663] = 32'b00000000000000000101001000100000;
assign LUT_1[61664] = 32'b00000000000000001000000000100100;
assign LUT_1[61665] = 32'b00000000000000000001010010100000;
assign LUT_1[61666] = 32'b00000000000000000011101110110101;
assign LUT_1[61667] = 32'b11111111111111111101000000110001;
assign LUT_1[61668] = 32'b00000000000000001111111001111011;
assign LUT_1[61669] = 32'b00000000000000001001001011110111;
assign LUT_1[61670] = 32'b00000000000000001011101000001100;
assign LUT_1[61671] = 32'b00000000000000000100111010001000;
assign LUT_1[61672] = 32'b00000000000000000111001110011001;
assign LUT_1[61673] = 32'b00000000000000000000100000010101;
assign LUT_1[61674] = 32'b00000000000000000010111100101010;
assign LUT_1[61675] = 32'b11111111111111111100001110100110;
assign LUT_1[61676] = 32'b00000000000000001111000111110000;
assign LUT_1[61677] = 32'b00000000000000001000011001101100;
assign LUT_1[61678] = 32'b00000000000000001010110110000001;
assign LUT_1[61679] = 32'b00000000000000000100000111111101;
assign LUT_1[61680] = 32'b00000000000000001001111100000110;
assign LUT_1[61681] = 32'b00000000000000000011001110000010;
assign LUT_1[61682] = 32'b00000000000000000101101010010111;
assign LUT_1[61683] = 32'b11111111111111111110111100010011;
assign LUT_1[61684] = 32'b00000000000000010001110101011101;
assign LUT_1[61685] = 32'b00000000000000001011000111011001;
assign LUT_1[61686] = 32'b00000000000000001101100011101110;
assign LUT_1[61687] = 32'b00000000000000000110110101101010;
assign LUT_1[61688] = 32'b00000000000000001001001001111011;
assign LUT_1[61689] = 32'b00000000000000000010011011110111;
assign LUT_1[61690] = 32'b00000000000000000100111000001100;
assign LUT_1[61691] = 32'b11111111111111111110001010001000;
assign LUT_1[61692] = 32'b00000000000000010001000011010010;
assign LUT_1[61693] = 32'b00000000000000001010010101001110;
assign LUT_1[61694] = 32'b00000000000000001100110001100011;
assign LUT_1[61695] = 32'b00000000000000000110000011011111;
assign LUT_1[61696] = 32'b11111111111111111111111100000110;
assign LUT_1[61697] = 32'b11111111111111111001001110000010;
assign LUT_1[61698] = 32'b11111111111111111011101010010111;
assign LUT_1[61699] = 32'b11111111111111110100111100010011;
assign LUT_1[61700] = 32'b00000000000000000111110101011101;
assign LUT_1[61701] = 32'b00000000000000000001000111011001;
assign LUT_1[61702] = 32'b00000000000000000011100011101110;
assign LUT_1[61703] = 32'b11111111111111111100110101101010;
assign LUT_1[61704] = 32'b11111111111111111111001001111011;
assign LUT_1[61705] = 32'b11111111111111111000011011110111;
assign LUT_1[61706] = 32'b11111111111111111010111000001100;
assign LUT_1[61707] = 32'b11111111111111110100001010001000;
assign LUT_1[61708] = 32'b00000000000000000111000011010010;
assign LUT_1[61709] = 32'b00000000000000000000010101001110;
assign LUT_1[61710] = 32'b00000000000000000010110001100011;
assign LUT_1[61711] = 32'b11111111111111111100000011011111;
assign LUT_1[61712] = 32'b00000000000000000001110111101000;
assign LUT_1[61713] = 32'b11111111111111111011001001100100;
assign LUT_1[61714] = 32'b11111111111111111101100101111001;
assign LUT_1[61715] = 32'b11111111111111110110110111110101;
assign LUT_1[61716] = 32'b00000000000000001001110000111111;
assign LUT_1[61717] = 32'b00000000000000000011000010111011;
assign LUT_1[61718] = 32'b00000000000000000101011111010000;
assign LUT_1[61719] = 32'b11111111111111111110110001001100;
assign LUT_1[61720] = 32'b00000000000000000001000101011101;
assign LUT_1[61721] = 32'b11111111111111111010010111011001;
assign LUT_1[61722] = 32'b11111111111111111100110011101110;
assign LUT_1[61723] = 32'b11111111111111110110000101101010;
assign LUT_1[61724] = 32'b00000000000000001000111110110100;
assign LUT_1[61725] = 32'b00000000000000000010010000110000;
assign LUT_1[61726] = 32'b00000000000000000100101101000101;
assign LUT_1[61727] = 32'b11111111111111111101111111000001;
assign LUT_1[61728] = 32'b00000000000000000000110111000101;
assign LUT_1[61729] = 32'b11111111111111111010001001000001;
assign LUT_1[61730] = 32'b11111111111111111100100101010110;
assign LUT_1[61731] = 32'b11111111111111110101110111010010;
assign LUT_1[61732] = 32'b00000000000000001000110000011100;
assign LUT_1[61733] = 32'b00000000000000000010000010011000;
assign LUT_1[61734] = 32'b00000000000000000100011110101101;
assign LUT_1[61735] = 32'b11111111111111111101110000101001;
assign LUT_1[61736] = 32'b00000000000000000000000100111010;
assign LUT_1[61737] = 32'b11111111111111111001010110110110;
assign LUT_1[61738] = 32'b11111111111111111011110011001011;
assign LUT_1[61739] = 32'b11111111111111110101000101000111;
assign LUT_1[61740] = 32'b00000000000000000111111110010001;
assign LUT_1[61741] = 32'b00000000000000000001010000001101;
assign LUT_1[61742] = 32'b00000000000000000011101100100010;
assign LUT_1[61743] = 32'b11111111111111111100111110011110;
assign LUT_1[61744] = 32'b00000000000000000010110010100111;
assign LUT_1[61745] = 32'b11111111111111111100000100100011;
assign LUT_1[61746] = 32'b11111111111111111110100000111000;
assign LUT_1[61747] = 32'b11111111111111110111110010110100;
assign LUT_1[61748] = 32'b00000000000000001010101011111110;
assign LUT_1[61749] = 32'b00000000000000000011111101111010;
assign LUT_1[61750] = 32'b00000000000000000110011010001111;
assign LUT_1[61751] = 32'b11111111111111111111101100001011;
assign LUT_1[61752] = 32'b00000000000000000010000000011100;
assign LUT_1[61753] = 32'b11111111111111111011010010011000;
assign LUT_1[61754] = 32'b11111111111111111101101110101101;
assign LUT_1[61755] = 32'b11111111111111110111000000101001;
assign LUT_1[61756] = 32'b00000000000000001001111001110011;
assign LUT_1[61757] = 32'b00000000000000000011001011101111;
assign LUT_1[61758] = 32'b00000000000000000101101000000100;
assign LUT_1[61759] = 32'b11111111111111111110111010000000;
assign LUT_1[61760] = 32'b00000000000000000001111001101110;
assign LUT_1[61761] = 32'b11111111111111111011001011101010;
assign LUT_1[61762] = 32'b11111111111111111101100111111111;
assign LUT_1[61763] = 32'b11111111111111110110111001111011;
assign LUT_1[61764] = 32'b00000000000000001001110011000101;
assign LUT_1[61765] = 32'b00000000000000000011000101000001;
assign LUT_1[61766] = 32'b00000000000000000101100001010110;
assign LUT_1[61767] = 32'b11111111111111111110110011010010;
assign LUT_1[61768] = 32'b00000000000000000001000111100011;
assign LUT_1[61769] = 32'b11111111111111111010011001011111;
assign LUT_1[61770] = 32'b11111111111111111100110101110100;
assign LUT_1[61771] = 32'b11111111111111110110000111110000;
assign LUT_1[61772] = 32'b00000000000000001001000000111010;
assign LUT_1[61773] = 32'b00000000000000000010010010110110;
assign LUT_1[61774] = 32'b00000000000000000100101111001011;
assign LUT_1[61775] = 32'b11111111111111111110000001000111;
assign LUT_1[61776] = 32'b00000000000000000011110101010000;
assign LUT_1[61777] = 32'b11111111111111111101000111001100;
assign LUT_1[61778] = 32'b11111111111111111111100011100001;
assign LUT_1[61779] = 32'b11111111111111111000110101011101;
assign LUT_1[61780] = 32'b00000000000000001011101110100111;
assign LUT_1[61781] = 32'b00000000000000000101000000100011;
assign LUT_1[61782] = 32'b00000000000000000111011100111000;
assign LUT_1[61783] = 32'b00000000000000000000101110110100;
assign LUT_1[61784] = 32'b00000000000000000011000011000101;
assign LUT_1[61785] = 32'b11111111111111111100010101000001;
assign LUT_1[61786] = 32'b11111111111111111110110001010110;
assign LUT_1[61787] = 32'b11111111111111111000000011010010;
assign LUT_1[61788] = 32'b00000000000000001010111100011100;
assign LUT_1[61789] = 32'b00000000000000000100001110011000;
assign LUT_1[61790] = 32'b00000000000000000110101010101101;
assign LUT_1[61791] = 32'b11111111111111111111111100101001;
assign LUT_1[61792] = 32'b00000000000000000010110100101101;
assign LUT_1[61793] = 32'b11111111111111111100000110101001;
assign LUT_1[61794] = 32'b11111111111111111110100010111110;
assign LUT_1[61795] = 32'b11111111111111110111110100111010;
assign LUT_1[61796] = 32'b00000000000000001010101110000100;
assign LUT_1[61797] = 32'b00000000000000000100000000000000;
assign LUT_1[61798] = 32'b00000000000000000110011100010101;
assign LUT_1[61799] = 32'b11111111111111111111101110010001;
assign LUT_1[61800] = 32'b00000000000000000010000010100010;
assign LUT_1[61801] = 32'b11111111111111111011010100011110;
assign LUT_1[61802] = 32'b11111111111111111101110000110011;
assign LUT_1[61803] = 32'b11111111111111110111000010101111;
assign LUT_1[61804] = 32'b00000000000000001001111011111001;
assign LUT_1[61805] = 32'b00000000000000000011001101110101;
assign LUT_1[61806] = 32'b00000000000000000101101010001010;
assign LUT_1[61807] = 32'b11111111111111111110111100000110;
assign LUT_1[61808] = 32'b00000000000000000100110000001111;
assign LUT_1[61809] = 32'b11111111111111111110000010001011;
assign LUT_1[61810] = 32'b00000000000000000000011110100000;
assign LUT_1[61811] = 32'b11111111111111111001110000011100;
assign LUT_1[61812] = 32'b00000000000000001100101001100110;
assign LUT_1[61813] = 32'b00000000000000000101111011100010;
assign LUT_1[61814] = 32'b00000000000000001000010111110111;
assign LUT_1[61815] = 32'b00000000000000000001101001110011;
assign LUT_1[61816] = 32'b00000000000000000011111110000100;
assign LUT_1[61817] = 32'b11111111111111111101010000000000;
assign LUT_1[61818] = 32'b11111111111111111111101100010101;
assign LUT_1[61819] = 32'b11111111111111111000111110010001;
assign LUT_1[61820] = 32'b00000000000000001011110111011011;
assign LUT_1[61821] = 32'b00000000000000000101001001010111;
assign LUT_1[61822] = 32'b00000000000000000111100101101100;
assign LUT_1[61823] = 32'b00000000000000000000110111101000;
assign LUT_1[61824] = 32'b00000000000000000010111100001001;
assign LUT_1[61825] = 32'b11111111111111111100001110000101;
assign LUT_1[61826] = 32'b11111111111111111110101010011010;
assign LUT_1[61827] = 32'b11111111111111110111111100010110;
assign LUT_1[61828] = 32'b00000000000000001010110101100000;
assign LUT_1[61829] = 32'b00000000000000000100000111011100;
assign LUT_1[61830] = 32'b00000000000000000110100011110001;
assign LUT_1[61831] = 32'b11111111111111111111110101101101;
assign LUT_1[61832] = 32'b00000000000000000010001001111110;
assign LUT_1[61833] = 32'b11111111111111111011011011111010;
assign LUT_1[61834] = 32'b11111111111111111101111000001111;
assign LUT_1[61835] = 32'b11111111111111110111001010001011;
assign LUT_1[61836] = 32'b00000000000000001010000011010101;
assign LUT_1[61837] = 32'b00000000000000000011010101010001;
assign LUT_1[61838] = 32'b00000000000000000101110001100110;
assign LUT_1[61839] = 32'b11111111111111111111000011100010;
assign LUT_1[61840] = 32'b00000000000000000100110111101011;
assign LUT_1[61841] = 32'b11111111111111111110001001100111;
assign LUT_1[61842] = 32'b00000000000000000000100101111100;
assign LUT_1[61843] = 32'b11111111111111111001110111111000;
assign LUT_1[61844] = 32'b00000000000000001100110001000010;
assign LUT_1[61845] = 32'b00000000000000000110000010111110;
assign LUT_1[61846] = 32'b00000000000000001000011111010011;
assign LUT_1[61847] = 32'b00000000000000000001110001001111;
assign LUT_1[61848] = 32'b00000000000000000100000101100000;
assign LUT_1[61849] = 32'b11111111111111111101010111011100;
assign LUT_1[61850] = 32'b11111111111111111111110011110001;
assign LUT_1[61851] = 32'b11111111111111111001000101101101;
assign LUT_1[61852] = 32'b00000000000000001011111110110111;
assign LUT_1[61853] = 32'b00000000000000000101010000110011;
assign LUT_1[61854] = 32'b00000000000000000111101101001000;
assign LUT_1[61855] = 32'b00000000000000000000111111000100;
assign LUT_1[61856] = 32'b00000000000000000011110111001000;
assign LUT_1[61857] = 32'b11111111111111111101001001000100;
assign LUT_1[61858] = 32'b11111111111111111111100101011001;
assign LUT_1[61859] = 32'b11111111111111111000110111010101;
assign LUT_1[61860] = 32'b00000000000000001011110000011111;
assign LUT_1[61861] = 32'b00000000000000000101000010011011;
assign LUT_1[61862] = 32'b00000000000000000111011110110000;
assign LUT_1[61863] = 32'b00000000000000000000110000101100;
assign LUT_1[61864] = 32'b00000000000000000011000100111101;
assign LUT_1[61865] = 32'b11111111111111111100010110111001;
assign LUT_1[61866] = 32'b11111111111111111110110011001110;
assign LUT_1[61867] = 32'b11111111111111111000000101001010;
assign LUT_1[61868] = 32'b00000000000000001010111110010100;
assign LUT_1[61869] = 32'b00000000000000000100010000010000;
assign LUT_1[61870] = 32'b00000000000000000110101100100101;
assign LUT_1[61871] = 32'b11111111111111111111111110100001;
assign LUT_1[61872] = 32'b00000000000000000101110010101010;
assign LUT_1[61873] = 32'b11111111111111111111000100100110;
assign LUT_1[61874] = 32'b00000000000000000001100000111011;
assign LUT_1[61875] = 32'b11111111111111111010110010110111;
assign LUT_1[61876] = 32'b00000000000000001101101100000001;
assign LUT_1[61877] = 32'b00000000000000000110111101111101;
assign LUT_1[61878] = 32'b00000000000000001001011010010010;
assign LUT_1[61879] = 32'b00000000000000000010101100001110;
assign LUT_1[61880] = 32'b00000000000000000101000000011111;
assign LUT_1[61881] = 32'b11111111111111111110010010011011;
assign LUT_1[61882] = 32'b00000000000000000000101110110000;
assign LUT_1[61883] = 32'b11111111111111111010000000101100;
assign LUT_1[61884] = 32'b00000000000000001100111001110110;
assign LUT_1[61885] = 32'b00000000000000000110001011110010;
assign LUT_1[61886] = 32'b00000000000000001000101000000111;
assign LUT_1[61887] = 32'b00000000000000000001111010000011;
assign LUT_1[61888] = 32'b00000000000000000100111001110001;
assign LUT_1[61889] = 32'b11111111111111111110001011101101;
assign LUT_1[61890] = 32'b00000000000000000000101000000010;
assign LUT_1[61891] = 32'b11111111111111111001111001111110;
assign LUT_1[61892] = 32'b00000000000000001100110011001000;
assign LUT_1[61893] = 32'b00000000000000000110000101000100;
assign LUT_1[61894] = 32'b00000000000000001000100001011001;
assign LUT_1[61895] = 32'b00000000000000000001110011010101;
assign LUT_1[61896] = 32'b00000000000000000100000111100110;
assign LUT_1[61897] = 32'b11111111111111111101011001100010;
assign LUT_1[61898] = 32'b11111111111111111111110101110111;
assign LUT_1[61899] = 32'b11111111111111111001000111110011;
assign LUT_1[61900] = 32'b00000000000000001100000000111101;
assign LUT_1[61901] = 32'b00000000000000000101010010111001;
assign LUT_1[61902] = 32'b00000000000000000111101111001110;
assign LUT_1[61903] = 32'b00000000000000000001000001001010;
assign LUT_1[61904] = 32'b00000000000000000110110101010011;
assign LUT_1[61905] = 32'b00000000000000000000000111001111;
assign LUT_1[61906] = 32'b00000000000000000010100011100100;
assign LUT_1[61907] = 32'b11111111111111111011110101100000;
assign LUT_1[61908] = 32'b00000000000000001110101110101010;
assign LUT_1[61909] = 32'b00000000000000001000000000100110;
assign LUT_1[61910] = 32'b00000000000000001010011100111011;
assign LUT_1[61911] = 32'b00000000000000000011101110110111;
assign LUT_1[61912] = 32'b00000000000000000110000011001000;
assign LUT_1[61913] = 32'b11111111111111111111010101000100;
assign LUT_1[61914] = 32'b00000000000000000001110001011001;
assign LUT_1[61915] = 32'b11111111111111111011000011010101;
assign LUT_1[61916] = 32'b00000000000000001101111100011111;
assign LUT_1[61917] = 32'b00000000000000000111001110011011;
assign LUT_1[61918] = 32'b00000000000000001001101010110000;
assign LUT_1[61919] = 32'b00000000000000000010111100101100;
assign LUT_1[61920] = 32'b00000000000000000101110100110000;
assign LUT_1[61921] = 32'b11111111111111111111000110101100;
assign LUT_1[61922] = 32'b00000000000000000001100011000001;
assign LUT_1[61923] = 32'b11111111111111111010110100111101;
assign LUT_1[61924] = 32'b00000000000000001101101110000111;
assign LUT_1[61925] = 32'b00000000000000000111000000000011;
assign LUT_1[61926] = 32'b00000000000000001001011100011000;
assign LUT_1[61927] = 32'b00000000000000000010101110010100;
assign LUT_1[61928] = 32'b00000000000000000101000010100101;
assign LUT_1[61929] = 32'b11111111111111111110010100100001;
assign LUT_1[61930] = 32'b00000000000000000000110000110110;
assign LUT_1[61931] = 32'b11111111111111111010000010110010;
assign LUT_1[61932] = 32'b00000000000000001100111011111100;
assign LUT_1[61933] = 32'b00000000000000000110001101111000;
assign LUT_1[61934] = 32'b00000000000000001000101010001101;
assign LUT_1[61935] = 32'b00000000000000000001111100001001;
assign LUT_1[61936] = 32'b00000000000000000111110000010010;
assign LUT_1[61937] = 32'b00000000000000000001000010001110;
assign LUT_1[61938] = 32'b00000000000000000011011110100011;
assign LUT_1[61939] = 32'b11111111111111111100110000011111;
assign LUT_1[61940] = 32'b00000000000000001111101001101001;
assign LUT_1[61941] = 32'b00000000000000001000111011100101;
assign LUT_1[61942] = 32'b00000000000000001011010111111010;
assign LUT_1[61943] = 32'b00000000000000000100101001110110;
assign LUT_1[61944] = 32'b00000000000000000110111110000111;
assign LUT_1[61945] = 32'b00000000000000000000010000000011;
assign LUT_1[61946] = 32'b00000000000000000010101100011000;
assign LUT_1[61947] = 32'b11111111111111111011111110010100;
assign LUT_1[61948] = 32'b00000000000000001110110111011110;
assign LUT_1[61949] = 32'b00000000000000001000001001011010;
assign LUT_1[61950] = 32'b00000000000000001010100101101111;
assign LUT_1[61951] = 32'b00000000000000000011110111101011;
assign LUT_1[61952] = 32'b11111111111111111011110110010111;
assign LUT_1[61953] = 32'b11111111111111110101001000010011;
assign LUT_1[61954] = 32'b11111111111111110111100100101000;
assign LUT_1[61955] = 32'b11111111111111110000110110100100;
assign LUT_1[61956] = 32'b00000000000000000011101111101110;
assign LUT_1[61957] = 32'b11111111111111111101000001101010;
assign LUT_1[61958] = 32'b11111111111111111111011101111111;
assign LUT_1[61959] = 32'b11111111111111111000101111111011;
assign LUT_1[61960] = 32'b11111111111111111011000100001100;
assign LUT_1[61961] = 32'b11111111111111110100010110001000;
assign LUT_1[61962] = 32'b11111111111111110110110010011101;
assign LUT_1[61963] = 32'b11111111111111110000000100011001;
assign LUT_1[61964] = 32'b00000000000000000010111101100011;
assign LUT_1[61965] = 32'b11111111111111111100001111011111;
assign LUT_1[61966] = 32'b11111111111111111110101011110100;
assign LUT_1[61967] = 32'b11111111111111110111111101110000;
assign LUT_1[61968] = 32'b11111111111111111101110001111001;
assign LUT_1[61969] = 32'b11111111111111110111000011110101;
assign LUT_1[61970] = 32'b11111111111111111001100000001010;
assign LUT_1[61971] = 32'b11111111111111110010110010000110;
assign LUT_1[61972] = 32'b00000000000000000101101011010000;
assign LUT_1[61973] = 32'b11111111111111111110111101001100;
assign LUT_1[61974] = 32'b00000000000000000001011001100001;
assign LUT_1[61975] = 32'b11111111111111111010101011011101;
assign LUT_1[61976] = 32'b11111111111111111100111111101110;
assign LUT_1[61977] = 32'b11111111111111110110010001101010;
assign LUT_1[61978] = 32'b11111111111111111000101101111111;
assign LUT_1[61979] = 32'b11111111111111110001111111111011;
assign LUT_1[61980] = 32'b00000000000000000100111001000101;
assign LUT_1[61981] = 32'b11111111111111111110001011000001;
assign LUT_1[61982] = 32'b00000000000000000000100111010110;
assign LUT_1[61983] = 32'b11111111111111111001111001010010;
assign LUT_1[61984] = 32'b11111111111111111100110001010110;
assign LUT_1[61985] = 32'b11111111111111110110000011010010;
assign LUT_1[61986] = 32'b11111111111111111000011111100111;
assign LUT_1[61987] = 32'b11111111111111110001110001100011;
assign LUT_1[61988] = 32'b00000000000000000100101010101101;
assign LUT_1[61989] = 32'b11111111111111111101111100101001;
assign LUT_1[61990] = 32'b00000000000000000000011000111110;
assign LUT_1[61991] = 32'b11111111111111111001101010111010;
assign LUT_1[61992] = 32'b11111111111111111011111111001011;
assign LUT_1[61993] = 32'b11111111111111110101010001000111;
assign LUT_1[61994] = 32'b11111111111111110111101101011100;
assign LUT_1[61995] = 32'b11111111111111110000111111011000;
assign LUT_1[61996] = 32'b00000000000000000011111000100010;
assign LUT_1[61997] = 32'b11111111111111111101001010011110;
assign LUT_1[61998] = 32'b11111111111111111111100110110011;
assign LUT_1[61999] = 32'b11111111111111111000111000101111;
assign LUT_1[62000] = 32'b11111111111111111110101100111000;
assign LUT_1[62001] = 32'b11111111111111110111111110110100;
assign LUT_1[62002] = 32'b11111111111111111010011011001001;
assign LUT_1[62003] = 32'b11111111111111110011101101000101;
assign LUT_1[62004] = 32'b00000000000000000110100110001111;
assign LUT_1[62005] = 32'b11111111111111111111111000001011;
assign LUT_1[62006] = 32'b00000000000000000010010100100000;
assign LUT_1[62007] = 32'b11111111111111111011100110011100;
assign LUT_1[62008] = 32'b11111111111111111101111010101101;
assign LUT_1[62009] = 32'b11111111111111110111001100101001;
assign LUT_1[62010] = 32'b11111111111111111001101000111110;
assign LUT_1[62011] = 32'b11111111111111110010111010111010;
assign LUT_1[62012] = 32'b00000000000000000101110100000100;
assign LUT_1[62013] = 32'b11111111111111111111000110000000;
assign LUT_1[62014] = 32'b00000000000000000001100010010101;
assign LUT_1[62015] = 32'b11111111111111111010110100010001;
assign LUT_1[62016] = 32'b11111111111111111101110011111111;
assign LUT_1[62017] = 32'b11111111111111110111000101111011;
assign LUT_1[62018] = 32'b11111111111111111001100010010000;
assign LUT_1[62019] = 32'b11111111111111110010110100001100;
assign LUT_1[62020] = 32'b00000000000000000101101101010110;
assign LUT_1[62021] = 32'b11111111111111111110111111010010;
assign LUT_1[62022] = 32'b00000000000000000001011011100111;
assign LUT_1[62023] = 32'b11111111111111111010101101100011;
assign LUT_1[62024] = 32'b11111111111111111101000001110100;
assign LUT_1[62025] = 32'b11111111111111110110010011110000;
assign LUT_1[62026] = 32'b11111111111111111000110000000101;
assign LUT_1[62027] = 32'b11111111111111110010000010000001;
assign LUT_1[62028] = 32'b00000000000000000100111011001011;
assign LUT_1[62029] = 32'b11111111111111111110001101000111;
assign LUT_1[62030] = 32'b00000000000000000000101001011100;
assign LUT_1[62031] = 32'b11111111111111111001111011011000;
assign LUT_1[62032] = 32'b11111111111111111111101111100001;
assign LUT_1[62033] = 32'b11111111111111111001000001011101;
assign LUT_1[62034] = 32'b11111111111111111011011101110010;
assign LUT_1[62035] = 32'b11111111111111110100101111101110;
assign LUT_1[62036] = 32'b00000000000000000111101000111000;
assign LUT_1[62037] = 32'b00000000000000000000111010110100;
assign LUT_1[62038] = 32'b00000000000000000011010111001001;
assign LUT_1[62039] = 32'b11111111111111111100101001000101;
assign LUT_1[62040] = 32'b11111111111111111110111101010110;
assign LUT_1[62041] = 32'b11111111111111111000001111010010;
assign LUT_1[62042] = 32'b11111111111111111010101011100111;
assign LUT_1[62043] = 32'b11111111111111110011111101100011;
assign LUT_1[62044] = 32'b00000000000000000110110110101101;
assign LUT_1[62045] = 32'b00000000000000000000001000101001;
assign LUT_1[62046] = 32'b00000000000000000010100100111110;
assign LUT_1[62047] = 32'b11111111111111111011110110111010;
assign LUT_1[62048] = 32'b11111111111111111110101110111110;
assign LUT_1[62049] = 32'b11111111111111111000000000111010;
assign LUT_1[62050] = 32'b11111111111111111010011101001111;
assign LUT_1[62051] = 32'b11111111111111110011101111001011;
assign LUT_1[62052] = 32'b00000000000000000110101000010101;
assign LUT_1[62053] = 32'b11111111111111111111111010010001;
assign LUT_1[62054] = 32'b00000000000000000010010110100110;
assign LUT_1[62055] = 32'b11111111111111111011101000100010;
assign LUT_1[62056] = 32'b11111111111111111101111100110011;
assign LUT_1[62057] = 32'b11111111111111110111001110101111;
assign LUT_1[62058] = 32'b11111111111111111001101011000100;
assign LUT_1[62059] = 32'b11111111111111110010111101000000;
assign LUT_1[62060] = 32'b00000000000000000101110110001010;
assign LUT_1[62061] = 32'b11111111111111111111001000000110;
assign LUT_1[62062] = 32'b00000000000000000001100100011011;
assign LUT_1[62063] = 32'b11111111111111111010110110010111;
assign LUT_1[62064] = 32'b00000000000000000000101010100000;
assign LUT_1[62065] = 32'b11111111111111111001111100011100;
assign LUT_1[62066] = 32'b11111111111111111100011000110001;
assign LUT_1[62067] = 32'b11111111111111110101101010101101;
assign LUT_1[62068] = 32'b00000000000000001000100011110111;
assign LUT_1[62069] = 32'b00000000000000000001110101110011;
assign LUT_1[62070] = 32'b00000000000000000100010010001000;
assign LUT_1[62071] = 32'b11111111111111111101100100000100;
assign LUT_1[62072] = 32'b11111111111111111111111000010101;
assign LUT_1[62073] = 32'b11111111111111111001001010010001;
assign LUT_1[62074] = 32'b11111111111111111011100110100110;
assign LUT_1[62075] = 32'b11111111111111110100111000100010;
assign LUT_1[62076] = 32'b00000000000000000111110001101100;
assign LUT_1[62077] = 32'b00000000000000000001000011101000;
assign LUT_1[62078] = 32'b00000000000000000011011111111101;
assign LUT_1[62079] = 32'b11111111111111111100110001111001;
assign LUT_1[62080] = 32'b11111111111111111110110110011010;
assign LUT_1[62081] = 32'b11111111111111111000001000010110;
assign LUT_1[62082] = 32'b11111111111111111010100100101011;
assign LUT_1[62083] = 32'b11111111111111110011110110100111;
assign LUT_1[62084] = 32'b00000000000000000110101111110001;
assign LUT_1[62085] = 32'b00000000000000000000000001101101;
assign LUT_1[62086] = 32'b00000000000000000010011110000010;
assign LUT_1[62087] = 32'b11111111111111111011101111111110;
assign LUT_1[62088] = 32'b11111111111111111110000100001111;
assign LUT_1[62089] = 32'b11111111111111110111010110001011;
assign LUT_1[62090] = 32'b11111111111111111001110010100000;
assign LUT_1[62091] = 32'b11111111111111110011000100011100;
assign LUT_1[62092] = 32'b00000000000000000101111101100110;
assign LUT_1[62093] = 32'b11111111111111111111001111100010;
assign LUT_1[62094] = 32'b00000000000000000001101011110111;
assign LUT_1[62095] = 32'b11111111111111111010111101110011;
assign LUT_1[62096] = 32'b00000000000000000000110001111100;
assign LUT_1[62097] = 32'b11111111111111111010000011111000;
assign LUT_1[62098] = 32'b11111111111111111100100000001101;
assign LUT_1[62099] = 32'b11111111111111110101110010001001;
assign LUT_1[62100] = 32'b00000000000000001000101011010011;
assign LUT_1[62101] = 32'b00000000000000000001111101001111;
assign LUT_1[62102] = 32'b00000000000000000100011001100100;
assign LUT_1[62103] = 32'b11111111111111111101101011100000;
assign LUT_1[62104] = 32'b11111111111111111111111111110001;
assign LUT_1[62105] = 32'b11111111111111111001010001101101;
assign LUT_1[62106] = 32'b11111111111111111011101110000010;
assign LUT_1[62107] = 32'b11111111111111110100111111111110;
assign LUT_1[62108] = 32'b00000000000000000111111001001000;
assign LUT_1[62109] = 32'b00000000000000000001001011000100;
assign LUT_1[62110] = 32'b00000000000000000011100111011001;
assign LUT_1[62111] = 32'b11111111111111111100111001010101;
assign LUT_1[62112] = 32'b11111111111111111111110001011001;
assign LUT_1[62113] = 32'b11111111111111111001000011010101;
assign LUT_1[62114] = 32'b11111111111111111011011111101010;
assign LUT_1[62115] = 32'b11111111111111110100110001100110;
assign LUT_1[62116] = 32'b00000000000000000111101010110000;
assign LUT_1[62117] = 32'b00000000000000000000111100101100;
assign LUT_1[62118] = 32'b00000000000000000011011001000001;
assign LUT_1[62119] = 32'b11111111111111111100101010111101;
assign LUT_1[62120] = 32'b11111111111111111110111111001110;
assign LUT_1[62121] = 32'b11111111111111111000010001001010;
assign LUT_1[62122] = 32'b11111111111111111010101101011111;
assign LUT_1[62123] = 32'b11111111111111110011111111011011;
assign LUT_1[62124] = 32'b00000000000000000110111000100101;
assign LUT_1[62125] = 32'b00000000000000000000001010100001;
assign LUT_1[62126] = 32'b00000000000000000010100110110110;
assign LUT_1[62127] = 32'b11111111111111111011111000110010;
assign LUT_1[62128] = 32'b00000000000000000001101100111011;
assign LUT_1[62129] = 32'b11111111111111111010111110110111;
assign LUT_1[62130] = 32'b11111111111111111101011011001100;
assign LUT_1[62131] = 32'b11111111111111110110101101001000;
assign LUT_1[62132] = 32'b00000000000000001001100110010010;
assign LUT_1[62133] = 32'b00000000000000000010111000001110;
assign LUT_1[62134] = 32'b00000000000000000101010100100011;
assign LUT_1[62135] = 32'b11111111111111111110100110011111;
assign LUT_1[62136] = 32'b00000000000000000000111010110000;
assign LUT_1[62137] = 32'b11111111111111111010001100101100;
assign LUT_1[62138] = 32'b11111111111111111100101001000001;
assign LUT_1[62139] = 32'b11111111111111110101111010111101;
assign LUT_1[62140] = 32'b00000000000000001000110100000111;
assign LUT_1[62141] = 32'b00000000000000000010000110000011;
assign LUT_1[62142] = 32'b00000000000000000100100010011000;
assign LUT_1[62143] = 32'b11111111111111111101110100010100;
assign LUT_1[62144] = 32'b00000000000000000000110100000010;
assign LUT_1[62145] = 32'b11111111111111111010000101111110;
assign LUT_1[62146] = 32'b11111111111111111100100010010011;
assign LUT_1[62147] = 32'b11111111111111110101110100001111;
assign LUT_1[62148] = 32'b00000000000000001000101101011001;
assign LUT_1[62149] = 32'b00000000000000000001111111010101;
assign LUT_1[62150] = 32'b00000000000000000100011011101010;
assign LUT_1[62151] = 32'b11111111111111111101101101100110;
assign LUT_1[62152] = 32'b00000000000000000000000001110111;
assign LUT_1[62153] = 32'b11111111111111111001010011110011;
assign LUT_1[62154] = 32'b11111111111111111011110000001000;
assign LUT_1[62155] = 32'b11111111111111110101000010000100;
assign LUT_1[62156] = 32'b00000000000000000111111011001110;
assign LUT_1[62157] = 32'b00000000000000000001001101001010;
assign LUT_1[62158] = 32'b00000000000000000011101001011111;
assign LUT_1[62159] = 32'b11111111111111111100111011011011;
assign LUT_1[62160] = 32'b00000000000000000010101111100100;
assign LUT_1[62161] = 32'b11111111111111111100000001100000;
assign LUT_1[62162] = 32'b11111111111111111110011101110101;
assign LUT_1[62163] = 32'b11111111111111110111101111110001;
assign LUT_1[62164] = 32'b00000000000000001010101000111011;
assign LUT_1[62165] = 32'b00000000000000000011111010110111;
assign LUT_1[62166] = 32'b00000000000000000110010111001100;
assign LUT_1[62167] = 32'b11111111111111111111101001001000;
assign LUT_1[62168] = 32'b00000000000000000001111101011001;
assign LUT_1[62169] = 32'b11111111111111111011001111010101;
assign LUT_1[62170] = 32'b11111111111111111101101011101010;
assign LUT_1[62171] = 32'b11111111111111110110111101100110;
assign LUT_1[62172] = 32'b00000000000000001001110110110000;
assign LUT_1[62173] = 32'b00000000000000000011001000101100;
assign LUT_1[62174] = 32'b00000000000000000101100101000001;
assign LUT_1[62175] = 32'b11111111111111111110110110111101;
assign LUT_1[62176] = 32'b00000000000000000001101111000001;
assign LUT_1[62177] = 32'b11111111111111111011000000111101;
assign LUT_1[62178] = 32'b11111111111111111101011101010010;
assign LUT_1[62179] = 32'b11111111111111110110101111001110;
assign LUT_1[62180] = 32'b00000000000000001001101000011000;
assign LUT_1[62181] = 32'b00000000000000000010111010010100;
assign LUT_1[62182] = 32'b00000000000000000101010110101001;
assign LUT_1[62183] = 32'b11111111111111111110101000100101;
assign LUT_1[62184] = 32'b00000000000000000000111100110110;
assign LUT_1[62185] = 32'b11111111111111111010001110110010;
assign LUT_1[62186] = 32'b11111111111111111100101011000111;
assign LUT_1[62187] = 32'b11111111111111110101111101000011;
assign LUT_1[62188] = 32'b00000000000000001000110110001101;
assign LUT_1[62189] = 32'b00000000000000000010001000001001;
assign LUT_1[62190] = 32'b00000000000000000100100100011110;
assign LUT_1[62191] = 32'b11111111111111111101110110011010;
assign LUT_1[62192] = 32'b00000000000000000011101010100011;
assign LUT_1[62193] = 32'b11111111111111111100111100011111;
assign LUT_1[62194] = 32'b11111111111111111111011000110100;
assign LUT_1[62195] = 32'b11111111111111111000101010110000;
assign LUT_1[62196] = 32'b00000000000000001011100011111010;
assign LUT_1[62197] = 32'b00000000000000000100110101110110;
assign LUT_1[62198] = 32'b00000000000000000111010010001011;
assign LUT_1[62199] = 32'b00000000000000000000100100000111;
assign LUT_1[62200] = 32'b00000000000000000010111000011000;
assign LUT_1[62201] = 32'b11111111111111111100001010010100;
assign LUT_1[62202] = 32'b11111111111111111110100110101001;
assign LUT_1[62203] = 32'b11111111111111110111111000100101;
assign LUT_1[62204] = 32'b00000000000000001010110001101111;
assign LUT_1[62205] = 32'b00000000000000000100000011101011;
assign LUT_1[62206] = 32'b00000000000000000110100000000000;
assign LUT_1[62207] = 32'b11111111111111111111110001111100;
assign LUT_1[62208] = 32'b11111111111111111001101010100011;
assign LUT_1[62209] = 32'b11111111111111110010111100011111;
assign LUT_1[62210] = 32'b11111111111111110101011000110100;
assign LUT_1[62211] = 32'b11111111111111101110101010110000;
assign LUT_1[62212] = 32'b00000000000000000001100011111010;
assign LUT_1[62213] = 32'b11111111111111111010110101110110;
assign LUT_1[62214] = 32'b11111111111111111101010010001011;
assign LUT_1[62215] = 32'b11111111111111110110100100000111;
assign LUT_1[62216] = 32'b11111111111111111000111000011000;
assign LUT_1[62217] = 32'b11111111111111110010001010010100;
assign LUT_1[62218] = 32'b11111111111111110100100110101001;
assign LUT_1[62219] = 32'b11111111111111101101111000100101;
assign LUT_1[62220] = 32'b00000000000000000000110001101111;
assign LUT_1[62221] = 32'b11111111111111111010000011101011;
assign LUT_1[62222] = 32'b11111111111111111100100000000000;
assign LUT_1[62223] = 32'b11111111111111110101110001111100;
assign LUT_1[62224] = 32'b11111111111111111011100110000101;
assign LUT_1[62225] = 32'b11111111111111110100111000000001;
assign LUT_1[62226] = 32'b11111111111111110111010100010110;
assign LUT_1[62227] = 32'b11111111111111110000100110010010;
assign LUT_1[62228] = 32'b00000000000000000011011111011100;
assign LUT_1[62229] = 32'b11111111111111111100110001011000;
assign LUT_1[62230] = 32'b11111111111111111111001101101101;
assign LUT_1[62231] = 32'b11111111111111111000011111101001;
assign LUT_1[62232] = 32'b11111111111111111010110011111010;
assign LUT_1[62233] = 32'b11111111111111110100000101110110;
assign LUT_1[62234] = 32'b11111111111111110110100010001011;
assign LUT_1[62235] = 32'b11111111111111101111110100000111;
assign LUT_1[62236] = 32'b00000000000000000010101101010001;
assign LUT_1[62237] = 32'b11111111111111111011111111001101;
assign LUT_1[62238] = 32'b11111111111111111110011011100010;
assign LUT_1[62239] = 32'b11111111111111110111101101011110;
assign LUT_1[62240] = 32'b11111111111111111010100101100010;
assign LUT_1[62241] = 32'b11111111111111110011110111011110;
assign LUT_1[62242] = 32'b11111111111111110110010011110011;
assign LUT_1[62243] = 32'b11111111111111101111100101101111;
assign LUT_1[62244] = 32'b00000000000000000010011110111001;
assign LUT_1[62245] = 32'b11111111111111111011110000110101;
assign LUT_1[62246] = 32'b11111111111111111110001101001010;
assign LUT_1[62247] = 32'b11111111111111110111011111000110;
assign LUT_1[62248] = 32'b11111111111111111001110011010111;
assign LUT_1[62249] = 32'b11111111111111110011000101010011;
assign LUT_1[62250] = 32'b11111111111111110101100001101000;
assign LUT_1[62251] = 32'b11111111111111101110110011100100;
assign LUT_1[62252] = 32'b00000000000000000001101100101110;
assign LUT_1[62253] = 32'b11111111111111111010111110101010;
assign LUT_1[62254] = 32'b11111111111111111101011010111111;
assign LUT_1[62255] = 32'b11111111111111110110101100111011;
assign LUT_1[62256] = 32'b11111111111111111100100001000100;
assign LUT_1[62257] = 32'b11111111111111110101110011000000;
assign LUT_1[62258] = 32'b11111111111111111000001111010101;
assign LUT_1[62259] = 32'b11111111111111110001100001010001;
assign LUT_1[62260] = 32'b00000000000000000100011010011011;
assign LUT_1[62261] = 32'b11111111111111111101101100010111;
assign LUT_1[62262] = 32'b00000000000000000000001000101100;
assign LUT_1[62263] = 32'b11111111111111111001011010101000;
assign LUT_1[62264] = 32'b11111111111111111011101110111001;
assign LUT_1[62265] = 32'b11111111111111110101000000110101;
assign LUT_1[62266] = 32'b11111111111111110111011101001010;
assign LUT_1[62267] = 32'b11111111111111110000101111000110;
assign LUT_1[62268] = 32'b00000000000000000011101000010000;
assign LUT_1[62269] = 32'b11111111111111111100111010001100;
assign LUT_1[62270] = 32'b11111111111111111111010110100001;
assign LUT_1[62271] = 32'b11111111111111111000101000011101;
assign LUT_1[62272] = 32'b11111111111111111011101000001011;
assign LUT_1[62273] = 32'b11111111111111110100111010000111;
assign LUT_1[62274] = 32'b11111111111111110111010110011100;
assign LUT_1[62275] = 32'b11111111111111110000101000011000;
assign LUT_1[62276] = 32'b00000000000000000011100001100010;
assign LUT_1[62277] = 32'b11111111111111111100110011011110;
assign LUT_1[62278] = 32'b11111111111111111111001111110011;
assign LUT_1[62279] = 32'b11111111111111111000100001101111;
assign LUT_1[62280] = 32'b11111111111111111010110110000000;
assign LUT_1[62281] = 32'b11111111111111110100000111111100;
assign LUT_1[62282] = 32'b11111111111111110110100100010001;
assign LUT_1[62283] = 32'b11111111111111101111110110001101;
assign LUT_1[62284] = 32'b00000000000000000010101111010111;
assign LUT_1[62285] = 32'b11111111111111111100000001010011;
assign LUT_1[62286] = 32'b11111111111111111110011101101000;
assign LUT_1[62287] = 32'b11111111111111110111101111100100;
assign LUT_1[62288] = 32'b11111111111111111101100011101101;
assign LUT_1[62289] = 32'b11111111111111110110110101101001;
assign LUT_1[62290] = 32'b11111111111111111001010001111110;
assign LUT_1[62291] = 32'b11111111111111110010100011111010;
assign LUT_1[62292] = 32'b00000000000000000101011101000100;
assign LUT_1[62293] = 32'b11111111111111111110101111000000;
assign LUT_1[62294] = 32'b00000000000000000001001011010101;
assign LUT_1[62295] = 32'b11111111111111111010011101010001;
assign LUT_1[62296] = 32'b11111111111111111100110001100010;
assign LUT_1[62297] = 32'b11111111111111110110000011011110;
assign LUT_1[62298] = 32'b11111111111111111000011111110011;
assign LUT_1[62299] = 32'b11111111111111110001110001101111;
assign LUT_1[62300] = 32'b00000000000000000100101010111001;
assign LUT_1[62301] = 32'b11111111111111111101111100110101;
assign LUT_1[62302] = 32'b00000000000000000000011001001010;
assign LUT_1[62303] = 32'b11111111111111111001101011000110;
assign LUT_1[62304] = 32'b11111111111111111100100011001010;
assign LUT_1[62305] = 32'b11111111111111110101110101000110;
assign LUT_1[62306] = 32'b11111111111111111000010001011011;
assign LUT_1[62307] = 32'b11111111111111110001100011010111;
assign LUT_1[62308] = 32'b00000000000000000100011100100001;
assign LUT_1[62309] = 32'b11111111111111111101101110011101;
assign LUT_1[62310] = 32'b00000000000000000000001010110010;
assign LUT_1[62311] = 32'b11111111111111111001011100101110;
assign LUT_1[62312] = 32'b11111111111111111011110000111111;
assign LUT_1[62313] = 32'b11111111111111110101000010111011;
assign LUT_1[62314] = 32'b11111111111111110111011111010000;
assign LUT_1[62315] = 32'b11111111111111110000110001001100;
assign LUT_1[62316] = 32'b00000000000000000011101010010110;
assign LUT_1[62317] = 32'b11111111111111111100111100010010;
assign LUT_1[62318] = 32'b11111111111111111111011000100111;
assign LUT_1[62319] = 32'b11111111111111111000101010100011;
assign LUT_1[62320] = 32'b11111111111111111110011110101100;
assign LUT_1[62321] = 32'b11111111111111110111110000101000;
assign LUT_1[62322] = 32'b11111111111111111010001100111101;
assign LUT_1[62323] = 32'b11111111111111110011011110111001;
assign LUT_1[62324] = 32'b00000000000000000110011000000011;
assign LUT_1[62325] = 32'b11111111111111111111101001111111;
assign LUT_1[62326] = 32'b00000000000000000010000110010100;
assign LUT_1[62327] = 32'b11111111111111111011011000010000;
assign LUT_1[62328] = 32'b11111111111111111101101100100001;
assign LUT_1[62329] = 32'b11111111111111110110111110011101;
assign LUT_1[62330] = 32'b11111111111111111001011010110010;
assign LUT_1[62331] = 32'b11111111111111110010101100101110;
assign LUT_1[62332] = 32'b00000000000000000101100101111000;
assign LUT_1[62333] = 32'b11111111111111111110110111110100;
assign LUT_1[62334] = 32'b00000000000000000001010100001001;
assign LUT_1[62335] = 32'b11111111111111111010100110000101;
assign LUT_1[62336] = 32'b11111111111111111100101010100110;
assign LUT_1[62337] = 32'b11111111111111110101111100100010;
assign LUT_1[62338] = 32'b11111111111111111000011000110111;
assign LUT_1[62339] = 32'b11111111111111110001101010110011;
assign LUT_1[62340] = 32'b00000000000000000100100011111101;
assign LUT_1[62341] = 32'b11111111111111111101110101111001;
assign LUT_1[62342] = 32'b00000000000000000000010010001110;
assign LUT_1[62343] = 32'b11111111111111111001100100001010;
assign LUT_1[62344] = 32'b11111111111111111011111000011011;
assign LUT_1[62345] = 32'b11111111111111110101001010010111;
assign LUT_1[62346] = 32'b11111111111111110111100110101100;
assign LUT_1[62347] = 32'b11111111111111110000111000101000;
assign LUT_1[62348] = 32'b00000000000000000011110001110010;
assign LUT_1[62349] = 32'b11111111111111111101000011101110;
assign LUT_1[62350] = 32'b11111111111111111111100000000011;
assign LUT_1[62351] = 32'b11111111111111111000110001111111;
assign LUT_1[62352] = 32'b11111111111111111110100110001000;
assign LUT_1[62353] = 32'b11111111111111110111111000000100;
assign LUT_1[62354] = 32'b11111111111111111010010100011001;
assign LUT_1[62355] = 32'b11111111111111110011100110010101;
assign LUT_1[62356] = 32'b00000000000000000110011111011111;
assign LUT_1[62357] = 32'b11111111111111111111110001011011;
assign LUT_1[62358] = 32'b00000000000000000010001101110000;
assign LUT_1[62359] = 32'b11111111111111111011011111101100;
assign LUT_1[62360] = 32'b11111111111111111101110011111101;
assign LUT_1[62361] = 32'b11111111111111110111000101111001;
assign LUT_1[62362] = 32'b11111111111111111001100010001110;
assign LUT_1[62363] = 32'b11111111111111110010110100001010;
assign LUT_1[62364] = 32'b00000000000000000101101101010100;
assign LUT_1[62365] = 32'b11111111111111111110111111010000;
assign LUT_1[62366] = 32'b00000000000000000001011011100101;
assign LUT_1[62367] = 32'b11111111111111111010101101100001;
assign LUT_1[62368] = 32'b11111111111111111101100101100101;
assign LUT_1[62369] = 32'b11111111111111110110110111100001;
assign LUT_1[62370] = 32'b11111111111111111001010011110110;
assign LUT_1[62371] = 32'b11111111111111110010100101110010;
assign LUT_1[62372] = 32'b00000000000000000101011110111100;
assign LUT_1[62373] = 32'b11111111111111111110110000111000;
assign LUT_1[62374] = 32'b00000000000000000001001101001101;
assign LUT_1[62375] = 32'b11111111111111111010011111001001;
assign LUT_1[62376] = 32'b11111111111111111100110011011010;
assign LUT_1[62377] = 32'b11111111111111110110000101010110;
assign LUT_1[62378] = 32'b11111111111111111000100001101011;
assign LUT_1[62379] = 32'b11111111111111110001110011100111;
assign LUT_1[62380] = 32'b00000000000000000100101100110001;
assign LUT_1[62381] = 32'b11111111111111111101111110101101;
assign LUT_1[62382] = 32'b00000000000000000000011011000010;
assign LUT_1[62383] = 32'b11111111111111111001101100111110;
assign LUT_1[62384] = 32'b11111111111111111111100001000111;
assign LUT_1[62385] = 32'b11111111111111111000110011000011;
assign LUT_1[62386] = 32'b11111111111111111011001111011000;
assign LUT_1[62387] = 32'b11111111111111110100100001010100;
assign LUT_1[62388] = 32'b00000000000000000111011010011110;
assign LUT_1[62389] = 32'b00000000000000000000101100011010;
assign LUT_1[62390] = 32'b00000000000000000011001000101111;
assign LUT_1[62391] = 32'b11111111111111111100011010101011;
assign LUT_1[62392] = 32'b11111111111111111110101110111100;
assign LUT_1[62393] = 32'b11111111111111111000000000111000;
assign LUT_1[62394] = 32'b11111111111111111010011101001101;
assign LUT_1[62395] = 32'b11111111111111110011101111001001;
assign LUT_1[62396] = 32'b00000000000000000110101000010011;
assign LUT_1[62397] = 32'b11111111111111111111111010001111;
assign LUT_1[62398] = 32'b00000000000000000010010110100100;
assign LUT_1[62399] = 32'b11111111111111111011101000100000;
assign LUT_1[62400] = 32'b11111111111111111110101000001110;
assign LUT_1[62401] = 32'b11111111111111110111111010001010;
assign LUT_1[62402] = 32'b11111111111111111010010110011111;
assign LUT_1[62403] = 32'b11111111111111110011101000011011;
assign LUT_1[62404] = 32'b00000000000000000110100001100101;
assign LUT_1[62405] = 32'b11111111111111111111110011100001;
assign LUT_1[62406] = 32'b00000000000000000010001111110110;
assign LUT_1[62407] = 32'b11111111111111111011100001110010;
assign LUT_1[62408] = 32'b11111111111111111101110110000011;
assign LUT_1[62409] = 32'b11111111111111110111000111111111;
assign LUT_1[62410] = 32'b11111111111111111001100100010100;
assign LUT_1[62411] = 32'b11111111111111110010110110010000;
assign LUT_1[62412] = 32'b00000000000000000101101111011010;
assign LUT_1[62413] = 32'b11111111111111111111000001010110;
assign LUT_1[62414] = 32'b00000000000000000001011101101011;
assign LUT_1[62415] = 32'b11111111111111111010101111100111;
assign LUT_1[62416] = 32'b00000000000000000000100011110000;
assign LUT_1[62417] = 32'b11111111111111111001110101101100;
assign LUT_1[62418] = 32'b11111111111111111100010010000001;
assign LUT_1[62419] = 32'b11111111111111110101100011111101;
assign LUT_1[62420] = 32'b00000000000000001000011101000111;
assign LUT_1[62421] = 32'b00000000000000000001101111000011;
assign LUT_1[62422] = 32'b00000000000000000100001011011000;
assign LUT_1[62423] = 32'b11111111111111111101011101010100;
assign LUT_1[62424] = 32'b11111111111111111111110001100101;
assign LUT_1[62425] = 32'b11111111111111111001000011100001;
assign LUT_1[62426] = 32'b11111111111111111011011111110110;
assign LUT_1[62427] = 32'b11111111111111110100110001110010;
assign LUT_1[62428] = 32'b00000000000000000111101010111100;
assign LUT_1[62429] = 32'b00000000000000000000111100111000;
assign LUT_1[62430] = 32'b00000000000000000011011001001101;
assign LUT_1[62431] = 32'b11111111111111111100101011001001;
assign LUT_1[62432] = 32'b11111111111111111111100011001101;
assign LUT_1[62433] = 32'b11111111111111111000110101001001;
assign LUT_1[62434] = 32'b11111111111111111011010001011110;
assign LUT_1[62435] = 32'b11111111111111110100100011011010;
assign LUT_1[62436] = 32'b00000000000000000111011100100100;
assign LUT_1[62437] = 32'b00000000000000000000101110100000;
assign LUT_1[62438] = 32'b00000000000000000011001010110101;
assign LUT_1[62439] = 32'b11111111111111111100011100110001;
assign LUT_1[62440] = 32'b11111111111111111110110001000010;
assign LUT_1[62441] = 32'b11111111111111111000000010111110;
assign LUT_1[62442] = 32'b11111111111111111010011111010011;
assign LUT_1[62443] = 32'b11111111111111110011110001001111;
assign LUT_1[62444] = 32'b00000000000000000110101010011001;
assign LUT_1[62445] = 32'b11111111111111111111111100010101;
assign LUT_1[62446] = 32'b00000000000000000010011000101010;
assign LUT_1[62447] = 32'b11111111111111111011101010100110;
assign LUT_1[62448] = 32'b00000000000000000001011110101111;
assign LUT_1[62449] = 32'b11111111111111111010110000101011;
assign LUT_1[62450] = 32'b11111111111111111101001101000000;
assign LUT_1[62451] = 32'b11111111111111110110011110111100;
assign LUT_1[62452] = 32'b00000000000000001001011000000110;
assign LUT_1[62453] = 32'b00000000000000000010101010000010;
assign LUT_1[62454] = 32'b00000000000000000101000110010111;
assign LUT_1[62455] = 32'b11111111111111111110011000010011;
assign LUT_1[62456] = 32'b00000000000000000000101100100100;
assign LUT_1[62457] = 32'b11111111111111111001111110100000;
assign LUT_1[62458] = 32'b11111111111111111100011010110101;
assign LUT_1[62459] = 32'b11111111111111110101101100110001;
assign LUT_1[62460] = 32'b00000000000000001000100101111011;
assign LUT_1[62461] = 32'b00000000000000000001110111110111;
assign LUT_1[62462] = 32'b00000000000000000100010100001100;
assign LUT_1[62463] = 32'b11111111111111111101100110001000;
assign LUT_1[62464] = 32'b00000000000000001000011110101010;
assign LUT_1[62465] = 32'b00000000000000000001110000100110;
assign LUT_1[62466] = 32'b00000000000000000100001100111011;
assign LUT_1[62467] = 32'b11111111111111111101011110110111;
assign LUT_1[62468] = 32'b00000000000000010000011000000001;
assign LUT_1[62469] = 32'b00000000000000001001101001111101;
assign LUT_1[62470] = 32'b00000000000000001100000110010010;
assign LUT_1[62471] = 32'b00000000000000000101011000001110;
assign LUT_1[62472] = 32'b00000000000000000111101100011111;
assign LUT_1[62473] = 32'b00000000000000000000111110011011;
assign LUT_1[62474] = 32'b00000000000000000011011010110000;
assign LUT_1[62475] = 32'b11111111111111111100101100101100;
assign LUT_1[62476] = 32'b00000000000000001111100101110110;
assign LUT_1[62477] = 32'b00000000000000001000110111110010;
assign LUT_1[62478] = 32'b00000000000000001011010100000111;
assign LUT_1[62479] = 32'b00000000000000000100100110000011;
assign LUT_1[62480] = 32'b00000000000000001010011010001100;
assign LUT_1[62481] = 32'b00000000000000000011101100001000;
assign LUT_1[62482] = 32'b00000000000000000110001000011101;
assign LUT_1[62483] = 32'b11111111111111111111011010011001;
assign LUT_1[62484] = 32'b00000000000000010010010011100011;
assign LUT_1[62485] = 32'b00000000000000001011100101011111;
assign LUT_1[62486] = 32'b00000000000000001110000001110100;
assign LUT_1[62487] = 32'b00000000000000000111010011110000;
assign LUT_1[62488] = 32'b00000000000000001001101000000001;
assign LUT_1[62489] = 32'b00000000000000000010111001111101;
assign LUT_1[62490] = 32'b00000000000000000101010110010010;
assign LUT_1[62491] = 32'b11111111111111111110101000001110;
assign LUT_1[62492] = 32'b00000000000000010001100001011000;
assign LUT_1[62493] = 32'b00000000000000001010110011010100;
assign LUT_1[62494] = 32'b00000000000000001101001111101001;
assign LUT_1[62495] = 32'b00000000000000000110100001100101;
assign LUT_1[62496] = 32'b00000000000000001001011001101001;
assign LUT_1[62497] = 32'b00000000000000000010101011100101;
assign LUT_1[62498] = 32'b00000000000000000101000111111010;
assign LUT_1[62499] = 32'b11111111111111111110011001110110;
assign LUT_1[62500] = 32'b00000000000000010001010011000000;
assign LUT_1[62501] = 32'b00000000000000001010100100111100;
assign LUT_1[62502] = 32'b00000000000000001101000001010001;
assign LUT_1[62503] = 32'b00000000000000000110010011001101;
assign LUT_1[62504] = 32'b00000000000000001000100111011110;
assign LUT_1[62505] = 32'b00000000000000000001111001011010;
assign LUT_1[62506] = 32'b00000000000000000100010101101111;
assign LUT_1[62507] = 32'b11111111111111111101100111101011;
assign LUT_1[62508] = 32'b00000000000000010000100000110101;
assign LUT_1[62509] = 32'b00000000000000001001110010110001;
assign LUT_1[62510] = 32'b00000000000000001100001111000110;
assign LUT_1[62511] = 32'b00000000000000000101100001000010;
assign LUT_1[62512] = 32'b00000000000000001011010101001011;
assign LUT_1[62513] = 32'b00000000000000000100100111000111;
assign LUT_1[62514] = 32'b00000000000000000111000011011100;
assign LUT_1[62515] = 32'b00000000000000000000010101011000;
assign LUT_1[62516] = 32'b00000000000000010011001110100010;
assign LUT_1[62517] = 32'b00000000000000001100100000011110;
assign LUT_1[62518] = 32'b00000000000000001110111100110011;
assign LUT_1[62519] = 32'b00000000000000001000001110101111;
assign LUT_1[62520] = 32'b00000000000000001010100011000000;
assign LUT_1[62521] = 32'b00000000000000000011110100111100;
assign LUT_1[62522] = 32'b00000000000000000110010001010001;
assign LUT_1[62523] = 32'b11111111111111111111100011001101;
assign LUT_1[62524] = 32'b00000000000000010010011100010111;
assign LUT_1[62525] = 32'b00000000000000001011101110010011;
assign LUT_1[62526] = 32'b00000000000000001110001010101000;
assign LUT_1[62527] = 32'b00000000000000000111011100100100;
assign LUT_1[62528] = 32'b00000000000000001010011100010010;
assign LUT_1[62529] = 32'b00000000000000000011101110001110;
assign LUT_1[62530] = 32'b00000000000000000110001010100011;
assign LUT_1[62531] = 32'b11111111111111111111011100011111;
assign LUT_1[62532] = 32'b00000000000000010010010101101001;
assign LUT_1[62533] = 32'b00000000000000001011100111100101;
assign LUT_1[62534] = 32'b00000000000000001110000011111010;
assign LUT_1[62535] = 32'b00000000000000000111010101110110;
assign LUT_1[62536] = 32'b00000000000000001001101010000111;
assign LUT_1[62537] = 32'b00000000000000000010111100000011;
assign LUT_1[62538] = 32'b00000000000000000101011000011000;
assign LUT_1[62539] = 32'b11111111111111111110101010010100;
assign LUT_1[62540] = 32'b00000000000000010001100011011110;
assign LUT_1[62541] = 32'b00000000000000001010110101011010;
assign LUT_1[62542] = 32'b00000000000000001101010001101111;
assign LUT_1[62543] = 32'b00000000000000000110100011101011;
assign LUT_1[62544] = 32'b00000000000000001100010111110100;
assign LUT_1[62545] = 32'b00000000000000000101101001110000;
assign LUT_1[62546] = 32'b00000000000000001000000110000101;
assign LUT_1[62547] = 32'b00000000000000000001011000000001;
assign LUT_1[62548] = 32'b00000000000000010100010001001011;
assign LUT_1[62549] = 32'b00000000000000001101100011000111;
assign LUT_1[62550] = 32'b00000000000000001111111111011100;
assign LUT_1[62551] = 32'b00000000000000001001010001011000;
assign LUT_1[62552] = 32'b00000000000000001011100101101001;
assign LUT_1[62553] = 32'b00000000000000000100110111100101;
assign LUT_1[62554] = 32'b00000000000000000111010011111010;
assign LUT_1[62555] = 32'b00000000000000000000100101110110;
assign LUT_1[62556] = 32'b00000000000000010011011111000000;
assign LUT_1[62557] = 32'b00000000000000001100110000111100;
assign LUT_1[62558] = 32'b00000000000000001111001101010001;
assign LUT_1[62559] = 32'b00000000000000001000011111001101;
assign LUT_1[62560] = 32'b00000000000000001011010111010001;
assign LUT_1[62561] = 32'b00000000000000000100101001001101;
assign LUT_1[62562] = 32'b00000000000000000111000101100010;
assign LUT_1[62563] = 32'b00000000000000000000010111011110;
assign LUT_1[62564] = 32'b00000000000000010011010000101000;
assign LUT_1[62565] = 32'b00000000000000001100100010100100;
assign LUT_1[62566] = 32'b00000000000000001110111110111001;
assign LUT_1[62567] = 32'b00000000000000001000010000110101;
assign LUT_1[62568] = 32'b00000000000000001010100101000110;
assign LUT_1[62569] = 32'b00000000000000000011110111000010;
assign LUT_1[62570] = 32'b00000000000000000110010011010111;
assign LUT_1[62571] = 32'b11111111111111111111100101010011;
assign LUT_1[62572] = 32'b00000000000000010010011110011101;
assign LUT_1[62573] = 32'b00000000000000001011110000011001;
assign LUT_1[62574] = 32'b00000000000000001110001100101110;
assign LUT_1[62575] = 32'b00000000000000000111011110101010;
assign LUT_1[62576] = 32'b00000000000000001101010010110011;
assign LUT_1[62577] = 32'b00000000000000000110100100101111;
assign LUT_1[62578] = 32'b00000000000000001001000001000100;
assign LUT_1[62579] = 32'b00000000000000000010010011000000;
assign LUT_1[62580] = 32'b00000000000000010101001100001010;
assign LUT_1[62581] = 32'b00000000000000001110011110000110;
assign LUT_1[62582] = 32'b00000000000000010000111010011011;
assign LUT_1[62583] = 32'b00000000000000001010001100010111;
assign LUT_1[62584] = 32'b00000000000000001100100000101000;
assign LUT_1[62585] = 32'b00000000000000000101110010100100;
assign LUT_1[62586] = 32'b00000000000000001000001110111001;
assign LUT_1[62587] = 32'b00000000000000000001100000110101;
assign LUT_1[62588] = 32'b00000000000000010100011001111111;
assign LUT_1[62589] = 32'b00000000000000001101101011111011;
assign LUT_1[62590] = 32'b00000000000000010000001000010000;
assign LUT_1[62591] = 32'b00000000000000001001011010001100;
assign LUT_1[62592] = 32'b00000000000000001011011110101101;
assign LUT_1[62593] = 32'b00000000000000000100110000101001;
assign LUT_1[62594] = 32'b00000000000000000111001100111110;
assign LUT_1[62595] = 32'b00000000000000000000011110111010;
assign LUT_1[62596] = 32'b00000000000000010011011000000100;
assign LUT_1[62597] = 32'b00000000000000001100101010000000;
assign LUT_1[62598] = 32'b00000000000000001111000110010101;
assign LUT_1[62599] = 32'b00000000000000001000011000010001;
assign LUT_1[62600] = 32'b00000000000000001010101100100010;
assign LUT_1[62601] = 32'b00000000000000000011111110011110;
assign LUT_1[62602] = 32'b00000000000000000110011010110011;
assign LUT_1[62603] = 32'b11111111111111111111101100101111;
assign LUT_1[62604] = 32'b00000000000000010010100101111001;
assign LUT_1[62605] = 32'b00000000000000001011110111110101;
assign LUT_1[62606] = 32'b00000000000000001110010100001010;
assign LUT_1[62607] = 32'b00000000000000000111100110000110;
assign LUT_1[62608] = 32'b00000000000000001101011010001111;
assign LUT_1[62609] = 32'b00000000000000000110101100001011;
assign LUT_1[62610] = 32'b00000000000000001001001000100000;
assign LUT_1[62611] = 32'b00000000000000000010011010011100;
assign LUT_1[62612] = 32'b00000000000000010101010011100110;
assign LUT_1[62613] = 32'b00000000000000001110100101100010;
assign LUT_1[62614] = 32'b00000000000000010001000001110111;
assign LUT_1[62615] = 32'b00000000000000001010010011110011;
assign LUT_1[62616] = 32'b00000000000000001100101000000100;
assign LUT_1[62617] = 32'b00000000000000000101111010000000;
assign LUT_1[62618] = 32'b00000000000000001000010110010101;
assign LUT_1[62619] = 32'b00000000000000000001101000010001;
assign LUT_1[62620] = 32'b00000000000000010100100001011011;
assign LUT_1[62621] = 32'b00000000000000001101110011010111;
assign LUT_1[62622] = 32'b00000000000000010000001111101100;
assign LUT_1[62623] = 32'b00000000000000001001100001101000;
assign LUT_1[62624] = 32'b00000000000000001100011001101100;
assign LUT_1[62625] = 32'b00000000000000000101101011101000;
assign LUT_1[62626] = 32'b00000000000000001000000111111101;
assign LUT_1[62627] = 32'b00000000000000000001011001111001;
assign LUT_1[62628] = 32'b00000000000000010100010011000011;
assign LUT_1[62629] = 32'b00000000000000001101100100111111;
assign LUT_1[62630] = 32'b00000000000000010000000001010100;
assign LUT_1[62631] = 32'b00000000000000001001010011010000;
assign LUT_1[62632] = 32'b00000000000000001011100111100001;
assign LUT_1[62633] = 32'b00000000000000000100111001011101;
assign LUT_1[62634] = 32'b00000000000000000111010101110010;
assign LUT_1[62635] = 32'b00000000000000000000100111101110;
assign LUT_1[62636] = 32'b00000000000000010011100000111000;
assign LUT_1[62637] = 32'b00000000000000001100110010110100;
assign LUT_1[62638] = 32'b00000000000000001111001111001001;
assign LUT_1[62639] = 32'b00000000000000001000100001000101;
assign LUT_1[62640] = 32'b00000000000000001110010101001110;
assign LUT_1[62641] = 32'b00000000000000000111100111001010;
assign LUT_1[62642] = 32'b00000000000000001010000011011111;
assign LUT_1[62643] = 32'b00000000000000000011010101011011;
assign LUT_1[62644] = 32'b00000000000000010110001110100101;
assign LUT_1[62645] = 32'b00000000000000001111100000100001;
assign LUT_1[62646] = 32'b00000000000000010001111100110110;
assign LUT_1[62647] = 32'b00000000000000001011001110110010;
assign LUT_1[62648] = 32'b00000000000000001101100011000011;
assign LUT_1[62649] = 32'b00000000000000000110110100111111;
assign LUT_1[62650] = 32'b00000000000000001001010001010100;
assign LUT_1[62651] = 32'b00000000000000000010100011010000;
assign LUT_1[62652] = 32'b00000000000000010101011100011010;
assign LUT_1[62653] = 32'b00000000000000001110101110010110;
assign LUT_1[62654] = 32'b00000000000000010001001010101011;
assign LUT_1[62655] = 32'b00000000000000001010011100100111;
assign LUT_1[62656] = 32'b00000000000000001101011100010101;
assign LUT_1[62657] = 32'b00000000000000000110101110010001;
assign LUT_1[62658] = 32'b00000000000000001001001010100110;
assign LUT_1[62659] = 32'b00000000000000000010011100100010;
assign LUT_1[62660] = 32'b00000000000000010101010101101100;
assign LUT_1[62661] = 32'b00000000000000001110100111101000;
assign LUT_1[62662] = 32'b00000000000000010001000011111101;
assign LUT_1[62663] = 32'b00000000000000001010010101111001;
assign LUT_1[62664] = 32'b00000000000000001100101010001010;
assign LUT_1[62665] = 32'b00000000000000000101111100000110;
assign LUT_1[62666] = 32'b00000000000000001000011000011011;
assign LUT_1[62667] = 32'b00000000000000000001101010010111;
assign LUT_1[62668] = 32'b00000000000000010100100011100001;
assign LUT_1[62669] = 32'b00000000000000001101110101011101;
assign LUT_1[62670] = 32'b00000000000000010000010001110010;
assign LUT_1[62671] = 32'b00000000000000001001100011101110;
assign LUT_1[62672] = 32'b00000000000000001111010111110111;
assign LUT_1[62673] = 32'b00000000000000001000101001110011;
assign LUT_1[62674] = 32'b00000000000000001011000110001000;
assign LUT_1[62675] = 32'b00000000000000000100011000000100;
assign LUT_1[62676] = 32'b00000000000000010111010001001110;
assign LUT_1[62677] = 32'b00000000000000010000100011001010;
assign LUT_1[62678] = 32'b00000000000000010010111111011111;
assign LUT_1[62679] = 32'b00000000000000001100010001011011;
assign LUT_1[62680] = 32'b00000000000000001110100101101100;
assign LUT_1[62681] = 32'b00000000000000000111110111101000;
assign LUT_1[62682] = 32'b00000000000000001010010011111101;
assign LUT_1[62683] = 32'b00000000000000000011100101111001;
assign LUT_1[62684] = 32'b00000000000000010110011111000011;
assign LUT_1[62685] = 32'b00000000000000001111110000111111;
assign LUT_1[62686] = 32'b00000000000000010010001101010100;
assign LUT_1[62687] = 32'b00000000000000001011011111010000;
assign LUT_1[62688] = 32'b00000000000000001110010111010100;
assign LUT_1[62689] = 32'b00000000000000000111101001010000;
assign LUT_1[62690] = 32'b00000000000000001010000101100101;
assign LUT_1[62691] = 32'b00000000000000000011010111100001;
assign LUT_1[62692] = 32'b00000000000000010110010000101011;
assign LUT_1[62693] = 32'b00000000000000001111100010100111;
assign LUT_1[62694] = 32'b00000000000000010001111110111100;
assign LUT_1[62695] = 32'b00000000000000001011010000111000;
assign LUT_1[62696] = 32'b00000000000000001101100101001001;
assign LUT_1[62697] = 32'b00000000000000000110110111000101;
assign LUT_1[62698] = 32'b00000000000000001001010011011010;
assign LUT_1[62699] = 32'b00000000000000000010100101010110;
assign LUT_1[62700] = 32'b00000000000000010101011110100000;
assign LUT_1[62701] = 32'b00000000000000001110110000011100;
assign LUT_1[62702] = 32'b00000000000000010001001100110001;
assign LUT_1[62703] = 32'b00000000000000001010011110101101;
assign LUT_1[62704] = 32'b00000000000000010000010010110110;
assign LUT_1[62705] = 32'b00000000000000001001100100110010;
assign LUT_1[62706] = 32'b00000000000000001100000001000111;
assign LUT_1[62707] = 32'b00000000000000000101010011000011;
assign LUT_1[62708] = 32'b00000000000000011000001100001101;
assign LUT_1[62709] = 32'b00000000000000010001011110001001;
assign LUT_1[62710] = 32'b00000000000000010011111010011110;
assign LUT_1[62711] = 32'b00000000000000001101001100011010;
assign LUT_1[62712] = 32'b00000000000000001111100000101011;
assign LUT_1[62713] = 32'b00000000000000001000110010100111;
assign LUT_1[62714] = 32'b00000000000000001011001110111100;
assign LUT_1[62715] = 32'b00000000000000000100100000111000;
assign LUT_1[62716] = 32'b00000000000000010111011010000010;
assign LUT_1[62717] = 32'b00000000000000010000101011111110;
assign LUT_1[62718] = 32'b00000000000000010011001000010011;
assign LUT_1[62719] = 32'b00000000000000001100011010001111;
assign LUT_1[62720] = 32'b00000000000000000110010010110110;
assign LUT_1[62721] = 32'b11111111111111111111100100110010;
assign LUT_1[62722] = 32'b00000000000000000010000001000111;
assign LUT_1[62723] = 32'b11111111111111111011010011000011;
assign LUT_1[62724] = 32'b00000000000000001110001100001101;
assign LUT_1[62725] = 32'b00000000000000000111011110001001;
assign LUT_1[62726] = 32'b00000000000000001001111010011110;
assign LUT_1[62727] = 32'b00000000000000000011001100011010;
assign LUT_1[62728] = 32'b00000000000000000101100000101011;
assign LUT_1[62729] = 32'b11111111111111111110110010100111;
assign LUT_1[62730] = 32'b00000000000000000001001110111100;
assign LUT_1[62731] = 32'b11111111111111111010100000111000;
assign LUT_1[62732] = 32'b00000000000000001101011010000010;
assign LUT_1[62733] = 32'b00000000000000000110101011111110;
assign LUT_1[62734] = 32'b00000000000000001001001000010011;
assign LUT_1[62735] = 32'b00000000000000000010011010001111;
assign LUT_1[62736] = 32'b00000000000000001000001110011000;
assign LUT_1[62737] = 32'b00000000000000000001100000010100;
assign LUT_1[62738] = 32'b00000000000000000011111100101001;
assign LUT_1[62739] = 32'b11111111111111111101001110100101;
assign LUT_1[62740] = 32'b00000000000000010000000111101111;
assign LUT_1[62741] = 32'b00000000000000001001011001101011;
assign LUT_1[62742] = 32'b00000000000000001011110110000000;
assign LUT_1[62743] = 32'b00000000000000000101000111111100;
assign LUT_1[62744] = 32'b00000000000000000111011100001101;
assign LUT_1[62745] = 32'b00000000000000000000101110001001;
assign LUT_1[62746] = 32'b00000000000000000011001010011110;
assign LUT_1[62747] = 32'b11111111111111111100011100011010;
assign LUT_1[62748] = 32'b00000000000000001111010101100100;
assign LUT_1[62749] = 32'b00000000000000001000100111100000;
assign LUT_1[62750] = 32'b00000000000000001011000011110101;
assign LUT_1[62751] = 32'b00000000000000000100010101110001;
assign LUT_1[62752] = 32'b00000000000000000111001101110101;
assign LUT_1[62753] = 32'b00000000000000000000011111110001;
assign LUT_1[62754] = 32'b00000000000000000010111100000110;
assign LUT_1[62755] = 32'b11111111111111111100001110000010;
assign LUT_1[62756] = 32'b00000000000000001111000111001100;
assign LUT_1[62757] = 32'b00000000000000001000011001001000;
assign LUT_1[62758] = 32'b00000000000000001010110101011101;
assign LUT_1[62759] = 32'b00000000000000000100000111011001;
assign LUT_1[62760] = 32'b00000000000000000110011011101010;
assign LUT_1[62761] = 32'b11111111111111111111101101100110;
assign LUT_1[62762] = 32'b00000000000000000010001001111011;
assign LUT_1[62763] = 32'b11111111111111111011011011110111;
assign LUT_1[62764] = 32'b00000000000000001110010101000001;
assign LUT_1[62765] = 32'b00000000000000000111100110111101;
assign LUT_1[62766] = 32'b00000000000000001010000011010010;
assign LUT_1[62767] = 32'b00000000000000000011010101001110;
assign LUT_1[62768] = 32'b00000000000000001001001001010111;
assign LUT_1[62769] = 32'b00000000000000000010011011010011;
assign LUT_1[62770] = 32'b00000000000000000100110111101000;
assign LUT_1[62771] = 32'b11111111111111111110001001100100;
assign LUT_1[62772] = 32'b00000000000000010001000010101110;
assign LUT_1[62773] = 32'b00000000000000001010010100101010;
assign LUT_1[62774] = 32'b00000000000000001100110000111111;
assign LUT_1[62775] = 32'b00000000000000000110000010111011;
assign LUT_1[62776] = 32'b00000000000000001000010111001100;
assign LUT_1[62777] = 32'b00000000000000000001101001001000;
assign LUT_1[62778] = 32'b00000000000000000100000101011101;
assign LUT_1[62779] = 32'b11111111111111111101010111011001;
assign LUT_1[62780] = 32'b00000000000000010000010000100011;
assign LUT_1[62781] = 32'b00000000000000001001100010011111;
assign LUT_1[62782] = 32'b00000000000000001011111110110100;
assign LUT_1[62783] = 32'b00000000000000000101010000110000;
assign LUT_1[62784] = 32'b00000000000000001000010000011110;
assign LUT_1[62785] = 32'b00000000000000000001100010011010;
assign LUT_1[62786] = 32'b00000000000000000011111110101111;
assign LUT_1[62787] = 32'b11111111111111111101010000101011;
assign LUT_1[62788] = 32'b00000000000000010000001001110101;
assign LUT_1[62789] = 32'b00000000000000001001011011110001;
assign LUT_1[62790] = 32'b00000000000000001011111000000110;
assign LUT_1[62791] = 32'b00000000000000000101001010000010;
assign LUT_1[62792] = 32'b00000000000000000111011110010011;
assign LUT_1[62793] = 32'b00000000000000000000110000001111;
assign LUT_1[62794] = 32'b00000000000000000011001100100100;
assign LUT_1[62795] = 32'b11111111111111111100011110100000;
assign LUT_1[62796] = 32'b00000000000000001111010111101010;
assign LUT_1[62797] = 32'b00000000000000001000101001100110;
assign LUT_1[62798] = 32'b00000000000000001011000101111011;
assign LUT_1[62799] = 32'b00000000000000000100010111110111;
assign LUT_1[62800] = 32'b00000000000000001010001100000000;
assign LUT_1[62801] = 32'b00000000000000000011011101111100;
assign LUT_1[62802] = 32'b00000000000000000101111010010001;
assign LUT_1[62803] = 32'b11111111111111111111001100001101;
assign LUT_1[62804] = 32'b00000000000000010010000101010111;
assign LUT_1[62805] = 32'b00000000000000001011010111010011;
assign LUT_1[62806] = 32'b00000000000000001101110011101000;
assign LUT_1[62807] = 32'b00000000000000000111000101100100;
assign LUT_1[62808] = 32'b00000000000000001001011001110101;
assign LUT_1[62809] = 32'b00000000000000000010101011110001;
assign LUT_1[62810] = 32'b00000000000000000101001000000110;
assign LUT_1[62811] = 32'b11111111111111111110011010000010;
assign LUT_1[62812] = 32'b00000000000000010001010011001100;
assign LUT_1[62813] = 32'b00000000000000001010100101001000;
assign LUT_1[62814] = 32'b00000000000000001101000001011101;
assign LUT_1[62815] = 32'b00000000000000000110010011011001;
assign LUT_1[62816] = 32'b00000000000000001001001011011101;
assign LUT_1[62817] = 32'b00000000000000000010011101011001;
assign LUT_1[62818] = 32'b00000000000000000100111001101110;
assign LUT_1[62819] = 32'b11111111111111111110001011101010;
assign LUT_1[62820] = 32'b00000000000000010001000100110100;
assign LUT_1[62821] = 32'b00000000000000001010010110110000;
assign LUT_1[62822] = 32'b00000000000000001100110011000101;
assign LUT_1[62823] = 32'b00000000000000000110000101000001;
assign LUT_1[62824] = 32'b00000000000000001000011001010010;
assign LUT_1[62825] = 32'b00000000000000000001101011001110;
assign LUT_1[62826] = 32'b00000000000000000100000111100011;
assign LUT_1[62827] = 32'b11111111111111111101011001011111;
assign LUT_1[62828] = 32'b00000000000000010000010010101001;
assign LUT_1[62829] = 32'b00000000000000001001100100100101;
assign LUT_1[62830] = 32'b00000000000000001100000000111010;
assign LUT_1[62831] = 32'b00000000000000000101010010110110;
assign LUT_1[62832] = 32'b00000000000000001011000110111111;
assign LUT_1[62833] = 32'b00000000000000000100011000111011;
assign LUT_1[62834] = 32'b00000000000000000110110101010000;
assign LUT_1[62835] = 32'b00000000000000000000000111001100;
assign LUT_1[62836] = 32'b00000000000000010011000000010110;
assign LUT_1[62837] = 32'b00000000000000001100010010010010;
assign LUT_1[62838] = 32'b00000000000000001110101110100111;
assign LUT_1[62839] = 32'b00000000000000001000000000100011;
assign LUT_1[62840] = 32'b00000000000000001010010100110100;
assign LUT_1[62841] = 32'b00000000000000000011100110110000;
assign LUT_1[62842] = 32'b00000000000000000110000011000101;
assign LUT_1[62843] = 32'b11111111111111111111010101000001;
assign LUT_1[62844] = 32'b00000000000000010010001110001011;
assign LUT_1[62845] = 32'b00000000000000001011100000000111;
assign LUT_1[62846] = 32'b00000000000000001101111100011100;
assign LUT_1[62847] = 32'b00000000000000000111001110011000;
assign LUT_1[62848] = 32'b00000000000000001001010010111001;
assign LUT_1[62849] = 32'b00000000000000000010100100110101;
assign LUT_1[62850] = 32'b00000000000000000101000001001010;
assign LUT_1[62851] = 32'b11111111111111111110010011000110;
assign LUT_1[62852] = 32'b00000000000000010001001100010000;
assign LUT_1[62853] = 32'b00000000000000001010011110001100;
assign LUT_1[62854] = 32'b00000000000000001100111010100001;
assign LUT_1[62855] = 32'b00000000000000000110001100011101;
assign LUT_1[62856] = 32'b00000000000000001000100000101110;
assign LUT_1[62857] = 32'b00000000000000000001110010101010;
assign LUT_1[62858] = 32'b00000000000000000100001110111111;
assign LUT_1[62859] = 32'b11111111111111111101100000111011;
assign LUT_1[62860] = 32'b00000000000000010000011010000101;
assign LUT_1[62861] = 32'b00000000000000001001101100000001;
assign LUT_1[62862] = 32'b00000000000000001100001000010110;
assign LUT_1[62863] = 32'b00000000000000000101011010010010;
assign LUT_1[62864] = 32'b00000000000000001011001110011011;
assign LUT_1[62865] = 32'b00000000000000000100100000010111;
assign LUT_1[62866] = 32'b00000000000000000110111100101100;
assign LUT_1[62867] = 32'b00000000000000000000001110101000;
assign LUT_1[62868] = 32'b00000000000000010011000111110010;
assign LUT_1[62869] = 32'b00000000000000001100011001101110;
assign LUT_1[62870] = 32'b00000000000000001110110110000011;
assign LUT_1[62871] = 32'b00000000000000001000000111111111;
assign LUT_1[62872] = 32'b00000000000000001010011100010000;
assign LUT_1[62873] = 32'b00000000000000000011101110001100;
assign LUT_1[62874] = 32'b00000000000000000110001010100001;
assign LUT_1[62875] = 32'b11111111111111111111011100011101;
assign LUT_1[62876] = 32'b00000000000000010010010101100111;
assign LUT_1[62877] = 32'b00000000000000001011100111100011;
assign LUT_1[62878] = 32'b00000000000000001110000011111000;
assign LUT_1[62879] = 32'b00000000000000000111010101110100;
assign LUT_1[62880] = 32'b00000000000000001010001101111000;
assign LUT_1[62881] = 32'b00000000000000000011011111110100;
assign LUT_1[62882] = 32'b00000000000000000101111100001001;
assign LUT_1[62883] = 32'b11111111111111111111001110000101;
assign LUT_1[62884] = 32'b00000000000000010010000111001111;
assign LUT_1[62885] = 32'b00000000000000001011011001001011;
assign LUT_1[62886] = 32'b00000000000000001101110101100000;
assign LUT_1[62887] = 32'b00000000000000000111000111011100;
assign LUT_1[62888] = 32'b00000000000000001001011011101101;
assign LUT_1[62889] = 32'b00000000000000000010101101101001;
assign LUT_1[62890] = 32'b00000000000000000101001001111110;
assign LUT_1[62891] = 32'b11111111111111111110011011111010;
assign LUT_1[62892] = 32'b00000000000000010001010101000100;
assign LUT_1[62893] = 32'b00000000000000001010100111000000;
assign LUT_1[62894] = 32'b00000000000000001101000011010101;
assign LUT_1[62895] = 32'b00000000000000000110010101010001;
assign LUT_1[62896] = 32'b00000000000000001100001001011010;
assign LUT_1[62897] = 32'b00000000000000000101011011010110;
assign LUT_1[62898] = 32'b00000000000000000111110111101011;
assign LUT_1[62899] = 32'b00000000000000000001001001100111;
assign LUT_1[62900] = 32'b00000000000000010100000010110001;
assign LUT_1[62901] = 32'b00000000000000001101010100101101;
assign LUT_1[62902] = 32'b00000000000000001111110001000010;
assign LUT_1[62903] = 32'b00000000000000001001000010111110;
assign LUT_1[62904] = 32'b00000000000000001011010111001111;
assign LUT_1[62905] = 32'b00000000000000000100101001001011;
assign LUT_1[62906] = 32'b00000000000000000111000101100000;
assign LUT_1[62907] = 32'b00000000000000000000010111011100;
assign LUT_1[62908] = 32'b00000000000000010011010000100110;
assign LUT_1[62909] = 32'b00000000000000001100100010100010;
assign LUT_1[62910] = 32'b00000000000000001110111110110111;
assign LUT_1[62911] = 32'b00000000000000001000010000110011;
assign LUT_1[62912] = 32'b00000000000000001011010000100001;
assign LUT_1[62913] = 32'b00000000000000000100100010011101;
assign LUT_1[62914] = 32'b00000000000000000110111110110010;
assign LUT_1[62915] = 32'b00000000000000000000010000101110;
assign LUT_1[62916] = 32'b00000000000000010011001001111000;
assign LUT_1[62917] = 32'b00000000000000001100011011110100;
assign LUT_1[62918] = 32'b00000000000000001110111000001001;
assign LUT_1[62919] = 32'b00000000000000001000001010000101;
assign LUT_1[62920] = 32'b00000000000000001010011110010110;
assign LUT_1[62921] = 32'b00000000000000000011110000010010;
assign LUT_1[62922] = 32'b00000000000000000110001100100111;
assign LUT_1[62923] = 32'b11111111111111111111011110100011;
assign LUT_1[62924] = 32'b00000000000000010010010111101101;
assign LUT_1[62925] = 32'b00000000000000001011101001101001;
assign LUT_1[62926] = 32'b00000000000000001110000101111110;
assign LUT_1[62927] = 32'b00000000000000000111010111111010;
assign LUT_1[62928] = 32'b00000000000000001101001100000011;
assign LUT_1[62929] = 32'b00000000000000000110011101111111;
assign LUT_1[62930] = 32'b00000000000000001000111010010100;
assign LUT_1[62931] = 32'b00000000000000000010001100010000;
assign LUT_1[62932] = 32'b00000000000000010101000101011010;
assign LUT_1[62933] = 32'b00000000000000001110010111010110;
assign LUT_1[62934] = 32'b00000000000000010000110011101011;
assign LUT_1[62935] = 32'b00000000000000001010000101100111;
assign LUT_1[62936] = 32'b00000000000000001100011001111000;
assign LUT_1[62937] = 32'b00000000000000000101101011110100;
assign LUT_1[62938] = 32'b00000000000000001000001000001001;
assign LUT_1[62939] = 32'b00000000000000000001011010000101;
assign LUT_1[62940] = 32'b00000000000000010100010011001111;
assign LUT_1[62941] = 32'b00000000000000001101100101001011;
assign LUT_1[62942] = 32'b00000000000000010000000001100000;
assign LUT_1[62943] = 32'b00000000000000001001010011011100;
assign LUT_1[62944] = 32'b00000000000000001100001011100000;
assign LUT_1[62945] = 32'b00000000000000000101011101011100;
assign LUT_1[62946] = 32'b00000000000000000111111001110001;
assign LUT_1[62947] = 32'b00000000000000000001001011101101;
assign LUT_1[62948] = 32'b00000000000000010100000100110111;
assign LUT_1[62949] = 32'b00000000000000001101010110110011;
assign LUT_1[62950] = 32'b00000000000000001111110011001000;
assign LUT_1[62951] = 32'b00000000000000001001000101000100;
assign LUT_1[62952] = 32'b00000000000000001011011001010101;
assign LUT_1[62953] = 32'b00000000000000000100101011010001;
assign LUT_1[62954] = 32'b00000000000000000111000111100110;
assign LUT_1[62955] = 32'b00000000000000000000011001100010;
assign LUT_1[62956] = 32'b00000000000000010011010010101100;
assign LUT_1[62957] = 32'b00000000000000001100100100101000;
assign LUT_1[62958] = 32'b00000000000000001111000000111101;
assign LUT_1[62959] = 32'b00000000000000001000010010111001;
assign LUT_1[62960] = 32'b00000000000000001110000111000010;
assign LUT_1[62961] = 32'b00000000000000000111011000111110;
assign LUT_1[62962] = 32'b00000000000000001001110101010011;
assign LUT_1[62963] = 32'b00000000000000000011000111001111;
assign LUT_1[62964] = 32'b00000000000000010110000000011001;
assign LUT_1[62965] = 32'b00000000000000001111010010010101;
assign LUT_1[62966] = 32'b00000000000000010001101110101010;
assign LUT_1[62967] = 32'b00000000000000001011000000100110;
assign LUT_1[62968] = 32'b00000000000000001101010100110111;
assign LUT_1[62969] = 32'b00000000000000000110100110110011;
assign LUT_1[62970] = 32'b00000000000000001001000011001000;
assign LUT_1[62971] = 32'b00000000000000000010010101000100;
assign LUT_1[62972] = 32'b00000000000000010101001110001110;
assign LUT_1[62973] = 32'b00000000000000001110100000001010;
assign LUT_1[62974] = 32'b00000000000000010000111100011111;
assign LUT_1[62975] = 32'b00000000000000001010001110011011;
assign LUT_1[62976] = 32'b00000000000000000010001101000111;
assign LUT_1[62977] = 32'b11111111111111111011011111000011;
assign LUT_1[62978] = 32'b11111111111111111101111011011000;
assign LUT_1[62979] = 32'b11111111111111110111001101010100;
assign LUT_1[62980] = 32'b00000000000000001010000110011110;
assign LUT_1[62981] = 32'b00000000000000000011011000011010;
assign LUT_1[62982] = 32'b00000000000000000101110100101111;
assign LUT_1[62983] = 32'b11111111111111111111000110101011;
assign LUT_1[62984] = 32'b00000000000000000001011010111100;
assign LUT_1[62985] = 32'b11111111111111111010101100111000;
assign LUT_1[62986] = 32'b11111111111111111101001001001101;
assign LUT_1[62987] = 32'b11111111111111110110011011001001;
assign LUT_1[62988] = 32'b00000000000000001001010100010011;
assign LUT_1[62989] = 32'b00000000000000000010100110001111;
assign LUT_1[62990] = 32'b00000000000000000101000010100100;
assign LUT_1[62991] = 32'b11111111111111111110010100100000;
assign LUT_1[62992] = 32'b00000000000000000100001000101001;
assign LUT_1[62993] = 32'b11111111111111111101011010100101;
assign LUT_1[62994] = 32'b11111111111111111111110110111010;
assign LUT_1[62995] = 32'b11111111111111111001001000110110;
assign LUT_1[62996] = 32'b00000000000000001100000010000000;
assign LUT_1[62997] = 32'b00000000000000000101010011111100;
assign LUT_1[62998] = 32'b00000000000000000111110000010001;
assign LUT_1[62999] = 32'b00000000000000000001000010001101;
assign LUT_1[63000] = 32'b00000000000000000011010110011110;
assign LUT_1[63001] = 32'b11111111111111111100101000011010;
assign LUT_1[63002] = 32'b11111111111111111111000100101111;
assign LUT_1[63003] = 32'b11111111111111111000010110101011;
assign LUT_1[63004] = 32'b00000000000000001011001111110101;
assign LUT_1[63005] = 32'b00000000000000000100100001110001;
assign LUT_1[63006] = 32'b00000000000000000110111110000110;
assign LUT_1[63007] = 32'b00000000000000000000010000000010;
assign LUT_1[63008] = 32'b00000000000000000011001000000110;
assign LUT_1[63009] = 32'b11111111111111111100011010000010;
assign LUT_1[63010] = 32'b11111111111111111110110110010111;
assign LUT_1[63011] = 32'b11111111111111111000001000010011;
assign LUT_1[63012] = 32'b00000000000000001011000001011101;
assign LUT_1[63013] = 32'b00000000000000000100010011011001;
assign LUT_1[63014] = 32'b00000000000000000110101111101110;
assign LUT_1[63015] = 32'b00000000000000000000000001101010;
assign LUT_1[63016] = 32'b00000000000000000010010101111011;
assign LUT_1[63017] = 32'b11111111111111111011100111110111;
assign LUT_1[63018] = 32'b11111111111111111110000100001100;
assign LUT_1[63019] = 32'b11111111111111110111010110001000;
assign LUT_1[63020] = 32'b00000000000000001010001111010010;
assign LUT_1[63021] = 32'b00000000000000000011100001001110;
assign LUT_1[63022] = 32'b00000000000000000101111101100011;
assign LUT_1[63023] = 32'b11111111111111111111001111011111;
assign LUT_1[63024] = 32'b00000000000000000101000011101000;
assign LUT_1[63025] = 32'b11111111111111111110010101100100;
assign LUT_1[63026] = 32'b00000000000000000000110001111001;
assign LUT_1[63027] = 32'b11111111111111111010000011110101;
assign LUT_1[63028] = 32'b00000000000000001100111100111111;
assign LUT_1[63029] = 32'b00000000000000000110001110111011;
assign LUT_1[63030] = 32'b00000000000000001000101011010000;
assign LUT_1[63031] = 32'b00000000000000000001111101001100;
assign LUT_1[63032] = 32'b00000000000000000100010001011101;
assign LUT_1[63033] = 32'b11111111111111111101100011011001;
assign LUT_1[63034] = 32'b11111111111111111111111111101110;
assign LUT_1[63035] = 32'b11111111111111111001010001101010;
assign LUT_1[63036] = 32'b00000000000000001100001010110100;
assign LUT_1[63037] = 32'b00000000000000000101011100110000;
assign LUT_1[63038] = 32'b00000000000000000111111001000101;
assign LUT_1[63039] = 32'b00000000000000000001001011000001;
assign LUT_1[63040] = 32'b00000000000000000100001010101111;
assign LUT_1[63041] = 32'b11111111111111111101011100101011;
assign LUT_1[63042] = 32'b11111111111111111111111001000000;
assign LUT_1[63043] = 32'b11111111111111111001001010111100;
assign LUT_1[63044] = 32'b00000000000000001100000100000110;
assign LUT_1[63045] = 32'b00000000000000000101010110000010;
assign LUT_1[63046] = 32'b00000000000000000111110010010111;
assign LUT_1[63047] = 32'b00000000000000000001000100010011;
assign LUT_1[63048] = 32'b00000000000000000011011000100100;
assign LUT_1[63049] = 32'b11111111111111111100101010100000;
assign LUT_1[63050] = 32'b11111111111111111111000110110101;
assign LUT_1[63051] = 32'b11111111111111111000011000110001;
assign LUT_1[63052] = 32'b00000000000000001011010001111011;
assign LUT_1[63053] = 32'b00000000000000000100100011110111;
assign LUT_1[63054] = 32'b00000000000000000111000000001100;
assign LUT_1[63055] = 32'b00000000000000000000010010001000;
assign LUT_1[63056] = 32'b00000000000000000110000110010001;
assign LUT_1[63057] = 32'b11111111111111111111011000001101;
assign LUT_1[63058] = 32'b00000000000000000001110100100010;
assign LUT_1[63059] = 32'b11111111111111111011000110011110;
assign LUT_1[63060] = 32'b00000000000000001101111111101000;
assign LUT_1[63061] = 32'b00000000000000000111010001100100;
assign LUT_1[63062] = 32'b00000000000000001001101101111001;
assign LUT_1[63063] = 32'b00000000000000000010111111110101;
assign LUT_1[63064] = 32'b00000000000000000101010100000110;
assign LUT_1[63065] = 32'b11111111111111111110100110000010;
assign LUT_1[63066] = 32'b00000000000000000001000010010111;
assign LUT_1[63067] = 32'b11111111111111111010010100010011;
assign LUT_1[63068] = 32'b00000000000000001101001101011101;
assign LUT_1[63069] = 32'b00000000000000000110011111011001;
assign LUT_1[63070] = 32'b00000000000000001000111011101110;
assign LUT_1[63071] = 32'b00000000000000000010001101101010;
assign LUT_1[63072] = 32'b00000000000000000101000101101110;
assign LUT_1[63073] = 32'b11111111111111111110010111101010;
assign LUT_1[63074] = 32'b00000000000000000000110011111111;
assign LUT_1[63075] = 32'b11111111111111111010000101111011;
assign LUT_1[63076] = 32'b00000000000000001100111111000101;
assign LUT_1[63077] = 32'b00000000000000000110010001000001;
assign LUT_1[63078] = 32'b00000000000000001000101101010110;
assign LUT_1[63079] = 32'b00000000000000000001111111010010;
assign LUT_1[63080] = 32'b00000000000000000100010011100011;
assign LUT_1[63081] = 32'b11111111111111111101100101011111;
assign LUT_1[63082] = 32'b00000000000000000000000001110100;
assign LUT_1[63083] = 32'b11111111111111111001010011110000;
assign LUT_1[63084] = 32'b00000000000000001100001100111010;
assign LUT_1[63085] = 32'b00000000000000000101011110110110;
assign LUT_1[63086] = 32'b00000000000000000111111011001011;
assign LUT_1[63087] = 32'b00000000000000000001001101000111;
assign LUT_1[63088] = 32'b00000000000000000111000001010000;
assign LUT_1[63089] = 32'b00000000000000000000010011001100;
assign LUT_1[63090] = 32'b00000000000000000010101111100001;
assign LUT_1[63091] = 32'b11111111111111111100000001011101;
assign LUT_1[63092] = 32'b00000000000000001110111010100111;
assign LUT_1[63093] = 32'b00000000000000001000001100100011;
assign LUT_1[63094] = 32'b00000000000000001010101000111000;
assign LUT_1[63095] = 32'b00000000000000000011111010110100;
assign LUT_1[63096] = 32'b00000000000000000110001111000101;
assign LUT_1[63097] = 32'b11111111111111111111100001000001;
assign LUT_1[63098] = 32'b00000000000000000001111101010110;
assign LUT_1[63099] = 32'b11111111111111111011001111010010;
assign LUT_1[63100] = 32'b00000000000000001110001000011100;
assign LUT_1[63101] = 32'b00000000000000000111011010011000;
assign LUT_1[63102] = 32'b00000000000000001001110110101101;
assign LUT_1[63103] = 32'b00000000000000000011001000101001;
assign LUT_1[63104] = 32'b00000000000000000101001101001010;
assign LUT_1[63105] = 32'b11111111111111111110011111000110;
assign LUT_1[63106] = 32'b00000000000000000000111011011011;
assign LUT_1[63107] = 32'b11111111111111111010001101010111;
assign LUT_1[63108] = 32'b00000000000000001101000110100001;
assign LUT_1[63109] = 32'b00000000000000000110011000011101;
assign LUT_1[63110] = 32'b00000000000000001000110100110010;
assign LUT_1[63111] = 32'b00000000000000000010000110101110;
assign LUT_1[63112] = 32'b00000000000000000100011010111111;
assign LUT_1[63113] = 32'b11111111111111111101101100111011;
assign LUT_1[63114] = 32'b00000000000000000000001001010000;
assign LUT_1[63115] = 32'b11111111111111111001011011001100;
assign LUT_1[63116] = 32'b00000000000000001100010100010110;
assign LUT_1[63117] = 32'b00000000000000000101100110010010;
assign LUT_1[63118] = 32'b00000000000000001000000010100111;
assign LUT_1[63119] = 32'b00000000000000000001010100100011;
assign LUT_1[63120] = 32'b00000000000000000111001000101100;
assign LUT_1[63121] = 32'b00000000000000000000011010101000;
assign LUT_1[63122] = 32'b00000000000000000010110110111101;
assign LUT_1[63123] = 32'b11111111111111111100001000111001;
assign LUT_1[63124] = 32'b00000000000000001111000010000011;
assign LUT_1[63125] = 32'b00000000000000001000010011111111;
assign LUT_1[63126] = 32'b00000000000000001010110000010100;
assign LUT_1[63127] = 32'b00000000000000000100000010010000;
assign LUT_1[63128] = 32'b00000000000000000110010110100001;
assign LUT_1[63129] = 32'b11111111111111111111101000011101;
assign LUT_1[63130] = 32'b00000000000000000010000100110010;
assign LUT_1[63131] = 32'b11111111111111111011010110101110;
assign LUT_1[63132] = 32'b00000000000000001110001111111000;
assign LUT_1[63133] = 32'b00000000000000000111100001110100;
assign LUT_1[63134] = 32'b00000000000000001001111110001001;
assign LUT_1[63135] = 32'b00000000000000000011010000000101;
assign LUT_1[63136] = 32'b00000000000000000110001000001001;
assign LUT_1[63137] = 32'b11111111111111111111011010000101;
assign LUT_1[63138] = 32'b00000000000000000001110110011010;
assign LUT_1[63139] = 32'b11111111111111111011001000010110;
assign LUT_1[63140] = 32'b00000000000000001110000001100000;
assign LUT_1[63141] = 32'b00000000000000000111010011011100;
assign LUT_1[63142] = 32'b00000000000000001001101111110001;
assign LUT_1[63143] = 32'b00000000000000000011000001101101;
assign LUT_1[63144] = 32'b00000000000000000101010101111110;
assign LUT_1[63145] = 32'b11111111111111111110100111111010;
assign LUT_1[63146] = 32'b00000000000000000001000100001111;
assign LUT_1[63147] = 32'b11111111111111111010010110001011;
assign LUT_1[63148] = 32'b00000000000000001101001111010101;
assign LUT_1[63149] = 32'b00000000000000000110100001010001;
assign LUT_1[63150] = 32'b00000000000000001000111101100110;
assign LUT_1[63151] = 32'b00000000000000000010001111100010;
assign LUT_1[63152] = 32'b00000000000000001000000011101011;
assign LUT_1[63153] = 32'b00000000000000000001010101100111;
assign LUT_1[63154] = 32'b00000000000000000011110001111100;
assign LUT_1[63155] = 32'b11111111111111111101000011111000;
assign LUT_1[63156] = 32'b00000000000000001111111101000010;
assign LUT_1[63157] = 32'b00000000000000001001001110111110;
assign LUT_1[63158] = 32'b00000000000000001011101011010011;
assign LUT_1[63159] = 32'b00000000000000000100111101001111;
assign LUT_1[63160] = 32'b00000000000000000111010001100000;
assign LUT_1[63161] = 32'b00000000000000000000100011011100;
assign LUT_1[63162] = 32'b00000000000000000010111111110001;
assign LUT_1[63163] = 32'b11111111111111111100010001101101;
assign LUT_1[63164] = 32'b00000000000000001111001010110111;
assign LUT_1[63165] = 32'b00000000000000001000011100110011;
assign LUT_1[63166] = 32'b00000000000000001010111001001000;
assign LUT_1[63167] = 32'b00000000000000000100001011000100;
assign LUT_1[63168] = 32'b00000000000000000111001010110010;
assign LUT_1[63169] = 32'b00000000000000000000011100101110;
assign LUT_1[63170] = 32'b00000000000000000010111001000011;
assign LUT_1[63171] = 32'b11111111111111111100001010111111;
assign LUT_1[63172] = 32'b00000000000000001111000100001001;
assign LUT_1[63173] = 32'b00000000000000001000010110000101;
assign LUT_1[63174] = 32'b00000000000000001010110010011010;
assign LUT_1[63175] = 32'b00000000000000000100000100010110;
assign LUT_1[63176] = 32'b00000000000000000110011000100111;
assign LUT_1[63177] = 32'b11111111111111111111101010100011;
assign LUT_1[63178] = 32'b00000000000000000010000110111000;
assign LUT_1[63179] = 32'b11111111111111111011011000110100;
assign LUT_1[63180] = 32'b00000000000000001110010001111110;
assign LUT_1[63181] = 32'b00000000000000000111100011111010;
assign LUT_1[63182] = 32'b00000000000000001010000000001111;
assign LUT_1[63183] = 32'b00000000000000000011010010001011;
assign LUT_1[63184] = 32'b00000000000000001001000110010100;
assign LUT_1[63185] = 32'b00000000000000000010011000010000;
assign LUT_1[63186] = 32'b00000000000000000100110100100101;
assign LUT_1[63187] = 32'b11111111111111111110000110100001;
assign LUT_1[63188] = 32'b00000000000000010000111111101011;
assign LUT_1[63189] = 32'b00000000000000001010010001100111;
assign LUT_1[63190] = 32'b00000000000000001100101101111100;
assign LUT_1[63191] = 32'b00000000000000000101111111111000;
assign LUT_1[63192] = 32'b00000000000000001000010100001001;
assign LUT_1[63193] = 32'b00000000000000000001100110000101;
assign LUT_1[63194] = 32'b00000000000000000100000010011010;
assign LUT_1[63195] = 32'b11111111111111111101010100010110;
assign LUT_1[63196] = 32'b00000000000000010000001101100000;
assign LUT_1[63197] = 32'b00000000000000001001011111011100;
assign LUT_1[63198] = 32'b00000000000000001011111011110001;
assign LUT_1[63199] = 32'b00000000000000000101001101101101;
assign LUT_1[63200] = 32'b00000000000000001000000101110001;
assign LUT_1[63201] = 32'b00000000000000000001010111101101;
assign LUT_1[63202] = 32'b00000000000000000011110100000010;
assign LUT_1[63203] = 32'b11111111111111111101000101111110;
assign LUT_1[63204] = 32'b00000000000000001111111111001000;
assign LUT_1[63205] = 32'b00000000000000001001010001000100;
assign LUT_1[63206] = 32'b00000000000000001011101101011001;
assign LUT_1[63207] = 32'b00000000000000000100111111010101;
assign LUT_1[63208] = 32'b00000000000000000111010011100110;
assign LUT_1[63209] = 32'b00000000000000000000100101100010;
assign LUT_1[63210] = 32'b00000000000000000011000001110111;
assign LUT_1[63211] = 32'b11111111111111111100010011110011;
assign LUT_1[63212] = 32'b00000000000000001111001100111101;
assign LUT_1[63213] = 32'b00000000000000001000011110111001;
assign LUT_1[63214] = 32'b00000000000000001010111011001110;
assign LUT_1[63215] = 32'b00000000000000000100001101001010;
assign LUT_1[63216] = 32'b00000000000000001010000001010011;
assign LUT_1[63217] = 32'b00000000000000000011010011001111;
assign LUT_1[63218] = 32'b00000000000000000101101111100100;
assign LUT_1[63219] = 32'b11111111111111111111000001100000;
assign LUT_1[63220] = 32'b00000000000000010001111010101010;
assign LUT_1[63221] = 32'b00000000000000001011001100100110;
assign LUT_1[63222] = 32'b00000000000000001101101000111011;
assign LUT_1[63223] = 32'b00000000000000000110111010110111;
assign LUT_1[63224] = 32'b00000000000000001001001111001000;
assign LUT_1[63225] = 32'b00000000000000000010100001000100;
assign LUT_1[63226] = 32'b00000000000000000100111101011001;
assign LUT_1[63227] = 32'b11111111111111111110001111010101;
assign LUT_1[63228] = 32'b00000000000000010001001000011111;
assign LUT_1[63229] = 32'b00000000000000001010011010011011;
assign LUT_1[63230] = 32'b00000000000000001100110110110000;
assign LUT_1[63231] = 32'b00000000000000000110001000101100;
assign LUT_1[63232] = 32'b00000000000000000000000001010011;
assign LUT_1[63233] = 32'b11111111111111111001010011001111;
assign LUT_1[63234] = 32'b11111111111111111011101111100100;
assign LUT_1[63235] = 32'b11111111111111110101000001100000;
assign LUT_1[63236] = 32'b00000000000000000111111010101010;
assign LUT_1[63237] = 32'b00000000000000000001001100100110;
assign LUT_1[63238] = 32'b00000000000000000011101000111011;
assign LUT_1[63239] = 32'b11111111111111111100111010110111;
assign LUT_1[63240] = 32'b11111111111111111111001111001000;
assign LUT_1[63241] = 32'b11111111111111111000100001000100;
assign LUT_1[63242] = 32'b11111111111111111010111101011001;
assign LUT_1[63243] = 32'b11111111111111110100001111010101;
assign LUT_1[63244] = 32'b00000000000000000111001000011111;
assign LUT_1[63245] = 32'b00000000000000000000011010011011;
assign LUT_1[63246] = 32'b00000000000000000010110110110000;
assign LUT_1[63247] = 32'b11111111111111111100001000101100;
assign LUT_1[63248] = 32'b00000000000000000001111100110101;
assign LUT_1[63249] = 32'b11111111111111111011001110110001;
assign LUT_1[63250] = 32'b11111111111111111101101011000110;
assign LUT_1[63251] = 32'b11111111111111110110111101000010;
assign LUT_1[63252] = 32'b00000000000000001001110110001100;
assign LUT_1[63253] = 32'b00000000000000000011001000001000;
assign LUT_1[63254] = 32'b00000000000000000101100100011101;
assign LUT_1[63255] = 32'b11111111111111111110110110011001;
assign LUT_1[63256] = 32'b00000000000000000001001010101010;
assign LUT_1[63257] = 32'b11111111111111111010011100100110;
assign LUT_1[63258] = 32'b11111111111111111100111000111011;
assign LUT_1[63259] = 32'b11111111111111110110001010110111;
assign LUT_1[63260] = 32'b00000000000000001001000100000001;
assign LUT_1[63261] = 32'b00000000000000000010010101111101;
assign LUT_1[63262] = 32'b00000000000000000100110010010010;
assign LUT_1[63263] = 32'b11111111111111111110000100001110;
assign LUT_1[63264] = 32'b00000000000000000000111100010010;
assign LUT_1[63265] = 32'b11111111111111111010001110001110;
assign LUT_1[63266] = 32'b11111111111111111100101010100011;
assign LUT_1[63267] = 32'b11111111111111110101111100011111;
assign LUT_1[63268] = 32'b00000000000000001000110101101001;
assign LUT_1[63269] = 32'b00000000000000000010000111100101;
assign LUT_1[63270] = 32'b00000000000000000100100011111010;
assign LUT_1[63271] = 32'b11111111111111111101110101110110;
assign LUT_1[63272] = 32'b00000000000000000000001010000111;
assign LUT_1[63273] = 32'b11111111111111111001011100000011;
assign LUT_1[63274] = 32'b11111111111111111011111000011000;
assign LUT_1[63275] = 32'b11111111111111110101001010010100;
assign LUT_1[63276] = 32'b00000000000000001000000011011110;
assign LUT_1[63277] = 32'b00000000000000000001010101011010;
assign LUT_1[63278] = 32'b00000000000000000011110001101111;
assign LUT_1[63279] = 32'b11111111111111111101000011101011;
assign LUT_1[63280] = 32'b00000000000000000010110111110100;
assign LUT_1[63281] = 32'b11111111111111111100001001110000;
assign LUT_1[63282] = 32'b11111111111111111110100110000101;
assign LUT_1[63283] = 32'b11111111111111110111111000000001;
assign LUT_1[63284] = 32'b00000000000000001010110001001011;
assign LUT_1[63285] = 32'b00000000000000000100000011000111;
assign LUT_1[63286] = 32'b00000000000000000110011111011100;
assign LUT_1[63287] = 32'b11111111111111111111110001011000;
assign LUT_1[63288] = 32'b00000000000000000010000101101001;
assign LUT_1[63289] = 32'b11111111111111111011010111100101;
assign LUT_1[63290] = 32'b11111111111111111101110011111010;
assign LUT_1[63291] = 32'b11111111111111110111000101110110;
assign LUT_1[63292] = 32'b00000000000000001001111111000000;
assign LUT_1[63293] = 32'b00000000000000000011010000111100;
assign LUT_1[63294] = 32'b00000000000000000101101101010001;
assign LUT_1[63295] = 32'b11111111111111111110111111001101;
assign LUT_1[63296] = 32'b00000000000000000001111110111011;
assign LUT_1[63297] = 32'b11111111111111111011010000110111;
assign LUT_1[63298] = 32'b11111111111111111101101101001100;
assign LUT_1[63299] = 32'b11111111111111110110111111001000;
assign LUT_1[63300] = 32'b00000000000000001001111000010010;
assign LUT_1[63301] = 32'b00000000000000000011001010001110;
assign LUT_1[63302] = 32'b00000000000000000101100110100011;
assign LUT_1[63303] = 32'b11111111111111111110111000011111;
assign LUT_1[63304] = 32'b00000000000000000001001100110000;
assign LUT_1[63305] = 32'b11111111111111111010011110101100;
assign LUT_1[63306] = 32'b11111111111111111100111011000001;
assign LUT_1[63307] = 32'b11111111111111110110001100111101;
assign LUT_1[63308] = 32'b00000000000000001001000110000111;
assign LUT_1[63309] = 32'b00000000000000000010011000000011;
assign LUT_1[63310] = 32'b00000000000000000100110100011000;
assign LUT_1[63311] = 32'b11111111111111111110000110010100;
assign LUT_1[63312] = 32'b00000000000000000011111010011101;
assign LUT_1[63313] = 32'b11111111111111111101001100011001;
assign LUT_1[63314] = 32'b11111111111111111111101000101110;
assign LUT_1[63315] = 32'b11111111111111111000111010101010;
assign LUT_1[63316] = 32'b00000000000000001011110011110100;
assign LUT_1[63317] = 32'b00000000000000000101000101110000;
assign LUT_1[63318] = 32'b00000000000000000111100010000101;
assign LUT_1[63319] = 32'b00000000000000000000110100000001;
assign LUT_1[63320] = 32'b00000000000000000011001000010010;
assign LUT_1[63321] = 32'b11111111111111111100011010001110;
assign LUT_1[63322] = 32'b11111111111111111110110110100011;
assign LUT_1[63323] = 32'b11111111111111111000001000011111;
assign LUT_1[63324] = 32'b00000000000000001011000001101001;
assign LUT_1[63325] = 32'b00000000000000000100010011100101;
assign LUT_1[63326] = 32'b00000000000000000110101111111010;
assign LUT_1[63327] = 32'b00000000000000000000000001110110;
assign LUT_1[63328] = 32'b00000000000000000010111001111010;
assign LUT_1[63329] = 32'b11111111111111111100001011110110;
assign LUT_1[63330] = 32'b11111111111111111110101000001011;
assign LUT_1[63331] = 32'b11111111111111110111111010000111;
assign LUT_1[63332] = 32'b00000000000000001010110011010001;
assign LUT_1[63333] = 32'b00000000000000000100000101001101;
assign LUT_1[63334] = 32'b00000000000000000110100001100010;
assign LUT_1[63335] = 32'b11111111111111111111110011011110;
assign LUT_1[63336] = 32'b00000000000000000010000111101111;
assign LUT_1[63337] = 32'b11111111111111111011011001101011;
assign LUT_1[63338] = 32'b11111111111111111101110110000000;
assign LUT_1[63339] = 32'b11111111111111110111000111111100;
assign LUT_1[63340] = 32'b00000000000000001010000001000110;
assign LUT_1[63341] = 32'b00000000000000000011010011000010;
assign LUT_1[63342] = 32'b00000000000000000101101111010111;
assign LUT_1[63343] = 32'b11111111111111111111000001010011;
assign LUT_1[63344] = 32'b00000000000000000100110101011100;
assign LUT_1[63345] = 32'b11111111111111111110000111011000;
assign LUT_1[63346] = 32'b00000000000000000000100011101101;
assign LUT_1[63347] = 32'b11111111111111111001110101101001;
assign LUT_1[63348] = 32'b00000000000000001100101110110011;
assign LUT_1[63349] = 32'b00000000000000000110000000101111;
assign LUT_1[63350] = 32'b00000000000000001000011101000100;
assign LUT_1[63351] = 32'b00000000000000000001101111000000;
assign LUT_1[63352] = 32'b00000000000000000100000011010001;
assign LUT_1[63353] = 32'b11111111111111111101010101001101;
assign LUT_1[63354] = 32'b11111111111111111111110001100010;
assign LUT_1[63355] = 32'b11111111111111111001000011011110;
assign LUT_1[63356] = 32'b00000000000000001011111100101000;
assign LUT_1[63357] = 32'b00000000000000000101001110100100;
assign LUT_1[63358] = 32'b00000000000000000111101010111001;
assign LUT_1[63359] = 32'b00000000000000000000111100110101;
assign LUT_1[63360] = 32'b00000000000000000011000001010110;
assign LUT_1[63361] = 32'b11111111111111111100010011010010;
assign LUT_1[63362] = 32'b11111111111111111110101111100111;
assign LUT_1[63363] = 32'b11111111111111111000000001100011;
assign LUT_1[63364] = 32'b00000000000000001010111010101101;
assign LUT_1[63365] = 32'b00000000000000000100001100101001;
assign LUT_1[63366] = 32'b00000000000000000110101000111110;
assign LUT_1[63367] = 32'b11111111111111111111111010111010;
assign LUT_1[63368] = 32'b00000000000000000010001111001011;
assign LUT_1[63369] = 32'b11111111111111111011100001000111;
assign LUT_1[63370] = 32'b11111111111111111101111101011100;
assign LUT_1[63371] = 32'b11111111111111110111001111011000;
assign LUT_1[63372] = 32'b00000000000000001010001000100010;
assign LUT_1[63373] = 32'b00000000000000000011011010011110;
assign LUT_1[63374] = 32'b00000000000000000101110110110011;
assign LUT_1[63375] = 32'b11111111111111111111001000101111;
assign LUT_1[63376] = 32'b00000000000000000100111100111000;
assign LUT_1[63377] = 32'b11111111111111111110001110110100;
assign LUT_1[63378] = 32'b00000000000000000000101011001001;
assign LUT_1[63379] = 32'b11111111111111111001111101000101;
assign LUT_1[63380] = 32'b00000000000000001100110110001111;
assign LUT_1[63381] = 32'b00000000000000000110001000001011;
assign LUT_1[63382] = 32'b00000000000000001000100100100000;
assign LUT_1[63383] = 32'b00000000000000000001110110011100;
assign LUT_1[63384] = 32'b00000000000000000100001010101101;
assign LUT_1[63385] = 32'b11111111111111111101011100101001;
assign LUT_1[63386] = 32'b11111111111111111111111000111110;
assign LUT_1[63387] = 32'b11111111111111111001001010111010;
assign LUT_1[63388] = 32'b00000000000000001100000100000100;
assign LUT_1[63389] = 32'b00000000000000000101010110000000;
assign LUT_1[63390] = 32'b00000000000000000111110010010101;
assign LUT_1[63391] = 32'b00000000000000000001000100010001;
assign LUT_1[63392] = 32'b00000000000000000011111100010101;
assign LUT_1[63393] = 32'b11111111111111111101001110010001;
assign LUT_1[63394] = 32'b11111111111111111111101010100110;
assign LUT_1[63395] = 32'b11111111111111111000111100100010;
assign LUT_1[63396] = 32'b00000000000000001011110101101100;
assign LUT_1[63397] = 32'b00000000000000000101000111101000;
assign LUT_1[63398] = 32'b00000000000000000111100011111101;
assign LUT_1[63399] = 32'b00000000000000000000110101111001;
assign LUT_1[63400] = 32'b00000000000000000011001010001010;
assign LUT_1[63401] = 32'b11111111111111111100011100000110;
assign LUT_1[63402] = 32'b11111111111111111110111000011011;
assign LUT_1[63403] = 32'b11111111111111111000001010010111;
assign LUT_1[63404] = 32'b00000000000000001011000011100001;
assign LUT_1[63405] = 32'b00000000000000000100010101011101;
assign LUT_1[63406] = 32'b00000000000000000110110001110010;
assign LUT_1[63407] = 32'b00000000000000000000000011101110;
assign LUT_1[63408] = 32'b00000000000000000101110111110111;
assign LUT_1[63409] = 32'b11111111111111111111001001110011;
assign LUT_1[63410] = 32'b00000000000000000001100110001000;
assign LUT_1[63411] = 32'b11111111111111111010111000000100;
assign LUT_1[63412] = 32'b00000000000000001101110001001110;
assign LUT_1[63413] = 32'b00000000000000000111000011001010;
assign LUT_1[63414] = 32'b00000000000000001001011111011111;
assign LUT_1[63415] = 32'b00000000000000000010110001011011;
assign LUT_1[63416] = 32'b00000000000000000101000101101100;
assign LUT_1[63417] = 32'b11111111111111111110010111101000;
assign LUT_1[63418] = 32'b00000000000000000000110011111101;
assign LUT_1[63419] = 32'b11111111111111111010000101111001;
assign LUT_1[63420] = 32'b00000000000000001100111111000011;
assign LUT_1[63421] = 32'b00000000000000000110010000111111;
assign LUT_1[63422] = 32'b00000000000000001000101101010100;
assign LUT_1[63423] = 32'b00000000000000000001111111010000;
assign LUT_1[63424] = 32'b00000000000000000100111110111110;
assign LUT_1[63425] = 32'b11111111111111111110010000111010;
assign LUT_1[63426] = 32'b00000000000000000000101101001111;
assign LUT_1[63427] = 32'b11111111111111111001111111001011;
assign LUT_1[63428] = 32'b00000000000000001100111000010101;
assign LUT_1[63429] = 32'b00000000000000000110001010010001;
assign LUT_1[63430] = 32'b00000000000000001000100110100110;
assign LUT_1[63431] = 32'b00000000000000000001111000100010;
assign LUT_1[63432] = 32'b00000000000000000100001100110011;
assign LUT_1[63433] = 32'b11111111111111111101011110101111;
assign LUT_1[63434] = 32'b11111111111111111111111011000100;
assign LUT_1[63435] = 32'b11111111111111111001001101000000;
assign LUT_1[63436] = 32'b00000000000000001100000110001010;
assign LUT_1[63437] = 32'b00000000000000000101011000000110;
assign LUT_1[63438] = 32'b00000000000000000111110100011011;
assign LUT_1[63439] = 32'b00000000000000000001000110010111;
assign LUT_1[63440] = 32'b00000000000000000110111010100000;
assign LUT_1[63441] = 32'b00000000000000000000001100011100;
assign LUT_1[63442] = 32'b00000000000000000010101000110001;
assign LUT_1[63443] = 32'b11111111111111111011111010101101;
assign LUT_1[63444] = 32'b00000000000000001110110011110111;
assign LUT_1[63445] = 32'b00000000000000001000000101110011;
assign LUT_1[63446] = 32'b00000000000000001010100010001000;
assign LUT_1[63447] = 32'b00000000000000000011110100000100;
assign LUT_1[63448] = 32'b00000000000000000110001000010101;
assign LUT_1[63449] = 32'b11111111111111111111011010010001;
assign LUT_1[63450] = 32'b00000000000000000001110110100110;
assign LUT_1[63451] = 32'b11111111111111111011001000100010;
assign LUT_1[63452] = 32'b00000000000000001110000001101100;
assign LUT_1[63453] = 32'b00000000000000000111010011101000;
assign LUT_1[63454] = 32'b00000000000000001001101111111101;
assign LUT_1[63455] = 32'b00000000000000000011000001111001;
assign LUT_1[63456] = 32'b00000000000000000101111001111101;
assign LUT_1[63457] = 32'b11111111111111111111001011111001;
assign LUT_1[63458] = 32'b00000000000000000001101000001110;
assign LUT_1[63459] = 32'b11111111111111111010111010001010;
assign LUT_1[63460] = 32'b00000000000000001101110011010100;
assign LUT_1[63461] = 32'b00000000000000000111000101010000;
assign LUT_1[63462] = 32'b00000000000000001001100001100101;
assign LUT_1[63463] = 32'b00000000000000000010110011100001;
assign LUT_1[63464] = 32'b00000000000000000101000111110010;
assign LUT_1[63465] = 32'b11111111111111111110011001101110;
assign LUT_1[63466] = 32'b00000000000000000000110110000011;
assign LUT_1[63467] = 32'b11111111111111111010000111111111;
assign LUT_1[63468] = 32'b00000000000000001101000001001001;
assign LUT_1[63469] = 32'b00000000000000000110010011000101;
assign LUT_1[63470] = 32'b00000000000000001000101111011010;
assign LUT_1[63471] = 32'b00000000000000000010000001010110;
assign LUT_1[63472] = 32'b00000000000000000111110101011111;
assign LUT_1[63473] = 32'b00000000000000000001000111011011;
assign LUT_1[63474] = 32'b00000000000000000011100011110000;
assign LUT_1[63475] = 32'b11111111111111111100110101101100;
assign LUT_1[63476] = 32'b00000000000000001111101110110110;
assign LUT_1[63477] = 32'b00000000000000001001000000110010;
assign LUT_1[63478] = 32'b00000000000000001011011101000111;
assign LUT_1[63479] = 32'b00000000000000000100101111000011;
assign LUT_1[63480] = 32'b00000000000000000111000011010100;
assign LUT_1[63481] = 32'b00000000000000000000010101010000;
assign LUT_1[63482] = 32'b00000000000000000010110001100101;
assign LUT_1[63483] = 32'b11111111111111111100000011100001;
assign LUT_1[63484] = 32'b00000000000000001110111100101011;
assign LUT_1[63485] = 32'b00000000000000001000001110100111;
assign LUT_1[63486] = 32'b00000000000000001010101010111100;
assign LUT_1[63487] = 32'b00000000000000000011111100111000;
assign LUT_1[63488] = 32'b00000000000000000011001001110101;
assign LUT_1[63489] = 32'b11111111111111111100011011110001;
assign LUT_1[63490] = 32'b11111111111111111110111000000110;
assign LUT_1[63491] = 32'b11111111111111111000001010000010;
assign LUT_1[63492] = 32'b00000000000000001011000011001100;
assign LUT_1[63493] = 32'b00000000000000000100010101001000;
assign LUT_1[63494] = 32'b00000000000000000110110001011101;
assign LUT_1[63495] = 32'b00000000000000000000000011011001;
assign LUT_1[63496] = 32'b00000000000000000010010111101010;
assign LUT_1[63497] = 32'b11111111111111111011101001100110;
assign LUT_1[63498] = 32'b11111111111111111110000101111011;
assign LUT_1[63499] = 32'b11111111111111110111010111110111;
assign LUT_1[63500] = 32'b00000000000000001010010001000001;
assign LUT_1[63501] = 32'b00000000000000000011100010111101;
assign LUT_1[63502] = 32'b00000000000000000101111111010010;
assign LUT_1[63503] = 32'b11111111111111111111010001001110;
assign LUT_1[63504] = 32'b00000000000000000101000101010111;
assign LUT_1[63505] = 32'b11111111111111111110010111010011;
assign LUT_1[63506] = 32'b00000000000000000000110011101000;
assign LUT_1[63507] = 32'b11111111111111111010000101100100;
assign LUT_1[63508] = 32'b00000000000000001100111110101110;
assign LUT_1[63509] = 32'b00000000000000000110010000101010;
assign LUT_1[63510] = 32'b00000000000000001000101100111111;
assign LUT_1[63511] = 32'b00000000000000000001111110111011;
assign LUT_1[63512] = 32'b00000000000000000100010011001100;
assign LUT_1[63513] = 32'b11111111111111111101100101001000;
assign LUT_1[63514] = 32'b00000000000000000000000001011101;
assign LUT_1[63515] = 32'b11111111111111111001010011011001;
assign LUT_1[63516] = 32'b00000000000000001100001100100011;
assign LUT_1[63517] = 32'b00000000000000000101011110011111;
assign LUT_1[63518] = 32'b00000000000000000111111010110100;
assign LUT_1[63519] = 32'b00000000000000000001001100110000;
assign LUT_1[63520] = 32'b00000000000000000100000100110100;
assign LUT_1[63521] = 32'b11111111111111111101010110110000;
assign LUT_1[63522] = 32'b11111111111111111111110011000101;
assign LUT_1[63523] = 32'b11111111111111111001000101000001;
assign LUT_1[63524] = 32'b00000000000000001011111110001011;
assign LUT_1[63525] = 32'b00000000000000000101010000000111;
assign LUT_1[63526] = 32'b00000000000000000111101100011100;
assign LUT_1[63527] = 32'b00000000000000000000111110011000;
assign LUT_1[63528] = 32'b00000000000000000011010010101001;
assign LUT_1[63529] = 32'b11111111111111111100100100100101;
assign LUT_1[63530] = 32'b11111111111111111111000000111010;
assign LUT_1[63531] = 32'b11111111111111111000010010110110;
assign LUT_1[63532] = 32'b00000000000000001011001100000000;
assign LUT_1[63533] = 32'b00000000000000000100011101111100;
assign LUT_1[63534] = 32'b00000000000000000110111010010001;
assign LUT_1[63535] = 32'b00000000000000000000001100001101;
assign LUT_1[63536] = 32'b00000000000000000110000000010110;
assign LUT_1[63537] = 32'b11111111111111111111010010010010;
assign LUT_1[63538] = 32'b00000000000000000001101110100111;
assign LUT_1[63539] = 32'b11111111111111111011000000100011;
assign LUT_1[63540] = 32'b00000000000000001101111001101101;
assign LUT_1[63541] = 32'b00000000000000000111001011101001;
assign LUT_1[63542] = 32'b00000000000000001001100111111110;
assign LUT_1[63543] = 32'b00000000000000000010111001111010;
assign LUT_1[63544] = 32'b00000000000000000101001110001011;
assign LUT_1[63545] = 32'b11111111111111111110100000000111;
assign LUT_1[63546] = 32'b00000000000000000000111100011100;
assign LUT_1[63547] = 32'b11111111111111111010001110011000;
assign LUT_1[63548] = 32'b00000000000000001101000111100010;
assign LUT_1[63549] = 32'b00000000000000000110011001011110;
assign LUT_1[63550] = 32'b00000000000000001000110101110011;
assign LUT_1[63551] = 32'b00000000000000000010000111101111;
assign LUT_1[63552] = 32'b00000000000000000101000111011101;
assign LUT_1[63553] = 32'b11111111111111111110011001011001;
assign LUT_1[63554] = 32'b00000000000000000000110101101110;
assign LUT_1[63555] = 32'b11111111111111111010000111101010;
assign LUT_1[63556] = 32'b00000000000000001101000000110100;
assign LUT_1[63557] = 32'b00000000000000000110010010110000;
assign LUT_1[63558] = 32'b00000000000000001000101111000101;
assign LUT_1[63559] = 32'b00000000000000000010000001000001;
assign LUT_1[63560] = 32'b00000000000000000100010101010010;
assign LUT_1[63561] = 32'b11111111111111111101100111001110;
assign LUT_1[63562] = 32'b00000000000000000000000011100011;
assign LUT_1[63563] = 32'b11111111111111111001010101011111;
assign LUT_1[63564] = 32'b00000000000000001100001110101001;
assign LUT_1[63565] = 32'b00000000000000000101100000100101;
assign LUT_1[63566] = 32'b00000000000000000111111100111010;
assign LUT_1[63567] = 32'b00000000000000000001001110110110;
assign LUT_1[63568] = 32'b00000000000000000111000010111111;
assign LUT_1[63569] = 32'b00000000000000000000010100111011;
assign LUT_1[63570] = 32'b00000000000000000010110001010000;
assign LUT_1[63571] = 32'b11111111111111111100000011001100;
assign LUT_1[63572] = 32'b00000000000000001110111100010110;
assign LUT_1[63573] = 32'b00000000000000001000001110010010;
assign LUT_1[63574] = 32'b00000000000000001010101010100111;
assign LUT_1[63575] = 32'b00000000000000000011111100100011;
assign LUT_1[63576] = 32'b00000000000000000110010000110100;
assign LUT_1[63577] = 32'b11111111111111111111100010110000;
assign LUT_1[63578] = 32'b00000000000000000001111111000101;
assign LUT_1[63579] = 32'b11111111111111111011010001000001;
assign LUT_1[63580] = 32'b00000000000000001110001010001011;
assign LUT_1[63581] = 32'b00000000000000000111011100000111;
assign LUT_1[63582] = 32'b00000000000000001001111000011100;
assign LUT_1[63583] = 32'b00000000000000000011001010011000;
assign LUT_1[63584] = 32'b00000000000000000110000010011100;
assign LUT_1[63585] = 32'b11111111111111111111010100011000;
assign LUT_1[63586] = 32'b00000000000000000001110000101101;
assign LUT_1[63587] = 32'b11111111111111111011000010101001;
assign LUT_1[63588] = 32'b00000000000000001101111011110011;
assign LUT_1[63589] = 32'b00000000000000000111001101101111;
assign LUT_1[63590] = 32'b00000000000000001001101010000100;
assign LUT_1[63591] = 32'b00000000000000000010111100000000;
assign LUT_1[63592] = 32'b00000000000000000101010000010001;
assign LUT_1[63593] = 32'b11111111111111111110100010001101;
assign LUT_1[63594] = 32'b00000000000000000000111110100010;
assign LUT_1[63595] = 32'b11111111111111111010010000011110;
assign LUT_1[63596] = 32'b00000000000000001101001001101000;
assign LUT_1[63597] = 32'b00000000000000000110011011100100;
assign LUT_1[63598] = 32'b00000000000000001000110111111001;
assign LUT_1[63599] = 32'b00000000000000000010001001110101;
assign LUT_1[63600] = 32'b00000000000000000111111101111110;
assign LUT_1[63601] = 32'b00000000000000000001001111111010;
assign LUT_1[63602] = 32'b00000000000000000011101100001111;
assign LUT_1[63603] = 32'b11111111111111111100111110001011;
assign LUT_1[63604] = 32'b00000000000000001111110111010101;
assign LUT_1[63605] = 32'b00000000000000001001001001010001;
assign LUT_1[63606] = 32'b00000000000000001011100101100110;
assign LUT_1[63607] = 32'b00000000000000000100110111100010;
assign LUT_1[63608] = 32'b00000000000000000111001011110011;
assign LUT_1[63609] = 32'b00000000000000000000011101101111;
assign LUT_1[63610] = 32'b00000000000000000010111010000100;
assign LUT_1[63611] = 32'b11111111111111111100001100000000;
assign LUT_1[63612] = 32'b00000000000000001111000101001010;
assign LUT_1[63613] = 32'b00000000000000001000010111000110;
assign LUT_1[63614] = 32'b00000000000000001010110011011011;
assign LUT_1[63615] = 32'b00000000000000000100000101010111;
assign LUT_1[63616] = 32'b00000000000000000110001001111000;
assign LUT_1[63617] = 32'b11111111111111111111011011110100;
assign LUT_1[63618] = 32'b00000000000000000001111000001001;
assign LUT_1[63619] = 32'b11111111111111111011001010000101;
assign LUT_1[63620] = 32'b00000000000000001110000011001111;
assign LUT_1[63621] = 32'b00000000000000000111010101001011;
assign LUT_1[63622] = 32'b00000000000000001001110001100000;
assign LUT_1[63623] = 32'b00000000000000000011000011011100;
assign LUT_1[63624] = 32'b00000000000000000101010111101101;
assign LUT_1[63625] = 32'b11111111111111111110101001101001;
assign LUT_1[63626] = 32'b00000000000000000001000101111110;
assign LUT_1[63627] = 32'b11111111111111111010010111111010;
assign LUT_1[63628] = 32'b00000000000000001101010001000100;
assign LUT_1[63629] = 32'b00000000000000000110100011000000;
assign LUT_1[63630] = 32'b00000000000000001000111111010101;
assign LUT_1[63631] = 32'b00000000000000000010010001010001;
assign LUT_1[63632] = 32'b00000000000000001000000101011010;
assign LUT_1[63633] = 32'b00000000000000000001010111010110;
assign LUT_1[63634] = 32'b00000000000000000011110011101011;
assign LUT_1[63635] = 32'b11111111111111111101000101100111;
assign LUT_1[63636] = 32'b00000000000000001111111110110001;
assign LUT_1[63637] = 32'b00000000000000001001010000101101;
assign LUT_1[63638] = 32'b00000000000000001011101101000010;
assign LUT_1[63639] = 32'b00000000000000000100111110111110;
assign LUT_1[63640] = 32'b00000000000000000111010011001111;
assign LUT_1[63641] = 32'b00000000000000000000100101001011;
assign LUT_1[63642] = 32'b00000000000000000011000001100000;
assign LUT_1[63643] = 32'b11111111111111111100010011011100;
assign LUT_1[63644] = 32'b00000000000000001111001100100110;
assign LUT_1[63645] = 32'b00000000000000001000011110100010;
assign LUT_1[63646] = 32'b00000000000000001010111010110111;
assign LUT_1[63647] = 32'b00000000000000000100001100110011;
assign LUT_1[63648] = 32'b00000000000000000111000100110111;
assign LUT_1[63649] = 32'b00000000000000000000010110110011;
assign LUT_1[63650] = 32'b00000000000000000010110011001000;
assign LUT_1[63651] = 32'b11111111111111111100000101000100;
assign LUT_1[63652] = 32'b00000000000000001110111110001110;
assign LUT_1[63653] = 32'b00000000000000001000010000001010;
assign LUT_1[63654] = 32'b00000000000000001010101100011111;
assign LUT_1[63655] = 32'b00000000000000000011111110011011;
assign LUT_1[63656] = 32'b00000000000000000110010010101100;
assign LUT_1[63657] = 32'b11111111111111111111100100101000;
assign LUT_1[63658] = 32'b00000000000000000010000000111101;
assign LUT_1[63659] = 32'b11111111111111111011010010111001;
assign LUT_1[63660] = 32'b00000000000000001110001100000011;
assign LUT_1[63661] = 32'b00000000000000000111011101111111;
assign LUT_1[63662] = 32'b00000000000000001001111010010100;
assign LUT_1[63663] = 32'b00000000000000000011001100010000;
assign LUT_1[63664] = 32'b00000000000000001001000000011001;
assign LUT_1[63665] = 32'b00000000000000000010010010010101;
assign LUT_1[63666] = 32'b00000000000000000100101110101010;
assign LUT_1[63667] = 32'b11111111111111111110000000100110;
assign LUT_1[63668] = 32'b00000000000000010000111001110000;
assign LUT_1[63669] = 32'b00000000000000001010001011101100;
assign LUT_1[63670] = 32'b00000000000000001100101000000001;
assign LUT_1[63671] = 32'b00000000000000000101111001111101;
assign LUT_1[63672] = 32'b00000000000000001000001110001110;
assign LUT_1[63673] = 32'b00000000000000000001100000001010;
assign LUT_1[63674] = 32'b00000000000000000011111100011111;
assign LUT_1[63675] = 32'b11111111111111111101001110011011;
assign LUT_1[63676] = 32'b00000000000000010000000111100101;
assign LUT_1[63677] = 32'b00000000000000001001011001100001;
assign LUT_1[63678] = 32'b00000000000000001011110101110110;
assign LUT_1[63679] = 32'b00000000000000000101000111110010;
assign LUT_1[63680] = 32'b00000000000000001000000111100000;
assign LUT_1[63681] = 32'b00000000000000000001011001011100;
assign LUT_1[63682] = 32'b00000000000000000011110101110001;
assign LUT_1[63683] = 32'b11111111111111111101000111101101;
assign LUT_1[63684] = 32'b00000000000000010000000000110111;
assign LUT_1[63685] = 32'b00000000000000001001010010110011;
assign LUT_1[63686] = 32'b00000000000000001011101111001000;
assign LUT_1[63687] = 32'b00000000000000000101000001000100;
assign LUT_1[63688] = 32'b00000000000000000111010101010101;
assign LUT_1[63689] = 32'b00000000000000000000100111010001;
assign LUT_1[63690] = 32'b00000000000000000011000011100110;
assign LUT_1[63691] = 32'b11111111111111111100010101100010;
assign LUT_1[63692] = 32'b00000000000000001111001110101100;
assign LUT_1[63693] = 32'b00000000000000001000100000101000;
assign LUT_1[63694] = 32'b00000000000000001010111100111101;
assign LUT_1[63695] = 32'b00000000000000000100001110111001;
assign LUT_1[63696] = 32'b00000000000000001010000011000010;
assign LUT_1[63697] = 32'b00000000000000000011010100111110;
assign LUT_1[63698] = 32'b00000000000000000101110001010011;
assign LUT_1[63699] = 32'b11111111111111111111000011001111;
assign LUT_1[63700] = 32'b00000000000000010001111100011001;
assign LUT_1[63701] = 32'b00000000000000001011001110010101;
assign LUT_1[63702] = 32'b00000000000000001101101010101010;
assign LUT_1[63703] = 32'b00000000000000000110111100100110;
assign LUT_1[63704] = 32'b00000000000000001001010000110111;
assign LUT_1[63705] = 32'b00000000000000000010100010110011;
assign LUT_1[63706] = 32'b00000000000000000100111111001000;
assign LUT_1[63707] = 32'b11111111111111111110010001000100;
assign LUT_1[63708] = 32'b00000000000000010001001010001110;
assign LUT_1[63709] = 32'b00000000000000001010011100001010;
assign LUT_1[63710] = 32'b00000000000000001100111000011111;
assign LUT_1[63711] = 32'b00000000000000000110001010011011;
assign LUT_1[63712] = 32'b00000000000000001001000010011111;
assign LUT_1[63713] = 32'b00000000000000000010010100011011;
assign LUT_1[63714] = 32'b00000000000000000100110000110000;
assign LUT_1[63715] = 32'b11111111111111111110000010101100;
assign LUT_1[63716] = 32'b00000000000000010000111011110110;
assign LUT_1[63717] = 32'b00000000000000001010001101110010;
assign LUT_1[63718] = 32'b00000000000000001100101010000111;
assign LUT_1[63719] = 32'b00000000000000000101111100000011;
assign LUT_1[63720] = 32'b00000000000000001000010000010100;
assign LUT_1[63721] = 32'b00000000000000000001100010010000;
assign LUT_1[63722] = 32'b00000000000000000011111110100101;
assign LUT_1[63723] = 32'b11111111111111111101010000100001;
assign LUT_1[63724] = 32'b00000000000000010000001001101011;
assign LUT_1[63725] = 32'b00000000000000001001011011100111;
assign LUT_1[63726] = 32'b00000000000000001011110111111100;
assign LUT_1[63727] = 32'b00000000000000000101001001111000;
assign LUT_1[63728] = 32'b00000000000000001010111110000001;
assign LUT_1[63729] = 32'b00000000000000000100001111111101;
assign LUT_1[63730] = 32'b00000000000000000110101100010010;
assign LUT_1[63731] = 32'b11111111111111111111111110001110;
assign LUT_1[63732] = 32'b00000000000000010010110111011000;
assign LUT_1[63733] = 32'b00000000000000001100001001010100;
assign LUT_1[63734] = 32'b00000000000000001110100101101001;
assign LUT_1[63735] = 32'b00000000000000000111110111100101;
assign LUT_1[63736] = 32'b00000000000000001010001011110110;
assign LUT_1[63737] = 32'b00000000000000000011011101110010;
assign LUT_1[63738] = 32'b00000000000000000101111010000111;
assign LUT_1[63739] = 32'b11111111111111111111001100000011;
assign LUT_1[63740] = 32'b00000000000000010010000101001101;
assign LUT_1[63741] = 32'b00000000000000001011010111001001;
assign LUT_1[63742] = 32'b00000000000000001101110011011110;
assign LUT_1[63743] = 32'b00000000000000000111000101011010;
assign LUT_1[63744] = 32'b00000000000000000000111110000001;
assign LUT_1[63745] = 32'b11111111111111111010001111111101;
assign LUT_1[63746] = 32'b11111111111111111100101100010010;
assign LUT_1[63747] = 32'b11111111111111110101111110001110;
assign LUT_1[63748] = 32'b00000000000000001000110111011000;
assign LUT_1[63749] = 32'b00000000000000000010001001010100;
assign LUT_1[63750] = 32'b00000000000000000100100101101001;
assign LUT_1[63751] = 32'b11111111111111111101110111100101;
assign LUT_1[63752] = 32'b00000000000000000000001011110110;
assign LUT_1[63753] = 32'b11111111111111111001011101110010;
assign LUT_1[63754] = 32'b11111111111111111011111010000111;
assign LUT_1[63755] = 32'b11111111111111110101001100000011;
assign LUT_1[63756] = 32'b00000000000000001000000101001101;
assign LUT_1[63757] = 32'b00000000000000000001010111001001;
assign LUT_1[63758] = 32'b00000000000000000011110011011110;
assign LUT_1[63759] = 32'b11111111111111111101000101011010;
assign LUT_1[63760] = 32'b00000000000000000010111001100011;
assign LUT_1[63761] = 32'b11111111111111111100001011011111;
assign LUT_1[63762] = 32'b11111111111111111110100111110100;
assign LUT_1[63763] = 32'b11111111111111110111111001110000;
assign LUT_1[63764] = 32'b00000000000000001010110010111010;
assign LUT_1[63765] = 32'b00000000000000000100000100110110;
assign LUT_1[63766] = 32'b00000000000000000110100001001011;
assign LUT_1[63767] = 32'b11111111111111111111110011000111;
assign LUT_1[63768] = 32'b00000000000000000010000111011000;
assign LUT_1[63769] = 32'b11111111111111111011011001010100;
assign LUT_1[63770] = 32'b11111111111111111101110101101001;
assign LUT_1[63771] = 32'b11111111111111110111000111100101;
assign LUT_1[63772] = 32'b00000000000000001010000000101111;
assign LUT_1[63773] = 32'b00000000000000000011010010101011;
assign LUT_1[63774] = 32'b00000000000000000101101111000000;
assign LUT_1[63775] = 32'b11111111111111111111000000111100;
assign LUT_1[63776] = 32'b00000000000000000001111001000000;
assign LUT_1[63777] = 32'b11111111111111111011001010111100;
assign LUT_1[63778] = 32'b11111111111111111101100111010001;
assign LUT_1[63779] = 32'b11111111111111110110111001001101;
assign LUT_1[63780] = 32'b00000000000000001001110010010111;
assign LUT_1[63781] = 32'b00000000000000000011000100010011;
assign LUT_1[63782] = 32'b00000000000000000101100000101000;
assign LUT_1[63783] = 32'b11111111111111111110110010100100;
assign LUT_1[63784] = 32'b00000000000000000001000110110101;
assign LUT_1[63785] = 32'b11111111111111111010011000110001;
assign LUT_1[63786] = 32'b11111111111111111100110101000110;
assign LUT_1[63787] = 32'b11111111111111110110000111000010;
assign LUT_1[63788] = 32'b00000000000000001001000000001100;
assign LUT_1[63789] = 32'b00000000000000000010010010001000;
assign LUT_1[63790] = 32'b00000000000000000100101110011101;
assign LUT_1[63791] = 32'b11111111111111111110000000011001;
assign LUT_1[63792] = 32'b00000000000000000011110100100010;
assign LUT_1[63793] = 32'b11111111111111111101000110011110;
assign LUT_1[63794] = 32'b11111111111111111111100010110011;
assign LUT_1[63795] = 32'b11111111111111111000110100101111;
assign LUT_1[63796] = 32'b00000000000000001011101101111001;
assign LUT_1[63797] = 32'b00000000000000000100111111110101;
assign LUT_1[63798] = 32'b00000000000000000111011100001010;
assign LUT_1[63799] = 32'b00000000000000000000101110000110;
assign LUT_1[63800] = 32'b00000000000000000011000010010111;
assign LUT_1[63801] = 32'b11111111111111111100010100010011;
assign LUT_1[63802] = 32'b11111111111111111110110000101000;
assign LUT_1[63803] = 32'b11111111111111111000000010100100;
assign LUT_1[63804] = 32'b00000000000000001010111011101110;
assign LUT_1[63805] = 32'b00000000000000000100001101101010;
assign LUT_1[63806] = 32'b00000000000000000110101001111111;
assign LUT_1[63807] = 32'b11111111111111111111111011111011;
assign LUT_1[63808] = 32'b00000000000000000010111011101001;
assign LUT_1[63809] = 32'b11111111111111111100001101100101;
assign LUT_1[63810] = 32'b11111111111111111110101001111010;
assign LUT_1[63811] = 32'b11111111111111110111111011110110;
assign LUT_1[63812] = 32'b00000000000000001010110101000000;
assign LUT_1[63813] = 32'b00000000000000000100000110111100;
assign LUT_1[63814] = 32'b00000000000000000110100011010001;
assign LUT_1[63815] = 32'b11111111111111111111110101001101;
assign LUT_1[63816] = 32'b00000000000000000010001001011110;
assign LUT_1[63817] = 32'b11111111111111111011011011011010;
assign LUT_1[63818] = 32'b11111111111111111101110111101111;
assign LUT_1[63819] = 32'b11111111111111110111001001101011;
assign LUT_1[63820] = 32'b00000000000000001010000010110101;
assign LUT_1[63821] = 32'b00000000000000000011010100110001;
assign LUT_1[63822] = 32'b00000000000000000101110001000110;
assign LUT_1[63823] = 32'b11111111111111111111000011000010;
assign LUT_1[63824] = 32'b00000000000000000100110111001011;
assign LUT_1[63825] = 32'b11111111111111111110001001000111;
assign LUT_1[63826] = 32'b00000000000000000000100101011100;
assign LUT_1[63827] = 32'b11111111111111111001110111011000;
assign LUT_1[63828] = 32'b00000000000000001100110000100010;
assign LUT_1[63829] = 32'b00000000000000000110000010011110;
assign LUT_1[63830] = 32'b00000000000000001000011110110011;
assign LUT_1[63831] = 32'b00000000000000000001110000101111;
assign LUT_1[63832] = 32'b00000000000000000100000101000000;
assign LUT_1[63833] = 32'b11111111111111111101010110111100;
assign LUT_1[63834] = 32'b11111111111111111111110011010001;
assign LUT_1[63835] = 32'b11111111111111111001000101001101;
assign LUT_1[63836] = 32'b00000000000000001011111110010111;
assign LUT_1[63837] = 32'b00000000000000000101010000010011;
assign LUT_1[63838] = 32'b00000000000000000111101100101000;
assign LUT_1[63839] = 32'b00000000000000000000111110100100;
assign LUT_1[63840] = 32'b00000000000000000011110110101000;
assign LUT_1[63841] = 32'b11111111111111111101001000100100;
assign LUT_1[63842] = 32'b11111111111111111111100100111001;
assign LUT_1[63843] = 32'b11111111111111111000110110110101;
assign LUT_1[63844] = 32'b00000000000000001011101111111111;
assign LUT_1[63845] = 32'b00000000000000000101000001111011;
assign LUT_1[63846] = 32'b00000000000000000111011110010000;
assign LUT_1[63847] = 32'b00000000000000000000110000001100;
assign LUT_1[63848] = 32'b00000000000000000011000100011101;
assign LUT_1[63849] = 32'b11111111111111111100010110011001;
assign LUT_1[63850] = 32'b11111111111111111110110010101110;
assign LUT_1[63851] = 32'b11111111111111111000000100101010;
assign LUT_1[63852] = 32'b00000000000000001010111101110100;
assign LUT_1[63853] = 32'b00000000000000000100001111110000;
assign LUT_1[63854] = 32'b00000000000000000110101100000101;
assign LUT_1[63855] = 32'b11111111111111111111111110000001;
assign LUT_1[63856] = 32'b00000000000000000101110010001010;
assign LUT_1[63857] = 32'b11111111111111111111000100000110;
assign LUT_1[63858] = 32'b00000000000000000001100000011011;
assign LUT_1[63859] = 32'b11111111111111111010110010010111;
assign LUT_1[63860] = 32'b00000000000000001101101011100001;
assign LUT_1[63861] = 32'b00000000000000000110111101011101;
assign LUT_1[63862] = 32'b00000000000000001001011001110010;
assign LUT_1[63863] = 32'b00000000000000000010101011101110;
assign LUT_1[63864] = 32'b00000000000000000100111111111111;
assign LUT_1[63865] = 32'b11111111111111111110010001111011;
assign LUT_1[63866] = 32'b00000000000000000000101110010000;
assign LUT_1[63867] = 32'b11111111111111111010000000001100;
assign LUT_1[63868] = 32'b00000000000000001100111001010110;
assign LUT_1[63869] = 32'b00000000000000000110001011010010;
assign LUT_1[63870] = 32'b00000000000000001000100111100111;
assign LUT_1[63871] = 32'b00000000000000000001111001100011;
assign LUT_1[63872] = 32'b00000000000000000011111110000100;
assign LUT_1[63873] = 32'b11111111111111111101010000000000;
assign LUT_1[63874] = 32'b11111111111111111111101100010101;
assign LUT_1[63875] = 32'b11111111111111111000111110010001;
assign LUT_1[63876] = 32'b00000000000000001011110111011011;
assign LUT_1[63877] = 32'b00000000000000000101001001010111;
assign LUT_1[63878] = 32'b00000000000000000111100101101100;
assign LUT_1[63879] = 32'b00000000000000000000110111101000;
assign LUT_1[63880] = 32'b00000000000000000011001011111001;
assign LUT_1[63881] = 32'b11111111111111111100011101110101;
assign LUT_1[63882] = 32'b11111111111111111110111010001010;
assign LUT_1[63883] = 32'b11111111111111111000001100000110;
assign LUT_1[63884] = 32'b00000000000000001011000101010000;
assign LUT_1[63885] = 32'b00000000000000000100010111001100;
assign LUT_1[63886] = 32'b00000000000000000110110011100001;
assign LUT_1[63887] = 32'b00000000000000000000000101011101;
assign LUT_1[63888] = 32'b00000000000000000101111001100110;
assign LUT_1[63889] = 32'b11111111111111111111001011100010;
assign LUT_1[63890] = 32'b00000000000000000001100111110111;
assign LUT_1[63891] = 32'b11111111111111111010111001110011;
assign LUT_1[63892] = 32'b00000000000000001101110010111101;
assign LUT_1[63893] = 32'b00000000000000000111000100111001;
assign LUT_1[63894] = 32'b00000000000000001001100001001110;
assign LUT_1[63895] = 32'b00000000000000000010110011001010;
assign LUT_1[63896] = 32'b00000000000000000101000111011011;
assign LUT_1[63897] = 32'b11111111111111111110011001010111;
assign LUT_1[63898] = 32'b00000000000000000000110101101100;
assign LUT_1[63899] = 32'b11111111111111111010000111101000;
assign LUT_1[63900] = 32'b00000000000000001101000000110010;
assign LUT_1[63901] = 32'b00000000000000000110010010101110;
assign LUT_1[63902] = 32'b00000000000000001000101111000011;
assign LUT_1[63903] = 32'b00000000000000000010000000111111;
assign LUT_1[63904] = 32'b00000000000000000100111001000011;
assign LUT_1[63905] = 32'b11111111111111111110001010111111;
assign LUT_1[63906] = 32'b00000000000000000000100111010100;
assign LUT_1[63907] = 32'b11111111111111111001111001010000;
assign LUT_1[63908] = 32'b00000000000000001100110010011010;
assign LUT_1[63909] = 32'b00000000000000000110000100010110;
assign LUT_1[63910] = 32'b00000000000000001000100000101011;
assign LUT_1[63911] = 32'b00000000000000000001110010100111;
assign LUT_1[63912] = 32'b00000000000000000100000110111000;
assign LUT_1[63913] = 32'b11111111111111111101011000110100;
assign LUT_1[63914] = 32'b11111111111111111111110101001001;
assign LUT_1[63915] = 32'b11111111111111111001000111000101;
assign LUT_1[63916] = 32'b00000000000000001100000000001111;
assign LUT_1[63917] = 32'b00000000000000000101010010001011;
assign LUT_1[63918] = 32'b00000000000000000111101110100000;
assign LUT_1[63919] = 32'b00000000000000000001000000011100;
assign LUT_1[63920] = 32'b00000000000000000110110100100101;
assign LUT_1[63921] = 32'b00000000000000000000000110100001;
assign LUT_1[63922] = 32'b00000000000000000010100010110110;
assign LUT_1[63923] = 32'b11111111111111111011110100110010;
assign LUT_1[63924] = 32'b00000000000000001110101101111100;
assign LUT_1[63925] = 32'b00000000000000000111111111111000;
assign LUT_1[63926] = 32'b00000000000000001010011100001101;
assign LUT_1[63927] = 32'b00000000000000000011101110001001;
assign LUT_1[63928] = 32'b00000000000000000110000010011010;
assign LUT_1[63929] = 32'b11111111111111111111010100010110;
assign LUT_1[63930] = 32'b00000000000000000001110000101011;
assign LUT_1[63931] = 32'b11111111111111111011000010100111;
assign LUT_1[63932] = 32'b00000000000000001101111011110001;
assign LUT_1[63933] = 32'b00000000000000000111001101101101;
assign LUT_1[63934] = 32'b00000000000000001001101010000010;
assign LUT_1[63935] = 32'b00000000000000000010111011111110;
assign LUT_1[63936] = 32'b00000000000000000101111011101100;
assign LUT_1[63937] = 32'b11111111111111111111001101101000;
assign LUT_1[63938] = 32'b00000000000000000001101001111101;
assign LUT_1[63939] = 32'b11111111111111111010111011111001;
assign LUT_1[63940] = 32'b00000000000000001101110101000011;
assign LUT_1[63941] = 32'b00000000000000000111000110111111;
assign LUT_1[63942] = 32'b00000000000000001001100011010100;
assign LUT_1[63943] = 32'b00000000000000000010110101010000;
assign LUT_1[63944] = 32'b00000000000000000101001001100001;
assign LUT_1[63945] = 32'b11111111111111111110011011011101;
assign LUT_1[63946] = 32'b00000000000000000000110111110010;
assign LUT_1[63947] = 32'b11111111111111111010001001101110;
assign LUT_1[63948] = 32'b00000000000000001101000010111000;
assign LUT_1[63949] = 32'b00000000000000000110010100110100;
assign LUT_1[63950] = 32'b00000000000000001000110001001001;
assign LUT_1[63951] = 32'b00000000000000000010000011000101;
assign LUT_1[63952] = 32'b00000000000000000111110111001110;
assign LUT_1[63953] = 32'b00000000000000000001001001001010;
assign LUT_1[63954] = 32'b00000000000000000011100101011111;
assign LUT_1[63955] = 32'b11111111111111111100110111011011;
assign LUT_1[63956] = 32'b00000000000000001111110000100101;
assign LUT_1[63957] = 32'b00000000000000001001000010100001;
assign LUT_1[63958] = 32'b00000000000000001011011110110110;
assign LUT_1[63959] = 32'b00000000000000000100110000110010;
assign LUT_1[63960] = 32'b00000000000000000111000101000011;
assign LUT_1[63961] = 32'b00000000000000000000010110111111;
assign LUT_1[63962] = 32'b00000000000000000010110011010100;
assign LUT_1[63963] = 32'b11111111111111111100000101010000;
assign LUT_1[63964] = 32'b00000000000000001110111110011010;
assign LUT_1[63965] = 32'b00000000000000001000010000010110;
assign LUT_1[63966] = 32'b00000000000000001010101100101011;
assign LUT_1[63967] = 32'b00000000000000000011111110100111;
assign LUT_1[63968] = 32'b00000000000000000110110110101011;
assign LUT_1[63969] = 32'b00000000000000000000001000100111;
assign LUT_1[63970] = 32'b00000000000000000010100100111100;
assign LUT_1[63971] = 32'b11111111111111111011110110111000;
assign LUT_1[63972] = 32'b00000000000000001110110000000010;
assign LUT_1[63973] = 32'b00000000000000001000000001111110;
assign LUT_1[63974] = 32'b00000000000000001010011110010011;
assign LUT_1[63975] = 32'b00000000000000000011110000001111;
assign LUT_1[63976] = 32'b00000000000000000110000100100000;
assign LUT_1[63977] = 32'b11111111111111111111010110011100;
assign LUT_1[63978] = 32'b00000000000000000001110010110001;
assign LUT_1[63979] = 32'b11111111111111111011000100101101;
assign LUT_1[63980] = 32'b00000000000000001101111101110111;
assign LUT_1[63981] = 32'b00000000000000000111001111110011;
assign LUT_1[63982] = 32'b00000000000000001001101100001000;
assign LUT_1[63983] = 32'b00000000000000000010111110000100;
assign LUT_1[63984] = 32'b00000000000000001000110010001101;
assign LUT_1[63985] = 32'b00000000000000000010000100001001;
assign LUT_1[63986] = 32'b00000000000000000100100000011110;
assign LUT_1[63987] = 32'b11111111111111111101110010011010;
assign LUT_1[63988] = 32'b00000000000000010000101011100100;
assign LUT_1[63989] = 32'b00000000000000001001111101100000;
assign LUT_1[63990] = 32'b00000000000000001100011001110101;
assign LUT_1[63991] = 32'b00000000000000000101101011110001;
assign LUT_1[63992] = 32'b00000000000000001000000000000010;
assign LUT_1[63993] = 32'b00000000000000000001010001111110;
assign LUT_1[63994] = 32'b00000000000000000011101110010011;
assign LUT_1[63995] = 32'b11111111111111111101000000001111;
assign LUT_1[63996] = 32'b00000000000000001111111001011001;
assign LUT_1[63997] = 32'b00000000000000001001001011010101;
assign LUT_1[63998] = 32'b00000000000000001011100111101010;
assign LUT_1[63999] = 32'b00000000000000000100111001100110;
assign LUT_1[64000] = 32'b11111111111111111100111000010010;
assign LUT_1[64001] = 32'b11111111111111110110001010001110;
assign LUT_1[64002] = 32'b11111111111111111000100110100011;
assign LUT_1[64003] = 32'b11111111111111110001111000011111;
assign LUT_1[64004] = 32'b00000000000000000100110001101001;
assign LUT_1[64005] = 32'b11111111111111111110000011100101;
assign LUT_1[64006] = 32'b00000000000000000000011111111010;
assign LUT_1[64007] = 32'b11111111111111111001110001110110;
assign LUT_1[64008] = 32'b11111111111111111100000110000111;
assign LUT_1[64009] = 32'b11111111111111110101011000000011;
assign LUT_1[64010] = 32'b11111111111111110111110100011000;
assign LUT_1[64011] = 32'b11111111111111110001000110010100;
assign LUT_1[64012] = 32'b00000000000000000011111111011110;
assign LUT_1[64013] = 32'b11111111111111111101010001011010;
assign LUT_1[64014] = 32'b11111111111111111111101101101111;
assign LUT_1[64015] = 32'b11111111111111111000111111101011;
assign LUT_1[64016] = 32'b11111111111111111110110011110100;
assign LUT_1[64017] = 32'b11111111111111111000000101110000;
assign LUT_1[64018] = 32'b11111111111111111010100010000101;
assign LUT_1[64019] = 32'b11111111111111110011110100000001;
assign LUT_1[64020] = 32'b00000000000000000110101101001011;
assign LUT_1[64021] = 32'b11111111111111111111111111000111;
assign LUT_1[64022] = 32'b00000000000000000010011011011100;
assign LUT_1[64023] = 32'b11111111111111111011101101011000;
assign LUT_1[64024] = 32'b11111111111111111110000001101001;
assign LUT_1[64025] = 32'b11111111111111110111010011100101;
assign LUT_1[64026] = 32'b11111111111111111001101111111010;
assign LUT_1[64027] = 32'b11111111111111110011000001110110;
assign LUT_1[64028] = 32'b00000000000000000101111011000000;
assign LUT_1[64029] = 32'b11111111111111111111001100111100;
assign LUT_1[64030] = 32'b00000000000000000001101001010001;
assign LUT_1[64031] = 32'b11111111111111111010111011001101;
assign LUT_1[64032] = 32'b11111111111111111101110011010001;
assign LUT_1[64033] = 32'b11111111111111110111000101001101;
assign LUT_1[64034] = 32'b11111111111111111001100001100010;
assign LUT_1[64035] = 32'b11111111111111110010110011011110;
assign LUT_1[64036] = 32'b00000000000000000101101100101000;
assign LUT_1[64037] = 32'b11111111111111111110111110100100;
assign LUT_1[64038] = 32'b00000000000000000001011010111001;
assign LUT_1[64039] = 32'b11111111111111111010101100110101;
assign LUT_1[64040] = 32'b11111111111111111101000001000110;
assign LUT_1[64041] = 32'b11111111111111110110010011000010;
assign LUT_1[64042] = 32'b11111111111111111000101111010111;
assign LUT_1[64043] = 32'b11111111111111110010000001010011;
assign LUT_1[64044] = 32'b00000000000000000100111010011101;
assign LUT_1[64045] = 32'b11111111111111111110001100011001;
assign LUT_1[64046] = 32'b00000000000000000000101000101110;
assign LUT_1[64047] = 32'b11111111111111111001111010101010;
assign LUT_1[64048] = 32'b11111111111111111111101110110011;
assign LUT_1[64049] = 32'b11111111111111111001000000101111;
assign LUT_1[64050] = 32'b11111111111111111011011101000100;
assign LUT_1[64051] = 32'b11111111111111110100101111000000;
assign LUT_1[64052] = 32'b00000000000000000111101000001010;
assign LUT_1[64053] = 32'b00000000000000000000111010000110;
assign LUT_1[64054] = 32'b00000000000000000011010110011011;
assign LUT_1[64055] = 32'b11111111111111111100101000010111;
assign LUT_1[64056] = 32'b11111111111111111110111100101000;
assign LUT_1[64057] = 32'b11111111111111111000001110100100;
assign LUT_1[64058] = 32'b11111111111111111010101010111001;
assign LUT_1[64059] = 32'b11111111111111110011111100110101;
assign LUT_1[64060] = 32'b00000000000000000110110101111111;
assign LUT_1[64061] = 32'b00000000000000000000000111111011;
assign LUT_1[64062] = 32'b00000000000000000010100100010000;
assign LUT_1[64063] = 32'b11111111111111111011110110001100;
assign LUT_1[64064] = 32'b11111111111111111110110101111010;
assign LUT_1[64065] = 32'b11111111111111111000000111110110;
assign LUT_1[64066] = 32'b11111111111111111010100100001011;
assign LUT_1[64067] = 32'b11111111111111110011110110000111;
assign LUT_1[64068] = 32'b00000000000000000110101111010001;
assign LUT_1[64069] = 32'b00000000000000000000000001001101;
assign LUT_1[64070] = 32'b00000000000000000010011101100010;
assign LUT_1[64071] = 32'b11111111111111111011101111011110;
assign LUT_1[64072] = 32'b11111111111111111110000011101111;
assign LUT_1[64073] = 32'b11111111111111110111010101101011;
assign LUT_1[64074] = 32'b11111111111111111001110010000000;
assign LUT_1[64075] = 32'b11111111111111110011000011111100;
assign LUT_1[64076] = 32'b00000000000000000101111101000110;
assign LUT_1[64077] = 32'b11111111111111111111001111000010;
assign LUT_1[64078] = 32'b00000000000000000001101011010111;
assign LUT_1[64079] = 32'b11111111111111111010111101010011;
assign LUT_1[64080] = 32'b00000000000000000000110001011100;
assign LUT_1[64081] = 32'b11111111111111111010000011011000;
assign LUT_1[64082] = 32'b11111111111111111100011111101101;
assign LUT_1[64083] = 32'b11111111111111110101110001101001;
assign LUT_1[64084] = 32'b00000000000000001000101010110011;
assign LUT_1[64085] = 32'b00000000000000000001111100101111;
assign LUT_1[64086] = 32'b00000000000000000100011001000100;
assign LUT_1[64087] = 32'b11111111111111111101101011000000;
assign LUT_1[64088] = 32'b11111111111111111111111111010001;
assign LUT_1[64089] = 32'b11111111111111111001010001001101;
assign LUT_1[64090] = 32'b11111111111111111011101101100010;
assign LUT_1[64091] = 32'b11111111111111110100111111011110;
assign LUT_1[64092] = 32'b00000000000000000111111000101000;
assign LUT_1[64093] = 32'b00000000000000000001001010100100;
assign LUT_1[64094] = 32'b00000000000000000011100110111001;
assign LUT_1[64095] = 32'b11111111111111111100111000110101;
assign LUT_1[64096] = 32'b11111111111111111111110000111001;
assign LUT_1[64097] = 32'b11111111111111111001000010110101;
assign LUT_1[64098] = 32'b11111111111111111011011111001010;
assign LUT_1[64099] = 32'b11111111111111110100110001000110;
assign LUT_1[64100] = 32'b00000000000000000111101010010000;
assign LUT_1[64101] = 32'b00000000000000000000111100001100;
assign LUT_1[64102] = 32'b00000000000000000011011000100001;
assign LUT_1[64103] = 32'b11111111111111111100101010011101;
assign LUT_1[64104] = 32'b11111111111111111110111110101110;
assign LUT_1[64105] = 32'b11111111111111111000010000101010;
assign LUT_1[64106] = 32'b11111111111111111010101100111111;
assign LUT_1[64107] = 32'b11111111111111110011111110111011;
assign LUT_1[64108] = 32'b00000000000000000110111000000101;
assign LUT_1[64109] = 32'b00000000000000000000001010000001;
assign LUT_1[64110] = 32'b00000000000000000010100110010110;
assign LUT_1[64111] = 32'b11111111111111111011111000010010;
assign LUT_1[64112] = 32'b00000000000000000001101100011011;
assign LUT_1[64113] = 32'b11111111111111111010111110010111;
assign LUT_1[64114] = 32'b11111111111111111101011010101100;
assign LUT_1[64115] = 32'b11111111111111110110101100101000;
assign LUT_1[64116] = 32'b00000000000000001001100101110010;
assign LUT_1[64117] = 32'b00000000000000000010110111101110;
assign LUT_1[64118] = 32'b00000000000000000101010100000011;
assign LUT_1[64119] = 32'b11111111111111111110100101111111;
assign LUT_1[64120] = 32'b00000000000000000000111010010000;
assign LUT_1[64121] = 32'b11111111111111111010001100001100;
assign LUT_1[64122] = 32'b11111111111111111100101000100001;
assign LUT_1[64123] = 32'b11111111111111110101111010011101;
assign LUT_1[64124] = 32'b00000000000000001000110011100111;
assign LUT_1[64125] = 32'b00000000000000000010000101100011;
assign LUT_1[64126] = 32'b00000000000000000100100001111000;
assign LUT_1[64127] = 32'b11111111111111111101110011110100;
assign LUT_1[64128] = 32'b11111111111111111111111000010101;
assign LUT_1[64129] = 32'b11111111111111111001001010010001;
assign LUT_1[64130] = 32'b11111111111111111011100110100110;
assign LUT_1[64131] = 32'b11111111111111110100111000100010;
assign LUT_1[64132] = 32'b00000000000000000111110001101100;
assign LUT_1[64133] = 32'b00000000000000000001000011101000;
assign LUT_1[64134] = 32'b00000000000000000011011111111101;
assign LUT_1[64135] = 32'b11111111111111111100110001111001;
assign LUT_1[64136] = 32'b11111111111111111111000110001010;
assign LUT_1[64137] = 32'b11111111111111111000011000000110;
assign LUT_1[64138] = 32'b11111111111111111010110100011011;
assign LUT_1[64139] = 32'b11111111111111110100000110010111;
assign LUT_1[64140] = 32'b00000000000000000110111111100001;
assign LUT_1[64141] = 32'b00000000000000000000010001011101;
assign LUT_1[64142] = 32'b00000000000000000010101101110010;
assign LUT_1[64143] = 32'b11111111111111111011111111101110;
assign LUT_1[64144] = 32'b00000000000000000001110011110111;
assign LUT_1[64145] = 32'b11111111111111111011000101110011;
assign LUT_1[64146] = 32'b11111111111111111101100010001000;
assign LUT_1[64147] = 32'b11111111111111110110110100000100;
assign LUT_1[64148] = 32'b00000000000000001001101101001110;
assign LUT_1[64149] = 32'b00000000000000000010111111001010;
assign LUT_1[64150] = 32'b00000000000000000101011011011111;
assign LUT_1[64151] = 32'b11111111111111111110101101011011;
assign LUT_1[64152] = 32'b00000000000000000001000001101100;
assign LUT_1[64153] = 32'b11111111111111111010010011101000;
assign LUT_1[64154] = 32'b11111111111111111100101111111101;
assign LUT_1[64155] = 32'b11111111111111110110000001111001;
assign LUT_1[64156] = 32'b00000000000000001000111011000011;
assign LUT_1[64157] = 32'b00000000000000000010001100111111;
assign LUT_1[64158] = 32'b00000000000000000100101001010100;
assign LUT_1[64159] = 32'b11111111111111111101111011010000;
assign LUT_1[64160] = 32'b00000000000000000000110011010100;
assign LUT_1[64161] = 32'b11111111111111111010000101010000;
assign LUT_1[64162] = 32'b11111111111111111100100001100101;
assign LUT_1[64163] = 32'b11111111111111110101110011100001;
assign LUT_1[64164] = 32'b00000000000000001000101100101011;
assign LUT_1[64165] = 32'b00000000000000000001111110100111;
assign LUT_1[64166] = 32'b00000000000000000100011010111100;
assign LUT_1[64167] = 32'b11111111111111111101101100111000;
assign LUT_1[64168] = 32'b00000000000000000000000001001001;
assign LUT_1[64169] = 32'b11111111111111111001010011000101;
assign LUT_1[64170] = 32'b11111111111111111011101111011010;
assign LUT_1[64171] = 32'b11111111111111110101000001010110;
assign LUT_1[64172] = 32'b00000000000000000111111010100000;
assign LUT_1[64173] = 32'b00000000000000000001001100011100;
assign LUT_1[64174] = 32'b00000000000000000011101000110001;
assign LUT_1[64175] = 32'b11111111111111111100111010101101;
assign LUT_1[64176] = 32'b00000000000000000010101110110110;
assign LUT_1[64177] = 32'b11111111111111111100000000110010;
assign LUT_1[64178] = 32'b11111111111111111110011101000111;
assign LUT_1[64179] = 32'b11111111111111110111101111000011;
assign LUT_1[64180] = 32'b00000000000000001010101000001101;
assign LUT_1[64181] = 32'b00000000000000000011111010001001;
assign LUT_1[64182] = 32'b00000000000000000110010110011110;
assign LUT_1[64183] = 32'b11111111111111111111101000011010;
assign LUT_1[64184] = 32'b00000000000000000001111100101011;
assign LUT_1[64185] = 32'b11111111111111111011001110100111;
assign LUT_1[64186] = 32'b11111111111111111101101010111100;
assign LUT_1[64187] = 32'b11111111111111110110111100111000;
assign LUT_1[64188] = 32'b00000000000000001001110110000010;
assign LUT_1[64189] = 32'b00000000000000000011000111111110;
assign LUT_1[64190] = 32'b00000000000000000101100100010011;
assign LUT_1[64191] = 32'b11111111111111111110110110001111;
assign LUT_1[64192] = 32'b00000000000000000001110101111101;
assign LUT_1[64193] = 32'b11111111111111111011000111111001;
assign LUT_1[64194] = 32'b11111111111111111101100100001110;
assign LUT_1[64195] = 32'b11111111111111110110110110001010;
assign LUT_1[64196] = 32'b00000000000000001001101111010100;
assign LUT_1[64197] = 32'b00000000000000000011000001010000;
assign LUT_1[64198] = 32'b00000000000000000101011101100101;
assign LUT_1[64199] = 32'b11111111111111111110101111100001;
assign LUT_1[64200] = 32'b00000000000000000001000011110010;
assign LUT_1[64201] = 32'b11111111111111111010010101101110;
assign LUT_1[64202] = 32'b11111111111111111100110010000011;
assign LUT_1[64203] = 32'b11111111111111110110000011111111;
assign LUT_1[64204] = 32'b00000000000000001000111101001001;
assign LUT_1[64205] = 32'b00000000000000000010001111000101;
assign LUT_1[64206] = 32'b00000000000000000100101011011010;
assign LUT_1[64207] = 32'b11111111111111111101111101010110;
assign LUT_1[64208] = 32'b00000000000000000011110001011111;
assign LUT_1[64209] = 32'b11111111111111111101000011011011;
assign LUT_1[64210] = 32'b11111111111111111111011111110000;
assign LUT_1[64211] = 32'b11111111111111111000110001101100;
assign LUT_1[64212] = 32'b00000000000000001011101010110110;
assign LUT_1[64213] = 32'b00000000000000000100111100110010;
assign LUT_1[64214] = 32'b00000000000000000111011001000111;
assign LUT_1[64215] = 32'b00000000000000000000101011000011;
assign LUT_1[64216] = 32'b00000000000000000010111111010100;
assign LUT_1[64217] = 32'b11111111111111111100010001010000;
assign LUT_1[64218] = 32'b11111111111111111110101101100101;
assign LUT_1[64219] = 32'b11111111111111110111111111100001;
assign LUT_1[64220] = 32'b00000000000000001010111000101011;
assign LUT_1[64221] = 32'b00000000000000000100001010100111;
assign LUT_1[64222] = 32'b00000000000000000110100110111100;
assign LUT_1[64223] = 32'b11111111111111111111111000111000;
assign LUT_1[64224] = 32'b00000000000000000010110000111100;
assign LUT_1[64225] = 32'b11111111111111111100000010111000;
assign LUT_1[64226] = 32'b11111111111111111110011111001101;
assign LUT_1[64227] = 32'b11111111111111110111110001001001;
assign LUT_1[64228] = 32'b00000000000000001010101010010011;
assign LUT_1[64229] = 32'b00000000000000000011111100001111;
assign LUT_1[64230] = 32'b00000000000000000110011000100100;
assign LUT_1[64231] = 32'b11111111111111111111101010100000;
assign LUT_1[64232] = 32'b00000000000000000001111110110001;
assign LUT_1[64233] = 32'b11111111111111111011010000101101;
assign LUT_1[64234] = 32'b11111111111111111101101101000010;
assign LUT_1[64235] = 32'b11111111111111110110111110111110;
assign LUT_1[64236] = 32'b00000000000000001001111000001000;
assign LUT_1[64237] = 32'b00000000000000000011001010000100;
assign LUT_1[64238] = 32'b00000000000000000101100110011001;
assign LUT_1[64239] = 32'b11111111111111111110111000010101;
assign LUT_1[64240] = 32'b00000000000000000100101100011110;
assign LUT_1[64241] = 32'b11111111111111111101111110011010;
assign LUT_1[64242] = 32'b00000000000000000000011010101111;
assign LUT_1[64243] = 32'b11111111111111111001101100101011;
assign LUT_1[64244] = 32'b00000000000000001100100101110101;
assign LUT_1[64245] = 32'b00000000000000000101110111110001;
assign LUT_1[64246] = 32'b00000000000000001000010100000110;
assign LUT_1[64247] = 32'b00000000000000000001100110000010;
assign LUT_1[64248] = 32'b00000000000000000011111010010011;
assign LUT_1[64249] = 32'b11111111111111111101001100001111;
assign LUT_1[64250] = 32'b11111111111111111111101000100100;
assign LUT_1[64251] = 32'b11111111111111111000111010100000;
assign LUT_1[64252] = 32'b00000000000000001011110011101010;
assign LUT_1[64253] = 32'b00000000000000000101000101100110;
assign LUT_1[64254] = 32'b00000000000000000111100001111011;
assign LUT_1[64255] = 32'b00000000000000000000110011110111;
assign LUT_1[64256] = 32'b11111111111111111010101100011110;
assign LUT_1[64257] = 32'b11111111111111110011111110011010;
assign LUT_1[64258] = 32'b11111111111111110110011010101111;
assign LUT_1[64259] = 32'b11111111111111101111101100101011;
assign LUT_1[64260] = 32'b00000000000000000010100101110101;
assign LUT_1[64261] = 32'b11111111111111111011110111110001;
assign LUT_1[64262] = 32'b11111111111111111110010100000110;
assign LUT_1[64263] = 32'b11111111111111110111100110000010;
assign LUT_1[64264] = 32'b11111111111111111001111010010011;
assign LUT_1[64265] = 32'b11111111111111110011001100001111;
assign LUT_1[64266] = 32'b11111111111111110101101000100100;
assign LUT_1[64267] = 32'b11111111111111101110111010100000;
assign LUT_1[64268] = 32'b00000000000000000001110011101010;
assign LUT_1[64269] = 32'b11111111111111111011000101100110;
assign LUT_1[64270] = 32'b11111111111111111101100001111011;
assign LUT_1[64271] = 32'b11111111111111110110110011110111;
assign LUT_1[64272] = 32'b11111111111111111100101000000000;
assign LUT_1[64273] = 32'b11111111111111110101111001111100;
assign LUT_1[64274] = 32'b11111111111111111000010110010001;
assign LUT_1[64275] = 32'b11111111111111110001101000001101;
assign LUT_1[64276] = 32'b00000000000000000100100001010111;
assign LUT_1[64277] = 32'b11111111111111111101110011010011;
assign LUT_1[64278] = 32'b00000000000000000000001111101000;
assign LUT_1[64279] = 32'b11111111111111111001100001100100;
assign LUT_1[64280] = 32'b11111111111111111011110101110101;
assign LUT_1[64281] = 32'b11111111111111110101000111110001;
assign LUT_1[64282] = 32'b11111111111111110111100100000110;
assign LUT_1[64283] = 32'b11111111111111110000110110000010;
assign LUT_1[64284] = 32'b00000000000000000011101111001100;
assign LUT_1[64285] = 32'b11111111111111111101000001001000;
assign LUT_1[64286] = 32'b11111111111111111111011101011101;
assign LUT_1[64287] = 32'b11111111111111111000101111011001;
assign LUT_1[64288] = 32'b11111111111111111011100111011101;
assign LUT_1[64289] = 32'b11111111111111110100111001011001;
assign LUT_1[64290] = 32'b11111111111111110111010101101110;
assign LUT_1[64291] = 32'b11111111111111110000100111101010;
assign LUT_1[64292] = 32'b00000000000000000011100000110100;
assign LUT_1[64293] = 32'b11111111111111111100110010110000;
assign LUT_1[64294] = 32'b11111111111111111111001111000101;
assign LUT_1[64295] = 32'b11111111111111111000100001000001;
assign LUT_1[64296] = 32'b11111111111111111010110101010010;
assign LUT_1[64297] = 32'b11111111111111110100000111001110;
assign LUT_1[64298] = 32'b11111111111111110110100011100011;
assign LUT_1[64299] = 32'b11111111111111101111110101011111;
assign LUT_1[64300] = 32'b00000000000000000010101110101001;
assign LUT_1[64301] = 32'b11111111111111111100000000100101;
assign LUT_1[64302] = 32'b11111111111111111110011100111010;
assign LUT_1[64303] = 32'b11111111111111110111101110110110;
assign LUT_1[64304] = 32'b11111111111111111101100010111111;
assign LUT_1[64305] = 32'b11111111111111110110110100111011;
assign LUT_1[64306] = 32'b11111111111111111001010001010000;
assign LUT_1[64307] = 32'b11111111111111110010100011001100;
assign LUT_1[64308] = 32'b00000000000000000101011100010110;
assign LUT_1[64309] = 32'b11111111111111111110101110010010;
assign LUT_1[64310] = 32'b00000000000000000001001010100111;
assign LUT_1[64311] = 32'b11111111111111111010011100100011;
assign LUT_1[64312] = 32'b11111111111111111100110000110100;
assign LUT_1[64313] = 32'b11111111111111110110000010110000;
assign LUT_1[64314] = 32'b11111111111111111000011111000101;
assign LUT_1[64315] = 32'b11111111111111110001110001000001;
assign LUT_1[64316] = 32'b00000000000000000100101010001011;
assign LUT_1[64317] = 32'b11111111111111111101111100000111;
assign LUT_1[64318] = 32'b00000000000000000000011000011100;
assign LUT_1[64319] = 32'b11111111111111111001101010011000;
assign LUT_1[64320] = 32'b11111111111111111100101010000110;
assign LUT_1[64321] = 32'b11111111111111110101111100000010;
assign LUT_1[64322] = 32'b11111111111111111000011000010111;
assign LUT_1[64323] = 32'b11111111111111110001101010010011;
assign LUT_1[64324] = 32'b00000000000000000100100011011101;
assign LUT_1[64325] = 32'b11111111111111111101110101011001;
assign LUT_1[64326] = 32'b00000000000000000000010001101110;
assign LUT_1[64327] = 32'b11111111111111111001100011101010;
assign LUT_1[64328] = 32'b11111111111111111011110111111011;
assign LUT_1[64329] = 32'b11111111111111110101001001110111;
assign LUT_1[64330] = 32'b11111111111111110111100110001100;
assign LUT_1[64331] = 32'b11111111111111110000111000001000;
assign LUT_1[64332] = 32'b00000000000000000011110001010010;
assign LUT_1[64333] = 32'b11111111111111111101000011001110;
assign LUT_1[64334] = 32'b11111111111111111111011111100011;
assign LUT_1[64335] = 32'b11111111111111111000110001011111;
assign LUT_1[64336] = 32'b11111111111111111110100101101000;
assign LUT_1[64337] = 32'b11111111111111110111110111100100;
assign LUT_1[64338] = 32'b11111111111111111010010011111001;
assign LUT_1[64339] = 32'b11111111111111110011100101110101;
assign LUT_1[64340] = 32'b00000000000000000110011110111111;
assign LUT_1[64341] = 32'b11111111111111111111110000111011;
assign LUT_1[64342] = 32'b00000000000000000010001101010000;
assign LUT_1[64343] = 32'b11111111111111111011011111001100;
assign LUT_1[64344] = 32'b11111111111111111101110011011101;
assign LUT_1[64345] = 32'b11111111111111110111000101011001;
assign LUT_1[64346] = 32'b11111111111111111001100001101110;
assign LUT_1[64347] = 32'b11111111111111110010110011101010;
assign LUT_1[64348] = 32'b00000000000000000101101100110100;
assign LUT_1[64349] = 32'b11111111111111111110111110110000;
assign LUT_1[64350] = 32'b00000000000000000001011011000101;
assign LUT_1[64351] = 32'b11111111111111111010101101000001;
assign LUT_1[64352] = 32'b11111111111111111101100101000101;
assign LUT_1[64353] = 32'b11111111111111110110110111000001;
assign LUT_1[64354] = 32'b11111111111111111001010011010110;
assign LUT_1[64355] = 32'b11111111111111110010100101010010;
assign LUT_1[64356] = 32'b00000000000000000101011110011100;
assign LUT_1[64357] = 32'b11111111111111111110110000011000;
assign LUT_1[64358] = 32'b00000000000000000001001100101101;
assign LUT_1[64359] = 32'b11111111111111111010011110101001;
assign LUT_1[64360] = 32'b11111111111111111100110010111010;
assign LUT_1[64361] = 32'b11111111111111110110000100110110;
assign LUT_1[64362] = 32'b11111111111111111000100001001011;
assign LUT_1[64363] = 32'b11111111111111110001110011000111;
assign LUT_1[64364] = 32'b00000000000000000100101100010001;
assign LUT_1[64365] = 32'b11111111111111111101111110001101;
assign LUT_1[64366] = 32'b00000000000000000000011010100010;
assign LUT_1[64367] = 32'b11111111111111111001101100011110;
assign LUT_1[64368] = 32'b11111111111111111111100000100111;
assign LUT_1[64369] = 32'b11111111111111111000110010100011;
assign LUT_1[64370] = 32'b11111111111111111011001110111000;
assign LUT_1[64371] = 32'b11111111111111110100100000110100;
assign LUT_1[64372] = 32'b00000000000000000111011001111110;
assign LUT_1[64373] = 32'b00000000000000000000101011111010;
assign LUT_1[64374] = 32'b00000000000000000011001000001111;
assign LUT_1[64375] = 32'b11111111111111111100011010001011;
assign LUT_1[64376] = 32'b11111111111111111110101110011100;
assign LUT_1[64377] = 32'b11111111111111111000000000011000;
assign LUT_1[64378] = 32'b11111111111111111010011100101101;
assign LUT_1[64379] = 32'b11111111111111110011101110101001;
assign LUT_1[64380] = 32'b00000000000000000110100111110011;
assign LUT_1[64381] = 32'b11111111111111111111111001101111;
assign LUT_1[64382] = 32'b00000000000000000010010110000100;
assign LUT_1[64383] = 32'b11111111111111111011101000000000;
assign LUT_1[64384] = 32'b11111111111111111101101100100001;
assign LUT_1[64385] = 32'b11111111111111110110111110011101;
assign LUT_1[64386] = 32'b11111111111111111001011010110010;
assign LUT_1[64387] = 32'b11111111111111110010101100101110;
assign LUT_1[64388] = 32'b00000000000000000101100101111000;
assign LUT_1[64389] = 32'b11111111111111111110110111110100;
assign LUT_1[64390] = 32'b00000000000000000001010100001001;
assign LUT_1[64391] = 32'b11111111111111111010100110000101;
assign LUT_1[64392] = 32'b11111111111111111100111010010110;
assign LUT_1[64393] = 32'b11111111111111110110001100010010;
assign LUT_1[64394] = 32'b11111111111111111000101000100111;
assign LUT_1[64395] = 32'b11111111111111110001111010100011;
assign LUT_1[64396] = 32'b00000000000000000100110011101101;
assign LUT_1[64397] = 32'b11111111111111111110000101101001;
assign LUT_1[64398] = 32'b00000000000000000000100001111110;
assign LUT_1[64399] = 32'b11111111111111111001110011111010;
assign LUT_1[64400] = 32'b11111111111111111111101000000011;
assign LUT_1[64401] = 32'b11111111111111111000111001111111;
assign LUT_1[64402] = 32'b11111111111111111011010110010100;
assign LUT_1[64403] = 32'b11111111111111110100101000010000;
assign LUT_1[64404] = 32'b00000000000000000111100001011010;
assign LUT_1[64405] = 32'b00000000000000000000110011010110;
assign LUT_1[64406] = 32'b00000000000000000011001111101011;
assign LUT_1[64407] = 32'b11111111111111111100100001100111;
assign LUT_1[64408] = 32'b11111111111111111110110101111000;
assign LUT_1[64409] = 32'b11111111111111111000000111110100;
assign LUT_1[64410] = 32'b11111111111111111010100100001001;
assign LUT_1[64411] = 32'b11111111111111110011110110000101;
assign LUT_1[64412] = 32'b00000000000000000110101111001111;
assign LUT_1[64413] = 32'b00000000000000000000000001001011;
assign LUT_1[64414] = 32'b00000000000000000010011101100000;
assign LUT_1[64415] = 32'b11111111111111111011101111011100;
assign LUT_1[64416] = 32'b11111111111111111110100111100000;
assign LUT_1[64417] = 32'b11111111111111110111111001011100;
assign LUT_1[64418] = 32'b11111111111111111010010101110001;
assign LUT_1[64419] = 32'b11111111111111110011100111101101;
assign LUT_1[64420] = 32'b00000000000000000110100000110111;
assign LUT_1[64421] = 32'b11111111111111111111110010110011;
assign LUT_1[64422] = 32'b00000000000000000010001111001000;
assign LUT_1[64423] = 32'b11111111111111111011100001000100;
assign LUT_1[64424] = 32'b11111111111111111101110101010101;
assign LUT_1[64425] = 32'b11111111111111110111000111010001;
assign LUT_1[64426] = 32'b11111111111111111001100011100110;
assign LUT_1[64427] = 32'b11111111111111110010110101100010;
assign LUT_1[64428] = 32'b00000000000000000101101110101100;
assign LUT_1[64429] = 32'b11111111111111111111000000101000;
assign LUT_1[64430] = 32'b00000000000000000001011100111101;
assign LUT_1[64431] = 32'b11111111111111111010101110111001;
assign LUT_1[64432] = 32'b00000000000000000000100011000010;
assign LUT_1[64433] = 32'b11111111111111111001110100111110;
assign LUT_1[64434] = 32'b11111111111111111100010001010011;
assign LUT_1[64435] = 32'b11111111111111110101100011001111;
assign LUT_1[64436] = 32'b00000000000000001000011100011001;
assign LUT_1[64437] = 32'b00000000000000000001101110010101;
assign LUT_1[64438] = 32'b00000000000000000100001010101010;
assign LUT_1[64439] = 32'b11111111111111111101011100100110;
assign LUT_1[64440] = 32'b11111111111111111111110000110111;
assign LUT_1[64441] = 32'b11111111111111111001000010110011;
assign LUT_1[64442] = 32'b11111111111111111011011111001000;
assign LUT_1[64443] = 32'b11111111111111110100110001000100;
assign LUT_1[64444] = 32'b00000000000000000111101010001110;
assign LUT_1[64445] = 32'b00000000000000000000111100001010;
assign LUT_1[64446] = 32'b00000000000000000011011000011111;
assign LUT_1[64447] = 32'b11111111111111111100101010011011;
assign LUT_1[64448] = 32'b11111111111111111111101010001001;
assign LUT_1[64449] = 32'b11111111111111111000111100000101;
assign LUT_1[64450] = 32'b11111111111111111011011000011010;
assign LUT_1[64451] = 32'b11111111111111110100101010010110;
assign LUT_1[64452] = 32'b00000000000000000111100011100000;
assign LUT_1[64453] = 32'b00000000000000000000110101011100;
assign LUT_1[64454] = 32'b00000000000000000011010001110001;
assign LUT_1[64455] = 32'b11111111111111111100100011101101;
assign LUT_1[64456] = 32'b11111111111111111110110111111110;
assign LUT_1[64457] = 32'b11111111111111111000001001111010;
assign LUT_1[64458] = 32'b11111111111111111010100110001111;
assign LUT_1[64459] = 32'b11111111111111110011111000001011;
assign LUT_1[64460] = 32'b00000000000000000110110001010101;
assign LUT_1[64461] = 32'b00000000000000000000000011010001;
assign LUT_1[64462] = 32'b00000000000000000010011111100110;
assign LUT_1[64463] = 32'b11111111111111111011110001100010;
assign LUT_1[64464] = 32'b00000000000000000001100101101011;
assign LUT_1[64465] = 32'b11111111111111111010110111100111;
assign LUT_1[64466] = 32'b11111111111111111101010011111100;
assign LUT_1[64467] = 32'b11111111111111110110100101111000;
assign LUT_1[64468] = 32'b00000000000000001001011111000010;
assign LUT_1[64469] = 32'b00000000000000000010110000111110;
assign LUT_1[64470] = 32'b00000000000000000101001101010011;
assign LUT_1[64471] = 32'b11111111111111111110011111001111;
assign LUT_1[64472] = 32'b00000000000000000000110011100000;
assign LUT_1[64473] = 32'b11111111111111111010000101011100;
assign LUT_1[64474] = 32'b11111111111111111100100001110001;
assign LUT_1[64475] = 32'b11111111111111110101110011101101;
assign LUT_1[64476] = 32'b00000000000000001000101100110111;
assign LUT_1[64477] = 32'b00000000000000000001111110110011;
assign LUT_1[64478] = 32'b00000000000000000100011011001000;
assign LUT_1[64479] = 32'b11111111111111111101101101000100;
assign LUT_1[64480] = 32'b00000000000000000000100101001000;
assign LUT_1[64481] = 32'b11111111111111111001110111000100;
assign LUT_1[64482] = 32'b11111111111111111100010011011001;
assign LUT_1[64483] = 32'b11111111111111110101100101010101;
assign LUT_1[64484] = 32'b00000000000000001000011110011111;
assign LUT_1[64485] = 32'b00000000000000000001110000011011;
assign LUT_1[64486] = 32'b00000000000000000100001100110000;
assign LUT_1[64487] = 32'b11111111111111111101011110101100;
assign LUT_1[64488] = 32'b11111111111111111111110010111101;
assign LUT_1[64489] = 32'b11111111111111111001000100111001;
assign LUT_1[64490] = 32'b11111111111111111011100001001110;
assign LUT_1[64491] = 32'b11111111111111110100110011001010;
assign LUT_1[64492] = 32'b00000000000000000111101100010100;
assign LUT_1[64493] = 32'b00000000000000000000111110010000;
assign LUT_1[64494] = 32'b00000000000000000011011010100101;
assign LUT_1[64495] = 32'b11111111111111111100101100100001;
assign LUT_1[64496] = 32'b00000000000000000010100000101010;
assign LUT_1[64497] = 32'b11111111111111111011110010100110;
assign LUT_1[64498] = 32'b11111111111111111110001110111011;
assign LUT_1[64499] = 32'b11111111111111110111100000110111;
assign LUT_1[64500] = 32'b00000000000000001010011010000001;
assign LUT_1[64501] = 32'b00000000000000000011101011111101;
assign LUT_1[64502] = 32'b00000000000000000110001000010010;
assign LUT_1[64503] = 32'b11111111111111111111011010001110;
assign LUT_1[64504] = 32'b00000000000000000001101110011111;
assign LUT_1[64505] = 32'b11111111111111111011000000011011;
assign LUT_1[64506] = 32'b11111111111111111101011100110000;
assign LUT_1[64507] = 32'b11111111111111110110101110101100;
assign LUT_1[64508] = 32'b00000000000000001001100111110110;
assign LUT_1[64509] = 32'b00000000000000000010111001110010;
assign LUT_1[64510] = 32'b00000000000000000101010110000111;
assign LUT_1[64511] = 32'b11111111111111111110101000000011;
assign LUT_1[64512] = 32'b00000000000000001001100000100101;
assign LUT_1[64513] = 32'b00000000000000000010110010100001;
assign LUT_1[64514] = 32'b00000000000000000101001110110110;
assign LUT_1[64515] = 32'b11111111111111111110100000110010;
assign LUT_1[64516] = 32'b00000000000000010001011001111100;
assign LUT_1[64517] = 32'b00000000000000001010101011111000;
assign LUT_1[64518] = 32'b00000000000000001101001000001101;
assign LUT_1[64519] = 32'b00000000000000000110011010001001;
assign LUT_1[64520] = 32'b00000000000000001000101110011010;
assign LUT_1[64521] = 32'b00000000000000000010000000010110;
assign LUT_1[64522] = 32'b00000000000000000100011100101011;
assign LUT_1[64523] = 32'b11111111111111111101101110100111;
assign LUT_1[64524] = 32'b00000000000000010000100111110001;
assign LUT_1[64525] = 32'b00000000000000001001111001101101;
assign LUT_1[64526] = 32'b00000000000000001100010110000010;
assign LUT_1[64527] = 32'b00000000000000000101100111111110;
assign LUT_1[64528] = 32'b00000000000000001011011100000111;
assign LUT_1[64529] = 32'b00000000000000000100101110000011;
assign LUT_1[64530] = 32'b00000000000000000111001010011000;
assign LUT_1[64531] = 32'b00000000000000000000011100010100;
assign LUT_1[64532] = 32'b00000000000000010011010101011110;
assign LUT_1[64533] = 32'b00000000000000001100100111011010;
assign LUT_1[64534] = 32'b00000000000000001111000011101111;
assign LUT_1[64535] = 32'b00000000000000001000010101101011;
assign LUT_1[64536] = 32'b00000000000000001010101001111100;
assign LUT_1[64537] = 32'b00000000000000000011111011111000;
assign LUT_1[64538] = 32'b00000000000000000110011000001101;
assign LUT_1[64539] = 32'b11111111111111111111101010001001;
assign LUT_1[64540] = 32'b00000000000000010010100011010011;
assign LUT_1[64541] = 32'b00000000000000001011110101001111;
assign LUT_1[64542] = 32'b00000000000000001110010001100100;
assign LUT_1[64543] = 32'b00000000000000000111100011100000;
assign LUT_1[64544] = 32'b00000000000000001010011011100100;
assign LUT_1[64545] = 32'b00000000000000000011101101100000;
assign LUT_1[64546] = 32'b00000000000000000110001001110101;
assign LUT_1[64547] = 32'b11111111111111111111011011110001;
assign LUT_1[64548] = 32'b00000000000000010010010100111011;
assign LUT_1[64549] = 32'b00000000000000001011100110110111;
assign LUT_1[64550] = 32'b00000000000000001110000011001100;
assign LUT_1[64551] = 32'b00000000000000000111010101001000;
assign LUT_1[64552] = 32'b00000000000000001001101001011001;
assign LUT_1[64553] = 32'b00000000000000000010111011010101;
assign LUT_1[64554] = 32'b00000000000000000101010111101010;
assign LUT_1[64555] = 32'b11111111111111111110101001100110;
assign LUT_1[64556] = 32'b00000000000000010001100010110000;
assign LUT_1[64557] = 32'b00000000000000001010110100101100;
assign LUT_1[64558] = 32'b00000000000000001101010001000001;
assign LUT_1[64559] = 32'b00000000000000000110100010111101;
assign LUT_1[64560] = 32'b00000000000000001100010111000110;
assign LUT_1[64561] = 32'b00000000000000000101101001000010;
assign LUT_1[64562] = 32'b00000000000000001000000101010111;
assign LUT_1[64563] = 32'b00000000000000000001010111010011;
assign LUT_1[64564] = 32'b00000000000000010100010000011101;
assign LUT_1[64565] = 32'b00000000000000001101100010011001;
assign LUT_1[64566] = 32'b00000000000000001111111110101110;
assign LUT_1[64567] = 32'b00000000000000001001010000101010;
assign LUT_1[64568] = 32'b00000000000000001011100100111011;
assign LUT_1[64569] = 32'b00000000000000000100110110110111;
assign LUT_1[64570] = 32'b00000000000000000111010011001100;
assign LUT_1[64571] = 32'b00000000000000000000100101001000;
assign LUT_1[64572] = 32'b00000000000000010011011110010010;
assign LUT_1[64573] = 32'b00000000000000001100110000001110;
assign LUT_1[64574] = 32'b00000000000000001111001100100011;
assign LUT_1[64575] = 32'b00000000000000001000011110011111;
assign LUT_1[64576] = 32'b00000000000000001011011110001101;
assign LUT_1[64577] = 32'b00000000000000000100110000001001;
assign LUT_1[64578] = 32'b00000000000000000111001100011110;
assign LUT_1[64579] = 32'b00000000000000000000011110011010;
assign LUT_1[64580] = 32'b00000000000000010011010111100100;
assign LUT_1[64581] = 32'b00000000000000001100101001100000;
assign LUT_1[64582] = 32'b00000000000000001111000101110101;
assign LUT_1[64583] = 32'b00000000000000001000010111110001;
assign LUT_1[64584] = 32'b00000000000000001010101100000010;
assign LUT_1[64585] = 32'b00000000000000000011111101111110;
assign LUT_1[64586] = 32'b00000000000000000110011010010011;
assign LUT_1[64587] = 32'b11111111111111111111101100001111;
assign LUT_1[64588] = 32'b00000000000000010010100101011001;
assign LUT_1[64589] = 32'b00000000000000001011110111010101;
assign LUT_1[64590] = 32'b00000000000000001110010011101010;
assign LUT_1[64591] = 32'b00000000000000000111100101100110;
assign LUT_1[64592] = 32'b00000000000000001101011001101111;
assign LUT_1[64593] = 32'b00000000000000000110101011101011;
assign LUT_1[64594] = 32'b00000000000000001001001000000000;
assign LUT_1[64595] = 32'b00000000000000000010011001111100;
assign LUT_1[64596] = 32'b00000000000000010101010011000110;
assign LUT_1[64597] = 32'b00000000000000001110100101000010;
assign LUT_1[64598] = 32'b00000000000000010001000001010111;
assign LUT_1[64599] = 32'b00000000000000001010010011010011;
assign LUT_1[64600] = 32'b00000000000000001100100111100100;
assign LUT_1[64601] = 32'b00000000000000000101111001100000;
assign LUT_1[64602] = 32'b00000000000000001000010101110101;
assign LUT_1[64603] = 32'b00000000000000000001100111110001;
assign LUT_1[64604] = 32'b00000000000000010100100000111011;
assign LUT_1[64605] = 32'b00000000000000001101110010110111;
assign LUT_1[64606] = 32'b00000000000000010000001111001100;
assign LUT_1[64607] = 32'b00000000000000001001100001001000;
assign LUT_1[64608] = 32'b00000000000000001100011001001100;
assign LUT_1[64609] = 32'b00000000000000000101101011001000;
assign LUT_1[64610] = 32'b00000000000000001000000111011101;
assign LUT_1[64611] = 32'b00000000000000000001011001011001;
assign LUT_1[64612] = 32'b00000000000000010100010010100011;
assign LUT_1[64613] = 32'b00000000000000001101100100011111;
assign LUT_1[64614] = 32'b00000000000000010000000000110100;
assign LUT_1[64615] = 32'b00000000000000001001010010110000;
assign LUT_1[64616] = 32'b00000000000000001011100111000001;
assign LUT_1[64617] = 32'b00000000000000000100111000111101;
assign LUT_1[64618] = 32'b00000000000000000111010101010010;
assign LUT_1[64619] = 32'b00000000000000000000100111001110;
assign LUT_1[64620] = 32'b00000000000000010011100000011000;
assign LUT_1[64621] = 32'b00000000000000001100110010010100;
assign LUT_1[64622] = 32'b00000000000000001111001110101001;
assign LUT_1[64623] = 32'b00000000000000001000100000100101;
assign LUT_1[64624] = 32'b00000000000000001110010100101110;
assign LUT_1[64625] = 32'b00000000000000000111100110101010;
assign LUT_1[64626] = 32'b00000000000000001010000010111111;
assign LUT_1[64627] = 32'b00000000000000000011010100111011;
assign LUT_1[64628] = 32'b00000000000000010110001110000101;
assign LUT_1[64629] = 32'b00000000000000001111100000000001;
assign LUT_1[64630] = 32'b00000000000000010001111100010110;
assign LUT_1[64631] = 32'b00000000000000001011001110010010;
assign LUT_1[64632] = 32'b00000000000000001101100010100011;
assign LUT_1[64633] = 32'b00000000000000000110110100011111;
assign LUT_1[64634] = 32'b00000000000000001001010000110100;
assign LUT_1[64635] = 32'b00000000000000000010100010110000;
assign LUT_1[64636] = 32'b00000000000000010101011011111010;
assign LUT_1[64637] = 32'b00000000000000001110101101110110;
assign LUT_1[64638] = 32'b00000000000000010001001010001011;
assign LUT_1[64639] = 32'b00000000000000001010011100000111;
assign LUT_1[64640] = 32'b00000000000000001100100000101000;
assign LUT_1[64641] = 32'b00000000000000000101110010100100;
assign LUT_1[64642] = 32'b00000000000000001000001110111001;
assign LUT_1[64643] = 32'b00000000000000000001100000110101;
assign LUT_1[64644] = 32'b00000000000000010100011001111111;
assign LUT_1[64645] = 32'b00000000000000001101101011111011;
assign LUT_1[64646] = 32'b00000000000000010000001000010000;
assign LUT_1[64647] = 32'b00000000000000001001011010001100;
assign LUT_1[64648] = 32'b00000000000000001011101110011101;
assign LUT_1[64649] = 32'b00000000000000000101000000011001;
assign LUT_1[64650] = 32'b00000000000000000111011100101110;
assign LUT_1[64651] = 32'b00000000000000000000101110101010;
assign LUT_1[64652] = 32'b00000000000000010011100111110100;
assign LUT_1[64653] = 32'b00000000000000001100111001110000;
assign LUT_1[64654] = 32'b00000000000000001111010110000101;
assign LUT_1[64655] = 32'b00000000000000001000101000000001;
assign LUT_1[64656] = 32'b00000000000000001110011100001010;
assign LUT_1[64657] = 32'b00000000000000000111101110000110;
assign LUT_1[64658] = 32'b00000000000000001010001010011011;
assign LUT_1[64659] = 32'b00000000000000000011011100010111;
assign LUT_1[64660] = 32'b00000000000000010110010101100001;
assign LUT_1[64661] = 32'b00000000000000001111100111011101;
assign LUT_1[64662] = 32'b00000000000000010010000011110010;
assign LUT_1[64663] = 32'b00000000000000001011010101101110;
assign LUT_1[64664] = 32'b00000000000000001101101001111111;
assign LUT_1[64665] = 32'b00000000000000000110111011111011;
assign LUT_1[64666] = 32'b00000000000000001001011000010000;
assign LUT_1[64667] = 32'b00000000000000000010101010001100;
assign LUT_1[64668] = 32'b00000000000000010101100011010110;
assign LUT_1[64669] = 32'b00000000000000001110110101010010;
assign LUT_1[64670] = 32'b00000000000000010001010001100111;
assign LUT_1[64671] = 32'b00000000000000001010100011100011;
assign LUT_1[64672] = 32'b00000000000000001101011011100111;
assign LUT_1[64673] = 32'b00000000000000000110101101100011;
assign LUT_1[64674] = 32'b00000000000000001001001001111000;
assign LUT_1[64675] = 32'b00000000000000000010011011110100;
assign LUT_1[64676] = 32'b00000000000000010101010100111110;
assign LUT_1[64677] = 32'b00000000000000001110100110111010;
assign LUT_1[64678] = 32'b00000000000000010001000011001111;
assign LUT_1[64679] = 32'b00000000000000001010010101001011;
assign LUT_1[64680] = 32'b00000000000000001100101001011100;
assign LUT_1[64681] = 32'b00000000000000000101111011011000;
assign LUT_1[64682] = 32'b00000000000000001000010111101101;
assign LUT_1[64683] = 32'b00000000000000000001101001101001;
assign LUT_1[64684] = 32'b00000000000000010100100010110011;
assign LUT_1[64685] = 32'b00000000000000001101110100101111;
assign LUT_1[64686] = 32'b00000000000000010000010001000100;
assign LUT_1[64687] = 32'b00000000000000001001100011000000;
assign LUT_1[64688] = 32'b00000000000000001111010111001001;
assign LUT_1[64689] = 32'b00000000000000001000101001000101;
assign LUT_1[64690] = 32'b00000000000000001011000101011010;
assign LUT_1[64691] = 32'b00000000000000000100010111010110;
assign LUT_1[64692] = 32'b00000000000000010111010000100000;
assign LUT_1[64693] = 32'b00000000000000010000100010011100;
assign LUT_1[64694] = 32'b00000000000000010010111110110001;
assign LUT_1[64695] = 32'b00000000000000001100010000101101;
assign LUT_1[64696] = 32'b00000000000000001110100100111110;
assign LUT_1[64697] = 32'b00000000000000000111110110111010;
assign LUT_1[64698] = 32'b00000000000000001010010011001111;
assign LUT_1[64699] = 32'b00000000000000000011100101001011;
assign LUT_1[64700] = 32'b00000000000000010110011110010101;
assign LUT_1[64701] = 32'b00000000000000001111110000010001;
assign LUT_1[64702] = 32'b00000000000000010010001100100110;
assign LUT_1[64703] = 32'b00000000000000001011011110100010;
assign LUT_1[64704] = 32'b00000000000000001110011110010000;
assign LUT_1[64705] = 32'b00000000000000000111110000001100;
assign LUT_1[64706] = 32'b00000000000000001010001100100001;
assign LUT_1[64707] = 32'b00000000000000000011011110011101;
assign LUT_1[64708] = 32'b00000000000000010110010111100111;
assign LUT_1[64709] = 32'b00000000000000001111101001100011;
assign LUT_1[64710] = 32'b00000000000000010010000101111000;
assign LUT_1[64711] = 32'b00000000000000001011010111110100;
assign LUT_1[64712] = 32'b00000000000000001101101100000101;
assign LUT_1[64713] = 32'b00000000000000000110111110000001;
assign LUT_1[64714] = 32'b00000000000000001001011010010110;
assign LUT_1[64715] = 32'b00000000000000000010101100010010;
assign LUT_1[64716] = 32'b00000000000000010101100101011100;
assign LUT_1[64717] = 32'b00000000000000001110110111011000;
assign LUT_1[64718] = 32'b00000000000000010001010011101101;
assign LUT_1[64719] = 32'b00000000000000001010100101101001;
assign LUT_1[64720] = 32'b00000000000000010000011001110010;
assign LUT_1[64721] = 32'b00000000000000001001101011101110;
assign LUT_1[64722] = 32'b00000000000000001100001000000011;
assign LUT_1[64723] = 32'b00000000000000000101011001111111;
assign LUT_1[64724] = 32'b00000000000000011000010011001001;
assign LUT_1[64725] = 32'b00000000000000010001100101000101;
assign LUT_1[64726] = 32'b00000000000000010100000001011010;
assign LUT_1[64727] = 32'b00000000000000001101010011010110;
assign LUT_1[64728] = 32'b00000000000000001111100111100111;
assign LUT_1[64729] = 32'b00000000000000001000111001100011;
assign LUT_1[64730] = 32'b00000000000000001011010101111000;
assign LUT_1[64731] = 32'b00000000000000000100100111110100;
assign LUT_1[64732] = 32'b00000000000000010111100000111110;
assign LUT_1[64733] = 32'b00000000000000010000110010111010;
assign LUT_1[64734] = 32'b00000000000000010011001111001111;
assign LUT_1[64735] = 32'b00000000000000001100100001001011;
assign LUT_1[64736] = 32'b00000000000000001111011001001111;
assign LUT_1[64737] = 32'b00000000000000001000101011001011;
assign LUT_1[64738] = 32'b00000000000000001011000111100000;
assign LUT_1[64739] = 32'b00000000000000000100011001011100;
assign LUT_1[64740] = 32'b00000000000000010111010010100110;
assign LUT_1[64741] = 32'b00000000000000010000100100100010;
assign LUT_1[64742] = 32'b00000000000000010011000000110111;
assign LUT_1[64743] = 32'b00000000000000001100010010110011;
assign LUT_1[64744] = 32'b00000000000000001110100111000100;
assign LUT_1[64745] = 32'b00000000000000000111111001000000;
assign LUT_1[64746] = 32'b00000000000000001010010101010101;
assign LUT_1[64747] = 32'b00000000000000000011100111010001;
assign LUT_1[64748] = 32'b00000000000000010110100000011011;
assign LUT_1[64749] = 32'b00000000000000001111110010010111;
assign LUT_1[64750] = 32'b00000000000000010010001110101100;
assign LUT_1[64751] = 32'b00000000000000001011100000101000;
assign LUT_1[64752] = 32'b00000000000000010001010100110001;
assign LUT_1[64753] = 32'b00000000000000001010100110101101;
assign LUT_1[64754] = 32'b00000000000000001101000011000010;
assign LUT_1[64755] = 32'b00000000000000000110010100111110;
assign LUT_1[64756] = 32'b00000000000000011001001110001000;
assign LUT_1[64757] = 32'b00000000000000010010100000000100;
assign LUT_1[64758] = 32'b00000000000000010100111100011001;
assign LUT_1[64759] = 32'b00000000000000001110001110010101;
assign LUT_1[64760] = 32'b00000000000000010000100010100110;
assign LUT_1[64761] = 32'b00000000000000001001110100100010;
assign LUT_1[64762] = 32'b00000000000000001100010000110111;
assign LUT_1[64763] = 32'b00000000000000000101100010110011;
assign LUT_1[64764] = 32'b00000000000000011000011011111101;
assign LUT_1[64765] = 32'b00000000000000010001101101111001;
assign LUT_1[64766] = 32'b00000000000000010100001010001110;
assign LUT_1[64767] = 32'b00000000000000001101011100001010;
assign LUT_1[64768] = 32'b00000000000000000111010100110001;
assign LUT_1[64769] = 32'b00000000000000000000100110101101;
assign LUT_1[64770] = 32'b00000000000000000011000011000010;
assign LUT_1[64771] = 32'b11111111111111111100010100111110;
assign LUT_1[64772] = 32'b00000000000000001111001110001000;
assign LUT_1[64773] = 32'b00000000000000001000100000000100;
assign LUT_1[64774] = 32'b00000000000000001010111100011001;
assign LUT_1[64775] = 32'b00000000000000000100001110010101;
assign LUT_1[64776] = 32'b00000000000000000110100010100110;
assign LUT_1[64777] = 32'b11111111111111111111110100100010;
assign LUT_1[64778] = 32'b00000000000000000010010000110111;
assign LUT_1[64779] = 32'b11111111111111111011100010110011;
assign LUT_1[64780] = 32'b00000000000000001110011011111101;
assign LUT_1[64781] = 32'b00000000000000000111101101111001;
assign LUT_1[64782] = 32'b00000000000000001010001010001110;
assign LUT_1[64783] = 32'b00000000000000000011011100001010;
assign LUT_1[64784] = 32'b00000000000000001001010000010011;
assign LUT_1[64785] = 32'b00000000000000000010100010001111;
assign LUT_1[64786] = 32'b00000000000000000100111110100100;
assign LUT_1[64787] = 32'b11111111111111111110010000100000;
assign LUT_1[64788] = 32'b00000000000000010001001001101010;
assign LUT_1[64789] = 32'b00000000000000001010011011100110;
assign LUT_1[64790] = 32'b00000000000000001100110111111011;
assign LUT_1[64791] = 32'b00000000000000000110001001110111;
assign LUT_1[64792] = 32'b00000000000000001000011110001000;
assign LUT_1[64793] = 32'b00000000000000000001110000000100;
assign LUT_1[64794] = 32'b00000000000000000100001100011001;
assign LUT_1[64795] = 32'b11111111111111111101011110010101;
assign LUT_1[64796] = 32'b00000000000000010000010111011111;
assign LUT_1[64797] = 32'b00000000000000001001101001011011;
assign LUT_1[64798] = 32'b00000000000000001100000101110000;
assign LUT_1[64799] = 32'b00000000000000000101010111101100;
assign LUT_1[64800] = 32'b00000000000000001000001111110000;
assign LUT_1[64801] = 32'b00000000000000000001100001101100;
assign LUT_1[64802] = 32'b00000000000000000011111110000001;
assign LUT_1[64803] = 32'b11111111111111111101001111111101;
assign LUT_1[64804] = 32'b00000000000000010000001001000111;
assign LUT_1[64805] = 32'b00000000000000001001011011000011;
assign LUT_1[64806] = 32'b00000000000000001011110111011000;
assign LUT_1[64807] = 32'b00000000000000000101001001010100;
assign LUT_1[64808] = 32'b00000000000000000111011101100101;
assign LUT_1[64809] = 32'b00000000000000000000101111100001;
assign LUT_1[64810] = 32'b00000000000000000011001011110110;
assign LUT_1[64811] = 32'b11111111111111111100011101110010;
assign LUT_1[64812] = 32'b00000000000000001111010110111100;
assign LUT_1[64813] = 32'b00000000000000001000101000111000;
assign LUT_1[64814] = 32'b00000000000000001011000101001101;
assign LUT_1[64815] = 32'b00000000000000000100010111001001;
assign LUT_1[64816] = 32'b00000000000000001010001011010010;
assign LUT_1[64817] = 32'b00000000000000000011011101001110;
assign LUT_1[64818] = 32'b00000000000000000101111001100011;
assign LUT_1[64819] = 32'b11111111111111111111001011011111;
assign LUT_1[64820] = 32'b00000000000000010010000100101001;
assign LUT_1[64821] = 32'b00000000000000001011010110100101;
assign LUT_1[64822] = 32'b00000000000000001101110010111010;
assign LUT_1[64823] = 32'b00000000000000000111000100110110;
assign LUT_1[64824] = 32'b00000000000000001001011001000111;
assign LUT_1[64825] = 32'b00000000000000000010101011000011;
assign LUT_1[64826] = 32'b00000000000000000101000111011000;
assign LUT_1[64827] = 32'b11111111111111111110011001010100;
assign LUT_1[64828] = 32'b00000000000000010001010010011110;
assign LUT_1[64829] = 32'b00000000000000001010100100011010;
assign LUT_1[64830] = 32'b00000000000000001101000000101111;
assign LUT_1[64831] = 32'b00000000000000000110010010101011;
assign LUT_1[64832] = 32'b00000000000000001001010010011001;
assign LUT_1[64833] = 32'b00000000000000000010100100010101;
assign LUT_1[64834] = 32'b00000000000000000101000000101010;
assign LUT_1[64835] = 32'b11111111111111111110010010100110;
assign LUT_1[64836] = 32'b00000000000000010001001011110000;
assign LUT_1[64837] = 32'b00000000000000001010011101101100;
assign LUT_1[64838] = 32'b00000000000000001100111010000001;
assign LUT_1[64839] = 32'b00000000000000000110001011111101;
assign LUT_1[64840] = 32'b00000000000000001000100000001110;
assign LUT_1[64841] = 32'b00000000000000000001110010001010;
assign LUT_1[64842] = 32'b00000000000000000100001110011111;
assign LUT_1[64843] = 32'b11111111111111111101100000011011;
assign LUT_1[64844] = 32'b00000000000000010000011001100101;
assign LUT_1[64845] = 32'b00000000000000001001101011100001;
assign LUT_1[64846] = 32'b00000000000000001100000111110110;
assign LUT_1[64847] = 32'b00000000000000000101011001110010;
assign LUT_1[64848] = 32'b00000000000000001011001101111011;
assign LUT_1[64849] = 32'b00000000000000000100011111110111;
assign LUT_1[64850] = 32'b00000000000000000110111100001100;
assign LUT_1[64851] = 32'b00000000000000000000001110001000;
assign LUT_1[64852] = 32'b00000000000000010011000111010010;
assign LUT_1[64853] = 32'b00000000000000001100011001001110;
assign LUT_1[64854] = 32'b00000000000000001110110101100011;
assign LUT_1[64855] = 32'b00000000000000001000000111011111;
assign LUT_1[64856] = 32'b00000000000000001010011011110000;
assign LUT_1[64857] = 32'b00000000000000000011101101101100;
assign LUT_1[64858] = 32'b00000000000000000110001010000001;
assign LUT_1[64859] = 32'b11111111111111111111011011111101;
assign LUT_1[64860] = 32'b00000000000000010010010101000111;
assign LUT_1[64861] = 32'b00000000000000001011100111000011;
assign LUT_1[64862] = 32'b00000000000000001110000011011000;
assign LUT_1[64863] = 32'b00000000000000000111010101010100;
assign LUT_1[64864] = 32'b00000000000000001010001101011000;
assign LUT_1[64865] = 32'b00000000000000000011011111010100;
assign LUT_1[64866] = 32'b00000000000000000101111011101001;
assign LUT_1[64867] = 32'b11111111111111111111001101100101;
assign LUT_1[64868] = 32'b00000000000000010010000110101111;
assign LUT_1[64869] = 32'b00000000000000001011011000101011;
assign LUT_1[64870] = 32'b00000000000000001101110101000000;
assign LUT_1[64871] = 32'b00000000000000000111000110111100;
assign LUT_1[64872] = 32'b00000000000000001001011011001101;
assign LUT_1[64873] = 32'b00000000000000000010101101001001;
assign LUT_1[64874] = 32'b00000000000000000101001001011110;
assign LUT_1[64875] = 32'b11111111111111111110011011011010;
assign LUT_1[64876] = 32'b00000000000000010001010100100100;
assign LUT_1[64877] = 32'b00000000000000001010100110100000;
assign LUT_1[64878] = 32'b00000000000000001101000010110101;
assign LUT_1[64879] = 32'b00000000000000000110010100110001;
assign LUT_1[64880] = 32'b00000000000000001100001000111010;
assign LUT_1[64881] = 32'b00000000000000000101011010110110;
assign LUT_1[64882] = 32'b00000000000000000111110111001011;
assign LUT_1[64883] = 32'b00000000000000000001001001000111;
assign LUT_1[64884] = 32'b00000000000000010100000010010001;
assign LUT_1[64885] = 32'b00000000000000001101010100001101;
assign LUT_1[64886] = 32'b00000000000000001111110000100010;
assign LUT_1[64887] = 32'b00000000000000001001000010011110;
assign LUT_1[64888] = 32'b00000000000000001011010110101111;
assign LUT_1[64889] = 32'b00000000000000000100101000101011;
assign LUT_1[64890] = 32'b00000000000000000111000101000000;
assign LUT_1[64891] = 32'b00000000000000000000010110111100;
assign LUT_1[64892] = 32'b00000000000000010011010000000110;
assign LUT_1[64893] = 32'b00000000000000001100100010000010;
assign LUT_1[64894] = 32'b00000000000000001110111110010111;
assign LUT_1[64895] = 32'b00000000000000001000010000010011;
assign LUT_1[64896] = 32'b00000000000000001010010100110100;
assign LUT_1[64897] = 32'b00000000000000000011100110110000;
assign LUT_1[64898] = 32'b00000000000000000110000011000101;
assign LUT_1[64899] = 32'b11111111111111111111010101000001;
assign LUT_1[64900] = 32'b00000000000000010010001110001011;
assign LUT_1[64901] = 32'b00000000000000001011100000000111;
assign LUT_1[64902] = 32'b00000000000000001101111100011100;
assign LUT_1[64903] = 32'b00000000000000000111001110011000;
assign LUT_1[64904] = 32'b00000000000000001001100010101001;
assign LUT_1[64905] = 32'b00000000000000000010110100100101;
assign LUT_1[64906] = 32'b00000000000000000101010000111010;
assign LUT_1[64907] = 32'b11111111111111111110100010110110;
assign LUT_1[64908] = 32'b00000000000000010001011100000000;
assign LUT_1[64909] = 32'b00000000000000001010101101111100;
assign LUT_1[64910] = 32'b00000000000000001101001010010001;
assign LUT_1[64911] = 32'b00000000000000000110011100001101;
assign LUT_1[64912] = 32'b00000000000000001100010000010110;
assign LUT_1[64913] = 32'b00000000000000000101100010010010;
assign LUT_1[64914] = 32'b00000000000000000111111110100111;
assign LUT_1[64915] = 32'b00000000000000000001010000100011;
assign LUT_1[64916] = 32'b00000000000000010100001001101101;
assign LUT_1[64917] = 32'b00000000000000001101011011101001;
assign LUT_1[64918] = 32'b00000000000000001111110111111110;
assign LUT_1[64919] = 32'b00000000000000001001001001111010;
assign LUT_1[64920] = 32'b00000000000000001011011110001011;
assign LUT_1[64921] = 32'b00000000000000000100110000000111;
assign LUT_1[64922] = 32'b00000000000000000111001100011100;
assign LUT_1[64923] = 32'b00000000000000000000011110011000;
assign LUT_1[64924] = 32'b00000000000000010011010111100010;
assign LUT_1[64925] = 32'b00000000000000001100101001011110;
assign LUT_1[64926] = 32'b00000000000000001111000101110011;
assign LUT_1[64927] = 32'b00000000000000001000010111101111;
assign LUT_1[64928] = 32'b00000000000000001011001111110011;
assign LUT_1[64929] = 32'b00000000000000000100100001101111;
assign LUT_1[64930] = 32'b00000000000000000110111110000100;
assign LUT_1[64931] = 32'b00000000000000000000010000000000;
assign LUT_1[64932] = 32'b00000000000000010011001001001010;
assign LUT_1[64933] = 32'b00000000000000001100011011000110;
assign LUT_1[64934] = 32'b00000000000000001110110111011011;
assign LUT_1[64935] = 32'b00000000000000001000001001010111;
assign LUT_1[64936] = 32'b00000000000000001010011101101000;
assign LUT_1[64937] = 32'b00000000000000000011101111100100;
assign LUT_1[64938] = 32'b00000000000000000110001011111001;
assign LUT_1[64939] = 32'b11111111111111111111011101110101;
assign LUT_1[64940] = 32'b00000000000000010010010110111111;
assign LUT_1[64941] = 32'b00000000000000001011101000111011;
assign LUT_1[64942] = 32'b00000000000000001110000101010000;
assign LUT_1[64943] = 32'b00000000000000000111010111001100;
assign LUT_1[64944] = 32'b00000000000000001101001011010101;
assign LUT_1[64945] = 32'b00000000000000000110011101010001;
assign LUT_1[64946] = 32'b00000000000000001000111001100110;
assign LUT_1[64947] = 32'b00000000000000000010001011100010;
assign LUT_1[64948] = 32'b00000000000000010101000100101100;
assign LUT_1[64949] = 32'b00000000000000001110010110101000;
assign LUT_1[64950] = 32'b00000000000000010000110010111101;
assign LUT_1[64951] = 32'b00000000000000001010000100111001;
assign LUT_1[64952] = 32'b00000000000000001100011001001010;
assign LUT_1[64953] = 32'b00000000000000000101101011000110;
assign LUT_1[64954] = 32'b00000000000000001000000111011011;
assign LUT_1[64955] = 32'b00000000000000000001011001010111;
assign LUT_1[64956] = 32'b00000000000000010100010010100001;
assign LUT_1[64957] = 32'b00000000000000001101100100011101;
assign LUT_1[64958] = 32'b00000000000000010000000000110010;
assign LUT_1[64959] = 32'b00000000000000001001010010101110;
assign LUT_1[64960] = 32'b00000000000000001100010010011100;
assign LUT_1[64961] = 32'b00000000000000000101100100011000;
assign LUT_1[64962] = 32'b00000000000000001000000000101101;
assign LUT_1[64963] = 32'b00000000000000000001010010101001;
assign LUT_1[64964] = 32'b00000000000000010100001011110011;
assign LUT_1[64965] = 32'b00000000000000001101011101101111;
assign LUT_1[64966] = 32'b00000000000000001111111010000100;
assign LUT_1[64967] = 32'b00000000000000001001001100000000;
assign LUT_1[64968] = 32'b00000000000000001011100000010001;
assign LUT_1[64969] = 32'b00000000000000000100110010001101;
assign LUT_1[64970] = 32'b00000000000000000111001110100010;
assign LUT_1[64971] = 32'b00000000000000000000100000011110;
assign LUT_1[64972] = 32'b00000000000000010011011001101000;
assign LUT_1[64973] = 32'b00000000000000001100101011100100;
assign LUT_1[64974] = 32'b00000000000000001111000111111001;
assign LUT_1[64975] = 32'b00000000000000001000011001110101;
assign LUT_1[64976] = 32'b00000000000000001110001101111110;
assign LUT_1[64977] = 32'b00000000000000000111011111111010;
assign LUT_1[64978] = 32'b00000000000000001001111100001111;
assign LUT_1[64979] = 32'b00000000000000000011001110001011;
assign LUT_1[64980] = 32'b00000000000000010110000111010101;
assign LUT_1[64981] = 32'b00000000000000001111011001010001;
assign LUT_1[64982] = 32'b00000000000000010001110101100110;
assign LUT_1[64983] = 32'b00000000000000001011000111100010;
assign LUT_1[64984] = 32'b00000000000000001101011011110011;
assign LUT_1[64985] = 32'b00000000000000000110101101101111;
assign LUT_1[64986] = 32'b00000000000000001001001010000100;
assign LUT_1[64987] = 32'b00000000000000000010011100000000;
assign LUT_1[64988] = 32'b00000000000000010101010101001010;
assign LUT_1[64989] = 32'b00000000000000001110100111000110;
assign LUT_1[64990] = 32'b00000000000000010001000011011011;
assign LUT_1[64991] = 32'b00000000000000001010010101010111;
assign LUT_1[64992] = 32'b00000000000000001101001101011011;
assign LUT_1[64993] = 32'b00000000000000000110011111010111;
assign LUT_1[64994] = 32'b00000000000000001000111011101100;
assign LUT_1[64995] = 32'b00000000000000000010001101101000;
assign LUT_1[64996] = 32'b00000000000000010101000110110010;
assign LUT_1[64997] = 32'b00000000000000001110011000101110;
assign LUT_1[64998] = 32'b00000000000000010000110101000011;
assign LUT_1[64999] = 32'b00000000000000001010000110111111;
assign LUT_1[65000] = 32'b00000000000000001100011011010000;
assign LUT_1[65001] = 32'b00000000000000000101101101001100;
assign LUT_1[65002] = 32'b00000000000000001000001001100001;
assign LUT_1[65003] = 32'b00000000000000000001011011011101;
assign LUT_1[65004] = 32'b00000000000000010100010100100111;
assign LUT_1[65005] = 32'b00000000000000001101100110100011;
assign LUT_1[65006] = 32'b00000000000000010000000010111000;
assign LUT_1[65007] = 32'b00000000000000001001010100110100;
assign LUT_1[65008] = 32'b00000000000000001111001000111101;
assign LUT_1[65009] = 32'b00000000000000001000011010111001;
assign LUT_1[65010] = 32'b00000000000000001010110111001110;
assign LUT_1[65011] = 32'b00000000000000000100001001001010;
assign LUT_1[65012] = 32'b00000000000000010111000010010100;
assign LUT_1[65013] = 32'b00000000000000010000010100010000;
assign LUT_1[65014] = 32'b00000000000000010010110000100101;
assign LUT_1[65015] = 32'b00000000000000001100000010100001;
assign LUT_1[65016] = 32'b00000000000000001110010110110010;
assign LUT_1[65017] = 32'b00000000000000000111101000101110;
assign LUT_1[65018] = 32'b00000000000000001010000101000011;
assign LUT_1[65019] = 32'b00000000000000000011010110111111;
assign LUT_1[65020] = 32'b00000000000000010110010000001001;
assign LUT_1[65021] = 32'b00000000000000001111100010000101;
assign LUT_1[65022] = 32'b00000000000000010001111110011010;
assign LUT_1[65023] = 32'b00000000000000001011010000010110;
assign LUT_1[65024] = 32'b00000000000000000011001111000010;
assign LUT_1[65025] = 32'b11111111111111111100100000111110;
assign LUT_1[65026] = 32'b11111111111111111110111101010011;
assign LUT_1[65027] = 32'b11111111111111111000001111001111;
assign LUT_1[65028] = 32'b00000000000000001011001000011001;
assign LUT_1[65029] = 32'b00000000000000000100011010010101;
assign LUT_1[65030] = 32'b00000000000000000110110110101010;
assign LUT_1[65031] = 32'b00000000000000000000001000100110;
assign LUT_1[65032] = 32'b00000000000000000010011100110111;
assign LUT_1[65033] = 32'b11111111111111111011101110110011;
assign LUT_1[65034] = 32'b11111111111111111110001011001000;
assign LUT_1[65035] = 32'b11111111111111110111011101000100;
assign LUT_1[65036] = 32'b00000000000000001010010110001110;
assign LUT_1[65037] = 32'b00000000000000000011101000001010;
assign LUT_1[65038] = 32'b00000000000000000110000100011111;
assign LUT_1[65039] = 32'b11111111111111111111010110011011;
assign LUT_1[65040] = 32'b00000000000000000101001010100100;
assign LUT_1[65041] = 32'b11111111111111111110011100100000;
assign LUT_1[65042] = 32'b00000000000000000000111000110101;
assign LUT_1[65043] = 32'b11111111111111111010001010110001;
assign LUT_1[65044] = 32'b00000000000000001101000011111011;
assign LUT_1[65045] = 32'b00000000000000000110010101110111;
assign LUT_1[65046] = 32'b00000000000000001000110010001100;
assign LUT_1[65047] = 32'b00000000000000000010000100001000;
assign LUT_1[65048] = 32'b00000000000000000100011000011001;
assign LUT_1[65049] = 32'b11111111111111111101101010010101;
assign LUT_1[65050] = 32'b00000000000000000000000110101010;
assign LUT_1[65051] = 32'b11111111111111111001011000100110;
assign LUT_1[65052] = 32'b00000000000000001100010001110000;
assign LUT_1[65053] = 32'b00000000000000000101100011101100;
assign LUT_1[65054] = 32'b00000000000000001000000000000001;
assign LUT_1[65055] = 32'b00000000000000000001010001111101;
assign LUT_1[65056] = 32'b00000000000000000100001010000001;
assign LUT_1[65057] = 32'b11111111111111111101011011111101;
assign LUT_1[65058] = 32'b11111111111111111111111000010010;
assign LUT_1[65059] = 32'b11111111111111111001001010001110;
assign LUT_1[65060] = 32'b00000000000000001100000011011000;
assign LUT_1[65061] = 32'b00000000000000000101010101010100;
assign LUT_1[65062] = 32'b00000000000000000111110001101001;
assign LUT_1[65063] = 32'b00000000000000000001000011100101;
assign LUT_1[65064] = 32'b00000000000000000011010111110110;
assign LUT_1[65065] = 32'b11111111111111111100101001110010;
assign LUT_1[65066] = 32'b11111111111111111111000110000111;
assign LUT_1[65067] = 32'b11111111111111111000011000000011;
assign LUT_1[65068] = 32'b00000000000000001011010001001101;
assign LUT_1[65069] = 32'b00000000000000000100100011001001;
assign LUT_1[65070] = 32'b00000000000000000110111111011110;
assign LUT_1[65071] = 32'b00000000000000000000010001011010;
assign LUT_1[65072] = 32'b00000000000000000110000101100011;
assign LUT_1[65073] = 32'b11111111111111111111010111011111;
assign LUT_1[65074] = 32'b00000000000000000001110011110100;
assign LUT_1[65075] = 32'b11111111111111111011000101110000;
assign LUT_1[65076] = 32'b00000000000000001101111110111010;
assign LUT_1[65077] = 32'b00000000000000000111010000110110;
assign LUT_1[65078] = 32'b00000000000000001001101101001011;
assign LUT_1[65079] = 32'b00000000000000000010111111000111;
assign LUT_1[65080] = 32'b00000000000000000101010011011000;
assign LUT_1[65081] = 32'b11111111111111111110100101010100;
assign LUT_1[65082] = 32'b00000000000000000001000001101001;
assign LUT_1[65083] = 32'b11111111111111111010010011100101;
assign LUT_1[65084] = 32'b00000000000000001101001100101111;
assign LUT_1[65085] = 32'b00000000000000000110011110101011;
assign LUT_1[65086] = 32'b00000000000000001000111011000000;
assign LUT_1[65087] = 32'b00000000000000000010001100111100;
assign LUT_1[65088] = 32'b00000000000000000101001100101010;
assign LUT_1[65089] = 32'b11111111111111111110011110100110;
assign LUT_1[65090] = 32'b00000000000000000000111010111011;
assign LUT_1[65091] = 32'b11111111111111111010001100110111;
assign LUT_1[65092] = 32'b00000000000000001101000110000001;
assign LUT_1[65093] = 32'b00000000000000000110010111111101;
assign LUT_1[65094] = 32'b00000000000000001000110100010010;
assign LUT_1[65095] = 32'b00000000000000000010000110001110;
assign LUT_1[65096] = 32'b00000000000000000100011010011111;
assign LUT_1[65097] = 32'b11111111111111111101101100011011;
assign LUT_1[65098] = 32'b00000000000000000000001000110000;
assign LUT_1[65099] = 32'b11111111111111111001011010101100;
assign LUT_1[65100] = 32'b00000000000000001100010011110110;
assign LUT_1[65101] = 32'b00000000000000000101100101110010;
assign LUT_1[65102] = 32'b00000000000000001000000010000111;
assign LUT_1[65103] = 32'b00000000000000000001010100000011;
assign LUT_1[65104] = 32'b00000000000000000111001000001100;
assign LUT_1[65105] = 32'b00000000000000000000011010001000;
assign LUT_1[65106] = 32'b00000000000000000010110110011101;
assign LUT_1[65107] = 32'b11111111111111111100001000011001;
assign LUT_1[65108] = 32'b00000000000000001111000001100011;
assign LUT_1[65109] = 32'b00000000000000001000010011011111;
assign LUT_1[65110] = 32'b00000000000000001010101111110100;
assign LUT_1[65111] = 32'b00000000000000000100000001110000;
assign LUT_1[65112] = 32'b00000000000000000110010110000001;
assign LUT_1[65113] = 32'b11111111111111111111100111111101;
assign LUT_1[65114] = 32'b00000000000000000010000100010010;
assign LUT_1[65115] = 32'b11111111111111111011010110001110;
assign LUT_1[65116] = 32'b00000000000000001110001111011000;
assign LUT_1[65117] = 32'b00000000000000000111100001010100;
assign LUT_1[65118] = 32'b00000000000000001001111101101001;
assign LUT_1[65119] = 32'b00000000000000000011001111100101;
assign LUT_1[65120] = 32'b00000000000000000110000111101001;
assign LUT_1[65121] = 32'b11111111111111111111011001100101;
assign LUT_1[65122] = 32'b00000000000000000001110101111010;
assign LUT_1[65123] = 32'b11111111111111111011000111110110;
assign LUT_1[65124] = 32'b00000000000000001110000001000000;
assign LUT_1[65125] = 32'b00000000000000000111010010111100;
assign LUT_1[65126] = 32'b00000000000000001001101111010001;
assign LUT_1[65127] = 32'b00000000000000000011000001001101;
assign LUT_1[65128] = 32'b00000000000000000101010101011110;
assign LUT_1[65129] = 32'b11111111111111111110100111011010;
assign LUT_1[65130] = 32'b00000000000000000001000011101111;
assign LUT_1[65131] = 32'b11111111111111111010010101101011;
assign LUT_1[65132] = 32'b00000000000000001101001110110101;
assign LUT_1[65133] = 32'b00000000000000000110100000110001;
assign LUT_1[65134] = 32'b00000000000000001000111101000110;
assign LUT_1[65135] = 32'b00000000000000000010001111000010;
assign LUT_1[65136] = 32'b00000000000000001000000011001011;
assign LUT_1[65137] = 32'b00000000000000000001010101000111;
assign LUT_1[65138] = 32'b00000000000000000011110001011100;
assign LUT_1[65139] = 32'b11111111111111111101000011011000;
assign LUT_1[65140] = 32'b00000000000000001111111100100010;
assign LUT_1[65141] = 32'b00000000000000001001001110011110;
assign LUT_1[65142] = 32'b00000000000000001011101010110011;
assign LUT_1[65143] = 32'b00000000000000000100111100101111;
assign LUT_1[65144] = 32'b00000000000000000111010001000000;
assign LUT_1[65145] = 32'b00000000000000000000100010111100;
assign LUT_1[65146] = 32'b00000000000000000010111111010001;
assign LUT_1[65147] = 32'b11111111111111111100010001001101;
assign LUT_1[65148] = 32'b00000000000000001111001010010111;
assign LUT_1[65149] = 32'b00000000000000001000011100010011;
assign LUT_1[65150] = 32'b00000000000000001010111000101000;
assign LUT_1[65151] = 32'b00000000000000000100001010100100;
assign LUT_1[65152] = 32'b00000000000000000110001111000101;
assign LUT_1[65153] = 32'b11111111111111111111100001000001;
assign LUT_1[65154] = 32'b00000000000000000001111101010110;
assign LUT_1[65155] = 32'b11111111111111111011001111010010;
assign LUT_1[65156] = 32'b00000000000000001110001000011100;
assign LUT_1[65157] = 32'b00000000000000000111011010011000;
assign LUT_1[65158] = 32'b00000000000000001001110110101101;
assign LUT_1[65159] = 32'b00000000000000000011001000101001;
assign LUT_1[65160] = 32'b00000000000000000101011100111010;
assign LUT_1[65161] = 32'b11111111111111111110101110110110;
assign LUT_1[65162] = 32'b00000000000000000001001011001011;
assign LUT_1[65163] = 32'b11111111111111111010011101000111;
assign LUT_1[65164] = 32'b00000000000000001101010110010001;
assign LUT_1[65165] = 32'b00000000000000000110101000001101;
assign LUT_1[65166] = 32'b00000000000000001001000100100010;
assign LUT_1[65167] = 32'b00000000000000000010010110011110;
assign LUT_1[65168] = 32'b00000000000000001000001010100111;
assign LUT_1[65169] = 32'b00000000000000000001011100100011;
assign LUT_1[65170] = 32'b00000000000000000011111000111000;
assign LUT_1[65171] = 32'b11111111111111111101001010110100;
assign LUT_1[65172] = 32'b00000000000000010000000011111110;
assign LUT_1[65173] = 32'b00000000000000001001010101111010;
assign LUT_1[65174] = 32'b00000000000000001011110010001111;
assign LUT_1[65175] = 32'b00000000000000000101000100001011;
assign LUT_1[65176] = 32'b00000000000000000111011000011100;
assign LUT_1[65177] = 32'b00000000000000000000101010011000;
assign LUT_1[65178] = 32'b00000000000000000011000110101101;
assign LUT_1[65179] = 32'b11111111111111111100011000101001;
assign LUT_1[65180] = 32'b00000000000000001111010001110011;
assign LUT_1[65181] = 32'b00000000000000001000100011101111;
assign LUT_1[65182] = 32'b00000000000000001011000000000100;
assign LUT_1[65183] = 32'b00000000000000000100010010000000;
assign LUT_1[65184] = 32'b00000000000000000111001010000100;
assign LUT_1[65185] = 32'b00000000000000000000011100000000;
assign LUT_1[65186] = 32'b00000000000000000010111000010101;
assign LUT_1[65187] = 32'b11111111111111111100001010010001;
assign LUT_1[65188] = 32'b00000000000000001111000011011011;
assign LUT_1[65189] = 32'b00000000000000001000010101010111;
assign LUT_1[65190] = 32'b00000000000000001010110001101100;
assign LUT_1[65191] = 32'b00000000000000000100000011101000;
assign LUT_1[65192] = 32'b00000000000000000110010111111001;
assign LUT_1[65193] = 32'b11111111111111111111101001110101;
assign LUT_1[65194] = 32'b00000000000000000010000110001010;
assign LUT_1[65195] = 32'b11111111111111111011011000000110;
assign LUT_1[65196] = 32'b00000000000000001110010001010000;
assign LUT_1[65197] = 32'b00000000000000000111100011001100;
assign LUT_1[65198] = 32'b00000000000000001001111111100001;
assign LUT_1[65199] = 32'b00000000000000000011010001011101;
assign LUT_1[65200] = 32'b00000000000000001001000101100110;
assign LUT_1[65201] = 32'b00000000000000000010010111100010;
assign LUT_1[65202] = 32'b00000000000000000100110011110111;
assign LUT_1[65203] = 32'b11111111111111111110000101110011;
assign LUT_1[65204] = 32'b00000000000000010000111110111101;
assign LUT_1[65205] = 32'b00000000000000001010010000111001;
assign LUT_1[65206] = 32'b00000000000000001100101101001110;
assign LUT_1[65207] = 32'b00000000000000000101111111001010;
assign LUT_1[65208] = 32'b00000000000000001000010011011011;
assign LUT_1[65209] = 32'b00000000000000000001100101010111;
assign LUT_1[65210] = 32'b00000000000000000100000001101100;
assign LUT_1[65211] = 32'b11111111111111111101010011101000;
assign LUT_1[65212] = 32'b00000000000000010000001100110010;
assign LUT_1[65213] = 32'b00000000000000001001011110101110;
assign LUT_1[65214] = 32'b00000000000000001011111011000011;
assign LUT_1[65215] = 32'b00000000000000000101001100111111;
assign LUT_1[65216] = 32'b00000000000000001000001100101101;
assign LUT_1[65217] = 32'b00000000000000000001011110101001;
assign LUT_1[65218] = 32'b00000000000000000011111010111110;
assign LUT_1[65219] = 32'b11111111111111111101001100111010;
assign LUT_1[65220] = 32'b00000000000000010000000110000100;
assign LUT_1[65221] = 32'b00000000000000001001011000000000;
assign LUT_1[65222] = 32'b00000000000000001011110100010101;
assign LUT_1[65223] = 32'b00000000000000000101000110010001;
assign LUT_1[65224] = 32'b00000000000000000111011010100010;
assign LUT_1[65225] = 32'b00000000000000000000101100011110;
assign LUT_1[65226] = 32'b00000000000000000011001000110011;
assign LUT_1[65227] = 32'b11111111111111111100011010101111;
assign LUT_1[65228] = 32'b00000000000000001111010011111001;
assign LUT_1[65229] = 32'b00000000000000001000100101110101;
assign LUT_1[65230] = 32'b00000000000000001011000010001010;
assign LUT_1[65231] = 32'b00000000000000000100010100000110;
assign LUT_1[65232] = 32'b00000000000000001010001000001111;
assign LUT_1[65233] = 32'b00000000000000000011011010001011;
assign LUT_1[65234] = 32'b00000000000000000101110110100000;
assign LUT_1[65235] = 32'b11111111111111111111001000011100;
assign LUT_1[65236] = 32'b00000000000000010010000001100110;
assign LUT_1[65237] = 32'b00000000000000001011010011100010;
assign LUT_1[65238] = 32'b00000000000000001101101111110111;
assign LUT_1[65239] = 32'b00000000000000000111000001110011;
assign LUT_1[65240] = 32'b00000000000000001001010110000100;
assign LUT_1[65241] = 32'b00000000000000000010101000000000;
assign LUT_1[65242] = 32'b00000000000000000101000100010101;
assign LUT_1[65243] = 32'b11111111111111111110010110010001;
assign LUT_1[65244] = 32'b00000000000000010001001111011011;
assign LUT_1[65245] = 32'b00000000000000001010100001010111;
assign LUT_1[65246] = 32'b00000000000000001100111101101100;
assign LUT_1[65247] = 32'b00000000000000000110001111101000;
assign LUT_1[65248] = 32'b00000000000000001001000111101100;
assign LUT_1[65249] = 32'b00000000000000000010011001101000;
assign LUT_1[65250] = 32'b00000000000000000100110101111101;
assign LUT_1[65251] = 32'b11111111111111111110000111111001;
assign LUT_1[65252] = 32'b00000000000000010001000001000011;
assign LUT_1[65253] = 32'b00000000000000001010010010111111;
assign LUT_1[65254] = 32'b00000000000000001100101111010100;
assign LUT_1[65255] = 32'b00000000000000000110000001010000;
assign LUT_1[65256] = 32'b00000000000000001000010101100001;
assign LUT_1[65257] = 32'b00000000000000000001100111011101;
assign LUT_1[65258] = 32'b00000000000000000100000011110010;
assign LUT_1[65259] = 32'b11111111111111111101010101101110;
assign LUT_1[65260] = 32'b00000000000000010000001110111000;
assign LUT_1[65261] = 32'b00000000000000001001100000110100;
assign LUT_1[65262] = 32'b00000000000000001011111101001001;
assign LUT_1[65263] = 32'b00000000000000000101001111000101;
assign LUT_1[65264] = 32'b00000000000000001011000011001110;
assign LUT_1[65265] = 32'b00000000000000000100010101001010;
assign LUT_1[65266] = 32'b00000000000000000110110001011111;
assign LUT_1[65267] = 32'b00000000000000000000000011011011;
assign LUT_1[65268] = 32'b00000000000000010010111100100101;
assign LUT_1[65269] = 32'b00000000000000001100001110100001;
assign LUT_1[65270] = 32'b00000000000000001110101010110110;
assign LUT_1[65271] = 32'b00000000000000000111111100110010;
assign LUT_1[65272] = 32'b00000000000000001010010001000011;
assign LUT_1[65273] = 32'b00000000000000000011100010111111;
assign LUT_1[65274] = 32'b00000000000000000101111111010100;
assign LUT_1[65275] = 32'b11111111111111111111010001010000;
assign LUT_1[65276] = 32'b00000000000000010010001010011010;
assign LUT_1[65277] = 32'b00000000000000001011011100010110;
assign LUT_1[65278] = 32'b00000000000000001101111000101011;
assign LUT_1[65279] = 32'b00000000000000000111001010100111;
assign LUT_1[65280] = 32'b00000000000000000001000011001110;
assign LUT_1[65281] = 32'b11111111111111111010010101001010;
assign LUT_1[65282] = 32'b11111111111111111100110001011111;
assign LUT_1[65283] = 32'b11111111111111110110000011011011;
assign LUT_1[65284] = 32'b00000000000000001000111100100101;
assign LUT_1[65285] = 32'b00000000000000000010001110100001;
assign LUT_1[65286] = 32'b00000000000000000100101010110110;
assign LUT_1[65287] = 32'b11111111111111111101111100110010;
assign LUT_1[65288] = 32'b00000000000000000000010001000011;
assign LUT_1[65289] = 32'b11111111111111111001100010111111;
assign LUT_1[65290] = 32'b11111111111111111011111111010100;
assign LUT_1[65291] = 32'b11111111111111110101010001010000;
assign LUT_1[65292] = 32'b00000000000000001000001010011010;
assign LUT_1[65293] = 32'b00000000000000000001011100010110;
assign LUT_1[65294] = 32'b00000000000000000011111000101011;
assign LUT_1[65295] = 32'b11111111111111111101001010100111;
assign LUT_1[65296] = 32'b00000000000000000010111110110000;
assign LUT_1[65297] = 32'b11111111111111111100010000101100;
assign LUT_1[65298] = 32'b11111111111111111110101101000001;
assign LUT_1[65299] = 32'b11111111111111110111111110111101;
assign LUT_1[65300] = 32'b00000000000000001010111000000111;
assign LUT_1[65301] = 32'b00000000000000000100001010000011;
assign LUT_1[65302] = 32'b00000000000000000110100110011000;
assign LUT_1[65303] = 32'b11111111111111111111111000010100;
assign LUT_1[65304] = 32'b00000000000000000010001100100101;
assign LUT_1[65305] = 32'b11111111111111111011011110100001;
assign LUT_1[65306] = 32'b11111111111111111101111010110110;
assign LUT_1[65307] = 32'b11111111111111110111001100110010;
assign LUT_1[65308] = 32'b00000000000000001010000101111100;
assign LUT_1[65309] = 32'b00000000000000000011010111111000;
assign LUT_1[65310] = 32'b00000000000000000101110100001101;
assign LUT_1[65311] = 32'b11111111111111111111000110001001;
assign LUT_1[65312] = 32'b00000000000000000001111110001101;
assign LUT_1[65313] = 32'b11111111111111111011010000001001;
assign LUT_1[65314] = 32'b11111111111111111101101100011110;
assign LUT_1[65315] = 32'b11111111111111110110111110011010;
assign LUT_1[65316] = 32'b00000000000000001001110111100100;
assign LUT_1[65317] = 32'b00000000000000000011001001100000;
assign LUT_1[65318] = 32'b00000000000000000101100101110101;
assign LUT_1[65319] = 32'b11111111111111111110110111110001;
assign LUT_1[65320] = 32'b00000000000000000001001100000010;
assign LUT_1[65321] = 32'b11111111111111111010011101111110;
assign LUT_1[65322] = 32'b11111111111111111100111010010011;
assign LUT_1[65323] = 32'b11111111111111110110001100001111;
assign LUT_1[65324] = 32'b00000000000000001001000101011001;
assign LUT_1[65325] = 32'b00000000000000000010010111010101;
assign LUT_1[65326] = 32'b00000000000000000100110011101010;
assign LUT_1[65327] = 32'b11111111111111111110000101100110;
assign LUT_1[65328] = 32'b00000000000000000011111001101111;
assign LUT_1[65329] = 32'b11111111111111111101001011101011;
assign LUT_1[65330] = 32'b11111111111111111111101000000000;
assign LUT_1[65331] = 32'b11111111111111111000111001111100;
assign LUT_1[65332] = 32'b00000000000000001011110011000110;
assign LUT_1[65333] = 32'b00000000000000000101000101000010;
assign LUT_1[65334] = 32'b00000000000000000111100001010111;
assign LUT_1[65335] = 32'b00000000000000000000110011010011;
assign LUT_1[65336] = 32'b00000000000000000011000111100100;
assign LUT_1[65337] = 32'b11111111111111111100011001100000;
assign LUT_1[65338] = 32'b11111111111111111110110101110101;
assign LUT_1[65339] = 32'b11111111111111111000000111110001;
assign LUT_1[65340] = 32'b00000000000000001011000000111011;
assign LUT_1[65341] = 32'b00000000000000000100010010110111;
assign LUT_1[65342] = 32'b00000000000000000110101111001100;
assign LUT_1[65343] = 32'b00000000000000000000000001001000;
assign LUT_1[65344] = 32'b00000000000000000011000000110110;
assign LUT_1[65345] = 32'b11111111111111111100010010110010;
assign LUT_1[65346] = 32'b11111111111111111110101111000111;
assign LUT_1[65347] = 32'b11111111111111111000000001000011;
assign LUT_1[65348] = 32'b00000000000000001010111010001101;
assign LUT_1[65349] = 32'b00000000000000000100001100001001;
assign LUT_1[65350] = 32'b00000000000000000110101000011110;
assign LUT_1[65351] = 32'b11111111111111111111111010011010;
assign LUT_1[65352] = 32'b00000000000000000010001110101011;
assign LUT_1[65353] = 32'b11111111111111111011100000100111;
assign LUT_1[65354] = 32'b11111111111111111101111100111100;
assign LUT_1[65355] = 32'b11111111111111110111001110111000;
assign LUT_1[65356] = 32'b00000000000000001010001000000010;
assign LUT_1[65357] = 32'b00000000000000000011011001111110;
assign LUT_1[65358] = 32'b00000000000000000101110110010011;
assign LUT_1[65359] = 32'b11111111111111111111001000001111;
assign LUT_1[65360] = 32'b00000000000000000100111100011000;
assign LUT_1[65361] = 32'b11111111111111111110001110010100;
assign LUT_1[65362] = 32'b00000000000000000000101010101001;
assign LUT_1[65363] = 32'b11111111111111111001111100100101;
assign LUT_1[65364] = 32'b00000000000000001100110101101111;
assign LUT_1[65365] = 32'b00000000000000000110000111101011;
assign LUT_1[65366] = 32'b00000000000000001000100100000000;
assign LUT_1[65367] = 32'b00000000000000000001110101111100;
assign LUT_1[65368] = 32'b00000000000000000100001010001101;
assign LUT_1[65369] = 32'b11111111111111111101011100001001;
assign LUT_1[65370] = 32'b11111111111111111111111000011110;
assign LUT_1[65371] = 32'b11111111111111111001001010011010;
assign LUT_1[65372] = 32'b00000000000000001100000011100100;
assign LUT_1[65373] = 32'b00000000000000000101010101100000;
assign LUT_1[65374] = 32'b00000000000000000111110001110101;
assign LUT_1[65375] = 32'b00000000000000000001000011110001;
assign LUT_1[65376] = 32'b00000000000000000011111011110101;
assign LUT_1[65377] = 32'b11111111111111111101001101110001;
assign LUT_1[65378] = 32'b11111111111111111111101010000110;
assign LUT_1[65379] = 32'b11111111111111111000111100000010;
assign LUT_1[65380] = 32'b00000000000000001011110101001100;
assign LUT_1[65381] = 32'b00000000000000000101000111001000;
assign LUT_1[65382] = 32'b00000000000000000111100011011101;
assign LUT_1[65383] = 32'b00000000000000000000110101011001;
assign LUT_1[65384] = 32'b00000000000000000011001001101010;
assign LUT_1[65385] = 32'b11111111111111111100011011100110;
assign LUT_1[65386] = 32'b11111111111111111110110111111011;
assign LUT_1[65387] = 32'b11111111111111111000001001110111;
assign LUT_1[65388] = 32'b00000000000000001011000011000001;
assign LUT_1[65389] = 32'b00000000000000000100010100111101;
assign LUT_1[65390] = 32'b00000000000000000110110001010010;
assign LUT_1[65391] = 32'b00000000000000000000000011001110;
assign LUT_1[65392] = 32'b00000000000000000101110111010111;
assign LUT_1[65393] = 32'b11111111111111111111001001010011;
assign LUT_1[65394] = 32'b00000000000000000001100101101000;
assign LUT_1[65395] = 32'b11111111111111111010110111100100;
assign LUT_1[65396] = 32'b00000000000000001101110000101110;
assign LUT_1[65397] = 32'b00000000000000000111000010101010;
assign LUT_1[65398] = 32'b00000000000000001001011110111111;
assign LUT_1[65399] = 32'b00000000000000000010110000111011;
assign LUT_1[65400] = 32'b00000000000000000101000101001100;
assign LUT_1[65401] = 32'b11111111111111111110010111001000;
assign LUT_1[65402] = 32'b00000000000000000000110011011101;
assign LUT_1[65403] = 32'b11111111111111111010000101011001;
assign LUT_1[65404] = 32'b00000000000000001100111110100011;
assign LUT_1[65405] = 32'b00000000000000000110010000011111;
assign LUT_1[65406] = 32'b00000000000000001000101100110100;
assign LUT_1[65407] = 32'b00000000000000000001111110110000;
assign LUT_1[65408] = 32'b00000000000000000100000011010001;
assign LUT_1[65409] = 32'b11111111111111111101010101001101;
assign LUT_1[65410] = 32'b11111111111111111111110001100010;
assign LUT_1[65411] = 32'b11111111111111111001000011011110;
assign LUT_1[65412] = 32'b00000000000000001011111100101000;
assign LUT_1[65413] = 32'b00000000000000000101001110100100;
assign LUT_1[65414] = 32'b00000000000000000111101010111001;
assign LUT_1[65415] = 32'b00000000000000000000111100110101;
assign LUT_1[65416] = 32'b00000000000000000011010001000110;
assign LUT_1[65417] = 32'b11111111111111111100100011000010;
assign LUT_1[65418] = 32'b11111111111111111110111111010111;
assign LUT_1[65419] = 32'b11111111111111111000010001010011;
assign LUT_1[65420] = 32'b00000000000000001011001010011101;
assign LUT_1[65421] = 32'b00000000000000000100011100011001;
assign LUT_1[65422] = 32'b00000000000000000110111000101110;
assign LUT_1[65423] = 32'b00000000000000000000001010101010;
assign LUT_1[65424] = 32'b00000000000000000101111110110011;
assign LUT_1[65425] = 32'b11111111111111111111010000101111;
assign LUT_1[65426] = 32'b00000000000000000001101101000100;
assign LUT_1[65427] = 32'b11111111111111111010111111000000;
assign LUT_1[65428] = 32'b00000000000000001101111000001010;
assign LUT_1[65429] = 32'b00000000000000000111001010000110;
assign LUT_1[65430] = 32'b00000000000000001001100110011011;
assign LUT_1[65431] = 32'b00000000000000000010111000010111;
assign LUT_1[65432] = 32'b00000000000000000101001100101000;
assign LUT_1[65433] = 32'b11111111111111111110011110100100;
assign LUT_1[65434] = 32'b00000000000000000000111010111001;
assign LUT_1[65435] = 32'b11111111111111111010001100110101;
assign LUT_1[65436] = 32'b00000000000000001101000101111111;
assign LUT_1[65437] = 32'b00000000000000000110010111111011;
assign LUT_1[65438] = 32'b00000000000000001000110100010000;
assign LUT_1[65439] = 32'b00000000000000000010000110001100;
assign LUT_1[65440] = 32'b00000000000000000100111110010000;
assign LUT_1[65441] = 32'b11111111111111111110010000001100;
assign LUT_1[65442] = 32'b00000000000000000000101100100001;
assign LUT_1[65443] = 32'b11111111111111111001111110011101;
assign LUT_1[65444] = 32'b00000000000000001100110111100111;
assign LUT_1[65445] = 32'b00000000000000000110001001100011;
assign LUT_1[65446] = 32'b00000000000000001000100101111000;
assign LUT_1[65447] = 32'b00000000000000000001110111110100;
assign LUT_1[65448] = 32'b00000000000000000100001100000101;
assign LUT_1[65449] = 32'b11111111111111111101011110000001;
assign LUT_1[65450] = 32'b11111111111111111111111010010110;
assign LUT_1[65451] = 32'b11111111111111111001001100010010;
assign LUT_1[65452] = 32'b00000000000000001100000101011100;
assign LUT_1[65453] = 32'b00000000000000000101010111011000;
assign LUT_1[65454] = 32'b00000000000000000111110011101101;
assign LUT_1[65455] = 32'b00000000000000000001000101101001;
assign LUT_1[65456] = 32'b00000000000000000110111001110010;
assign LUT_1[65457] = 32'b00000000000000000000001011101110;
assign LUT_1[65458] = 32'b00000000000000000010101000000011;
assign LUT_1[65459] = 32'b11111111111111111011111001111111;
assign LUT_1[65460] = 32'b00000000000000001110110011001001;
assign LUT_1[65461] = 32'b00000000000000001000000101000101;
assign LUT_1[65462] = 32'b00000000000000001010100001011010;
assign LUT_1[65463] = 32'b00000000000000000011110011010110;
assign LUT_1[65464] = 32'b00000000000000000110000111100111;
assign LUT_1[65465] = 32'b11111111111111111111011001100011;
assign LUT_1[65466] = 32'b00000000000000000001110101111000;
assign LUT_1[65467] = 32'b11111111111111111011000111110100;
assign LUT_1[65468] = 32'b00000000000000001110000000111110;
assign LUT_1[65469] = 32'b00000000000000000111010010111010;
assign LUT_1[65470] = 32'b00000000000000001001101111001111;
assign LUT_1[65471] = 32'b00000000000000000011000001001011;
assign LUT_1[65472] = 32'b00000000000000000110000000111001;
assign LUT_1[65473] = 32'b11111111111111111111010010110101;
assign LUT_1[65474] = 32'b00000000000000000001101111001010;
assign LUT_1[65475] = 32'b11111111111111111011000001000110;
assign LUT_1[65476] = 32'b00000000000000001101111010010000;
assign LUT_1[65477] = 32'b00000000000000000111001100001100;
assign LUT_1[65478] = 32'b00000000000000001001101000100001;
assign LUT_1[65479] = 32'b00000000000000000010111010011101;
assign LUT_1[65480] = 32'b00000000000000000101001110101110;
assign LUT_1[65481] = 32'b11111111111111111110100000101010;
assign LUT_1[65482] = 32'b00000000000000000000111100111111;
assign LUT_1[65483] = 32'b11111111111111111010001110111011;
assign LUT_1[65484] = 32'b00000000000000001101001000000101;
assign LUT_1[65485] = 32'b00000000000000000110011010000001;
assign LUT_1[65486] = 32'b00000000000000001000110110010110;
assign LUT_1[65487] = 32'b00000000000000000010001000010010;
assign LUT_1[65488] = 32'b00000000000000000111111100011011;
assign LUT_1[65489] = 32'b00000000000000000001001110010111;
assign LUT_1[65490] = 32'b00000000000000000011101010101100;
assign LUT_1[65491] = 32'b11111111111111111100111100101000;
assign LUT_1[65492] = 32'b00000000000000001111110101110010;
assign LUT_1[65493] = 32'b00000000000000001001000111101110;
assign LUT_1[65494] = 32'b00000000000000001011100100000011;
assign LUT_1[65495] = 32'b00000000000000000100110101111111;
assign LUT_1[65496] = 32'b00000000000000000111001010010000;
assign LUT_1[65497] = 32'b00000000000000000000011100001100;
assign LUT_1[65498] = 32'b00000000000000000010111000100001;
assign LUT_1[65499] = 32'b11111111111111111100001010011101;
assign LUT_1[65500] = 32'b00000000000000001111000011100111;
assign LUT_1[65501] = 32'b00000000000000001000010101100011;
assign LUT_1[65502] = 32'b00000000000000001010110001111000;
assign LUT_1[65503] = 32'b00000000000000000100000011110100;
assign LUT_1[65504] = 32'b00000000000000000110111011111000;
assign LUT_1[65505] = 32'b00000000000000000000001101110100;
assign LUT_1[65506] = 32'b00000000000000000010101010001001;
assign LUT_1[65507] = 32'b11111111111111111011111100000101;
assign LUT_1[65508] = 32'b00000000000000001110110101001111;
assign LUT_1[65509] = 32'b00000000000000001000000111001011;
assign LUT_1[65510] = 32'b00000000000000001010100011100000;
assign LUT_1[65511] = 32'b00000000000000000011110101011100;
assign LUT_1[65512] = 32'b00000000000000000110001001101101;
assign LUT_1[65513] = 32'b11111111111111111111011011101001;
assign LUT_1[65514] = 32'b00000000000000000001110111111110;
assign LUT_1[65515] = 32'b11111111111111111011001001111010;
assign LUT_1[65516] = 32'b00000000000000001110000011000100;
assign LUT_1[65517] = 32'b00000000000000000111010101000000;
assign LUT_1[65518] = 32'b00000000000000001001110001010101;
assign LUT_1[65519] = 32'b00000000000000000011000011010001;
assign LUT_1[65520] = 32'b00000000000000001000110111011010;
assign LUT_1[65521] = 32'b00000000000000000010001001010110;
assign LUT_1[65522] = 32'b00000000000000000100100101101011;
assign LUT_1[65523] = 32'b11111111111111111101110111100111;
assign LUT_1[65524] = 32'b00000000000000010000110000110001;
assign LUT_1[65525] = 32'b00000000000000001010000010101101;
assign LUT_1[65526] = 32'b00000000000000001100011111000010;
assign LUT_1[65527] = 32'b00000000000000000101110000111110;
assign LUT_1[65528] = 32'b00000000000000001000000101001111;
assign LUT_1[65529] = 32'b00000000000000000001010111001011;
assign LUT_1[65530] = 32'b00000000000000000011110011100000;
assign LUT_1[65531] = 32'b11111111111111111101000101011100;
assign LUT_1[65532] = 32'b00000000000000001111111110100110;
assign LUT_1[65533] = 32'b00000000000000001001010000100010;
assign LUT_1[65534] = 32'b00000000000000001011101100110111;
assign LUT_1[65535] = 32'b00000000000000000100111110110011;
endmodule
